module top (out,n29,n31,n38,n42,n48,n56,n57,n66,n73
        ,n78,n87,n88,n95,n104,n115,n116,n120,n126,n136
        ,n137,n142,n147,n152,n177,n184,n194,n215,n217,n222
        ,n231,n237,n238,n242,n248,n256,n257,n263,n277,n289
        ,n297,n305,n312,n313,n320,n332,n340,n349,n356,n396
        ,n404,n419,n441,n1343,n1359,n1375,n1381,n1392,n1547,n1554
        ,n1561,n1568,n1575,n1581,n1583,n1596,n1614,n1624,n1625,n1627
        ,n1628,n1630,n1631,n1633,n1634,n1636,n1637,n1640);
output out;
input n29;
input n31;
input n38;
input n42;
input n48;
input n56;
input n57;
input n66;
input n73;
input n78;
input n87;
input n88;
input n95;
input n104;
input n115;
input n116;
input n120;
input n126;
input n136;
input n137;
input n142;
input n147;
input n152;
input n177;
input n184;
input n194;
input n215;
input n217;
input n222;
input n231;
input n237;
input n238;
input n242;
input n248;
input n256;
input n257;
input n263;
input n277;
input n289;
input n297;
input n305;
input n312;
input n313;
input n320;
input n332;
input n340;
input n349;
input n356;
input n396;
input n404;
input n419;
input n441;
input n1343;
input n1359;
input n1375;
input n1381;
input n1392;
input n1547;
input n1554;
input n1561;
input n1568;
input n1575;
input n1581;
input n1583;
input n1596;
input n1614;
input n1624;
input n1625;
input n1627;
input n1628;
input n1630;
input n1631;
input n1633;
input n1634;
input n1636;
input n1637;
input n1640;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n239;
wire n240;
wire n241;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1582;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1626;
wire n1629;
wire n1632;
wire n1635;
wire n1638;
wire n1639;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
xor (out,n0,n1642);
nand (n0,n1,n1638);
or (n1,n2,n1618);
not (n2,n3);
nand (n3,n4,n1617);
or (n4,n5,n1346);
not (n5,n6);
or (n6,n7,n1344);
nor (n7,n8,n1343);
not (n8,n9);
nand (n9,n10,n1342);
or (n10,n11,n896);
not (n11,n12);
nand (n12,n13,n895);
or (n13,n14,n771);
xor (n14,n15,n686);
xor (n15,n16,n446);
xor (n16,n17,n360);
xor (n17,n18,n197);
xor (n18,n19,n159);
xor (n19,n20,n108);
or (n20,n21,n107);
and (n21,n22,n81);
xor (n22,n23,n50);
nand (n23,n24,n44);
or (n24,n25,n33);
not (n25,n26);
nor (n26,n27,n32);
and (n27,n28,n30);
not (n28,n29);
not (n30,n31);
and (n32,n31,n29);
not (n33,n34);
nor (n34,n35,n40);
nor (n35,n36,n39);
and (n36,n29,n37);
not (n37,n38);
nor (n39,n37,n29);
nand (n40,n41,n43);
or (n41,n37,n42);
nand (n43,n37,n42);
nand (n44,n45,n40);
nand (n45,n46,n49);
or (n46,n29,n47);
not (n47,n48);
nand (n49,n47,n29);
nand (n50,n51,n75);
or (n51,n52,n61);
not (n52,n53);
nand (n53,n54,n58);
not (n54,n55);
and (n55,n56,n57);
nand (n58,n59,n60);
not (n59,n57);
not (n60,n56);
nand (n61,n62,n69);
or (n62,n63,n67);
not (n63,n64);
nand (n64,n65,n57);
not (n65,n66);
not (n67,n68);
nand (n68,n59,n66);
not (n69,n70);
nand (n70,n71,n74);
or (n71,n72,n66);
not (n72,n73);
nand (n74,n72,n66);
nand (n75,n76,n70);
nand (n76,n77,n79);
or (n77,n57,n78);
not (n79,n80);
and (n80,n78,n57);
nand (n81,n82,n101);
or (n82,n83,n91);
not (n83,n84);
nor (n84,n85,n89);
and (n85,n86,n88);
not (n86,n87);
and (n89,n87,n90);
not (n90,n88);
not (n91,n92);
nor (n92,n93,n97);
nand (n93,n94,n96);
or (n94,n59,n95);
nand (n96,n59,n95);
nor (n97,n98,n99);
and (n98,n86,n95);
and (n99,n87,n100);
not (n100,n95);
nand (n101,n102,n93);
nand (n102,n103,n105);
or (n103,n104,n87);
not (n105,n106);
and (n106,n104,n87);
and (n107,n23,n50);
or (n108,n109,n158);
and (n109,n110,n154);
xor (n110,n111,n129);
nand (n111,n112,n123);
or (n112,n113,n117);
nand (n113,n114,n116);
not (n114,n115);
nor (n117,n118,n121);
and (n118,n119,n120);
not (n119,n116);
and (n121,n116,n122);
not (n122,n120);
or (n123,n124,n114);
nor (n124,n125,n127);
and (n125,n119,n126);
and (n127,n116,n128);
not (n128,n126);
nand (n129,n130,n149);
or (n130,n131,n144);
nand (n131,n132,n139);
not (n132,n133);
nand (n133,n134,n138);
or (n134,n135,n137);
not (n135,n136);
nand (n138,n135,n137);
nand (n139,n140,n143);
or (n140,n136,n141);
not (n141,n142);
nand (n143,n141,n136);
nor (n144,n145,n148);
and (n145,n146,n142);
not (n146,n147);
and (n148,n147,n141);
nand (n149,n150,n133);
nand (n150,n151,n153);
or (n151,n152,n141);
nand (n153,n141,n152);
nor (n154,n155,n157);
not (n155,n156);
and (n156,n40,n31);
nand (n157,n93,n88);
and (n158,n111,n129);
or (n159,n160,n196);
and (n160,n161,n172);
xor (n161,n162,n167);
nor (n162,n163,n28);
nor (n163,n164,n166);
nor (n164,n165,n42);
and (n165,n31,n38);
nor (n166,n31,n38);
and (n167,n168,n86);
nand (n168,n169,n170);
or (n169,n100,n88);
nand (n170,n171,n57);
or (n171,n90,n95);
nand (n172,n173,n187);
or (n173,n174,n181);
not (n174,n175);
nand (n175,n176,n179);
or (n176,n177,n178);
not (n178,n137);
or (n179,n137,n180);
not (n180,n177);
not (n181,n182);
nand (n182,n183,n185);
nand (n183,n184,n116,n178);
nand (n185,n186,n119,n137);
not (n186,n184);
nand (n187,n188,n191);
nand (n188,n189,n190);
or (n189,n186,n116);
nand (n190,n186,n116);
nand (n191,n192,n195);
or (n192,n193,n137);
not (n193,n194);
nand (n195,n137,n193);
and (n196,n162,n167);
xor (n197,n198,n281);
xor (n198,n199,n207);
nand (n199,n200,n202);
or (n200,n131,n201);
not (n201,n150);
or (n202,n132,n203);
not (n203,n204);
nand (n204,n205,n206);
or (n205,n180,n142);
nand (n206,n142,n180);
or (n207,n208,n280);
and (n208,n209,n251);
xor (n209,n210,n233);
nand (n210,n211,n228);
or (n211,n212,n219);
not (n212,n213);
nand (n213,n214,n218);
or (n214,n215,n216);
not (n216,n217);
nand (n218,n216,n215);
nand (n219,n220,n224);
nand (n220,n221,n223);
or (n221,n222,n216);
nand (n223,n216,n222);
not (n224,n225);
nand (n225,n226,n227);
or (n226,n141,n222);
nand (n227,n141,n222);
nand (n228,n225,n229);
nand (n229,n230,n232);
or (n230,n231,n216);
nand (n232,n216,n231);
nand (n233,n234,n245);
or (n234,n235,n239);
nand (n235,n236,n238);
not (n236,n237);
not (n239,n240);
nand (n240,n241,n243);
or (n241,n242,n238);
not (n243,n244);
and (n244,n242,n238);
nand (n245,n246,n237);
nand (n246,n247,n249);
or (n247,n248,n238);
not (n249,n250);
and (n250,n248,n238);
nand (n251,n252,n266);
or (n252,n253,n260);
not (n253,n254);
nand (n254,n255,n258);
or (n255,n256,n257);
not (n258,n259);
and (n259,n256,n257);
nor (n260,n261,n264);
and (n261,n262,n263);
not (n262,n238);
and (n264,n238,n265);
not (n265,n263);
or (n266,n267,n274);
nand (n267,n268,n260);
or (n268,n269,n272);
not (n269,n270);
nand (n270,n271,n263);
not (n271,n257);
not (n272,n273);
nand (n273,n257,n265);
not (n274,n275);
nand (n275,n276,n278);
or (n276,n277,n257);
not (n278,n279);
and (n279,n277,n257);
and (n280,n210,n233);
or (n281,n282,n359);
and (n282,n283,n334);
xor (n283,n284,n307);
nand (n284,n285,n302);
or (n285,n286,n293);
not (n286,n287);
nand (n287,n288,n291);
or (n288,n289,n290);
not (n290,n42);
or (n291,n292,n42);
not (n292,n289);
nand (n293,n294,n299);
not (n294,n295);
nand (n295,n296,n298);
or (n296,n216,n297);
nand (n298,n216,n297);
nand (n299,n300,n301);
or (n300,n297,n290);
nand (n301,n290,n297);
nand (n302,n295,n303);
nand (n303,n304,n306);
or (n304,n305,n290);
nand (n306,n290,n305);
nand (n307,n308,n326);
or (n308,n309,n316);
not (n309,n310);
nand (n310,n311,n314);
or (n311,n312,n313);
not (n314,n315);
and (n315,n312,n313);
nand (n316,n317,n322);
not (n317,n318);
nand (n318,n319,n321);
or (n319,n320,n271);
nand (n321,n271,n320);
nand (n322,n323,n325);
or (n323,n324,n313);
not (n324,n320);
nand (n325,n313,n324);
nand (n326,n327,n318);
not (n327,n328);
nor (n328,n329,n333);
and (n329,n330,n331);
not (n330,n313);
not (n331,n332);
and (n333,n313,n332);
nand (n334,n335,n352);
or (n335,n336,n345);
nand (n336,n337,n342);
not (n337,n338);
nand (n338,n339,n341);
or (n339,n330,n340);
nand (n341,n330,n340);
nand (n342,n343,n344);
or (n343,n340,n72);
nand (n344,n72,n340);
not (n345,n346);
nand (n346,n347,n350);
not (n347,n348);
and (n348,n349,n73);
nand (n350,n72,n351);
not (n351,n349);
or (n352,n337,n353);
not (n353,n354);
nor (n354,n355,n357);
and (n355,n356,n72);
and (n357,n358,n73);
not (n358,n356);
and (n359,n284,n307);
xor (n360,n361,n420);
xor (n361,n362,n387);
xor (n362,n363,n379);
xor (n363,n364,n372);
nand (n364,n365,n366);
or (n365,n353,n336);
nand (n366,n338,n367);
nand (n367,n368,n370);
not (n368,n369);
and (n369,n312,n73);
nand (n370,n72,n371);
not (n371,n312);
nand (n372,n373,n375);
or (n373,n374,n33);
not (n374,n45);
nand (n375,n376,n40);
nor (n376,n377,n378);
and (n377,n28,n292);
and (n378,n29,n289);
nand (n379,n380,n382);
or (n380,n381,n61);
not (n381,n76);
nand (n382,n70,n383);
nand (n383,n384,n385);
or (n384,n57,n349);
not (n385,n386);
and (n386,n349,n57);
xor (n387,n388,n415);
xor (n388,n389,n407);
nand (n389,n390,n406);
or (n390,n391,n399);
not (n391,n392);
nand (n392,n88,n393);
not (n393,n394);
nor (n394,n395,n397);
and (n395,n86,n396);
and (n397,n87,n398);
not (n398,n396);
nand (n399,n400,n31);
not (n400,n401);
nor (n401,n402,n405);
and (n402,n29,n403);
not (n403,n404);
and (n405,n28,n404);
nand (n406,n391,n399);
nand (n407,n408,n410);
or (n408,n91,n409);
not (n409,n102);
or (n410,n411,n412);
not (n411,n93);
nor (n412,n413,n414);
and (n413,n86,n60);
and (n414,n87,n56);
nand (n415,n416,n417);
or (n416,n113,n124);
or (n417,n418,n114);
xnor (n418,n419,n116);
xor (n420,n421,n436);
xor (n421,n422,n429);
nand (n422,n423,n425);
or (n423,n424,n181);
not (n424,n191);
nand (n425,n426,n188);
nand (n426,n427,n428);
or (n427,n122,n137);
nand (n428,n137,n122);
nand (n429,n430,n432);
or (n430,n431,n219);
not (n431,n229);
nand (n432,n433,n225);
nand (n433,n434,n435);
or (n434,n146,n217);
nand (n435,n217,n146);
nand (n436,n437,n444);
or (n437,n236,n438);
not (n438,n439);
nand (n439,n440,n442);
or (n440,n441,n238);
not (n442,n443);
and (n443,n441,n238);
or (n444,n445,n235);
not (n445,n246);
or (n446,n447,n685);
and (n447,n448,n528);
xor (n448,n449,n482);
xor (n449,n450,n481);
xor (n450,n451,n480);
or (n451,n452,n479);
and (n452,n453,n471);
xor (n453,n454,n463);
nand (n454,n455,n462);
or (n455,n456,n336);
not (n456,n457);
nand (n457,n458,n460);
not (n458,n459);
and (n459,n78,n73);
nand (n460,n461,n72);
not (n461,n78);
nand (n462,n346,n338);
nand (n463,n464,n470);
or (n464,n465,n61);
not (n465,n466);
nand (n466,n467,n468);
or (n467,n104,n57);
not (n468,n469);
and (n469,n104,n57);
nand (n470,n53,n70);
nand (n471,n472,n477);
or (n472,n473,n113);
not (n473,n474);
nor (n474,n475,n476);
and (n475,n193,n119);
and (n476,n194,n116);
nand (n477,n478,n115);
not (n478,n117);
and (n479,n454,n463);
xor (n480,n110,n154);
xor (n481,n209,n251);
xor (n482,n483,n486);
xor (n483,n484,n485);
xor (n484,n283,n334);
xor (n485,n22,n81);
or (n486,n487,n527);
and (n487,n488,n505);
xor (n488,n489,n496);
nand (n489,n490,n495);
or (n490,n131,n491);
nor (n491,n492,n493);
and (n492,n141,n231);
and (n493,n142,n494);
not (n494,n231);
or (n495,n132,n144);
nand (n496,n497,n498);
or (n497,n236,n239);
nand (n498,n499,n504);
not (n499,n500);
nor (n500,n501,n503);
and (n501,n262,n502);
not (n502,n256);
and (n503,n238,n256);
not (n504,n235);
or (n505,n506,n526);
and (n506,n507,n523);
xor (n507,n508,n515);
nand (n508,n509,n510);
or (n509,n114,n473);
nand (n510,n511,n514);
nor (n511,n512,n513);
and (n512,n177,n116);
and (n513,n180,n119);
not (n514,n113);
nand (n515,n516,n521);
or (n516,n517,n131);
not (n517,n518);
nand (n518,n519,n520);
or (n519,n215,n141);
nand (n520,n141,n215);
nand (n521,n522,n133);
not (n522,n491);
nor (n523,n524,n525);
nand (n524,n295,n31);
nand (n525,n70,n88);
and (n526,n508,n515);
and (n527,n489,n496);
or (n528,n529,n684);
and (n529,n530,n599);
xor (n530,n531,n598);
or (n531,n532,n597);
and (n532,n533,n568);
xor (n533,n534,n542);
nand (n534,n535,n541);
or (n535,n235,n536);
not (n536,n537);
nor (n537,n538,n539);
and (n538,n277,n262);
and (n539,n540,n238);
not (n540,n277);
or (n541,n500,n236);
or (n542,n543,n567);
and (n543,n544,n556);
xor (n544,n545,n549);
nand (n545,n546,n548);
or (n546,n547,n525);
not (n547,n524);
nand (n548,n547,n525);
nand (n549,n550,n555);
or (n550,n113,n551);
nor (n551,n552,n553);
and (n552,n152,n119);
and (n553,n554,n116);
not (n554,n152);
nand (n555,n511,n115);
nand (n556,n557,n562);
or (n557,n181,n558);
not (n558,n559);
nor (n559,n560,n561);
and (n560,n494,n178);
and (n561,n231,n137);
or (n562,n563,n564);
not (n563,n188);
nor (n564,n565,n566);
and (n565,n146,n137);
and (n566,n147,n178);
and (n567,n545,n549);
or (n568,n569,n596);
and (n569,n570,n585);
xor (n570,n571,n578);
nand (n571,n572,n577);
or (n572,n573,n131);
not (n573,n574);
nand (n574,n575,n576);
or (n575,n305,n141);
nand (n576,n141,n305);
nand (n577,n133,n518);
nand (n578,n579,n580);
or (n579,n236,n536);
nand (n580,n581,n504);
nand (n581,n582,n584);
not (n582,n583);
and (n583,n332,n238);
nand (n584,n331,n262);
nand (n585,n586,n591);
or (n586,n587,n267);
not (n587,n588);
nor (n588,n589,n590);
and (n589,n358,n257);
and (n590,n356,n271);
nand (n591,n592,n593);
not (n592,n260);
nor (n593,n594,n595);
and (n594,n371,n257);
and (n595,n312,n271);
and (n596,n571,n578);
and (n597,n534,n542);
xor (n598,n488,n505);
xor (n599,n600,n651);
xor (n600,n601,n629);
or (n601,n602,n628);
and (n602,n603,n622);
xor (n603,n604,n614);
nand (n604,n605,n610);
or (n605,n294,n606);
not (n606,n607);
nand (n607,n608,n609);
or (n608,n42,n47);
nand (n609,n42,n47);
nand (n610,n294,n611,n299);
nand (n611,n612,n613);
or (n612,n42,n30);
nand (n613,n30,n42);
nand (n614,n615,n621);
or (n615,n616,n336);
not (n616,n617);
nand (n617,n618,n619);
or (n618,n73,n56);
not (n619,n620);
and (n620,n56,n73);
nand (n621,n338,n457);
nand (n622,n623,n624);
or (n623,n465,n69);
or (n624,n61,n625);
nor (n625,n626,n627);
and (n626,n59,n90);
and (n627,n88,n57);
and (n628,n604,n614);
or (n629,n630,n650);
and (n630,n631,n644);
xor (n631,n632,n639);
nor (n632,n633,n290);
and (n633,n634,n637);
nand (n634,n635,n216);
not (n635,n636);
and (n636,n31,n297);
nand (n637,n30,n638);
not (n638,n297);
nor (n639,n640,n57);
nor (n640,n641,n643);
and (n641,n642,n73);
nand (n642,n88,n65);
and (n643,n90,n66);
nand (n644,n645,n646);
or (n645,n564,n181);
nand (n646,n647,n188);
nor (n647,n648,n649);
and (n648,n554,n178);
and (n649,n152,n137);
and (n650,n632,n639);
or (n651,n652,n683);
and (n652,n653,n673);
xor (n653,n654,n665);
nand (n654,n655,n660);
or (n655,n656,n219);
not (n656,n657);
nand (n657,n658,n659);
or (n658,n289,n216);
nand (n659,n216,n289);
nand (n660,n225,n661);
nand (n661,n662,n664);
or (n662,n663,n217);
not (n663,n305);
nand (n664,n217,n663);
nand (n665,n666,n668);
or (n666,n267,n667);
not (n667,n593);
nand (n668,n592,n669);
nand (n669,n670,n671);
or (n670,n332,n257);
not (n671,n672);
and (n672,n332,n257);
nand (n673,n674,n679);
or (n674,n675,n316);
not (n675,n676);
nor (n676,n677,n678);
and (n677,n351,n313);
and (n678,n349,n330);
nand (n679,n318,n680);
nor (n680,n681,n682);
and (n681,n356,n330);
and (n682,n358,n313);
and (n683,n654,n665);
and (n684,n531,n598);
and (n685,n449,n482);
xor (n686,n687,n738);
xor (n687,n688,n691);
or (n688,n689,n690);
and (n689,n483,n486);
and (n690,n484,n485);
or (n691,n692,n737);
and (n692,n693,n728);
xor (n693,n694,n697);
or (n694,n695,n696);
and (n695,n600,n651);
and (n696,n601,n629);
or (n697,n698,n727);
and (n698,n699,n714);
xor (n699,n700,n701);
xor (n700,n453,n471);
xor (n701,n702,n711);
xor (n702,n703,n707);
nand (n703,n704,n706);
or (n704,n705,n267);
not (n705,n669);
nand (n706,n592,n275);
nand (n707,n708,n710);
or (n708,n709,n316);
not (n709,n680);
nand (n710,n318,n310);
nand (n711,n712,n713);
or (n712,n606,n293);
nand (n713,n295,n287);
xor (n714,n715,n723);
xor (n715,n716,n720);
nand (n716,n717,n719);
or (n717,n718,n181);
not (n718,n647);
nand (n719,n188,n175);
nand (n720,n721,n722);
or (n721,n156,n157);
nand (n722,n157,n156);
nand (n723,n724,n726);
or (n724,n219,n725);
not (n725,n661);
or (n726,n224,n212);
and (n727,n700,n701);
xor (n728,n729,n734);
xor (n729,n730,n731);
xor (n730,n161,n172);
or (n731,n732,n733);
and (n732,n715,n723);
and (n733,n716,n720);
or (n734,n735,n736);
and (n735,n702,n711);
and (n736,n703,n707);
and (n737,n694,n697);
xor (n738,n739,n768);
xor (n739,n740,n765);
xor (n740,n741,n757);
xor (n741,n742,n749);
nand (n742,n743,n744);
or (n743,n253,n267);
nand (n744,n592,n745);
nand (n745,n746,n747);
or (n746,n242,n257);
not (n747,n748);
and (n748,n242,n257);
nand (n749,n750,n752);
or (n750,n751,n293);
not (n751,n303);
nand (n752,n295,n753);
nand (n753,n754,n756);
or (n754,n42,n755);
not (n755,n215);
nand (n756,n42,n755);
nand (n757,n758,n764);
or (n758,n759,n317);
not (n759,n760);
nand (n760,n761,n763);
not (n761,n762);
and (n762,n277,n313);
nand (n763,n330,n540);
or (n764,n316,n328);
or (n765,n766,n767);
and (n766,n729,n734);
and (n767,n730,n731);
or (n768,n769,n770);
and (n769,n450,n481);
and (n770,n451,n480);
or (n771,n772,n894);
and (n772,n773,n893);
xor (n773,n774,n775);
xor (n774,n693,n728);
or (n775,n776,n892);
and (n776,n777,n811);
xor (n777,n778,n810);
or (n778,n779,n809);
and (n779,n780,n808);
xor (n780,n781,n782);
xor (n781,n631,n644);
or (n782,n783,n807);
and (n783,n784,n799);
xor (n784,n785,n792);
nand (n785,n786,n791);
or (n786,n787,n219);
not (n787,n788);
nand (n788,n789,n790);
or (n789,n48,n216);
nand (n790,n216,n48);
nand (n791,n657,n225);
nand (n792,n793,n798);
or (n793,n794,n316);
not (n794,n795);
nor (n795,n796,n797);
and (n796,n461,n313);
and (n797,n78,n330);
nand (n798,n318,n676);
nand (n799,n800,n806);
or (n800,n801,n336);
not (n801,n802);
nor (n802,n803,n805);
and (n803,n804,n73);
not (n804,n104);
and (n805,n104,n72);
nand (n806,n338,n617);
and (n807,n785,n792);
xor (n808,n653,n673);
and (n809,n781,n782);
xor (n810,n699,n714);
or (n811,n812,n891);
and (n812,n813,n816);
xor (n813,n814,n815);
xor (n814,n507,n523);
xor (n815,n603,n622);
or (n816,n817,n890);
and (n817,n818,n864);
xor (n818,n819,n840);
or (n819,n820,n839);
and (n820,n821,n832);
xor (n821,n822,n829);
nand (n822,n823,n828);
or (n823,n824,n181);
not (n824,n825);
nand (n825,n826,n827);
or (n826,n755,n137);
nand (n827,n137,n755);
nand (n828,n559,n188);
nor (n829,n830,n831);
nand (n830,n225,n31);
nand (n831,n338,n88);
nand (n832,n833,n838);
or (n833,n834,n131);
not (n834,n835);
nand (n835,n836,n837);
or (n836,n289,n141);
nand (n837,n289,n141);
nand (n838,n133,n574);
and (n839,n822,n829);
or (n840,n841,n863);
and (n841,n842,n856);
xor (n842,n843,n850);
nor (n843,n844,n216);
and (n844,n845,n848);
nand (n845,n846,n141);
not (n846,n847);
and (n847,n31,n222);
nand (n848,n30,n849);
not (n849,n222);
nor (n850,n851,n73);
nor (n851,n852,n855);
and (n852,n853,n313);
nand (n853,n88,n854);
not (n854,n340);
nor (n855,n88,n854);
nand (n856,n857,n862);
or (n857,n858,n219);
not (n858,n859);
nor (n859,n860,n861);
and (n860,n216,n30);
and (n861,n31,n217);
nand (n862,n788,n225);
and (n863,n843,n850);
or (n864,n865,n889);
and (n865,n866,n882);
xor (n866,n867,n874);
nand (n867,n868,n873);
or (n868,n869,n316);
not (n869,n870);
nor (n870,n871,n872);
and (n871,n60,n313);
and (n872,n56,n330);
nand (n873,n318,n795);
nand (n874,n875,n876);
or (n875,n337,n801);
nand (n876,n877,n881);
not (n877,n878);
nor (n878,n879,n880);
and (n879,n90,n72);
and (n880,n88,n73);
not (n881,n336);
nand (n882,n883,n888);
or (n883,n113,n884);
not (n884,n885);
nand (n885,n886,n887);
or (n886,n147,n119);
nand (n887,n119,n147);
or (n888,n551,n114);
and (n889,n867,n874);
and (n890,n819,n840);
and (n891,n814,n815);
and (n892,n778,n810);
xor (n893,n448,n528);
and (n894,n774,n775);
nand (n895,n14,n771);
nor (n896,n897,n1341);
and (n897,n898,n1336);
nand (n898,n899,n1335);
or (n899,n900,n1001);
not (n900,n901);
or (n901,n902,n919);
xor (n902,n903,n918);
xor (n903,n904,n917);
or (n904,n905,n916);
and (n905,n906,n915);
xor (n906,n907,n908);
xor (n907,n533,n568);
or (n908,n909,n914);
and (n909,n910,n913);
xor (n910,n911,n912);
xor (n911,n570,n585);
xor (n912,n784,n799);
xor (n913,n544,n556);
and (n914,n911,n912);
xor (n915,n780,n808);
and (n916,n907,n908);
xor (n917,n530,n599);
xor (n918,n777,n811);
or (n919,n920,n1000);
and (n920,n921,n999);
xor (n921,n922,n923);
xor (n922,n813,n816);
or (n923,n924,n998);
and (n924,n925,n997);
xor (n925,n926,n966);
or (n926,n927,n965);
and (n927,n928,n943);
xor (n928,n929,n936);
nand (n929,n930,n934);
or (n930,n931,n235);
nor (n931,n932,n933);
and (n932,n262,n371);
and (n933,n238,n312);
or (n934,n935,n236);
not (n935,n581);
nand (n936,n937,n942);
or (n937,n938,n267);
not (n938,n939);
nor (n939,n940,n941);
and (n940,n351,n257);
and (n941,n349,n271);
nand (n942,n592,n588);
or (n943,n944,n964);
and (n944,n945,n957);
xor (n945,n946,n953);
nand (n946,n947,n952);
or (n947,n948,n113);
not (n948,n949);
nor (n949,n950,n951);
and (n950,n231,n116);
and (n951,n494,n119);
nand (n952,n885,n115);
nand (n953,n954,n956);
or (n954,n955,n831);
not (n955,n830);
nand (n956,n955,n831);
nand (n957,n958,n963);
or (n958,n959,n181);
not (n959,n960);
nor (n960,n961,n962);
and (n961,n663,n178);
and (n962,n305,n137);
or (n963,n563,n824);
and (n964,n946,n953);
and (n965,n929,n936);
or (n966,n967,n996);
and (n967,n968,n995);
xor (n968,n969,n970);
xor (n969,n842,n856);
or (n970,n971,n994);
and (n971,n972,n986);
xor (n972,n973,n979);
nand (n973,n974,n978);
or (n974,n975,n235);
or (n975,n976,n977);
and (n976,n356,n262);
and (n977,n358,n238);
or (n978,n931,n236);
nand (n979,n980,n985);
or (n980,n981,n131);
not (n981,n982);
nor (n982,n983,n984);
and (n983,n47,n141);
and (n984,n48,n142);
nand (n985,n835,n133);
nand (n986,n987,n993);
or (n987,n988,n267);
not (n988,n989);
nand (n989,n990,n991);
or (n990,n78,n257);
not (n991,n992);
and (n992,n78,n257);
nand (n993,n592,n939);
and (n994,n973,n979);
xor (n995,n866,n882);
and (n996,n969,n970);
xor (n997,n818,n864);
and (n998,n926,n966);
xor (n999,n906,n915);
and (n1000,n922,n923);
not (n1001,n1002);
nand (n1002,n1003,n1332,n1334);
nand (n1003,n1004,n1076,n1325);
nand (n1004,n1005,n1007);
not (n1005,n1006);
xor (n1006,n921,n999);
not (n1007,n1008);
or (n1008,n1009,n1075);
and (n1009,n1010,n1074);
xor (n1010,n1011,n1012);
xor (n1011,n910,n913);
or (n1012,n1013,n1073);
and (n1013,n1014,n1072);
xor (n1014,n1015,n1016);
xor (n1015,n821,n832);
or (n1016,n1017,n1071);
and (n1017,n1018,n1050);
xor (n1018,n1019,n1026);
nand (n1019,n1020,n1025);
or (n1020,n1021,n316);
not (n1021,n1022);
nor (n1022,n1023,n1024);
and (n1023,n804,n313);
and (n1024,n104,n330);
nand (n1025,n318,n870);
or (n1026,n1027,n1049);
and (n1027,n1028,n1040);
xor (n1028,n1029,n1036);
nand (n1029,n1030,n1035);
or (n1030,n1031,n181);
not (n1031,n1032);
nand (n1032,n1033,n1034);
or (n1033,n289,n178);
nand (n1034,n178,n289);
nand (n1035,n960,n188);
nor (n1036,n1037,n1039);
not (n1037,n1038);
and (n1038,n318,n88);
nand (n1039,n31,n133);
nand (n1040,n1041,n1047);
or (n1041,n235,n1042);
not (n1042,n1043);
nand (n1043,n1044,n1046);
not (n1044,n1045);
and (n1045,n349,n238);
nand (n1046,n262,n351);
nand (n1047,n1048,n237);
not (n1048,n975);
and (n1049,n1029,n1036);
or (n1050,n1051,n1070);
and (n1051,n1052,n1064);
xor (n1052,n1053,n1059);
nor (n1053,n1054,n141);
and (n1054,n1055,n1058);
nand (n1055,n1056,n178);
not (n1056,n1057);
and (n1057,n31,n136);
nand (n1058,n30,n135);
nor (n1059,n1060,n313);
nor (n1060,n1061,n1063);
and (n1061,n1062,n257);
nand (n1062,n88,n324);
and (n1063,n90,n320);
nand (n1064,n1065,n1066);
or (n1065,n114,n948);
nand (n1066,n1067,n514);
nor (n1067,n1068,n1069);
and (n1068,n215,n116);
and (n1069,n755,n119);
and (n1070,n1053,n1059);
and (n1071,n1019,n1026);
xor (n1072,n928,n943);
and (n1073,n1015,n1016);
xor (n1074,n925,n997);
and (n1075,n1011,n1012);
nand (n1076,n1077,n1324);
or (n1077,n1078,n1310);
not (n1078,n1079);
nand (n1079,n1080,n1309);
or (n1080,n1081,n1181);
not (n1081,n1082);
nand (n1082,n1083,n1145);
not (n1083,n1084);
xor (n1084,n1085,n1115);
xor (n1085,n1086,n1087);
xor (n1086,n1018,n1050);
or (n1087,n1088,n1114);
and (n1088,n1089,n1113);
xor (n1089,n1090,n1112);
or (n1090,n1091,n1111);
and (n1091,n1092,n1107);
xor (n1092,n1093,n1100);
nand (n1093,n1094,n1099);
or (n1094,n1095,n181);
not (n1095,n1096);
nand (n1096,n1097,n1098);
or (n1097,n48,n178);
nand (n1098,n178,n48);
nand (n1099,n1032,n188);
nand (n1100,n1101,n1102);
or (n1101,n236,n1042);
nand (n1102,n1103,n504);
nand (n1103,n1104,n1106);
not (n1104,n1105);
and (n1105,n78,n238);
nand (n1106,n262,n461);
nand (n1107,n1108,n1110);
or (n1108,n1109,n1037);
not (n1109,n1039);
or (n1110,n1038,n1039);
and (n1111,n1093,n1100);
xor (n1112,n1052,n1064);
xor (n1113,n1028,n1040);
and (n1114,n1090,n1112);
xor (n1115,n1116,n1144);
xor (n1116,n1117,n1143);
or (n1117,n1118,n1142);
and (n1118,n1119,n1134);
xor (n1119,n1120,n1127);
nand (n1120,n1121,n1126);
or (n1121,n1122,n131);
not (n1122,n1123);
nor (n1123,n1124,n1125);
and (n1124,n141,n30);
and (n1125,n31,n142);
nand (n1126,n982,n133);
nand (n1127,n1128,n1133);
or (n1128,n1129,n267);
not (n1129,n1130);
nor (n1130,n1131,n1132);
and (n1131,n56,n271);
and (n1132,n60,n257);
nand (n1133,n592,n989);
nand (n1134,n1135,n1141);
or (n1135,n1136,n316);
not (n1136,n1137);
nand (n1137,n1138,n1139);
or (n1138,n88,n313);
not (n1139,n1140);
and (n1140,n88,n313);
nand (n1141,n318,n1022);
and (n1142,n1120,n1127);
xor (n1143,n972,n986);
xor (n1144,n945,n957);
not (n1145,n1146);
or (n1146,n1147,n1180);
and (n1147,n1148,n1179);
xor (n1148,n1149,n1150);
xor (n1149,n1119,n1134);
or (n1150,n1151,n1178);
and (n1151,n1152,n1166);
xor (n1152,n1153,n1159);
nand (n1153,n1154,n1158);
or (n1154,n1155,n267);
nor (n1155,n1156,n1157);
and (n1156,n804,n271);
and (n1157,n104,n257);
nand (n1158,n1130,n592);
nand (n1159,n1160,n1165);
or (n1160,n113,n1161);
not (n1161,n1162);
nor (n1162,n1163,n1164);
and (n1163,n305,n116);
and (n1164,n663,n119);
nand (n1165,n1067,n115);
and (n1166,n1167,n1173);
nor (n1167,n1168,n178);
and (n1168,n1169,n1172);
nand (n1169,n1170,n119);
not (n1170,n1171);
and (n1171,n31,n184);
nand (n1172,n186,n30);
nor (n1173,n1174,n257);
and (n1174,n1175,n1177);
nand (n1175,n1176,n238);
or (n1176,n90,n263);
nand (n1177,n90,n263);
and (n1178,n1153,n1159);
xor (n1179,n1089,n1113);
and (n1180,n1149,n1150);
not (n1181,n1182);
nand (n1182,n1183,n1308);
or (n1183,n1184,n1300);
not (n1184,n1185);
nand (n1185,n1186,n1299);
or (n1186,n1187,n1258);
not (n1187,n1188);
nand (n1188,n1189,n1219);
not (n1189,n1190);
xor (n1190,n1191,n1218);
xor (n1191,n1192,n1217);
or (n1192,n1193,n1216);
and (n1193,n1194,n1210);
xor (n1194,n1195,n1202);
nand (n1195,n1196,n1201);
or (n1196,n1197,n181);
not (n1197,n1198);
nand (n1198,n1199,n1200);
or (n1199,n31,n178);
nand (n1200,n178,n31);
nand (n1201,n1096,n188);
nand (n1202,n1203,n1209);
or (n1203,n1204,n235);
not (n1204,n1205);
nand (n1205,n1206,n1208);
not (n1206,n1207);
and (n1207,n56,n238);
nand (n1208,n262,n60);
nand (n1209,n1103,n237);
nand (n1210,n1211,n1215);
or (n1211,n267,n1212);
nor (n1212,n1213,n1214);
and (n1213,n271,n90);
and (n1214,n88,n257);
or (n1215,n260,n1155);
and (n1216,n1195,n1202);
xor (n1217,n1092,n1107);
xor (n1218,n1152,n1166);
not (n1219,n1220);
or (n1220,n1221,n1257);
and (n1221,n1222,n1235);
xor (n1222,n1223,n1230);
nand (n1223,n1224,n1225);
or (n1224,n114,n1161);
or (n1225,n113,n1226);
not (n1226,n1227);
nor (n1227,n1228,n1229);
and (n1228,n289,n116);
and (n1229,n292,n119);
xor (n1230,n1231,n1232);
xor (n1231,n1167,n1173);
nor (n1232,n1233,n1234);
nand (n1233,n592,n88);
nand (n1234,n188,n31);
or (n1235,n1236,n1256);
and (n1236,n1237,n1249);
xor (n1237,n1238,n1245);
nand (n1238,n1239,n1244);
or (n1239,n113,n1240);
not (n1240,n1241);
nor (n1241,n1242,n1243);
and (n1242,n47,n119);
and (n1243,n48,n116);
nand (n1244,n1227,n115);
nand (n1245,n1246,n1248);
or (n1246,n1234,n1247);
not (n1247,n1233);
nand (n1248,n1247,n1234);
nand (n1249,n1250,n1255);
or (n1250,n235,n1251);
not (n1251,n1252);
nor (n1252,n1253,n1254);
and (n1253,n804,n238);
and (n1254,n104,n262);
nand (n1255,n1205,n237);
and (n1256,n1238,n1245);
and (n1257,n1223,n1230);
not (n1258,n1259);
nand (n1259,n1260,n1298);
or (n1260,n1261,n1264);
nor (n1261,n1262,n1263);
xor (n1262,n1222,n1235);
xor (n1263,n1194,n1210);
nor (n1264,n1265,n1296);
and (n1265,n1266,n1283);
nand (n1266,n1267,n1269);
not (n1267,n1268);
xor (n1268,n1237,n1249);
not (n1269,n1270);
or (n1270,n1271,n1282);
and (n1271,n1272,n1276);
xor (n1272,n1273,n1275);
nor (n1273,n1274,n119);
and (n1274,n31,n115);
and (n1275,n262,n90,n237);
nand (n1276,n1277,n1278);
or (n1277,n236,n1251);
nand (n1278,n1279,n504);
nor (n1279,n1280,n1281);
and (n1280,n90,n238);
and (n1281,n88,n262);
and (n1282,n1273,n1275);
or (n1283,n1284,n1295);
and (n1284,n1285,n1294);
xor (n1285,n1286,n1288);
and (n1286,n1274,n1287);
and (n1287,n88,n237);
nand (n1288,n1289,n1290);
or (n1289,n114,n1240);
nand (n1290,n1291,n514);
nand (n1291,n1292,n1293);
or (n1292,n119,n31);
or (n1293,n30,n116);
xor (n1294,n1272,n1276);
and (n1295,n1286,n1288);
not (n1296,n1297);
nand (n1297,n1268,n1270);
nand (n1298,n1262,n1263);
nand (n1299,n1190,n1220);
not (n1300,n1301);
nand (n1301,n1302,n1304);
not (n1302,n1303);
xor (n1303,n1148,n1179);
not (n1304,n1305);
or (n1305,n1306,n1307);
and (n1306,n1191,n1218);
and (n1307,n1192,n1217);
nand (n1308,n1303,n1305);
nand (n1309,n1084,n1146);
not (n1310,n1311);
nand (n1311,n1312,n1320);
not (n1312,n1313);
xor (n1313,n1314,n1319);
xor (n1314,n1315,n1318);
or (n1315,n1316,n1317);
and (n1316,n1116,n1144);
and (n1317,n1117,n1143);
xor (n1318,n968,n995);
xor (n1319,n1014,n1072);
not (n1320,n1321);
or (n1321,n1322,n1323);
and (n1322,n1085,n1115);
and (n1323,n1086,n1087);
nand (n1324,n1313,n1321);
nand (n1325,n1326,n1328);
not (n1326,n1327);
xor (n1327,n1010,n1074);
not (n1328,n1329);
or (n1329,n1330,n1331);
and (n1330,n1314,n1319);
and (n1331,n1315,n1318);
nand (n1332,n1004,n1333);
nor (n1333,n1326,n1328);
nand (n1334,n1006,n1008);
nand (n1335,n902,n919);
or (n1336,n1337,n1338);
xor (n1337,n773,n893);
or (n1338,n1339,n1340);
and (n1339,n903,n918);
and (n1340,n904,n917);
and (n1341,n1337,n1338);
nand (n1342,n11,n896);
nor (n1344,n1345,n9);
not (n1345,n1343);
not (n1346,n1347);
nand (n1347,n1348,n1615);
nand (n1348,n1349,n1607);
nand (n1349,n1350,n1605);
or (n1350,n1351,n1360);
not (n1351,n1352);
nand (n1352,n1353,n1359);
not (n1353,n1354);
nand (n1354,n1355,n1358);
or (n1355,n1356,n1001);
not (n1356,n1357);
nand (n1357,n901,n1335);
or (n1358,n1357,n1002);
not (n1360,n1361);
nand (n1361,n1362,n1603);
or (n1362,n1363,n1376);
not (n1363,n1364);
nand (n1364,n1365,n1375);
not (n1365,n1366);
nand (n1366,n1367,n1374);
or (n1367,n1368,n1373);
nand (n1368,n1369,n1372);
or (n1369,n1370,n1371);
not (n1370,n1325);
not (n1371,n1076);
not (n1372,n1333);
nand (n1373,n1004,n1334);
nand (n1374,n1373,n1368);
not (n1376,n1377);
nand (n1377,n1378,n1597);
or (n1378,n1379,n1386);
nor (n1379,n1380,n1382);
not (n1380,n1381);
nand (n1382,n1383,n1385);
or (n1383,n1076,n1384);
nand (n1384,n1325,n1372);
nand (n1385,n1384,n1076);
not (n1386,n1387);
and (n1387,n1388,n1592);
or (n1388,n1389,n1591);
and (n1389,n1390,n1398);
xor (n1390,n1391,n1393);
not (n1391,n1392);
nand (n1393,n1394,n1397);
or (n1394,n1181,n1395);
not (n1395,n1396);
nand (n1396,n1082,n1309);
or (n1397,n1182,n1396);
or (n1398,n1399,n1548,n1590);
and (n1399,n1400,n1546);
xor (n1400,n1401,n1516);
xor (n1401,n1402,n1458);
xor (n1402,n1403,n1125);
xor (n1403,n1404,n1456);
xor (n1404,n1405,n1455);
xor (n1405,n1406,n1446);
xor (n1406,n1407,n1445);
xor (n1407,n1408,n1431);
xor (n1408,n1409,n1430);
xor (n1409,n1410,n1412);
xor (n1410,n1411,n1068);
and (n1411,n231,n115);
or (n1412,n1413,n1415);
and (n1413,n1414,n1163);
and (n1414,n215,n115);
and (n1415,n1416,n1417);
xor (n1416,n1414,n1163);
or (n1417,n1418,n1420);
and (n1418,n1419,n1228);
and (n1419,n305,n115);
and (n1420,n1421,n1422);
xor (n1421,n1419,n1228);
or (n1422,n1423,n1425);
and (n1423,n1424,n1243);
and (n1424,n289,n115);
and (n1425,n1426,n1427);
xor (n1426,n1424,n1243);
and (n1427,n1428,n1429);
and (n1428,n48,n115);
and (n1429,n31,n116);
and (n1430,n305,n184);
or (n1431,n1432,n1435);
and (n1432,n1433,n1434);
xor (n1433,n1416,n1417);
and (n1434,n289,n184);
and (n1435,n1436,n1437);
xor (n1436,n1433,n1434);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1421,n1422);
and (n1440,n48,n184);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
and (n1443,n1444,n1171);
xor (n1444,n1426,n1427);
and (n1445,n289,n137);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1436,n1437);
and (n1449,n48,n137);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
and (n1452,n1453,n1454);
xor (n1453,n1442,n1443);
and (n1454,n31,n137);
and (n1455,n48,n136);
and (n1456,n1457,n1057);
xor (n1457,n1451,n1452);
not (n1458,n1459);
xor (n1459,n1460,n1140);
xor (n1460,n1461,n1513);
xor (n1461,n1462,n1512);
xor (n1462,n1463,n1505);
xor (n1463,n1464,n1504);
xor (n1464,n1465,n1489);
xor (n1465,n1466,n1488);
xor (n1466,n1467,n1469);
xor (n1467,n1468,n1045);
and (n1468,n356,n237);
or (n1469,n1470,n1472);
and (n1470,n1471,n1105);
and (n1471,n349,n237);
and (n1472,n1473,n1474);
xor (n1473,n1471,n1105);
or (n1474,n1475,n1477);
and (n1475,n1476,n1207);
and (n1476,n78,n237);
and (n1477,n1478,n1479);
xor (n1478,n1476,n1207);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
and (n1481,n56,n237);
and (n1482,n104,n238);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
and (n1485,n1486,n1487);
and (n1486,n104,n237);
and (n1487,n88,n238);
and (n1488,n78,n263);
or (n1489,n1490,n1493);
and (n1490,n1491,n1492);
xor (n1491,n1473,n1474);
and (n1492,n56,n263);
and (n1493,n1494,n1495);
xor (n1494,n1491,n1492);
or (n1495,n1496,n1499);
and (n1496,n1497,n1498);
xor (n1497,n1478,n1479);
and (n1498,n104,n263);
and (n1499,n1500,n1501);
xor (n1500,n1497,n1498);
and (n1501,n1502,n1503);
xor (n1502,n1484,n1485);
and (n1503,n88,n263);
and (n1504,n56,n257);
or (n1505,n1506,n1508);
and (n1506,n1507,n1157);
xor (n1507,n1494,n1495);
and (n1508,n1509,n1510);
xor (n1509,n1507,n1157);
and (n1510,n1511,n1214);
xor (n1511,n1500,n1501);
and (n1512,n104,n320);
and (n1513,n1514,n1515);
xor (n1514,n1509,n1510);
and (n1515,n88,n320);
or (n1516,n1517,n1521,n1545);
and (n1517,n1518,n1519);
xor (n1518,n1457,n1057);
not (n1519,n1520);
xor (n1520,n1514,n1515);
and (n1521,n1519,n1522);
or (n1522,n1523,n1527,n1544);
and (n1523,n1524,n1525);
xor (n1524,n1453,n1454);
not (n1525,n1526);
xor (n1526,n1511,n1214);
and (n1527,n1525,n1528);
or (n1528,n1529,n1533,n1543);
and (n1529,n1530,n1531);
xor (n1530,n1444,n1171);
not (n1531,n1532);
xor (n1532,n1502,n1503);
and (n1533,n1531,n1534);
or (n1534,n1535,n1539,n1542);
and (n1535,n1536,n1537);
xor (n1536,n1428,n1429);
not (n1537,n1538);
xor (n1538,n1486,n1487);
and (n1539,n1537,n1540);
or (n1540,n1274,n1541);
not (n1541,n1287);
and (n1542,n1536,n1540);
and (n1543,n1530,n1534);
and (n1544,n1524,n1528);
and (n1545,n1518,n1522);
not (n1546,n1547);
and (n1548,n1546,n1549);
or (n1549,n1550,n1555,n1589);
and (n1550,n1551,n1553);
xor (n1551,n1552,n1522);
xor (n1552,n1518,n1519);
not (n1553,n1554);
and (n1555,n1553,n1556);
or (n1556,n1557,n1562,n1588);
and (n1557,n1558,n1560);
xor (n1558,n1559,n1528);
xor (n1559,n1524,n1525);
not (n1560,n1561);
and (n1562,n1560,n1563);
or (n1563,n1564,n1569,n1587);
and (n1564,n1565,n1567);
xor (n1565,n1566,n1534);
xor (n1566,n1530,n1531);
not (n1567,n1568);
and (n1569,n1567,n1570);
or (n1570,n1571,n1576,n1586);
and (n1571,n1572,n1574);
xor (n1572,n1573,n1540);
xor (n1573,n1536,n1537);
not (n1574,n1575);
and (n1576,n1577,n1574);
or (n1577,n1578,n1585);
and (n1578,n1579,n1584);
xor (n1579,n1580,n1582);
not (n1580,n1581);
not (n1582,n1583);
xor (n1584,n1274,n1287);
and (n1585,n1582,n1580);
and (n1586,n1572,n1577);
and (n1587,n1565,n1570);
and (n1588,n1558,n1563);
and (n1589,n1551,n1556);
and (n1590,n1400,n1549);
and (n1591,n1391,n1393);
nand (n1592,n1593,n1596);
not (n1593,n1594);
xnor (n1594,n1079,n1595);
nand (n1595,n1311,n1324);
nor (n1597,n1598,n1601);
nor (n1598,n1379,n1599);
nand (n1599,n1600,n1594);
not (n1600,n1596);
nor (n1601,n1602,n1381);
not (n1602,n1382);
nand (n1603,n1604,n1366);
not (n1604,n1375);
nand (n1605,n1606,n1354);
not (n1606,n1359);
nand (n1607,n1608,n1614);
not (n1608,n1609);
nand (n1609,n1610,n1613);
or (n1610,n1611,n898);
nand (n1611,n1612,n1336);
not (n1612,n1341);
nand (n1613,n898,n1611);
nand (n1615,n1616,n1609);
not (n1616,n1614);
or (n1617,n1347,n6);
and (n1618,n1619,n1635);
not (n1619,n1620);
or (n1620,n1621,n1632);
or (n1621,n1622,n1629);
or (n1622,n1623,n1626);
xor (n1623,n1624,n1625);
xor (n1626,n1627,n1628);
xor (n1629,n1630,n1631);
xor (n1632,n1633,n1634);
xor (n1635,n1636,n1637);
or (n1638,n1639,n1641);
not (n1639,n1640);
not (n1641,n1618);
wire s0n1642,s1n1642,notn1642;
or (n1642,s0n1642,s1n1642);
not(notn1642,n1641);
and (s0n1642,notn1642,n1640);
and (s1n1642,n1641,n1643);
xor (n1643,n1644,n2336);
xor (n1644,n1645,n1345);
xor (n1645,n1646,n2290);
xor (n1646,n1647,n1972);
xor (n1647,n1648,n1971);
xor (n1648,n1649,n1969);
xor (n1649,n1650,n1968);
xor (n1650,n1651,n1960);
xor (n1651,n1652,n1959);
xor (n1652,n1653,n1944);
xor (n1653,n1654,n1943);
xor (n1654,n1655,n1923);
xor (n1655,n1656,n1922);
xor (n1656,n1657,n1896);
xor (n1657,n1658,n1895);
xor (n1658,n1659,n1863);
xor (n1659,n1660,n1862);
xor (n1660,n1661,n1826);
xor (n1661,n1662,n1825);
xor (n1662,n1663,n1786);
xor (n1663,n1664,n1785);
xor (n1664,n1665,n1749);
xor (n1665,n1666,n1748);
xor (n1666,n1667,n1709);
xor (n1667,n1668,n1708);
xor (n1668,n1669,n1672);
xor (n1669,n1670,n1671);
and (n1670,n419,n115);
and (n1671,n126,n116);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
and (n1674,n126,n115);
and (n1675,n120,n116);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1681);
and (n1679,n1680,n476);
and (n1680,n120,n115);
and (n1681,n1682,n1683);
xor (n1682,n1680,n476);
or (n1683,n1684,n1686);
and (n1684,n1685,n512);
and (n1685,n194,n115);
and (n1686,n1687,n1688);
xor (n1687,n1685,n512);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
and (n1690,n177,n115);
and (n1691,n152,n116);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
and (n1696,n152,n115);
and (n1697,n147,n116);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1703);
and (n1701,n1702,n950);
and (n1702,n147,n115);
and (n1703,n1704,n1705);
xor (n1704,n1702,n950);
or (n1705,n1706,n1707);
and (n1706,n1411,n1068);
and (n1707,n1410,n1412);
and (n1708,n120,n184);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1677,n1678);
and (n1712,n194,n184);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1682,n1683);
and (n1718,n177,n184);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1687,n1688);
and (n1724,n152,n184);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1693,n1694);
and (n1730,n147,n184);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1699,n1700);
and (n1736,n231,n184);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1704,n1705);
and (n1742,n215,n184);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
or (n1745,n1746,n1747);
and (n1746,n1409,n1430);
and (n1747,n1408,n1431);
and (n1748,n194,n137);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
xor (n1751,n1714,n1715);
and (n1752,n177,n137);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
or (n1755,n1756,n1758);
and (n1756,n1757,n649);
xor (n1757,n1720,n1721);
and (n1758,n1759,n1760);
xor (n1759,n1757,n649);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1726,n1727);
and (n1763,n147,n137);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
or (n1766,n1767,n1769);
and (n1767,n1768,n561);
xor (n1768,n1732,n1733);
and (n1769,n1770,n1771);
xor (n1770,n1768,n561);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1738,n1739);
and (n1774,n215,n137);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1780);
and (n1778,n1779,n962);
xor (n1779,n1744,n1745);
and (n1780,n1781,n1782);
xor (n1781,n1779,n962);
or (n1782,n1783,n1784);
and (n1783,n1407,n1445);
and (n1784,n1406,n1446);
and (n1785,n177,n136);
or (n1786,n1787,n1790);
and (n1787,n1788,n1789);
xor (n1788,n1754,n1755);
and (n1789,n152,n136);
and (n1790,n1791,n1792);
xor (n1791,n1788,n1789);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1759,n1760);
and (n1795,n147,n136);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1765,n1766);
and (n1801,n231,n136);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1770,n1771);
and (n1807,n215,n136);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1776,n1777);
and (n1813,n305,n136);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1781,n1782);
and (n1819,n289,n136);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
or (n1822,n1823,n1824);
and (n1823,n1405,n1455);
and (n1824,n1404,n1456);
and (n1825,n152,n142);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1791,n1792);
and (n1829,n147,n142);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1836);
and (n1833,n1834,n1835);
xor (n1834,n1797,n1798);
and (n1835,n231,n142);
and (n1836,n1837,n1838);
xor (n1837,n1834,n1835);
or (n1838,n1839,n1842);
and (n1839,n1840,n1841);
xor (n1840,n1803,n1804);
and (n1841,n215,n142);
and (n1842,n1843,n1844);
xor (n1843,n1840,n1841);
or (n1844,n1845,n1848);
and (n1845,n1846,n1847);
xor (n1846,n1809,n1810);
and (n1847,n305,n142);
and (n1848,n1849,n1850);
xor (n1849,n1846,n1847);
or (n1850,n1851,n1854);
and (n1851,n1852,n1853);
xor (n1852,n1815,n1816);
and (n1853,n289,n142);
and (n1854,n1855,n1856);
xor (n1855,n1852,n1853);
or (n1856,n1857,n1859);
and (n1857,n1858,n984);
xor (n1858,n1821,n1822);
and (n1859,n1860,n1861);
xor (n1860,n1858,n984);
and (n1861,n1403,n1125);
and (n1862,n147,n222);
or (n1863,n1864,n1867);
and (n1864,n1865,n1866);
xor (n1865,n1831,n1832);
and (n1866,n231,n222);
and (n1867,n1868,n1869);
xor (n1868,n1865,n1866);
or (n1869,n1870,n1873);
and (n1870,n1871,n1872);
xor (n1871,n1837,n1838);
and (n1872,n215,n222);
and (n1873,n1874,n1875);
xor (n1874,n1871,n1872);
or (n1875,n1876,n1879);
and (n1876,n1877,n1878);
xor (n1877,n1843,n1844);
and (n1878,n305,n222);
and (n1879,n1880,n1881);
xor (n1880,n1877,n1878);
or (n1881,n1882,n1885);
and (n1882,n1883,n1884);
xor (n1883,n1849,n1850);
and (n1884,n289,n222);
and (n1885,n1886,n1887);
xor (n1886,n1883,n1884);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
xor (n1889,n1855,n1856);
and (n1890,n48,n222);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
and (n1893,n1894,n847);
xor (n1894,n1860,n1861);
and (n1895,n231,n217);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1868,n1869);
and (n1899,n215,n217);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1874,n1875);
and (n1905,n305,n217);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
or (n1908,n1909,n1912);
and (n1909,n1910,n1911);
xor (n1910,n1880,n1881);
and (n1911,n289,n217);
and (n1912,n1913,n1914);
xor (n1913,n1910,n1911);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1886,n1887);
and (n1917,n48,n217);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
and (n1920,n1921,n861);
xor (n1921,n1892,n1893);
and (n1922,n215,n297);
or (n1923,n1924,n1927);
and (n1924,n1925,n1926);
xor (n1925,n1901,n1902);
and (n1926,n305,n297);
and (n1927,n1928,n1929);
xor (n1928,n1925,n1926);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1907,n1908);
and (n1932,n289,n297);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1913,n1914);
and (n1938,n48,n297);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
and (n1941,n1942,n636);
xor (n1942,n1919,n1920);
and (n1943,n305,n42);
or (n1944,n1945,n1948);
and (n1945,n1946,n1947);
xor (n1946,n1928,n1929);
and (n1947,n289,n42);
and (n1948,n1949,n1950);
xor (n1949,n1946,n1947);
or (n1950,n1951,n1954);
and (n1951,n1952,n1953);
xor (n1952,n1934,n1935);
and (n1953,n48,n42);
and (n1954,n1955,n1956);
xor (n1955,n1952,n1953);
and (n1956,n1957,n1958);
xor (n1957,n1940,n1941);
and (n1958,n31,n42);
and (n1959,n289,n38);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
xor (n1962,n1949,n1950);
and (n1963,n48,n38);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
and (n1966,n1967,n165);
xor (n1967,n1955,n1956);
and (n1968,n48,n29);
and (n1969,n1970,n32);
xor (n1970,n1965,n1966);
and (n1971,n31,n404);
not (n1972,n1973);
xor (n1973,n1974,n2289);
xor (n1974,n1975,n2286);
xor (n1975,n1976,n106);
xor (n1976,n1977,n2277);
xor (n1977,n1978,n2276);
xor (n1978,n1979,n2264);
xor (n1979,n1980,n80);
xor (n1980,n1981,n2243);
xor (n1981,n1982,n2242);
xor (n1982,n1983,n2219);
xor (n1983,n1984,n2218);
xor (n1984,n1985,n2185);
xor (n1985,n1986,n2184);
xor (n1986,n1987,n2148);
xor (n1987,n1988,n333);
xor (n1988,n1989,n2109);
xor (n1989,n1990,n2108);
xor (n1990,n1991,n2072);
xor (n1991,n1992,n259);
xor (n1992,n1993,n2033);
xor (n1993,n1994,n2032);
xor (n1994,n1995,n1997);
xor (n1995,n1996,n250);
and (n1996,n441,n237);
or (n1997,n1998,n2000);
and (n1998,n1999,n244);
and (n1999,n248,n237);
and (n2000,n2001,n2002);
xor (n2001,n1999,n244);
or (n2002,n2003,n2005);
and (n2003,n2004,n503);
and (n2004,n242,n237);
and (n2005,n2006,n2007);
xor (n2006,n2004,n503);
or (n2007,n2008,n2011);
and (n2008,n2009,n2010);
and (n2009,n256,n237);
and (n2010,n277,n238);
and (n2011,n2012,n2013);
xor (n2012,n2009,n2010);
or (n2013,n2014,n2016);
and (n2014,n2015,n583);
and (n2015,n277,n237);
and (n2016,n2017,n2018);
xor (n2017,n2015,n583);
or (n2018,n2019,n2021);
and (n2019,n2020,n933);
and (n2020,n332,n237);
and (n2021,n2022,n2023);
xor (n2022,n2020,n933);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
and (n2025,n312,n237);
and (n2026,n356,n238);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2031);
and (n2030,n1468,n1045);
and (n2031,n1467,n1469);
and (n2032,n242,n263);
or (n2033,n2034,n2037);
and (n2034,n2035,n2036);
xor (n2035,n2001,n2002);
and (n2036,n256,n263);
and (n2037,n2038,n2039);
xor (n2038,n2035,n2036);
or (n2039,n2040,n2043);
and (n2040,n2041,n2042);
xor (n2041,n2006,n2007);
and (n2042,n277,n263);
and (n2043,n2044,n2045);
xor (n2044,n2041,n2042);
or (n2045,n2046,n2049);
and (n2046,n2047,n2048);
xor (n2047,n2012,n2013);
and (n2048,n332,n263);
and (n2049,n2050,n2051);
xor (n2050,n2047,n2048);
or (n2051,n2052,n2055);
and (n2052,n2053,n2054);
xor (n2053,n2017,n2018);
and (n2054,n312,n263);
and (n2055,n2056,n2057);
xor (n2056,n2053,n2054);
or (n2057,n2058,n2061);
and (n2058,n2059,n2060);
xor (n2059,n2022,n2023);
and (n2060,n356,n263);
and (n2061,n2062,n2063);
xor (n2062,n2059,n2060);
or (n2063,n2064,n2067);
and (n2064,n2065,n2066);
xor (n2065,n2028,n2029);
and (n2066,n349,n263);
and (n2067,n2068,n2069);
xor (n2068,n2065,n2066);
or (n2069,n2070,n2071);
and (n2070,n1466,n1488);
and (n2071,n1465,n1489);
or (n2072,n2073,n2075);
and (n2073,n2074,n279);
xor (n2074,n2038,n2039);
and (n2075,n2076,n2077);
xor (n2076,n2074,n279);
or (n2077,n2078,n2080);
and (n2078,n2079,n672);
xor (n2079,n2044,n2045);
and (n2080,n2081,n2082);
xor (n2081,n2079,n672);
or (n2082,n2083,n2086);
and (n2083,n2084,n2085);
xor (n2084,n2050,n2051);
and (n2085,n312,n257);
and (n2086,n2087,n2088);
xor (n2087,n2084,n2085);
or (n2088,n2089,n2092);
and (n2089,n2090,n2091);
xor (n2090,n2056,n2057);
and (n2091,n356,n257);
and (n2092,n2093,n2094);
xor (n2093,n2090,n2091);
or (n2094,n2095,n2098);
and (n2095,n2096,n2097);
xor (n2096,n2062,n2063);
and (n2097,n349,n257);
and (n2098,n2099,n2100);
xor (n2099,n2096,n2097);
or (n2100,n2101,n2103);
and (n2101,n2102,n992);
xor (n2102,n2068,n2069);
and (n2103,n2104,n2105);
xor (n2104,n2102,n992);
or (n2105,n2106,n2107);
and (n2106,n1464,n1504);
and (n2107,n1463,n1505);
and (n2108,n277,n320);
or (n2109,n2110,n2113);
and (n2110,n2111,n2112);
xor (n2111,n2076,n2077);
and (n2112,n332,n320);
and (n2113,n2114,n2115);
xor (n2114,n2111,n2112);
or (n2115,n2116,n2119);
and (n2116,n2117,n2118);
xor (n2117,n2081,n2082);
and (n2118,n312,n320);
and (n2119,n2120,n2121);
xor (n2120,n2117,n2118);
or (n2121,n2122,n2125);
and (n2122,n2123,n2124);
xor (n2123,n2087,n2088);
and (n2124,n356,n320);
and (n2125,n2126,n2127);
xor (n2126,n2123,n2124);
or (n2127,n2128,n2131);
and (n2128,n2129,n2130);
xor (n2129,n2093,n2094);
and (n2130,n349,n320);
and (n2131,n2132,n2133);
xor (n2132,n2129,n2130);
or (n2133,n2134,n2137);
and (n2134,n2135,n2136);
xor (n2135,n2099,n2100);
and (n2136,n78,n320);
and (n2137,n2138,n2139);
xor (n2138,n2135,n2136);
or (n2139,n2140,n2143);
and (n2140,n2141,n2142);
xor (n2141,n2104,n2105);
and (n2142,n56,n320);
and (n2143,n2144,n2145);
xor (n2144,n2141,n2142);
or (n2145,n2146,n2147);
and (n2146,n1462,n1512);
and (n2147,n1461,n1513);
or (n2148,n2149,n2151);
and (n2149,n2150,n315);
xor (n2150,n2114,n2115);
and (n2151,n2152,n2153);
xor (n2152,n2150,n315);
or (n2153,n2154,n2157);
and (n2154,n2155,n2156);
xor (n2155,n2120,n2121);
and (n2156,n356,n313);
and (n2157,n2158,n2159);
xor (n2158,n2155,n2156);
or (n2159,n2160,n2163);
and (n2160,n2161,n2162);
xor (n2161,n2126,n2127);
and (n2162,n349,n313);
and (n2163,n2164,n2165);
xor (n2164,n2161,n2162);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2132,n2133);
and (n2168,n78,n313);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2138,n2139);
and (n2174,n56,n313);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
or (n2177,n2178,n2181);
and (n2178,n2179,n2180);
xor (n2179,n2144,n2145);
and (n2180,n104,n313);
and (n2181,n2182,n2183);
xor (n2182,n2179,n2180);
and (n2183,n1460,n1140);
and (n2184,n312,n340);
or (n2185,n2186,n2189);
and (n2186,n2187,n2188);
xor (n2187,n2152,n2153);
and (n2188,n356,n340);
and (n2189,n2190,n2191);
xor (n2190,n2187,n2188);
or (n2191,n2192,n2195);
and (n2192,n2193,n2194);
xor (n2193,n2158,n2159);
and (n2194,n349,n340);
and (n2195,n2196,n2197);
xor (n2196,n2193,n2194);
or (n2197,n2198,n2201);
and (n2198,n2199,n2200);
xor (n2199,n2164,n2165);
and (n2200,n78,n340);
and (n2201,n2202,n2203);
xor (n2202,n2199,n2200);
or (n2203,n2204,n2207);
and (n2204,n2205,n2206);
xor (n2205,n2170,n2171);
and (n2206,n56,n340);
and (n2207,n2208,n2209);
xor (n2208,n2205,n2206);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2176,n2177);
and (n2212,n104,n340);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
and (n2215,n2216,n2217);
xor (n2216,n2182,n2183);
and (n2217,n88,n340);
and (n2218,n356,n73);
or (n2219,n2220,n2222);
and (n2220,n2221,n348);
xor (n2221,n2190,n2191);
and (n2222,n2223,n2224);
xor (n2223,n2221,n348);
or (n2224,n2225,n2227);
and (n2225,n2226,n459);
xor (n2226,n2196,n2197);
and (n2227,n2228,n2229);
xor (n2228,n2226,n459);
or (n2229,n2230,n2232);
and (n2230,n2231,n620);
xor (n2231,n2202,n2203);
and (n2232,n2233,n2234);
xor (n2233,n2231,n620);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2208,n2209);
and (n2237,n104,n73);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
and (n2240,n2241,n880);
xor (n2241,n2214,n2215);
and (n2242,n349,n66);
or (n2243,n2244,n2247);
and (n2244,n2245,n2246);
xor (n2245,n2223,n2224);
and (n2246,n78,n66);
and (n2247,n2248,n2249);
xor (n2248,n2245,n2246);
or (n2249,n2250,n2253);
and (n2250,n2251,n2252);
xor (n2251,n2228,n2229);
and (n2252,n56,n66);
and (n2253,n2254,n2255);
xor (n2254,n2251,n2252);
or (n2255,n2256,n2259);
and (n2256,n2257,n2258);
xor (n2257,n2233,n2234);
and (n2258,n104,n66);
and (n2259,n2260,n2261);
xor (n2260,n2257,n2258);
and (n2261,n2262,n2263);
xor (n2262,n2239,n2240);
and (n2263,n88,n66);
or (n2264,n2265,n2267);
and (n2265,n2266,n55);
xor (n2266,n2248,n2249);
and (n2267,n2268,n2269);
xor (n2268,n2266,n55);
or (n2269,n2270,n2272);
and (n2270,n2271,n469);
xor (n2271,n2254,n2255);
and (n2272,n2273,n2274);
xor (n2273,n2271,n469);
and (n2274,n2275,n627);
xor (n2275,n2260,n2261);
and (n2276,n56,n95);
or (n2277,n2278,n2281);
and (n2278,n2279,n2280);
xor (n2279,n2268,n2269);
and (n2280,n104,n95);
and (n2281,n2282,n2283);
xor (n2282,n2279,n2280);
and (n2283,n2284,n2285);
xor (n2284,n2273,n2274);
and (n2285,n88,n95);
and (n2286,n2287,n2288);
xor (n2287,n2282,n2283);
and (n2288,n88,n87);
and (n2289,n88,n396);
or (n2290,n2291,n2295,n2335);
and (n2291,n2292,n2293);
xor (n2292,n1970,n32);
not (n2293,n2294);
xor (n2294,n2287,n2288);
and (n2295,n2293,n2296);
or (n2296,n2297,n2301,n2334);
and (n2297,n2298,n2299);
xor (n2298,n1967,n165);
not (n2299,n2300);
xor (n2300,n2284,n2285);
and (n2301,n2299,n2302);
or (n2302,n2303,n2307,n2333);
and (n2303,n2304,n2305);
xor (n2304,n1957,n1958);
not (n2305,n2306);
xor (n2306,n2275,n627);
and (n2307,n2305,n2308);
or (n2308,n2309,n2313,n2332);
and (n2309,n2310,n2311);
xor (n2310,n1942,n636);
not (n2311,n2312);
xor (n2312,n2262,n2263);
and (n2313,n2311,n2314);
or (n2314,n2315,n2319,n2331);
and (n2315,n2316,n2317);
xor (n2316,n1921,n861);
not (n2317,n2318);
xor (n2318,n2241,n880);
and (n2319,n2317,n2320);
or (n2320,n2321,n2325,n2330);
and (n2321,n2322,n2323);
xor (n2322,n1894,n847);
not (n2323,n2324);
xor (n2324,n2216,n2217);
and (n2325,n2323,n2326);
or (n2326,n2327,n2328,n2329);
and (n2327,n1402,n1458);
and (n2328,n1458,n1516);
and (n2329,n1402,n1516);
and (n2330,n2322,n2326);
and (n2331,n2316,n2320);
and (n2332,n2310,n2314);
and (n2333,n2304,n2308);
and (n2334,n2298,n2302);
and (n2335,n2292,n2296);
or (n2336,n2337,n2340,n2371);
and (n2337,n2338,n1616);
xor (n2338,n2339,n2296);
xor (n2339,n2292,n2293);
and (n2340,n1616,n2341);
or (n2341,n2342,n2345,n2370);
and (n2342,n2343,n1606);
xor (n2343,n2344,n2302);
xor (n2344,n2298,n2299);
and (n2345,n1606,n2346);
or (n2346,n2347,n2350,n2369);
and (n2347,n2348,n1604);
xor (n2348,n2349,n2308);
xor (n2349,n2304,n2305);
and (n2350,n1604,n2351);
or (n2351,n2352,n2355,n2368);
and (n2352,n2353,n1380);
xor (n2353,n2354,n2314);
xor (n2354,n2310,n2311);
and (n2355,n1380,n2356);
or (n2356,n2357,n2360,n2367);
and (n2357,n2358,n1600);
xor (n2358,n2359,n2320);
xor (n2359,n2316,n2317);
and (n2360,n1600,n2361);
or (n2361,n2362,n2365,n2366);
and (n2362,n2363,n1391);
xor (n2363,n2364,n2326);
xor (n2364,n2322,n2323);
and (n2365,n1391,n1398);
and (n2366,n2363,n1398);
and (n2367,n2358,n2361);
and (n2368,n2353,n2356);
and (n2369,n2348,n2351);
and (n2370,n2343,n2346);
and (n2371,n2338,n2341);
endmodule
