module top (out,n12,n17,n19,n20,n22,n26,n29,n35,n53
        ,n67,n68,n69,n70,n71,n72,n73,n74,n78,n79
        ,n80,n84,n86,n88,n125,n127,n128,n129,n140,n141
        ,n142,n143,n155,n156,n157,n158,n171,n172,n173,n174
        ,n180,n182,n183,n186,n188,n191,n193,n194,n195,n275
        ,n381,n384,n386,n540,n542,n543,n546,n549,n550,n551
        ,n552,n555,n557,n561,n572,n573,n590,n593,n595,n596
        ,n598,n602,n608,n611,n613,n615,n619,n622,n624,n626
        ,n630,n633,n635,n637,n639,n647,n650,n652,n654,n658
        ,n661,n663,n665,n669,n672,n674,n676,n680,n683,n685
        ,n687,n695,n698,n700,n702,n706,n709,n711,n713,n717
        ,n720,n722,n724,n728,n731,n733,n735,n744,n747,n749
        ,n751,n765,n768,n770,n772,n791,n794,n796,n798,n807
        ,n810,n812,n814,n828,n831,n833,n835,n858,n861,n863
        ,n865,n881,n884,n886,n888,n933,n936,n938,n940,n944
        ,n947,n949,n951,n955,n958,n960,n962,n966,n969,n971
        ,n973,n982,n985,n987,n989,n993,n996,n998,n1000,n1004
        ,n1007,n1009,n1011,n1015,n1018,n1020,n1022,n1030,n1033,n1035
        ,n1037,n1041,n1044,n1046,n1048,n1052,n1055,n1057,n1059,n1063
        ,n1066,n1068,n1070,n1295,n1298,n1300,n1302,n1311,n1314,n1316
        ,n1318,n1327,n1330,n1332,n1334,n1343,n1346,n1348,n1350,n1359
        ,n1362,n1364,n1366,n1375,n1378,n1380,n1382,n1392,n1395,n1397
        ,n1399,n1407,n1410,n1412,n1414,n1822,n1825,n1827,n1829,n1839
        ,n1842,n1844,n1846,n1856,n1859,n1861,n1863,n1881,n1884,n1886
        ,n1888,n1908,n1911,n1913,n1915,n1934,n1937,n1939,n1941,n1963
        ,n1966,n1968,n1970,n1982,n1985,n1987,n1989,n2159,n2162,n2164
        ,n2166,n2175,n2178,n2180,n2182,n2191,n2194,n2196,n2198,n2207
        ,n2210,n2212,n2214,n2223,n2226,n2228,n2230,n2239,n2242,n2244
        ,n2246,n2255,n2258,n2260,n2262,n2270,n2273,n2275,n2277);
output out;
input n12;
input n17;
input n19;
input n20;
input n22;
input n26;
input n29;
input n35;
input n53;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n78;
input n79;
input n80;
input n84;
input n86;
input n88;
input n125;
input n127;
input n128;
input n129;
input n140;
input n141;
input n142;
input n143;
input n155;
input n156;
input n157;
input n158;
input n171;
input n172;
input n173;
input n174;
input n180;
input n182;
input n183;
input n186;
input n188;
input n191;
input n193;
input n194;
input n195;
input n275;
input n381;
input n384;
input n386;
input n540;
input n542;
input n543;
input n546;
input n549;
input n550;
input n551;
input n552;
input n555;
input n557;
input n561;
input n572;
input n573;
input n590;
input n593;
input n595;
input n596;
input n598;
input n602;
input n608;
input n611;
input n613;
input n615;
input n619;
input n622;
input n624;
input n626;
input n630;
input n633;
input n635;
input n637;
input n639;
input n647;
input n650;
input n652;
input n654;
input n658;
input n661;
input n663;
input n665;
input n669;
input n672;
input n674;
input n676;
input n680;
input n683;
input n685;
input n687;
input n695;
input n698;
input n700;
input n702;
input n706;
input n709;
input n711;
input n713;
input n717;
input n720;
input n722;
input n724;
input n728;
input n731;
input n733;
input n735;
input n744;
input n747;
input n749;
input n751;
input n765;
input n768;
input n770;
input n772;
input n791;
input n794;
input n796;
input n798;
input n807;
input n810;
input n812;
input n814;
input n828;
input n831;
input n833;
input n835;
input n858;
input n861;
input n863;
input n865;
input n881;
input n884;
input n886;
input n888;
input n933;
input n936;
input n938;
input n940;
input n944;
input n947;
input n949;
input n951;
input n955;
input n958;
input n960;
input n962;
input n966;
input n969;
input n971;
input n973;
input n982;
input n985;
input n987;
input n989;
input n993;
input n996;
input n998;
input n1000;
input n1004;
input n1007;
input n1009;
input n1011;
input n1015;
input n1018;
input n1020;
input n1022;
input n1030;
input n1033;
input n1035;
input n1037;
input n1041;
input n1044;
input n1046;
input n1048;
input n1052;
input n1055;
input n1057;
input n1059;
input n1063;
input n1066;
input n1068;
input n1070;
input n1295;
input n1298;
input n1300;
input n1302;
input n1311;
input n1314;
input n1316;
input n1318;
input n1327;
input n1330;
input n1332;
input n1334;
input n1343;
input n1346;
input n1348;
input n1350;
input n1359;
input n1362;
input n1364;
input n1366;
input n1375;
input n1378;
input n1380;
input n1382;
input n1392;
input n1395;
input n1397;
input n1399;
input n1407;
input n1410;
input n1412;
input n1414;
input n1822;
input n1825;
input n1827;
input n1829;
input n1839;
input n1842;
input n1844;
input n1846;
input n1856;
input n1859;
input n1861;
input n1863;
input n1881;
input n1884;
input n1886;
input n1888;
input n1908;
input n1911;
input n1913;
input n1915;
input n1934;
input n1937;
input n1939;
input n1941;
input n1963;
input n1966;
input n1968;
input n1970;
input n1982;
input n1985;
input n1987;
input n1989;
input n2159;
input n2162;
input n2164;
input n2166;
input n2175;
input n2178;
input n2180;
input n2182;
input n2191;
input n2194;
input n2196;
input n2198;
input n2207;
input n2210;
input n2212;
input n2214;
input n2223;
input n2226;
input n2228;
input n2230;
input n2239;
input n2242;
input n2244;
input n2246;
input n2255;
input n2258;
input n2260;
input n2262;
input n2270;
input n2273;
input n2275;
input n2277;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n21;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n75;
wire n76;
wire n77;
wire n81;
wire n82;
wire n83;
wire n85;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n184;
wire n185;
wire n187;
wire n189;
wire n190;
wire n192;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n382;
wire n383;
wire n385;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n541;
wire n544;
wire n545;
wire n547;
wire n548;
wire n553;
wire n554;
wire n556;
wire n558;
wire n559;
wire n560;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n591;
wire n592;
wire n594;
wire n597;
wire n599;
wire n600;
wire n601;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n609;
wire n610;
wire n612;
wire n614;
wire n616;
wire n617;
wire n618;
wire n620;
wire n621;
wire n623;
wire n625;
wire n627;
wire n628;
wire n629;
wire n631;
wire n632;
wire n634;
wire n636;
wire n638;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n648;
wire n649;
wire n651;
wire n653;
wire n655;
wire n656;
wire n657;
wire n659;
wire n660;
wire n662;
wire n664;
wire n666;
wire n667;
wire n668;
wire n670;
wire n671;
wire n673;
wire n675;
wire n677;
wire n678;
wire n679;
wire n681;
wire n682;
wire n684;
wire n686;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n696;
wire n697;
wire n699;
wire n701;
wire n703;
wire n704;
wire n705;
wire n707;
wire n708;
wire n710;
wire n712;
wire n714;
wire n715;
wire n716;
wire n718;
wire n719;
wire n721;
wire n723;
wire n725;
wire n726;
wire n727;
wire n729;
wire n730;
wire n732;
wire n734;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n745;
wire n746;
wire n748;
wire n750;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n766;
wire n767;
wire n769;
wire n771;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n792;
wire n793;
wire n795;
wire n797;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n808;
wire n809;
wire n811;
wire n813;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n829;
wire n830;
wire n832;
wire n834;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n859;
wire n860;
wire n862;
wire n864;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n882;
wire n883;
wire n885;
wire n887;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n934;
wire n935;
wire n937;
wire n939;
wire n941;
wire n942;
wire n943;
wire n945;
wire n946;
wire n948;
wire n950;
wire n952;
wire n953;
wire n954;
wire n956;
wire n957;
wire n959;
wire n961;
wire n963;
wire n964;
wire n965;
wire n967;
wire n968;
wire n970;
wire n972;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n983;
wire n984;
wire n986;
wire n988;
wire n990;
wire n991;
wire n992;
wire n994;
wire n995;
wire n997;
wire n999;
wire n1001;
wire n1002;
wire n1003;
wire n1005;
wire n1006;
wire n1008;
wire n1010;
wire n1012;
wire n1013;
wire n1014;
wire n1016;
wire n1017;
wire n1019;
wire n1021;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1031;
wire n1032;
wire n1034;
wire n1036;
wire n1038;
wire n1039;
wire n1040;
wire n1042;
wire n1043;
wire n1045;
wire n1047;
wire n1049;
wire n1050;
wire n1051;
wire n1053;
wire n1054;
wire n1056;
wire n1058;
wire n1060;
wire n1061;
wire n1062;
wire n1064;
wire n1065;
wire n1067;
wire n1069;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1296;
wire n1297;
wire n1299;
wire n1301;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1312;
wire n1313;
wire n1315;
wire n1317;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1328;
wire n1329;
wire n1331;
wire n1333;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1344;
wire n1345;
wire n1347;
wire n1349;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1360;
wire n1361;
wire n1363;
wire n1365;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1376;
wire n1377;
wire n1379;
wire n1381;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1393;
wire n1394;
wire n1396;
wire n1398;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1408;
wire n1409;
wire n1411;
wire n1413;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1823;
wire n1824;
wire n1826;
wire n1828;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1840;
wire n1841;
wire n1843;
wire n1845;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1857;
wire n1858;
wire n1860;
wire n1862;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1882;
wire n1883;
wire n1885;
wire n1887;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1909;
wire n1910;
wire n1912;
wire n1914;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1935;
wire n1936;
wire n1938;
wire n1940;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1964;
wire n1965;
wire n1967;
wire n1969;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1983;
wire n1984;
wire n1986;
wire n1988;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2160;
wire n2161;
wire n2163;
wire n2165;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2176;
wire n2177;
wire n2179;
wire n2181;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2192;
wire n2193;
wire n2195;
wire n2197;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2208;
wire n2209;
wire n2211;
wire n2213;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2224;
wire n2225;
wire n2227;
wire n2229;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2240;
wire n2241;
wire n2243;
wire n2245;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2256;
wire n2257;
wire n2259;
wire n2261;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2271;
wire n2272;
wire n2274;
wire n2276;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
xor (out,n0,n2690);
xor (n0,n1,n2667);
xor (n1,n2,n2568);
xor (n2,n3,n1812);
xor (n3,n4,n1717);
xor (n4,n5,n1288);
xor (n5,n6,n1072);
wire s0n6,s1n6,notn6;
or (n6,s0n6,s1n6);
not(notn6,n926);
and (s0n6,notn6,1'b0);
and (s1n6,n926,n8);
xor (n8,n9,n737);
wire s0n9,s1n9,notn9;
or (n9,s0n9,s1n9);
not(notn9,n583);
and (s0n9,notn9,1'b0);
and (s1n9,n583,n10);
wire s0n10,s1n10,notn10;
or (n10,s0n10,s1n10);
not(notn10,n566);
and (s0n10,notn10,n11);
and (s1n10,n566,n553);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n13);
and (s0n11,notn11,1'b0);
and (s1n11,n13,n12);
and (n13,n14,n547);
and (n14,n15,n31);
or (n15,n16,n21,n25,n28);
and (n16,n17,n18);
and (n18,n19,n20);
and (n21,n22,n23);
and (n23,n24,n20);
not (n24,n19);
and (n25,n26,n27);
nor (n27,n24,n20);
and (n28,n29,n30);
nor (n30,n19,n20);
and (n31,n32,n546);
not (n32,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n545);
and (s0n33,notn33,n34);
and (s1n33,n545,1'b0);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n175);
and (s0n34,notn34,n35);
and (s1n34,n175,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n538);
and (s0n36,notn36,n37);
and (s1n36,n538,n512);
or (n37,n38,n480,n511,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n38,n39,n479);
or (n39,n40,n478);
or (n40,n41,n477);
or (n41,n42,n475);
or (n42,n43,n474);
or (n43,n44,n472);
or (n44,n45,n470);
nor (n45,n46,n395,n404,n416,n428,n439,n450,n461);
or (n46,1'b0,n47,n389,n393);
and (n47,n48,n388);
wire s0n48,s1n48,notn48;
or (n48,s0n48,s1n48);
not(notn48,n379);
and (s0n48,notn48,n49);
and (s1n48,n379,n287);
wire s0n49,s1n49,notn49;
or (n49,s0n49,s1n49);
not(notn49,n246);
and (s0n49,notn49,1'b0);
and (s1n49,n246,n50);
or (n50,n51,n227,n231,n235,n238,n241,n243,1'b0);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n200,n211,n221);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n89);
and (s0n55,notn55,n56);
and (s1n55,n89,1'b0);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n87);
and (s0n56,notn56,n57);
and (s1n56,n87,n85);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n81);
and (s0n57,notn57,n58);
and (s1n57,n81,n75);
wire s0n58,s1n58,notn58;
or (n58,s0n58,s1n58);
not(notn58,n74);
and (s0n58,notn58,n59);
and (s1n58,n74,1'b0);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n73);
and (s0n59,notn59,n60);
and (s1n59,n73,1'b1);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n72);
and (s0n60,notn60,n61);
and (s1n60,n72,1'b0);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n71);
and (s0n61,notn61,n62);
and (s1n61,n71,1'b1);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n70);
and (s0n62,notn62,n63);
and (s1n62,n70,1'b0);
wire s0n63,s1n63,notn63;
or (n63,s0n63,s1n63);
not(notn63,n69);
and (s0n63,notn63,n64);
and (s1n63,n69,1'b1);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n68);
and (s0n64,notn64,n65);
and (s1n64,n68,1'b0);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n67);
and (s0n65,notn65,n52);
and (s1n65,n67,1'b1);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n80);
and (s0n75,notn75,n76);
and (s1n75,n80,1'b0);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n79);
and (s0n76,notn76,n77);
and (s1n76,n79,1'b1);
not (n77,n78);
or (n81,n82,n84);
or (n82,n83,n78);
or (n83,n80,n79);
not (n85,n86);
or (n87,n86,n88);
not (n89,n90);
or (n90,n91,n198);
or (n91,n92,n196);
or (n92,n93,n190);
or (n93,n94,n189);
or (n94,n95,n185);
or (n95,n96,n184);
or (n96,n97,n179);
or (n97,n98,n178);
or (n98,n99,n177);
or (n99,n100,n175);
or (n100,n101,n169);
or (n101,n102,n168);
or (n102,n103,n167);
or (n103,n104,n166);
or (n104,n105,n165);
or (n105,n106,n164);
or (n106,n107,n163);
or (n107,n108,n162);
or (n108,n109,n159);
or (n109,n110,n153);
or (n110,n111,n152);
or (n111,n112,n151);
or (n112,n113,n150);
or (n113,n114,n149);
or (n114,n115,n148);
or (n115,n116,n146);
or (n116,n117,n144);
or (n117,n118,n138);
or (n118,n119,n137);
or (n119,n120,n136);
or (n120,n121,n135);
or (n121,n122,n134);
or (n122,n123,n132);
or (n123,n124,n130);
nor (n124,n125,n126,n128,n129);
not (n126,n127);
nor (n130,n125,n126,n131,n129);
not (n131,n128);
and (n132,n125,n127,n128,n133);
not (n133,n129);
and (n134,n125,n126,n128,n133);
nor (n135,n125,n127,n131,n129);
and (n136,n125,n126,n128,n129);
and (n137,n125,n127,n128,n129);
nor (n138,n139,n141,n142,n143);
not (n139,n140);
nor (n144,n139,n145,n142,n143);
not (n145,n141);
and (n146,n139,n141,n142,n147);
not (n147,n143);
and (n148,n140,n141,n142,n147);
and (n149,n140,n145,n142,n147);
and (n150,n139,n145,n142,n143);
and (n151,n140,n145,n142,n143);
and (n152,n140,n141,n142,n143);
nor (n153,n154,n156,n157,n158);
not (n154,n155);
and (n159,n155,n156,n160,n161);
not (n160,n157);
not (n161,n158);
and (n162,n154,n156,n160,n161);
and (n163,n155,n156,n157,n161);
nor (n164,n155,n156,n160,n161);
and (n165,n154,n156,n157,n158);
and (n166,n154,n156,n160,n158);
and (n167,n155,n156,n160,n158);
nor (n168,n154,n156,n157,n161);
nor (n169,n170,n172,n173,n174);
not (n170,n171);
nor (n175,n171,n176,n173,n174);
not (n176,n172);
and (n177,n170,n176,n173,n174);
and (n178,n171,n176,n173,n174);
nor (n179,n180,n181,n183);
not (n181,n182);
and (n184,n180,n182,n183);
and (n185,n186,n187);
not (n187,n188);
nor (n189,n186,n187);
nor (n190,n191,n192,n194,n195);
not (n192,n193);
and (n196,n191,n193,n194,n197);
not (n197,n195);
and (n198,n199,n192,n194,n197);
not (n199,n191);
wire s0n200,s1n200,notn200;
or (n200,s0n200,s1n200);
not(notn200,n89);
and (s0n200,notn200,n201);
and (s1n200,n89,1'b0);
wire s0n201,s1n201,notn201;
or (n201,s0n201,s1n201);
not(notn201,n87);
and (s0n201,notn201,n202);
and (s1n201,n87,1'b0);
wire s0n202,s1n202,notn202;
or (n202,s0n202,s1n202);
not(notn202,n81);
and (s0n202,notn202,n203);
and (s1n202,n81,n83);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n74);
and (s0n203,notn203,n204);
and (s1n203,n74,1'b1);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n73);
and (s0n204,notn204,n205);
and (s1n204,n73,1'b1);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n72);
and (s0n205,notn205,n206);
and (s1n205,n72,1'b0);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n71);
and (s0n206,notn206,n207);
and (s1n206,n71,1'b0);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n70);
and (s0n207,notn207,n208);
and (s1n207,n70,1'b1);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n69);
and (s0n208,notn208,n209);
and (s1n208,n69,1'b1);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n68);
and (s0n209,notn209,n210);
and (s1n209,n68,1'b0);
not (n210,n67);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n89);
and (s0n211,notn211,n212);
and (s1n211,n89,1'b0);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n87);
and (s0n212,notn212,n213);
and (s1n212,n87,1'b0);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n81);
and (s0n213,notn213,n214);
and (s1n213,n81,n220);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n74);
and (s0n214,notn214,n215);
and (s1n214,n74,1'b1);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n73);
and (s0n215,notn215,n216);
and (s1n215,n73,1'b1);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n72);
and (s0n216,notn216,n217);
and (s1n216,n72,1'b0);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n71);
and (s0n217,notn217,n218);
and (s1n217,n71,1'b0);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n70);
and (s0n218,notn218,n219);
and (s1n218,n70,1'b0);
not (n219,n69);
not (n220,n83);
not (n221,n222);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n89);
and (s0n222,notn222,n223);
and (s1n222,n89,1'b0);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n87);
and (s0n223,notn223,n224);
and (s1n223,n87,1'b0);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n81);
and (s0n224,notn224,n225);
and (s1n224,n81,1'b0);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n74);
and (s0n225,notn225,n226);
and (s1n225,n74,1'b0);
not (n226,n73);
and (n227,n228,n229);
not (n228,n68);
and (n229,n230,n200,n211,n221);
not (n230,n55);
and (n231,n232,n233);
not (n232,n70);
and (n233,n55,n234,n211,n221);
not (n234,n200);
and (n235,n236,n237);
not (n236,n72);
and (n237,n230,n234,n211,n221);
and (n238,n239,n240);
not (n239,n74);
nor (n240,n230,n234,n211,n222);
and (n241,n77,n242);
nor (n242,n55,n234,n211,n222);
and (n243,n244,n245);
not (n244,n80);
nor (n245,n230,n200,n211,n222);
or (n246,n247,n276);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n274);
and (s0n247,notn247,n248);
and (s1n247,n274,1'b0);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n273);
and (s0n248,notn248,n249);
and (s1n248,n273,n268);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n267);
and (s0n249,notn249,n250);
and (s1n249,n267,n256);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n255);
and (s0n250,notn250,n251);
and (s1n250,n255,n118);
or (n251,n252,n149);
or (n252,n253,n148);
or (n253,n254,n146);
or (n254,n138,n144);
or (n255,n125,n127,n128,n129);
or (n256,1'b0,1'b0,n257,n263,n265);
and (n257,n258,n261);
or (n258,1'b0,1'b0,n259,n179);
and (n259,n260,n182,n183);
not (n260,n180);
and (n261,n170,n176,n173,n262);
not (n262,n174);
and (n263,n186,n264);
and (n264,n171,n176,n173,n262);
or (n265,n266,n177);
or (n266,n169,n175);
or (n267,n171,n172,n173,n174);
or (n268,n269,n168);
or (n269,n270,n166);
or (n270,n271,n163);
or (n271,n272,n162);
or (n272,n153,n159);
or (n273,n155,n156,n157,n158);
not (n274,n275);
wire s0n276,s1n276,notn276;
or (n276,s0n276,s1n276);
not(notn276,n274);
and (s0n276,notn276,n277);
and (s1n276,n274,1'b0);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n273);
and (s0n277,notn277,n278);
and (s1n277,n273,n286);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n267);
and (s0n278,notn278,n279);
and (s1n278,n267,n282);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n255);
and (s0n279,notn279,n280);
and (s1n279,n255,1'b0);
or (n280,n281,n152);
or (n281,n150,n151);
or (n282,1'b0,n178,n283,n285,1'b0);
and (n283,n284,n261);
or (n284,1'b0,n184,n259,1'b0);
and (n285,n188,n264);
or (n286,n165,n167);
not (n287,n288);
nor (n288,n49,n289,n305,n325,n342,n356,n367,n375);
wire s0n289,s1n289,notn289;
or (n289,s0n289,s1n289);
not(notn289,n246);
and (s0n289,notn289,1'b0);
and (s1n289,n246,n290);
or (n290,n291,n293,n295,n297,n299,n301,n303,1'b0);
and (n291,n292,n54);
xnor (n292,n67,n53);
and (n293,n294,n229);
xnor (n294,n69,n68);
and (n295,n296,n233);
xnor (n296,n71,n70);
and (n297,n298,n237);
xnor (n298,n73,n72);
and (n299,n300,n240);
xnor (n300,n84,n74);
and (n301,n302,n242);
xnor (n302,n79,n78);
and (n303,n304,n245);
xnor (n304,n88,n80);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n246);
and (s0n305,notn305,1'b0);
and (s1n305,n246,n306);
or (n306,n307,n310,n313,n316,n319,n322,1'b0,1'b0);
and (n307,n308,n54);
xnor (n308,n68,n309);
or (n309,n67,n53);
and (n310,n311,n229);
xnor (n311,n70,n312);
or (n312,n69,n68);
and (n313,n314,n233);
xnor (n314,n72,n315);
or (n315,n71,n70);
and (n316,n317,n237);
xnor (n317,n74,n318);
or (n318,n73,n72);
and (n319,n320,n240);
xnor (n320,n78,n321);
or (n321,n84,n74);
and (n322,n323,n242);
xnor (n323,n80,n324);
or (n324,n79,n78);
wire s0n325,s1n325,notn325;
or (n325,s0n325,s1n325);
not(notn325,n246);
and (s0n325,notn325,1'b0);
and (s1n325,n246,n326);
or (n326,n327,n330,n333,n336,n339,1'b0,1'b0,1'b0);
and (n327,n328,n54);
xnor (n328,n69,n329);
or (n329,n68,n309);
and (n330,n331,n229);
xnor (n331,n71,n332);
or (n332,n70,n312);
and (n333,n334,n233);
xnor (n334,n73,n335);
or (n335,n72,n315);
and (n336,n337,n237);
xnor (n337,n84,n338);
or (n338,n74,n318);
and (n339,n340,n240);
xnor (n340,n79,n341);
or (n341,n78,n321);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n246);
and (s0n342,notn342,1'b0);
and (s1n342,n246,n343);
or (n343,n344,n347,n350,n353,1'b0,1'b0,1'b0,1'b0);
and (n344,n345,n54);
xnor (n345,n70,n346);
or (n346,n69,n329);
and (n347,n348,n229);
xnor (n348,n72,n349);
or (n349,n71,n332);
and (n350,n351,n233);
xnor (n351,n74,n352);
or (n352,n73,n335);
and (n353,n354,n237);
xnor (n354,n78,n355);
or (n355,n84,n338);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n246);
and (s0n356,notn356,1'b0);
and (s1n356,n246,n357);
or (n357,n358,n361,n364,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n358,n359,n54);
xnor (n359,n71,n360);
or (n360,n70,n346);
and (n361,n362,n229);
xnor (n362,n73,n363);
or (n363,n72,n349);
and (n364,n365,n233);
xnor (n365,n84,n366);
or (n366,n74,n352);
wire s0n367,s1n367,notn367;
or (n367,s0n367,s1n367);
not(notn367,n246);
and (s0n367,notn367,1'b0);
and (s1n367,n246,n368);
or (n368,n369,n372,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n369,n370,n54);
xnor (n370,n72,n371);
or (n371,n71,n360);
and (n372,n373,n229);
xnor (n373,n74,n374);
or (n374,n73,n363);
wire s0n375,s1n375,notn375;
or (n375,s0n375,s1n375);
not(notn375,n246);
and (s0n375,notn375,1'b0);
and (s1n375,n246,n376);
and (n376,n377,n54);
xnor (n377,n73,n378);
or (n378,n72,n371);
nor (n379,n380,n382,n385);
not (n380,n381);
not (n382,n383);
xor (n383,n384,n381);
xor (n385,n386,n387);
and (n387,n384,n381);
and (n388,n247,n276);
and (n389,n390,n391);
xor (n390,n289,n49);
nor (n391,n247,n392);
not (n392,n276);
and (n393,n49,n394);
and (n394,n247,n392);
not (n395,n396);
or (n396,1'b0,n397,n399,n403);
and (n397,n398,n388);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n379);
and (s0n398,notn398,n289);
and (s1n398,n379,1'b0);
and (n399,n400,n391);
xor (n400,n401,n402);
not (n401,n305);
not (n402,n289);
and (n403,n289,n394);
or (n404,1'b0,n405,n407,n415);
and (n405,n406,n388);
wire s0n406,s1n406,notn406;
or (n406,s0n406,s1n406);
not(notn406,n379);
and (s0n406,notn406,n305);
and (s1n406,n379,1'b0);
and (n407,n408,n391);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n49);
and (s0n408,notn408,n409);
and (s1n408,n49,n412);
xor (n409,n410,n411);
not (n410,n325);
and (n411,n401,n402);
xor (n412,n325,n413);
and (n413,n305,n414);
and (n414,n289,n49);
and (n415,n305,n394);
not (n416,n417);
or (n417,1'b0,n418,n420,n427);
and (n418,n419,n388);
wire s0n419,s1n419,notn419;
or (n419,s0n419,s1n419);
not(notn419,n379);
and (s0n419,notn419,n325);
and (s1n419,n379,1'b0);
and (n420,n421,n391);
wire s0n421,s1n421,notn421;
or (n421,s0n421,s1n421);
not(notn421,n49);
and (s0n421,notn421,n422);
and (s1n421,n49,n425);
xor (n422,n423,n424);
not (n423,n342);
and (n424,n410,n411);
xor (n425,n342,n426);
and (n426,n325,n413);
and (n427,n325,n394);
or (n428,1'b0,n429,n431,n438);
and (n429,n430,n388);
wire s0n430,s1n430,notn430;
or (n430,s0n430,s1n430);
not(notn430,n379);
and (s0n430,notn430,n342);
and (s1n430,n379,1'b0);
and (n431,n432,n391);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n49);
and (s0n432,notn432,n433);
and (s1n432,n49,n436);
xor (n433,n434,n435);
not (n434,n356);
and (n435,n423,n424);
xor (n436,n356,n437);
and (n437,n342,n426);
and (n438,n342,n394);
or (n439,1'b0,n440,n442,n449);
and (n440,n441,n388);
wire s0n441,s1n441,notn441;
or (n441,s0n441,s1n441);
not(notn441,n379);
and (s0n441,notn441,n356);
and (s1n441,n379,1'b0);
and (n442,n443,n391);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n49);
and (s0n443,notn443,n444);
and (s1n443,n49,n447);
xor (n444,n445,n446);
not (n445,n367);
and (n446,n434,n435);
xor (n447,n367,n448);
and (n448,n356,n437);
and (n449,n356,n394);
or (n450,1'b0,n451,n453,n460);
and (n451,n452,n388);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n379);
and (s0n452,notn452,n367);
and (s1n452,n379,1'b0);
and (n453,n454,n391);
wire s0n454,s1n454,notn454;
or (n454,s0n454,s1n454);
not(notn454,n49);
and (s0n454,notn454,n455);
and (s1n454,n49,n458);
xor (n455,n456,n457);
not (n456,n375);
and (n457,n445,n446);
xor (n458,n375,n459);
and (n459,n367,n448);
and (n460,n367,n394);
or (n461,1'b0,n462,n464,n469);
and (n462,n463,n388);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n379);
and (s0n463,notn463,n375);
and (s1n463,n379,1'b0);
and (n464,n465,n391);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n49);
and (s0n465,notn465,n466);
and (s1n465,n49,n468);
not (n466,n467);
and (n467,n456,n457);
and (n468,n375,n459);
and (n469,n375,n394);
nor (n470,n471,n395,n404,n416,n428,n439,n450,n461);
not (n471,n46);
nor (n472,n46,n396,n473,n416,n428,n439,n450,n461);
not (n473,n404);
nor (n474,n471,n396,n473,n416,n428,n439,n450,n461);
nor (n475,n46,n395,n473,n417,n476,n439,n450,n461);
not (n476,n428);
nor (n477,n471,n395,n473,n417,n476,n439,n450,n461);
nor (n478,n46,n396,n404,n416,n476,n439,n450,n461);
nor (n479,n471,n396,n404,n416,n476,n439,n450,n461);
or (n480,n481,n496);
or (n481,n482,n495);
or (n482,n483,n494);
or (n483,n484,n493);
or (n484,n485,n492);
or (n485,n486,n491);
or (n486,n487,n490);
or (n487,n488,n489);
nor (n488,n46,n395,n473,n417,n428,n439,n450,n461);
nor (n489,n471,n395,n473,n417,n428,n439,n450,n461);
nor (n490,n46,n396,n404,n416,n428,n439,n450,n461);
nor (n491,n471,n396,n404,n416,n428,n439,n450,n461);
nor (n492,n46,n395,n404,n417,n476,n439,n450,n461);
nor (n493,n471,n395,n404,n417,n476,n439,n450,n461);
nor (n494,n46,n396,n473,n417,n476,n439,n450,n461);
nor (n495,n471,n396,n473,n417,n476,n439,n450,n461);
or (n496,n497,n510);
or (n497,n498,n509);
or (n498,n499,n508);
or (n499,n500,n507);
or (n500,n501,n506);
or (n501,n502,n505);
or (n502,n503,n504);
nor (n503,n46,n395,n473,n416,n428,n439,n450,n461);
nor (n504,n471,n395,n473,n416,n428,n439,n450,n461);
nor (n505,n46,n396,n404,n417,n476,n439,n450,n461);
nor (n506,n471,n396,n404,n417,n476,n439,n450,n461);
nor (n507,n46,n395,n404,n416,n476,n439,n450,n461);
nor (n508,n471,n395,n404,n416,n476,n439,n450,n461);
nor (n509,n46,n396,n473,n416,n476,n439,n450,n461);
nor (n510,n471,n396,n473,n416,n476,n439,n450,n461);
nor (n511,n471,n396,n473,n417,n428,n439,n450,n461);
or (n512,1'b0,n513,n520,n527,n288);
or (n513,n514,n478);
or (n514,n515,n477);
or (n515,n516,n475);
or (n516,n517,n495);
or (n517,n518,n472);
or (n518,n519,n470);
or (n519,n491,n45);
or (n520,n521,n494);
or (n521,n522,n493);
or (n522,n523,n492);
or (n523,n524,n506);
or (n524,n525,n490);
or (n525,n526,n489);
or (n526,n511,n488);
or (n527,n528,n505);
or (n528,n529,n504);
or (n529,n530,n503);
or (n530,n531,n474);
or (n531,n532,n537);
or (n532,n533,n536);
or (n533,n534,n535);
nor (n534,n471,n396,n404,n417,n428,n439,n450,n461);
nor (n535,n46,n395,n404,n417,n428,n439,n450,n461);
nor (n536,n471,n395,n404,n417,n428,n439,n450,n461);
nor (n537,n46,n396,n473,n417,n428,n439,n450,n461);
or (n538,n539,n544);
nor (n539,n540,n541,n543);
not (n541,n542);
and (n544,n540,n542,n543);
nor (n545,n170,n176,n173,n174);
nor (n547,n548,n550,n551,n552);
not (n548,n549);
or (n553,1'b0,n554,n556,n560,n563);
and (n554,n555,n547);
and (n556,n557,n558);
nor (n558,n549,n559,n551,n552);
not (n559,n550);
and (n560,n561,n562);
nor (n562,n548,n559,n551,n552);
and (n563,n12,n564);
and (n564,n548,n559,n551,n565);
not (n565,n552);
and (n566,n31,n567);
not (n567,n568);
wire s0n568,s1n568,notn568;
or (n568,s0n568,s1n568);
not(notn568,n581);
and (s0n568,notn568,n14);
and (s1n568,n581,n569);
or (n569,n570,n574,n577,n579);
and (n570,n17,n571);
and (n571,n572,n573);
and (n574,n22,n575);
and (n575,n576,n573);
not (n576,n572);
and (n577,n26,n578);
nor (n578,n576,n573);
and (n579,n29,n580);
nor (n580,n572,n573);
and (n581,n32,n582);
not (n582,n546);
and (n583,n584,n640);
not (n584,n585);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n31);
and (s0n585,notn585,1'b0);
and (s1n585,n31,n586);
wire s0n586,s1n586,notn586;
or (n586,s0n586,s1n586);
not(notn586,n639);
and (s0n586,notn586,n587);
and (s1n586,n639,n630);
or (n587,n588,n606,n617,n628);
and (n588,n589,n18);
wire s0n589,s1n589,notn589;
or (n589,s0n589,s1n589);
not(notn589,n568);
and (s0n589,notn589,n590);
and (s1n589,n568,n591);
or (n591,n592,n597,n601,n604);
and (n592,n593,n594);
nor (n594,n595,n596);
and (n597,n598,n599);
nor (n599,n600,n596);
not (n600,n595);
and (n601,n602,n603);
and (n603,n600,n596);
and (n604,n590,n605);
and (n605,n595,n596);
and (n606,n607,n23);
wire s0n607,s1n607,notn607;
or (n607,s0n607,s1n607);
not(notn607,n568);
and (s0n607,notn607,n608);
and (s1n607,n568,n609);
or (n609,n610,n612,n614,n616);
and (n610,n611,n594);
and (n612,n613,n599);
and (n614,n615,n603);
and (n616,n608,n605);
and (n617,n618,n27);
wire s0n618,s1n618,notn618;
or (n618,s0n618,s1n618);
not(notn618,n568);
and (s0n618,notn618,n619);
and (s1n618,n568,n620);
or (n620,n621,n623,n625,n627);
and (n621,n622,n594);
and (n623,n624,n599);
and (n625,n626,n603);
and (n627,n619,n605);
and (n628,n629,n30);
wire s0n629,s1n629,notn629;
or (n629,s0n629,s1n629);
not(notn629,n568);
and (s0n629,notn629,n630);
and (s1n629,n568,n631);
or (n631,n632,n634,n636,n638);
and (n632,n633,n594);
and (n634,n635,n599);
and (n636,n637,n603);
and (n638,n630,n605);
and (n640,n641,n689);
not (n641,n642);
wire s0n642,s1n642,notn642;
or (n642,s0n642,s1n642);
not(notn642,n31);
and (s0n642,notn642,1'b0);
and (s1n642,n31,n643);
wire s0n643,s1n643,notn643;
or (n643,s0n643,s1n643);
not(notn643,n639);
and (s0n643,notn643,n644);
and (s1n643,n639,n680);
or (n644,n645,n656,n667,n678);
and (n645,n646,n18);
wire s0n646,s1n646,notn646;
or (n646,s0n646,s1n646);
not(notn646,n568);
and (s0n646,notn646,n647);
and (s1n646,n568,n648);
or (n648,n649,n651,n653,n655);
and (n649,n650,n594);
and (n651,n652,n599);
and (n653,n654,n603);
and (n655,n647,n605);
and (n656,n657,n23);
wire s0n657,s1n657,notn657;
or (n657,s0n657,s1n657);
not(notn657,n568);
and (s0n657,notn657,n658);
and (s1n657,n568,n659);
or (n659,n660,n662,n664,n666);
and (n660,n661,n594);
and (n662,n663,n599);
and (n664,n665,n603);
and (n666,n658,n605);
and (n667,n668,n27);
wire s0n668,s1n668,notn668;
or (n668,s0n668,s1n668);
not(notn668,n568);
and (s0n668,notn668,n669);
and (s1n668,n568,n670);
or (n670,n671,n673,n675,n677);
and (n671,n672,n594);
and (n673,n674,n599);
and (n675,n676,n603);
and (n677,n669,n605);
and (n678,n679,n30);
wire s0n679,s1n679,notn679;
or (n679,s0n679,s1n679);
not(notn679,n568);
and (s0n679,notn679,n680);
and (s1n679,n568,n681);
or (n681,n682,n684,n686,n688);
and (n682,n683,n594);
and (n684,n685,n599);
and (n686,n687,n603);
and (n688,n680,n605);
not (n689,n690);
wire s0n690,s1n690,notn690;
or (n690,s0n690,s1n690);
not(notn690,n31);
and (s0n690,notn690,1'b0);
and (s1n690,n31,n691);
wire s0n691,s1n691,notn691;
or (n691,s0n691,s1n691);
not(notn691,n639);
and (s0n691,notn691,n692);
and (s1n691,n639,n728);
or (n692,n693,n704,n715,n726);
and (n693,n694,n18);
wire s0n694,s1n694,notn694;
or (n694,s0n694,s1n694);
not(notn694,n568);
and (s0n694,notn694,n695);
and (s1n694,n568,n696);
or (n696,n697,n699,n701,n703);
and (n697,n698,n594);
and (n699,n700,n599);
and (n701,n702,n603);
and (n703,n695,n605);
and (n704,n705,n23);
wire s0n705,s1n705,notn705;
or (n705,s0n705,s1n705);
not(notn705,n568);
and (s0n705,notn705,n706);
and (s1n705,n568,n707);
or (n707,n708,n710,n712,n714);
and (n708,n709,n594);
and (n710,n711,n599);
and (n712,n713,n603);
and (n714,n706,n605);
and (n715,n716,n27);
wire s0n716,s1n716,notn716;
or (n716,s0n716,s1n716);
not(notn716,n568);
and (s0n716,notn716,n717);
and (s1n716,n568,n718);
or (n718,n719,n721,n723,n725);
and (n719,n720,n594);
and (n721,n722,n599);
and (n723,n724,n603);
and (n725,n717,n605);
and (n726,n727,n30);
wire s0n727,s1n727,notn727;
or (n727,s0n727,s1n727);
not(notn727,n568);
and (s0n727,notn727,n728);
and (s1n727,n568,n729);
or (n729,n730,n732,n734,n736);
and (n730,n731,n594);
and (n732,n733,n599);
and (n734,n735,n603);
and (n736,n728,n605);
or (n737,n738,n777);
and (n738,n739,n778);
xor (n739,n740,n755);
xor (n740,n741,n753);
wire s0n741,s1n741,notn741;
or (n741,s0n741,s1n741);
not(notn741,n583);
and (s0n741,notn741,1'b0);
and (s1n741,n583,n742);
wire s0n742,s1n742,notn742;
or (n742,s0n742,s1n742);
not(notn742,n566);
and (s0n742,notn742,n743);
and (s1n742,n566,n745);
wire s0n743,s1n743,notn743;
or (n743,s0n743,s1n743);
not(notn743,n13);
and (s0n743,notn743,1'b0);
and (s1n743,n13,n744);
or (n745,1'b0,n746,n748,n750,n752);
and (n746,n747,n547);
and (n748,n749,n558);
and (n750,n751,n562);
and (n752,n744,n564);
wire s0n753,s1n753,notn753;
or (n753,s0n753,s1n753);
not(notn753,n754);
and (s0n753,notn753,1'b0);
and (s1n753,n754,n10);
xor (n754,n584,n640);
or (n755,n756,n777);
and (n756,n757,n774);
xor (n757,n758,n759);
wire s0n758,s1n758,notn758;
or (n758,s0n758,s1n758);
not(notn758,n754);
and (s0n758,notn758,1'b0);
and (s1n758,n754,n742);
xor (n759,n760,n762);
wire s0n760,s1n760,notn760;
or (n760,s0n760,s1n760);
not(notn760,n761);
and (s0n760,notn760,1'b0);
and (s1n760,n761,n10);
xor (n761,n641,n689);
wire s0n762,s1n762,notn762;
or (n762,s0n762,s1n762);
not(notn762,n583);
and (s0n762,notn762,1'b0);
and (s1n762,n583,n763);
wire s0n763,s1n763,notn763;
or (n763,s0n763,s1n763);
not(notn763,n566);
and (s0n763,notn763,n764);
and (s1n763,n566,n766);
wire s0n764,s1n764,notn764;
or (n764,s0n764,s1n764);
not(notn764,n13);
and (s0n764,notn764,1'b0);
and (s1n764,n13,n765);
or (n766,1'b0,n767,n769,n771,n773);
and (n767,n768,n547);
and (n769,n770,n558);
and (n771,n772,n562);
and (n773,n765,n564);
and (n774,n775,n776);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n761);
and (s0n775,notn775,1'b0);
and (s1n775,n761,n742);
wire s0n776,s1n776,notn776;
or (n776,s0n776,s1n776);
not(notn776,n690);
and (s0n776,notn776,1'b0);
and (s1n776,n690,n10);
and (n777,n758,n759);
nand (n778,n779,n925);
or (n779,n780,n920);
nor (n780,n781,n919);
and (n781,n782,n908);
nand (n782,n783,n907);
or (n783,n784,n841);
not (n784,n785);
or (n785,n786,n819);
xor (n786,n787,n816);
xor (n787,n788,n800);
wire s0n788,s1n788,notn788;
or (n788,s0n788,s1n788);
not(notn788,n754);
and (s0n788,notn788,1'b0);
and (s1n788,n754,n789);
wire s0n789,s1n789,notn789;
or (n789,s0n789,s1n789);
not(notn789,n566);
and (s0n789,notn789,n790);
and (s1n789,n566,n792);
wire s0n790,s1n790,notn790;
or (n790,s0n790,s1n790);
not(notn790,n13);
and (s0n790,notn790,1'b0);
and (s1n790,n13,n791);
or (n792,1'b0,n793,n795,n797,n799);
and (n793,n794,n547);
and (n795,n796,n558);
and (n797,n798,n562);
and (n799,n791,n564);
xor (n800,n801,n804);
xor (n801,n802,n803);
wire s0n802,s1n802,notn802;
or (n802,s0n802,s1n802);
not(notn802,n761);
and (s0n802,notn802,1'b0);
and (s1n802,n761,n763);
wire s0n803,s1n803,notn803;
or (n803,s0n803,s1n803);
not(notn803,n690);
and (s0n803,notn803,1'b0);
and (s1n803,n690,n742);
wire s0n804,s1n804,notn804;
or (n804,s0n804,s1n804);
not(notn804,n583);
and (s0n804,notn804,1'b0);
and (s1n804,n583,n805);
wire s0n805,s1n805,notn805;
or (n805,s0n805,s1n805);
not(notn805,n566);
and (s0n805,notn805,n806);
and (s1n805,n566,n808);
wire s0n806,s1n806,notn806;
or (n806,s0n806,s1n806);
not(notn806,n13);
and (s0n806,notn806,1'b0);
and (s1n806,n13,n807);
or (n808,1'b0,n809,n811,n813,n815);
and (n809,n810,n547);
and (n811,n812,n558);
and (n813,n814,n562);
and (n815,n807,n564);
and (n816,n817,n818);
wire s0n817,s1n817,notn817;
or (n817,s0n817,s1n817);
not(notn817,n761);
and (s0n817,notn817,1'b0);
and (s1n817,n761,n789);
wire s0n818,s1n818,notn818;
or (n818,s0n818,s1n818);
not(notn818,n690);
and (s0n818,notn818,1'b0);
and (s1n818,n690,n763);
or (n819,n820,n840);
and (n820,n821,n837);
xor (n821,n822,n823);
wire s0n822,s1n822,notn822;
or (n822,s0n822,s1n822);
not(notn822,n754);
and (s0n822,notn822,1'b0);
and (s1n822,n754,n805);
xor (n823,n824,n825);
xor (n824,n817,n818);
wire s0n825,s1n825,notn825;
or (n825,s0n825,s1n825);
not(notn825,n583);
and (s0n825,notn825,1'b0);
and (s1n825,n583,n826);
wire s0n826,s1n826,notn826;
or (n826,s0n826,s1n826);
not(notn826,n566);
and (s0n826,notn826,n827);
and (s1n826,n566,n829);
wire s0n827,s1n827,notn827;
or (n827,s0n827,s1n827);
not(notn827,n13);
and (s0n827,notn827,1'b0);
and (s1n827,n13,n828);
or (n829,1'b0,n830,n832,n834,n836);
and (n830,n831,n547);
and (n832,n833,n558);
and (n834,n835,n562);
and (n836,n828,n564);
and (n837,n838,n839);
wire s0n838,s1n838,notn838;
or (n838,s0n838,s1n838);
not(notn838,n761);
and (s0n838,notn838,1'b0);
and (s1n838,n761,n805);
wire s0n839,s1n839,notn839;
or (n839,s0n839,s1n839);
not(notn839,n690);
and (s0n839,notn839,1'b0);
and (s1n839,n690,n789);
and (n840,n822,n823);
not (n841,n842);
nand (n842,n843,n903,n906);
nand (n843,n844,n868,n900);
or (n844,n845,n846);
xor (n845,n821,n837);
or (n846,n847,n867);
and (n847,n848,n853);
xor (n848,n849,n850);
wire s0n849,s1n849,notn849;
or (n849,s0n849,s1n849);
not(notn849,n754);
and (s0n849,notn849,1'b0);
and (s1n849,n754,n826);
and (n850,n851,n852);
wire s0n851,s1n851,notn851;
or (n851,s0n851,s1n851);
not(notn851,n761);
and (s0n851,notn851,1'b0);
and (s1n851,n761,n826);
wire s0n852,s1n852,notn852;
or (n852,s0n852,s1n852);
not(notn852,n690);
and (s0n852,notn852,1'b0);
and (s1n852,n690,n805);
xor (n853,n854,n855);
xor (n854,n838,n839);
wire s0n855,s1n855,notn855;
or (n855,s0n855,s1n855);
not(notn855,n583);
and (s0n855,notn855,1'b0);
and (s1n855,n583,n856);
wire s0n856,s1n856,notn856;
or (n856,s0n856,s1n856);
not(notn856,n566);
and (s0n856,notn856,n857);
and (s1n856,n566,n859);
wire s0n857,s1n857,notn857;
or (n857,s0n857,s1n857);
not(notn857,n13);
and (s0n857,notn857,1'b0);
and (s1n857,n13,n858);
or (n859,1'b0,n860,n862,n864,n866);
and (n860,n861,n547);
and (n862,n863,n558);
and (n864,n865,n562);
and (n866,n858,n564);
and (n867,n849,n850);
or (n868,n869,n899);
and (n869,n870,n894);
xor (n870,n871,n874);
and (n871,n872,n873);
wire s0n872,s1n872,notn872;
or (n872,s0n872,s1n872);
not(notn872,n761);
and (s0n872,notn872,1'b0);
and (s1n872,n761,n856);
wire s0n873,s1n873,notn873;
or (n873,s0n873,s1n873);
not(notn873,n690);
and (s0n873,notn873,1'b0);
and (s1n873,n690,n826);
or (n874,n875,n893);
and (n875,n876,n892);
xor (n876,n877,n891);
and (n877,n878,n890);
wire s0n878,s1n878,notn878;
or (n878,s0n878,s1n878);
not(notn878,n761);
and (s0n878,notn878,1'b0);
and (s1n878,n761,n879);
wire s0n879,s1n879,notn879;
or (n879,s0n879,s1n879);
not(notn879,n566);
and (s0n879,notn879,n880);
and (s1n879,n566,n882);
wire s0n880,s1n880,notn880;
or (n880,s0n880,s1n880);
not(notn880,n13);
and (s0n880,notn880,1'b0);
and (s1n880,n13,n881);
or (n882,1'b0,n883,n885,n887,n889);
and (n883,n884,n547);
and (n885,n886,n558);
and (n887,n888,n562);
and (n889,n881,n564);
wire s0n890,s1n890,notn890;
or (n890,s0n890,s1n890);
not(notn890,n690);
and (s0n890,notn890,1'b0);
and (s1n890,n690,n856);
wire s0n891,s1n891,notn891;
or (n891,s0n891,s1n891);
not(notn891,n754);
and (s0n891,notn891,1'b0);
and (s1n891,n754,n879);
xor (n892,n872,n873);
and (n893,n877,n891);
xor (n894,n895,n898);
xor (n895,n896,n897);
wire s0n896,s1n896,notn896;
or (n896,s0n896,s1n896);
not(notn896,n583);
and (s0n896,notn896,1'b0);
and (s1n896,n583,n879);
xor (n897,n851,n852);
wire s0n898,s1n898,notn898;
or (n898,s0n898,s1n898);
not(notn898,n754);
and (s0n898,notn898,1'b0);
and (s1n898,n754,n856);
and (n899,n871,n874);
or (n900,n901,n902);
xor (n901,n848,n853);
and (n902,n895,n898);
nand (n903,n904,n844);
not (n904,n905);
nand (n905,n901,n902);
nand (n906,n845,n846);
nand (n907,n786,n819);
or (n908,n909,n916);
xor (n909,n910,n915);
xor (n910,n911,n912);
wire s0n911,s1n911,notn911;
or (n911,s0n911,s1n911);
not(notn911,n754);
and (s0n911,notn911,1'b0);
and (s1n911,n754,n763);
xor (n912,n913,n914);
xor (n913,n775,n776);
wire s0n914,s1n914,notn914;
or (n914,s0n914,s1n914);
not(notn914,n583);
and (s0n914,notn914,1'b0);
and (s1n914,n583,n789);
and (n915,n802,n803);
or (n916,n917,n918);
and (n917,n787,n816);
and (n918,n788,n800);
and (n919,n909,n916);
nor (n920,n921,n924);
or (n921,n922,n923);
and (n922,n910,n915);
and (n923,n911,n912);
xor (n924,n757,n774);
nand (n925,n921,n924);
and (n926,n927,n975);
not (n927,n928);
wire s0n928,s1n928,notn928;
or (n928,s0n928,s1n928);
not(notn928,n31);
and (s0n928,notn928,1'b0);
and (s1n928,n31,n929);
wire s0n929,s1n929,notn929;
or (n929,s0n929,s1n929);
not(notn929,n639);
and (s0n929,notn929,n930);
and (s1n929,n639,n966);
or (n930,n931,n942,n953,n964);
and (n931,n932,n18);
wire s0n932,s1n932,notn932;
or (n932,s0n932,s1n932);
not(notn932,n568);
and (s0n932,notn932,n933);
and (s1n932,n568,n934);
or (n934,n935,n937,n939,n941);
and (n935,n936,n594);
and (n937,n938,n599);
and (n939,n940,n603);
and (n941,n933,n605);
and (n942,n943,n23);
wire s0n943,s1n943,notn943;
or (n943,s0n943,s1n943);
not(notn943,n568);
and (s0n943,notn943,n944);
and (s1n943,n568,n945);
or (n945,n946,n948,n950,n952);
and (n946,n947,n594);
and (n948,n949,n599);
and (n950,n951,n603);
and (n952,n944,n605);
and (n953,n954,n27);
wire s0n954,s1n954,notn954;
or (n954,s0n954,s1n954);
not(notn954,n568);
and (s0n954,notn954,n955);
and (s1n954,n568,n956);
or (n956,n957,n959,n961,n963);
and (n957,n958,n594);
and (n959,n960,n599);
and (n961,n962,n603);
and (n963,n955,n605);
and (n964,n965,n30);
wire s0n965,s1n965,notn965;
or (n965,s0n965,s1n965);
not(notn965,n568);
and (s0n965,notn965,n966);
and (s1n965,n568,n967);
or (n967,n968,n970,n972,n974);
and (n968,n969,n594);
and (n970,n971,n599);
and (n972,n973,n603);
and (n974,n966,n605);
and (n975,n976,n1024);
not (n976,n977);
wire s0n977,s1n977,notn977;
or (n977,s0n977,s1n977);
not(notn977,n31);
and (s0n977,notn977,1'b0);
and (s1n977,n31,n978);
wire s0n978,s1n978,notn978;
or (n978,s0n978,s1n978);
not(notn978,n639);
and (s0n978,notn978,n979);
and (s1n978,n639,n1015);
or (n979,n980,n991,n1002,n1013);
and (n980,n981,n18);
wire s0n981,s1n981,notn981;
or (n981,s0n981,s1n981);
not(notn981,n568);
and (s0n981,notn981,n982);
and (s1n981,n568,n983);
or (n983,n984,n986,n988,n990);
and (n984,n985,n594);
and (n986,n987,n599);
and (n988,n989,n603);
and (n990,n982,n605);
and (n991,n992,n23);
wire s0n992,s1n992,notn992;
or (n992,s0n992,s1n992);
not(notn992,n568);
and (s0n992,notn992,n993);
and (s1n992,n568,n994);
or (n994,n995,n997,n999,n1001);
and (n995,n996,n594);
and (n997,n998,n599);
and (n999,n1000,n603);
and (n1001,n993,n605);
and (n1002,n1003,n27);
wire s0n1003,s1n1003,notn1003;
or (n1003,s0n1003,s1n1003);
not(notn1003,n568);
and (s0n1003,notn1003,n1004);
and (s1n1003,n568,n1005);
or (n1005,n1006,n1008,n1010,n1012);
and (n1006,n1007,n594);
and (n1008,n1009,n599);
and (n1010,n1011,n603);
and (n1012,n1004,n605);
and (n1013,n1014,n30);
wire s0n1014,s1n1014,notn1014;
or (n1014,s0n1014,s1n1014);
not(notn1014,n568);
and (s0n1014,notn1014,n1015);
and (s1n1014,n568,n1016);
or (n1016,n1017,n1019,n1021,n1023);
and (n1017,n1018,n594);
and (n1019,n1020,n599);
and (n1021,n1022,n603);
and (n1023,n1015,n605);
not (n1024,n1025);
wire s0n1025,s1n1025,notn1025;
or (n1025,s0n1025,s1n1025);
not(notn1025,n31);
and (s0n1025,notn1025,1'b0);
and (s1n1025,n31,n1026);
wire s0n1026,s1n1026,notn1026;
or (n1026,s0n1026,s1n1026);
not(notn1026,n639);
and (s0n1026,notn1026,n1027);
and (s1n1026,n639,n1063);
or (n1027,n1028,n1039,n1050,n1061);
and (n1028,n1029,n18);
wire s0n1029,s1n1029,notn1029;
or (n1029,s0n1029,s1n1029);
not(notn1029,n568);
and (s0n1029,notn1029,n1030);
and (s1n1029,n568,n1031);
or (n1031,n1032,n1034,n1036,n1038);
and (n1032,n1033,n594);
and (n1034,n1035,n599);
and (n1036,n1037,n603);
and (n1038,n1030,n605);
and (n1039,n1040,n23);
wire s0n1040,s1n1040,notn1040;
or (n1040,s0n1040,s1n1040);
not(notn1040,n568);
and (s0n1040,notn1040,n1041);
and (s1n1040,n568,n1042);
or (n1042,n1043,n1045,n1047,n1049);
and (n1043,n1044,n594);
and (n1045,n1046,n599);
and (n1047,n1048,n603);
and (n1049,n1041,n605);
and (n1050,n1051,n27);
wire s0n1051,s1n1051,notn1051;
or (n1051,s0n1051,s1n1051);
not(notn1051,n568);
and (s0n1051,notn1051,n1052);
and (s1n1051,n568,n1053);
or (n1053,n1054,n1056,n1058,n1060);
and (n1054,n1055,n594);
and (n1056,n1057,n599);
and (n1058,n1059,n603);
and (n1060,n1052,n605);
and (n1061,n1062,n30);
wire s0n1062,s1n1062,notn1062;
or (n1062,s0n1062,s1n1062);
not(notn1062,n568);
and (s0n1062,notn1062,n1063);
and (s1n1062,n568,n1064);
or (n1064,n1065,n1067,n1069,n1071);
and (n1065,n1066,n594);
and (n1067,n1068,n599);
and (n1069,n1070,n603);
and (n1071,n1063,n605);
or (n1072,n1073,n1202,n1287);
and (n1073,n1074,n1079);
xor (n1074,n1075,n1077);
and (n1075,n1076,n926);
xor (n1076,n739,n778);
wire s0n1077,s1n1077,notn1077;
or (n1077,s0n1077,s1n1077);
not(notn1077,n1078);
and (s0n1077,notn1077,1'b0);
and (s1n1077,n1078,n8);
xor (n1078,n927,n975);
and (n1079,n1080,n1082);
wire s0n1080,s1n1080,notn1080;
or (n1080,s0n1080,s1n1080);
not(notn1080,n1081);
and (s0n1080,notn1080,1'b0);
and (s1n1080,n1081,n8);
xor (n1081,n976,n1024);
or (n1082,n1083,n1086,n1201);
and (n1083,n1084,n1085);
and (n1084,n1076,n1081);
wire s0n1085,s1n1085,notn1085;
or (n1085,s0n1085,s1n1085);
not(notn1085,n1025);
and (s0n1085,notn1085,1'b0);
and (s1n1085,n1025,n8);
and (n1086,n1085,n1087);
or (n1087,n1088,n1143,n1200);
and (n1088,n1089,n1142);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n1081);
and (s0n1089,notn1089,1'b0);
and (s1n1089,n1081,n1090);
xor (n1090,n1091,n1110);
xor (n1091,n1092,n1093);
xor (n1092,n762,n758);
xor (n1093,n760,n1094);
or (n1094,n774,n1095,n1109);
and (n1095,n776,n1096);
or (n1096,n915,n1097,n1108);
and (n1097,n803,n1098);
or (n1098,n816,n1099,n1107);
and (n1099,n818,n1100);
or (n1100,n837,n1101,n1106);
and (n1101,n839,n1102);
or (n1102,n850,n1103,n871);
and (n1103,n852,n1104);
or (n1104,n871,n1105,n877);
and (n1105,n873,n877);
and (n1106,n838,n1102);
and (n1107,n817,n1100);
and (n1108,n802,n1098);
and (n1109,n775,n1096);
or (n1110,n1111,n1114,n1141);
and (n1111,n1112,n1113);
xor (n1112,n914,n911);
xor (n1113,n913,n1096);
and (n1114,n1113,n1115);
or (n1115,n1116,n1119,n1140);
and (n1116,n1117,n1118);
xor (n1117,n804,n788);
xor (n1118,n801,n1098);
and (n1119,n1118,n1120);
or (n1120,n1121,n1124,n1139);
and (n1121,n1122,n1123);
xor (n1122,n825,n822);
xor (n1123,n824,n1100);
and (n1124,n1123,n1125);
or (n1125,n1126,n1129,n1138);
and (n1126,n1127,n1128);
xor (n1127,n855,n849);
xor (n1128,n854,n1102);
and (n1129,n1128,n1130);
or (n1130,n1131,n1134,n1137);
and (n1131,n1132,n1133);
xor (n1132,n896,n898);
xor (n1133,n897,n1104);
and (n1134,n1133,n1135);
and (n1135,n891,n1136);
xor (n1136,n892,n877);
and (n1137,n1132,n1135);
and (n1138,n1127,n1130);
and (n1139,n1122,n1125);
and (n1140,n1117,n1120);
and (n1141,n1112,n1115);
and (n1142,n1076,n1025);
and (n1143,n1142,n1144);
or (n1144,n1145,n1151,n1199);
and (n1145,n1146,n1150);
and (n1146,n1147,n1081);
xor (n1147,n1148,n782);
nor (n1148,n1149,n919);
not (n1149,n908);
wire s0n1150,s1n1150,notn1150;
or (n1150,s0n1150,s1n1150);
not(notn1150,n1025);
and (s0n1150,notn1150,1'b0);
and (s1n1150,n1025,n1090);
and (n1151,n1150,n1152);
or (n1152,n1153,n1158,n1198);
and (n1153,n1154,n1157);
and (n1154,n1155,n1081);
xnor (n1155,n842,n1156);
nand (n1156,n785,n907);
and (n1157,n1147,n1025);
and (n1158,n1157,n1159);
or (n1159,n1160,n1165,n1197);
and (n1160,n1161,n1164);
wire s0n1161,s1n1161,notn1161;
or (n1161,s0n1161,s1n1161);
not(notn1161,n1081);
and (s0n1161,notn1161,1'b0);
and (s1n1161,n1081,n1162);
xor (n1162,n1163,n1125);
xor (n1163,n1122,n1123);
and (n1164,n1155,n1025);
and (n1165,n1164,n1166);
or (n1166,n1167,n1172,n1196);
and (n1167,n1168,n1171);
wire s0n1168,s1n1168,notn1168;
or (n1168,s0n1168,s1n1168);
not(notn1168,n1081);
and (s0n1168,notn1168,1'b0);
and (s1n1168,n1081,n1169);
xor (n1169,n1170,n1130);
xor (n1170,n1127,n1128);
wire s0n1171,s1n1171,notn1171;
or (n1171,s0n1171,s1n1171);
not(notn1171,n1025);
and (s0n1171,notn1171,1'b0);
and (s1n1171,n1025,n1162);
and (n1172,n1171,n1173);
or (n1173,n1174,n1178,n1195);
and (n1174,n1175,n1177);
and (n1175,n1176,n1081);
xor (n1176,n870,n894);
wire s0n1177,s1n1177,notn1177;
or (n1177,s0n1177,s1n1177);
not(notn1177,n1025);
and (s0n1177,notn1177,1'b0);
and (s1n1177,n1025,n1169);
and (n1178,n1177,n1179);
or (n1179,n1180,n1184,n1186);
and (n1180,n1181,n1183);
and (n1181,n1182,n1081);
xor (n1182,n876,n892);
and (n1183,n1176,n1025);
and (n1184,n1183,n1185);
or (n1185,n1186,n1190,n1191);
and (n1186,n1187,n1189);
wire s0n1187,s1n1187,notn1187;
or (n1187,s0n1187,s1n1187);
not(notn1187,n1081);
and (s0n1187,notn1187,1'b0);
and (s1n1187,n1081,n1188);
xor (n1188,n878,n890);
and (n1189,n1182,n1025);
and (n1190,n1189,n1191);
and (n1191,n1192,n1194);
wire s0n1192,s1n1192,notn1192;
or (n1192,s0n1192,s1n1192);
not(notn1192,n1081);
and (s0n1192,notn1192,1'b0);
and (s1n1192,n1081,n1193);
wire s0n1193,s1n1193,notn1193;
or (n1193,s0n1193,s1n1193);
not(notn1193,n690);
and (s0n1193,notn1193,1'b0);
and (s1n1193,n690,n879);
wire s0n1194,s1n1194,notn1194;
or (n1194,s0n1194,s1n1194);
not(notn1194,n1025);
and (s0n1194,notn1194,1'b0);
and (s1n1194,n1025,n1188);
and (n1195,n1175,n1179);
and (n1196,n1168,n1173);
and (n1197,n1161,n1166);
and (n1198,n1154,n1159);
and (n1199,n1146,n1152);
and (n1200,n1089,n1144);
and (n1201,n1084,n1087);
and (n1202,n1079,n1203);
or (n1203,n1204,n1209,n1286);
and (n1204,n1205,n1208);
xor (n1205,n1206,n1207);
wire s0n1206,s1n1206,notn1206;
or (n1206,s0n1206,s1n1206);
not(notn1206,n926);
and (s0n1206,notn1206,1'b0);
and (s1n1206,n926,n1090);
and (n1207,n1076,n1078);
xor (n1208,n1080,n1082);
and (n1209,n1208,n1210);
or (n1210,n1211,n1217,n1285);
and (n1211,n1212,n1215);
xor (n1212,n1213,n1214);
and (n1213,n1147,n926);
wire s0n1214,s1n1214,notn1214;
or (n1214,s0n1214,s1n1214);
not(notn1214,n1078);
and (s0n1214,notn1214,1'b0);
and (s1n1214,n1078,n1090);
xor (n1215,n1216,n1087);
xor (n1216,n1084,n1085);
and (n1217,n1215,n1218);
or (n1218,n1219,n1225,n1284);
and (n1219,n1220,n1223);
xor (n1220,n1221,n1222);
and (n1221,n1155,n926);
and (n1222,n1147,n1078);
xor (n1223,n1224,n1144);
xor (n1224,n1089,n1142);
and (n1225,n1223,n1226);
or (n1226,n1227,n1233,n1283);
and (n1227,n1228,n1231);
xor (n1228,n1229,n1230);
wire s0n1229,s1n1229,notn1229;
or (n1229,s0n1229,s1n1229);
not(notn1229,n926);
and (s0n1229,notn1229,1'b0);
and (s1n1229,n926,n1162);
and (n1230,n1155,n1078);
xor (n1231,n1232,n1152);
xor (n1232,n1146,n1150);
and (n1233,n1231,n1234);
or (n1234,n1235,n1241,n1282);
and (n1235,n1236,n1239);
xor (n1236,n1237,n1238);
wire s0n1237,s1n1237,notn1237;
or (n1237,s0n1237,s1n1237);
not(notn1237,n926);
and (s0n1237,notn1237,1'b0);
and (s1n1237,n926,n1169);
wire s0n1238,s1n1238,notn1238;
or (n1238,s0n1238,s1n1238);
not(notn1238,n1078);
and (s0n1238,notn1238,1'b0);
and (s1n1238,n1078,n1162);
xor (n1239,n1240,n1159);
xor (n1240,n1154,n1157);
and (n1241,n1239,n1242);
or (n1242,n1243,n1249,n1281);
and (n1243,n1244,n1247);
xor (n1244,n1245,n1246);
and (n1245,n1176,n926);
wire s0n1246,s1n1246,notn1246;
or (n1246,s0n1246,s1n1246);
not(notn1246,n1078);
and (s0n1246,notn1246,1'b0);
and (s1n1246,n1078,n1169);
xor (n1247,n1248,n1166);
xor (n1248,n1161,n1164);
and (n1249,n1247,n1250);
or (n1250,n1251,n1257,n1280);
and (n1251,n1252,n1255);
xor (n1252,n1253,n1254);
and (n1253,n1182,n926);
and (n1254,n1176,n1078);
xor (n1255,n1256,n1173);
xor (n1256,n1168,n1171);
and (n1257,n1255,n1258);
or (n1258,n1259,n1265,n1279);
and (n1259,n1260,n1263);
xor (n1260,n1261,n1262);
wire s0n1261,s1n1261,notn1261;
or (n1261,s0n1261,s1n1261);
not(notn1261,n926);
and (s0n1261,notn1261,1'b0);
and (s1n1261,n926,n1188);
and (n1262,n1182,n1078);
xor (n1263,n1264,n1179);
xor (n1264,n1175,n1177);
and (n1265,n1263,n1266);
or (n1266,n1267,n1273,n1278);
and (n1267,n1268,n1271);
xor (n1268,n1269,n1270);
wire s0n1269,s1n1269,notn1269;
or (n1269,s0n1269,s1n1269);
not(notn1269,n926);
and (s0n1269,notn1269,1'b0);
and (s1n1269,n926,n1193);
wire s0n1270,s1n1270,notn1270;
or (n1270,s0n1270,s1n1270);
not(notn1270,n1078);
and (s0n1270,notn1270,1'b0);
and (s1n1270,n1078,n1188);
xor (n1271,n1272,n1185);
xor (n1272,n1181,n1183);
and (n1273,n1271,n1274);
and (n1274,n1275,n1276);
wire s0n1275,s1n1275,notn1275;
or (n1275,s0n1275,s1n1275);
not(notn1275,n1078);
and (s0n1275,notn1275,1'b0);
and (s1n1275,n1078,n1193);
xor (n1276,n1277,n1191);
xor (n1277,n1187,n1189);
and (n1278,n1268,n1274);
and (n1279,n1260,n1266);
and (n1280,n1252,n1258);
and (n1281,n1244,n1250);
and (n1282,n1236,n1242);
and (n1283,n1228,n1234);
and (n1284,n1220,n1226);
and (n1285,n1212,n1218);
and (n1286,n1205,n1210);
and (n1287,n1074,n1203);
xor (n1288,n1289,n1475);
wire s0n1289,s1n1289,notn1289;
or (n1289,s0n1289,s1n1289);
not(notn1289,n926);
and (s0n1289,notn1289,1'b0);
and (s1n1289,n926,n1290);
or (n1290,n1291,n1421,n1474);
and (n1291,n1292,n1304);
and (n1292,n585,n1293);
wire s0n1293,s1n1293,notn1293;
or (n1293,s0n1293,s1n1293);
not(notn1293,n566);
and (s0n1293,notn1293,n1294);
and (s1n1293,n566,n1296);
wire s0n1294,s1n1294,notn1294;
or (n1294,s0n1294,s1n1294);
not(notn1294,n13);
and (s0n1294,notn1294,1'b0);
and (s1n1294,n13,n1295);
or (n1296,1'b0,n1297,n1299,n1301,n1303);
and (n1297,n1298,n547);
and (n1299,n1300,n558);
and (n1301,n1302,n562);
and (n1303,n1295,n564);
and (n1304,n1305,n1306);
wire s0n1305,s1n1305,notn1305;
or (n1305,s0n1305,s1n1305);
not(notn1305,n642);
and (s0n1305,notn1305,1'b0);
and (s1n1305,n642,n1293);
or (n1306,n1307,n1321,n1420);
and (n1307,n1308,n1320);
wire s0n1308,s1n1308,notn1308;
or (n1308,s0n1308,s1n1308);
not(notn1308,n642);
and (s0n1308,notn1308,1'b0);
and (s1n1308,n642,n1309);
wire s0n1309,s1n1309,notn1309;
or (n1309,s0n1309,s1n1309);
not(notn1309,n566);
and (s0n1309,notn1309,n1310);
and (s1n1309,n566,n1312);
wire s0n1310,s1n1310,notn1310;
or (n1310,s0n1310,s1n1310);
not(notn1310,n13);
and (s0n1310,notn1310,1'b0);
and (s1n1310,n13,n1311);
or (n1312,1'b0,n1313,n1315,n1317,n1319);
and (n1313,n1314,n547);
and (n1315,n1316,n558);
and (n1317,n1318,n562);
and (n1319,n1311,n564);
wire s0n1320,s1n1320,notn1320;
or (n1320,s0n1320,s1n1320);
not(notn1320,n690);
and (s0n1320,notn1320,1'b0);
and (s1n1320,n690,n1293);
and (n1321,n1320,n1322);
or (n1322,n1323,n1337,n1419);
and (n1323,n1324,n1336);
wire s0n1324,s1n1324,notn1324;
or (n1324,s0n1324,s1n1324);
not(notn1324,n642);
and (s0n1324,notn1324,1'b0);
and (s1n1324,n642,n1325);
wire s0n1325,s1n1325,notn1325;
or (n1325,s0n1325,s1n1325);
not(notn1325,n566);
and (s0n1325,notn1325,n1326);
and (s1n1325,n566,n1328);
wire s0n1326,s1n1326,notn1326;
or (n1326,s0n1326,s1n1326);
not(notn1326,n13);
and (s0n1326,notn1326,1'b0);
and (s1n1326,n13,n1327);
or (n1328,1'b0,n1329,n1331,n1333,n1335);
and (n1329,n1330,n547);
and (n1331,n1332,n558);
and (n1333,n1334,n562);
and (n1335,n1327,n564);
wire s0n1336,s1n1336,notn1336;
or (n1336,s0n1336,s1n1336);
not(notn1336,n690);
and (s0n1336,notn1336,1'b0);
and (s1n1336,n690,n1309);
and (n1337,n1336,n1338);
or (n1338,n1339,n1353,n1418);
and (n1339,n1340,n1352);
wire s0n1340,s1n1340,notn1340;
or (n1340,s0n1340,s1n1340);
not(notn1340,n642);
and (s0n1340,notn1340,1'b0);
and (s1n1340,n642,n1341);
wire s0n1341,s1n1341,notn1341;
or (n1341,s0n1341,s1n1341);
not(notn1341,n566);
and (s0n1341,notn1341,n1342);
and (s1n1341,n566,n1344);
wire s0n1342,s1n1342,notn1342;
or (n1342,s0n1342,s1n1342);
not(notn1342,n13);
and (s0n1342,notn1342,1'b0);
and (s1n1342,n13,n1343);
or (n1344,1'b0,n1345,n1347,n1349,n1351);
and (n1345,n1346,n547);
and (n1347,n1348,n558);
and (n1349,n1350,n562);
and (n1351,n1343,n564);
wire s0n1352,s1n1352,notn1352;
or (n1352,s0n1352,s1n1352);
not(notn1352,n690);
and (s0n1352,notn1352,1'b0);
and (s1n1352,n690,n1325);
and (n1353,n1352,n1354);
or (n1354,n1355,n1369,n1417);
and (n1355,n1356,n1368);
wire s0n1356,s1n1356,notn1356;
or (n1356,s0n1356,s1n1356);
not(notn1356,n642);
and (s0n1356,notn1356,1'b0);
and (s1n1356,n642,n1357);
wire s0n1357,s1n1357,notn1357;
or (n1357,s0n1357,s1n1357);
not(notn1357,n566);
and (s0n1357,notn1357,n1358);
and (s1n1357,n566,n1360);
wire s0n1358,s1n1358,notn1358;
or (n1358,s0n1358,s1n1358);
not(notn1358,n13);
and (s0n1358,notn1358,1'b0);
and (s1n1358,n13,n1359);
or (n1360,1'b0,n1361,n1363,n1365,n1367);
and (n1361,n1362,n547);
and (n1363,n1364,n558);
and (n1365,n1366,n562);
and (n1367,n1359,n564);
wire s0n1368,s1n1368,notn1368;
or (n1368,s0n1368,s1n1368);
not(notn1368,n690);
and (s0n1368,notn1368,1'b0);
and (s1n1368,n690,n1341);
and (n1369,n1368,n1370);
or (n1370,n1371,n1385,n1387);
and (n1371,n1372,n1384);
wire s0n1372,s1n1372,notn1372;
or (n1372,s0n1372,s1n1372);
not(notn1372,n642);
and (s0n1372,notn1372,1'b0);
and (s1n1372,n642,n1373);
wire s0n1373,s1n1373,notn1373;
or (n1373,s0n1373,s1n1373);
not(notn1373,n566);
and (s0n1373,notn1373,n1374);
and (s1n1373,n566,n1376);
wire s0n1374,s1n1374,notn1374;
or (n1374,s0n1374,s1n1374);
not(notn1374,n13);
and (s0n1374,notn1374,1'b0);
and (s1n1374,n13,n1375);
or (n1376,1'b0,n1377,n1379,n1381,n1383);
and (n1377,n1378,n547);
and (n1379,n1380,n558);
and (n1381,n1382,n562);
and (n1383,n1375,n564);
wire s0n1384,s1n1384,notn1384;
or (n1384,s0n1384,s1n1384);
not(notn1384,n690);
and (s0n1384,notn1384,1'b0);
and (s1n1384,n690,n1357);
and (n1385,n1384,n1386);
or (n1386,n1387,n1402,n1403);
and (n1387,n1388,n1401);
not (n1388,n1389);
nand (n1389,n642,n1390);
wire s0n1390,s1n1390,notn1390;
or (n1390,s0n1390,s1n1390);
not(notn1390,n566);
and (s0n1390,notn1390,n1391);
and (s1n1390,n566,n1393);
wire s0n1391,s1n1391,notn1391;
or (n1391,s0n1391,s1n1391);
not(notn1391,n13);
and (s0n1391,notn1391,1'b0);
and (s1n1391,n13,n1392);
or (n1393,1'b0,n1394,n1396,n1398,n1400);
and (n1394,n1395,n547);
and (n1396,n1397,n558);
and (n1398,n1399,n562);
and (n1400,n1392,n564);
wire s0n1401,s1n1401,notn1401;
or (n1401,s0n1401,s1n1401);
not(notn1401,n690);
and (s0n1401,notn1401,1'b0);
and (s1n1401,n690,n1373);
and (n1402,n1401,n1403);
and (n1403,n1404,n1416);
wire s0n1404,s1n1404,notn1404;
or (n1404,s0n1404,s1n1404);
not(notn1404,n642);
and (s0n1404,notn1404,1'b0);
and (s1n1404,n642,n1405);
wire s0n1405,s1n1405,notn1405;
or (n1405,s0n1405,s1n1405);
not(notn1405,n566);
and (s0n1405,notn1405,n1406);
and (s1n1405,n566,n1408);
wire s0n1406,s1n1406,notn1406;
or (n1406,s0n1406,s1n1406);
not(notn1406,n13);
and (s0n1406,notn1406,1'b0);
and (s1n1406,n13,n1407);
or (n1408,1'b0,n1409,n1411,n1413,n1415);
and (n1409,n1410,n547);
and (n1411,n1412,n558);
and (n1413,n1414,n562);
and (n1415,n1407,n564);
wire s0n1416,s1n1416,notn1416;
or (n1416,s0n1416,s1n1416);
not(notn1416,n690);
and (s0n1416,notn1416,1'b0);
and (s1n1416,n690,n1390);
and (n1417,n1356,n1370);
and (n1418,n1340,n1354);
and (n1419,n1324,n1338);
and (n1420,n1308,n1322);
and (n1421,n1304,n1422);
or (n1422,n1423,n1427,n1473);
and (n1423,n1424,n1426);
not (n1424,n1425);
nand (n1425,n585,n1309);
xor (n1426,n1305,n1306);
and (n1427,n1426,n1428);
or (n1428,n1429,n1434,n1472);
and (n1429,n1430,n1432);
not (n1430,n1431);
nand (n1431,n585,n1325);
xor (n1432,n1433,n1322);
xor (n1433,n1308,n1320);
and (n1434,n1432,n1435);
or (n1435,n1436,n1441,n1471);
and (n1436,n1437,n1439);
not (n1437,n1438);
nand (n1438,n585,n1341);
xor (n1439,n1440,n1338);
xor (n1440,n1324,n1336);
and (n1441,n1439,n1442);
or (n1442,n1443,n1448,n1470);
and (n1443,n1444,n1446);
not (n1444,n1445);
nand (n1445,n585,n1357);
xor (n1446,n1447,n1354);
xor (n1447,n1340,n1352);
and (n1448,n1446,n1449);
or (n1449,n1450,n1455,n1469);
and (n1450,n1451,n1453);
not (n1451,n1452);
nand (n1452,n585,n1373);
xor (n1453,n1454,n1370);
xor (n1454,n1356,n1368);
and (n1455,n1453,n1456);
or (n1456,n1457,n1462,n1468);
and (n1457,n1458,n1460);
not (n1458,n1459);
nand (n1459,n585,n1390);
xor (n1460,n1461,n1386);
xor (n1461,n1372,n1384);
and (n1462,n1460,n1463);
and (n1463,n1464,n1466);
not (n1464,n1465);
nand (n1465,n585,n1405);
xor (n1466,n1467,n1403);
xor (n1467,n1388,n1401);
and (n1468,n1458,n1463);
and (n1469,n1451,n1456);
and (n1470,n1444,n1449);
and (n1471,n1437,n1442);
and (n1472,n1430,n1435);
and (n1473,n1424,n1428);
and (n1474,n1292,n1422);
or (n1475,n1476,n1631,n1716);
and (n1476,n1477,n1482);
xor (n1477,n1478,n1481);
wire s0n1478,s1n1478,notn1478;
or (n1478,s0n1478,s1n1478);
not(notn1478,n926);
and (s0n1478,notn1478,1'b0);
and (s1n1478,n926,n1479);
xor (n1479,n1480,n1422);
xor (n1480,n1292,n1304);
wire s0n1481,s1n1481,notn1481;
or (n1481,s0n1481,s1n1481);
not(notn1481,n1078);
and (s0n1481,notn1481,1'b0);
and (s1n1481,n1078,n1290);
and (n1482,n1483,n1484);
wire s0n1483,s1n1483,notn1483;
or (n1483,s0n1483,s1n1483);
not(notn1483,n1081);
and (s0n1483,notn1483,1'b0);
and (s1n1483,n1081,n1290);
or (n1484,n1485,n1488,n1630);
and (n1485,n1486,n1487);
wire s0n1486,s1n1486,notn1486;
or (n1486,s0n1486,s1n1486);
not(notn1486,n1081);
and (s0n1486,notn1486,1'b0);
and (s1n1486,n1081,n1479);
wire s0n1487,s1n1487,notn1487;
or (n1487,s0n1487,s1n1487);
not(notn1487,n1025);
and (s0n1487,notn1487,1'b0);
and (s1n1487,n1025,n1290);
and (n1488,n1487,n1489);
or (n1489,n1490,n1576,n1629);
and (n1490,n1491,n1575);
and (n1491,n1492,n1081);
xor (n1492,n1493,n1506);
xor (n1493,n1494,n1502);
nand (n1494,n1495,n1499);
or (n1495,n1496,n1498);
and (n1496,n1497,n1431);
not (n1497,n1320);
not (n1498,n1308);
or (n1499,n1500,n1501);
not (n1500,n1352);
not (n1501,n1292);
not (n1502,n1503);
xnor (n1503,n1504,n1505);
not (n1504,n1424);
not (n1505,n1305);
or (n1506,n1507,n1574);
and (n1507,n1508,n1520);
xor (n1508,n1509,n1514);
nor (n1509,n1510,n1512);
and (n1510,n1511,n1308);
xor (n1511,n1497,n1431);
and (n1512,n1513,n1498);
not (n1513,n1511);
nand (n1514,n1515,n1517,n1519);
or (n1515,n1431,n1516);
not (n1516,n1340);
or (n1517,n1438,n1518);
not (n1518,n1336);
not (n1519,n1323);
nand (n1520,n1521,n1573);
or (n1521,n1522,n1534);
not (n1522,n1523);
nand (n1523,n1524,n1526);
xor (n1524,n1440,n1525);
not (n1525,n1437);
not (n1526,n1527);
nand (n1527,n1528,n1531,n1533);
or (n1528,n1529,n1530);
not (n1529,n1384);
not (n1530,n1430);
or (n1531,n1525,n1532);
not (n1532,n1356);
not (n1533,n1339);
not (n1534,n1535);
or (n1535,n1536,n1572);
and (n1536,n1537,n1547);
xor (n1537,n1538,n1544);
nand (n1538,n1539,n1541,n1543);
or (n1539,n1438,n1540);
not (n1540,n1401);
or (n1541,n1445,n1542);
not (n1542,n1372);
not (n1543,n1355);
nand (n1544,n1545,n1546);
or (n1545,n1445,n1447);
nand (n1546,n1447,n1445);
or (n1547,n1548,n1571);
and (n1548,n1549,n1558);
xor (n1549,n1550,n1556);
nand (n1550,n1551,n1553,n1555);
not (n1551,n1552);
and (n1552,n1451,n1388);
or (n1553,n1445,n1554);
not (n1554,n1416);
not (n1555,n1371);
xnor (n1556,n1557,n1454);
not (n1557,n1451);
or (n1558,n1559,n1570);
and (n1559,n1560,n1566);
xor (n1560,n1561,n1562);
nor (n1561,n1465,n1540);
xnor (n1562,n1563,n1542);
nand (n1563,n1564,n1565);
or (n1564,n1458,n1529);
nand (n1565,n1458,n1529);
nand (n1566,n1567,n1569);
or (n1567,n1568,n1389);
xnor (n1568,n1540,n1465);
not (n1569,n1403);
and (n1570,n1561,n1562);
and (n1571,n1550,n1556);
and (n1572,n1538,n1544);
or (n1573,n1524,n1526);
and (n1574,n1509,n1514);
wire s0n1575,s1n1575,notn1575;
or (n1575,s0n1575,s1n1575);
not(notn1575,n1025);
and (s0n1575,notn1575,1'b0);
and (s1n1575,n1025,n1479);
and (n1576,n1575,n1577);
or (n1577,n1578,n1582,n1628);
and (n1578,n1579,n1581);
and (n1579,n1580,n1081);
xor (n1580,n1508,n1520);
wire s0n1581,s1n1581,notn1581;
or (n1581,s0n1581,s1n1581);
not(notn1581,n1025);
and (s0n1581,notn1581,1'b0);
and (s1n1581,n1025,n1492);
and (n1582,n1581,n1583);
or (n1583,n1584,n1589,n1627);
and (n1584,n1585,n1588);
wire s0n1585,s1n1585,notn1585;
or (n1585,s0n1585,s1n1585);
not(notn1585,n1081);
and (s0n1585,notn1585,1'b0);
and (s1n1585,n1081,n1586);
xor (n1586,n1587,n1442);
xor (n1587,n1437,n1439);
wire s0n1588,s1n1588,notn1588;
or (n1588,s0n1588,s1n1588);
not(notn1588,n1025);
and (s0n1588,notn1588,1'b0);
and (s1n1588,n1025,n1580);
and (n1589,n1588,n1590);
or (n1590,n1591,n1595,n1626);
and (n1591,n1592,n1594);
and (n1592,n1593,n1081);
xor (n1593,n1537,n1547);
wire s0n1594,s1n1594,notn1594;
or (n1594,s0n1594,s1n1594);
not(notn1594,n1025);
and (s0n1594,notn1594,1'b0);
and (s1n1594,n1025,n1586);
and (n1595,n1594,n1596);
or (n1596,n1597,n1601,n1625);
and (n1597,n1598,n1600);
and (n1598,n1599,n1081);
xor (n1599,n1549,n1558);
wire s0n1600,s1n1600,notn1600;
or (n1600,s0n1600,s1n1600);
not(notn1600,n1025);
and (s0n1600,notn1600,1'b0);
and (s1n1600,n1025,n1593);
and (n1601,n1600,n1602);
or (n1602,n1603,n1607,n1624);
and (n1603,n1604,n1606);
and (n1604,n1605,n1081);
xor (n1605,n1560,n1566);
wire s0n1606,s1n1606,notn1606;
or (n1606,s0n1606,s1n1606);
not(notn1606,n1025);
and (s0n1606,notn1606,1'b0);
and (s1n1606,n1025,n1599);
and (n1607,n1606,n1608);
or (n1608,n1609,n1613,n1615);
and (n1609,n1610,n1612);
wire s0n1610,s1n1610,notn1610;
or (n1610,s0n1610,s1n1610);
not(notn1610,n1081);
and (s0n1610,notn1610,1'b0);
and (s1n1610,n1081,n1611);
xor (n1611,n1464,n1466);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n1025);
and (s0n1612,notn1612,1'b0);
and (s1n1612,n1025,n1605);
and (n1613,n1612,n1614);
or (n1614,n1615,n1619,n1620);
and (n1615,n1616,n1618);
wire s0n1616,s1n1616,notn1616;
or (n1616,s0n1616,s1n1616);
not(notn1616,n1081);
and (s0n1616,notn1616,1'b0);
and (s1n1616,n1081,n1617);
xor (n1617,n1404,n1416);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n1025);
and (s0n1618,notn1618,1'b0);
and (s1n1618,n1025,n1611);
and (n1619,n1618,n1620);
and (n1620,n1621,n1623);
wire s0n1621,s1n1621,notn1621;
or (n1621,s0n1621,s1n1621);
not(notn1621,n1081);
and (s0n1621,notn1621,1'b0);
and (s1n1621,n1081,n1622);
wire s0n1622,s1n1622,notn1622;
or (n1622,s0n1622,s1n1622);
not(notn1622,n690);
and (s0n1622,notn1622,1'b0);
and (s1n1622,n690,n1405);
wire s0n1623,s1n1623,notn1623;
or (n1623,s0n1623,s1n1623);
not(notn1623,n1025);
and (s0n1623,notn1623,1'b0);
and (s1n1623,n1025,n1617);
and (n1624,n1604,n1608);
and (n1625,n1598,n1602);
and (n1626,n1592,n1596);
and (n1627,n1585,n1590);
and (n1628,n1579,n1583);
and (n1629,n1491,n1577);
and (n1630,n1486,n1489);
and (n1631,n1482,n1632);
or (n1632,n1633,n1638,n1715);
and (n1633,n1634,n1637);
xor (n1634,n1635,n1636);
and (n1635,n1492,n926);
wire s0n1636,s1n1636,notn1636;
or (n1636,s0n1636,s1n1636);
not(notn1636,n1078);
and (s0n1636,notn1636,1'b0);
and (s1n1636,n1078,n1479);
xor (n1637,n1483,n1484);
and (n1638,n1637,n1639);
or (n1639,n1640,n1646,n1714);
and (n1640,n1641,n1644);
xor (n1641,n1642,n1643);
and (n1642,n1580,n926);
and (n1643,n1492,n1078);
xor (n1644,n1645,n1489);
xor (n1645,n1486,n1487);
and (n1646,n1644,n1647);
or (n1647,n1648,n1654,n1713);
and (n1648,n1649,n1652);
xor (n1649,n1650,n1651);
wire s0n1650,s1n1650,notn1650;
or (n1650,s0n1650,s1n1650);
not(notn1650,n926);
and (s0n1650,notn1650,1'b0);
and (s1n1650,n926,n1586);
and (n1651,n1580,n1078);
xor (n1652,n1653,n1577);
xor (n1653,n1491,n1575);
and (n1654,n1652,n1655);
or (n1655,n1656,n1662,n1712);
and (n1656,n1657,n1660);
xor (n1657,n1658,n1659);
and (n1658,n1593,n926);
wire s0n1659,s1n1659,notn1659;
or (n1659,s0n1659,s1n1659);
not(notn1659,n1078);
and (s0n1659,notn1659,1'b0);
and (s1n1659,n1078,n1586);
xor (n1660,n1661,n1583);
xor (n1661,n1579,n1581);
and (n1662,n1660,n1663);
or (n1663,n1664,n1670,n1711);
and (n1664,n1665,n1668);
xor (n1665,n1666,n1667);
and (n1666,n1599,n926);
and (n1667,n1593,n1078);
xor (n1668,n1669,n1590);
xor (n1669,n1585,n1588);
and (n1670,n1668,n1671);
or (n1671,n1672,n1678,n1710);
and (n1672,n1673,n1676);
xor (n1673,n1674,n1675);
and (n1674,n1605,n926);
and (n1675,n1599,n1078);
xor (n1676,n1677,n1596);
xor (n1677,n1592,n1594);
and (n1678,n1676,n1679);
or (n1679,n1680,n1686,n1709);
and (n1680,n1681,n1684);
xor (n1681,n1682,n1683);
wire s0n1682,s1n1682,notn1682;
or (n1682,s0n1682,s1n1682);
not(notn1682,n926);
and (s0n1682,notn1682,1'b0);
and (s1n1682,n926,n1611);
and (n1683,n1605,n1078);
xor (n1684,n1685,n1602);
xor (n1685,n1598,n1600);
and (n1686,n1684,n1687);
or (n1687,n1688,n1694,n1708);
and (n1688,n1689,n1692);
xor (n1689,n1690,n1691);
and (n1690,n926,n1617);
wire s0n1691,s1n1691,notn1691;
or (n1691,s0n1691,s1n1691);
not(notn1691,n1078);
and (s0n1691,notn1691,1'b0);
and (s1n1691,n1078,n1611);
xor (n1692,n1693,n1608);
xor (n1693,n1604,n1606);
and (n1694,n1692,n1695);
or (n1695,n1696,n1702,n1707);
and (n1696,n1697,n1700);
xor (n1697,n1698,n1699);
wire s0n1698,s1n1698,notn1698;
or (n1698,s0n1698,s1n1698);
not(notn1698,n926);
and (s0n1698,notn1698,1'b0);
and (s1n1698,n926,n1622);
and (n1699,n1078,n1617);
xor (n1700,n1701,n1614);
xor (n1701,n1610,n1612);
and (n1702,n1700,n1703);
and (n1703,n1704,n1705);
wire s0n1704,s1n1704,notn1704;
or (n1704,s0n1704,s1n1704);
not(notn1704,n1078);
and (s0n1704,notn1704,1'b0);
and (s1n1704,n1078,n1622);
xor (n1705,n1706,n1620);
xor (n1706,n1616,n1618);
and (n1707,n1697,n1703);
and (n1708,n1689,n1695);
and (n1709,n1681,n1687);
and (n1710,n1673,n1679);
and (n1711,n1665,n1671);
and (n1712,n1657,n1663);
and (n1713,n1649,n1655);
and (n1714,n1641,n1647);
and (n1715,n1634,n1639);
and (n1716,n1477,n1632);
or (n1717,n1718,n1723,n1811);
and (n1718,n1719,n1721);
xor (n1719,n1720,n1203);
xor (n1720,n1074,n1079);
xor (n1721,n1722,n1632);
xor (n1722,n1477,n1482);
and (n1723,n1721,n1724);
or (n1724,n1725,n1730,n1810);
and (n1725,n1726,n1728);
xor (n1726,n1727,n1210);
xor (n1727,n1205,n1208);
xor (n1728,n1729,n1639);
xor (n1729,n1634,n1637);
and (n1730,n1728,n1731);
or (n1731,n1732,n1737,n1809);
and (n1732,n1733,n1735);
xor (n1733,n1734,n1218);
xor (n1734,n1212,n1215);
xor (n1735,n1736,n1647);
xor (n1736,n1641,n1644);
and (n1737,n1735,n1738);
or (n1738,n1739,n1744,n1808);
and (n1739,n1740,n1742);
xor (n1740,n1741,n1226);
xor (n1741,n1220,n1223);
xor (n1742,n1743,n1655);
xor (n1743,n1649,n1652);
and (n1744,n1742,n1745);
or (n1745,n1746,n1751,n1807);
and (n1746,n1747,n1749);
xor (n1747,n1748,n1234);
xor (n1748,n1228,n1231);
xor (n1749,n1750,n1663);
xor (n1750,n1657,n1660);
and (n1751,n1749,n1752);
or (n1752,n1753,n1758,n1806);
and (n1753,n1754,n1756);
xor (n1754,n1755,n1242);
xor (n1755,n1236,n1239);
xor (n1756,n1757,n1671);
xor (n1757,n1665,n1668);
and (n1758,n1756,n1759);
or (n1759,n1760,n1765,n1805);
and (n1760,n1761,n1763);
xor (n1761,n1762,n1250);
xor (n1762,n1244,n1247);
xor (n1763,n1764,n1679);
xor (n1764,n1673,n1676);
and (n1765,n1763,n1766);
or (n1766,n1767,n1772,n1804);
and (n1767,n1768,n1770);
xor (n1768,n1769,n1258);
xor (n1769,n1252,n1255);
xor (n1770,n1771,n1687);
xor (n1771,n1681,n1684);
and (n1772,n1770,n1773);
or (n1773,n1774,n1779,n1803);
and (n1774,n1775,n1777);
xor (n1775,n1776,n1266);
xor (n1776,n1260,n1263);
xor (n1777,n1778,n1695);
xor (n1778,n1689,n1692);
and (n1779,n1777,n1780);
or (n1780,n1781,n1786,n1802);
and (n1781,n1782,n1784);
xor (n1782,n1783,n1274);
xor (n1783,n1268,n1271);
xor (n1784,n1785,n1703);
xor (n1785,n1697,n1700);
and (n1786,n1784,n1787);
or (n1787,n1788,n1791,n1801);
and (n1788,n1789,n1790);
xor (n1789,n1275,n1276);
xor (n1790,n1704,n1705);
and (n1791,n1790,n1792);
or (n1792,n1793,n1796,n1800);
and (n1793,n1794,n1795);
xor (n1794,n1192,n1194);
xor (n1795,n1621,n1623);
and (n1796,n1795,n1797);
and (n1797,n1798,n1799);
wire s0n1798,s1n1798,notn1798;
or (n1798,s0n1798,s1n1798);
not(notn1798,n1025);
and (s0n1798,notn1798,1'b0);
and (s1n1798,n1025,n1193);
wire s0n1799,s1n1799,notn1799;
or (n1799,s0n1799,s1n1799);
not(notn1799,n1025);
and (s0n1799,notn1799,1'b0);
and (s1n1799,n1025,n1622);
and (n1800,n1794,n1797);
and (n1801,n1789,n1792);
and (n1802,n1782,n1787);
and (n1803,n1775,n1780);
and (n1804,n1768,n1773);
and (n1805,n1761,n1766);
and (n1806,n1754,n1759);
and (n1807,n1747,n1752);
and (n1808,n1740,n1745);
and (n1809,n1733,n1738);
and (n1810,n1726,n1731);
and (n1811,n1719,n1724);
xor (n1812,n1813,n2473);
xor (n1813,n1814,n2151);
or (n1814,n1815,n2083,n2150);
and (n1815,n1816,n2016);
and (n1816,n1817,n928);
xnor (n1817,n1818,n1831);
not (n1818,n1819);
and (n1819,n583,n1820);
wire s0n1820,s1n1820,notn1820;
or (n1820,s0n1820,s1n1820);
not(notn1820,n566);
and (s0n1820,notn1820,n1821);
and (s1n1820,n566,n1823);
wire s0n1821,s1n1821,notn1821;
or (n1821,s0n1821,s1n1821);
not(notn1821,n13);
and (s0n1821,notn1821,1'b0);
and (s1n1821,n13,n1822);
or (n1823,1'b0,n1824,n1826,n1828,n1830);
and (n1824,n1825,n547);
and (n1826,n1827,n558);
and (n1828,n1829,n562);
and (n1830,n1822,n564);
or (n1831,n1832,n1869);
and (n1832,n1833,n1870);
xor (n1833,n1834,n1848);
xor (n1834,n1835,n1836);
and (n1835,n754,n1820);
and (n1836,n583,n1837);
wire s0n1837,s1n1837,notn1837;
or (n1837,s0n1837,s1n1837);
not(notn1837,n566);
and (s0n1837,notn1837,n1838);
and (s1n1837,n566,n1840);
wire s0n1838,s1n1838,notn1838;
or (n1838,s0n1838,s1n1838);
not(notn1838,n13);
and (s0n1838,notn1838,1'b0);
and (s1n1838,n13,n1839);
or (n1840,1'b0,n1841,n1843,n1845,n1847);
and (n1841,n1842,n547);
and (n1843,n1844,n558);
and (n1845,n1846,n562);
and (n1847,n1839,n564);
or (n1848,n1849,n1869);
and (n1849,n1850,n1866);
xor (n1850,n1851,n1865);
xor (n1851,n1852,n1853);
and (n1852,n761,n1820);
and (n1853,n583,n1854);
wire s0n1854,s1n1854,notn1854;
or (n1854,s0n1854,s1n1854);
not(notn1854,n566);
and (s0n1854,notn1854,n1855);
and (s1n1854,n566,n1857);
wire s0n1855,s1n1855,notn1855;
or (n1855,s0n1855,s1n1855);
not(notn1855,n13);
and (s0n1855,notn1855,1'b0);
and (s1n1855,n13,n1856);
or (n1857,1'b0,n1858,n1860,n1862,n1864);
and (n1858,n1859,n547);
and (n1860,n1861,n558);
and (n1862,n1863,n562);
and (n1864,n1856,n564);
and (n1865,n754,n1837);
and (n1866,n1867,n1868);
and (n1867,n761,n1837);
wire s0n1868,s1n1868,notn1868;
or (n1868,s0n1868,s1n1868);
not(notn1868,n690);
and (s0n1868,notn1868,1'b0);
and (s1n1868,n690,n1820);
and (n1869,n1851,n1865);
or (n1870,n1871,n2015);
and (n1871,n1872,n1896);
xor (n1872,n1873,n1895);
or (n1873,n1874,n1894);
and (n1874,n1875,n1891);
xor (n1875,n1876,n1890);
xor (n1876,n1877,n1878);
xor (n1877,n1867,n1868);
and (n1878,n583,n1879);
wire s0n1879,s1n1879,notn1879;
or (n1879,s0n1879,s1n1879);
not(notn1879,n566);
and (s0n1879,notn1879,n1880);
and (s1n1879,n566,n1882);
wire s0n1880,s1n1880,notn1880;
or (n1880,s0n1880,s1n1880);
not(notn1880,n13);
and (s0n1880,notn1880,1'b0);
and (s1n1880,n13,n1881);
or (n1882,1'b0,n1883,n1885,n1887,n1889);
and (n1883,n1884,n547);
and (n1885,n1886,n558);
and (n1887,n1888,n562);
and (n1889,n1881,n564);
and (n1890,n754,n1854);
and (n1891,n1892,n1893);
wire s0n1892,s1n1892,notn1892;
or (n1892,s0n1892,s1n1892);
not(notn1892,n690);
and (s0n1892,notn1892,1'b0);
and (s1n1892,n690,n1837);
and (n1893,n761,n1854);
and (n1894,n1876,n1890);
xor (n1895,n1850,n1866);
or (n1896,n1897,n2014);
and (n1897,n1898,n1922);
xor (n1898,n1899,n1921);
or (n1899,n1900,n1920);
and (n1900,n1901,n1917);
xor (n1901,n1902,n1903);
and (n1902,n754,n1879);
xor (n1903,n1904,n1905);
xor (n1904,n1892,n1893);
and (n1905,n583,n1906);
wire s0n1906,s1n1906,notn1906;
or (n1906,s0n1906,s1n1906);
not(notn1906,n566);
and (s0n1906,notn1906,n1907);
and (s1n1906,n566,n1909);
wire s0n1907,s1n1907,notn1907;
or (n1907,s0n1907,s1n1907);
not(notn1907,n13);
and (s0n1907,notn1907,1'b0);
and (s1n1907,n13,n1908);
or (n1909,1'b0,n1910,n1912,n1914,n1916);
and (n1910,n1911,n547);
and (n1912,n1913,n558);
and (n1914,n1915,n562);
and (n1916,n1908,n564);
and (n1917,n1918,n1919);
wire s0n1918,s1n1918,notn1918;
or (n1918,s0n1918,s1n1918);
not(notn1918,n690);
and (s0n1918,notn1918,1'b0);
and (s1n1918,n690,n1854);
and (n1919,n761,n1879);
and (n1920,n1902,n1903);
xor (n1921,n1875,n1891);
or (n1922,n1923,n2013);
and (n1923,n1924,n1948);
xor (n1924,n1925,n1947);
or (n1925,n1926,n1946);
and (n1926,n1927,n1943);
xor (n1927,n1928,n1929);
and (n1928,n754,n1906);
xor (n1929,n1930,n1931);
xor (n1930,n1918,n1919);
and (n1931,n583,n1932);
wire s0n1932,s1n1932,notn1932;
or (n1932,s0n1932,s1n1932);
not(notn1932,n566);
and (s0n1932,notn1932,n1933);
and (s1n1932,n566,n1935);
wire s0n1933,s1n1933,notn1933;
or (n1933,s0n1933,s1n1933);
not(notn1933,n13);
and (s0n1933,notn1933,1'b0);
and (s1n1933,n13,n1934);
or (n1935,1'b0,n1936,n1938,n1940,n1942);
and (n1936,n1937,n547);
and (n1938,n1939,n558);
and (n1940,n1941,n562);
and (n1942,n1934,n564);
and (n1943,n1944,n1945);
and (n1944,n761,n1906);
wire s0n1945,s1n1945,notn1945;
or (n1945,s0n1945,s1n1945);
not(notn1945,n690);
and (s0n1945,notn1945,1'b0);
and (s1n1945,n690,n1879);
and (n1946,n1928,n1929);
xor (n1947,n1901,n1917);
or (n1948,n1949,n2012);
and (n1949,n1950,n1974);
xor (n1950,n1951,n1973);
or (n1951,n1952,n1972);
and (n1952,n1953,n1958);
xor (n1953,n1954,n1955);
and (n1954,n754,n1932);
and (n1955,n1956,n1957);
wire s0n1956,s1n1956,notn1956;
or (n1956,s0n1956,s1n1956);
not(notn1956,n690);
and (s0n1956,notn1956,1'b0);
and (s1n1956,n690,n1906);
and (n1957,n761,n1932);
xor (n1958,n1959,n1960);
xor (n1959,n1944,n1945);
and (n1960,n583,n1961);
wire s0n1961,s1n1961,notn1961;
or (n1961,s0n1961,s1n1961);
not(notn1961,n566);
and (s0n1961,notn1961,n1962);
and (s1n1961,n566,n1964);
wire s0n1962,s1n1962,notn1962;
or (n1962,s0n1962,s1n1962);
not(notn1962,n13);
and (s0n1962,notn1962,1'b0);
and (s1n1962,n13,n1963);
or (n1964,1'b0,n1965,n1967,n1969,n1971);
and (n1965,n1966,n547);
and (n1967,n1968,n558);
and (n1969,n1970,n562);
and (n1971,n1963,n564);
and (n1972,n1954,n1955);
xor (n1973,n1927,n1943);
or (n1974,n1975,n2011);
and (n1975,n1976,n1994);
xor (n1976,n1977,n1993);
and (n1977,n1978,n1992);
xor (n1978,n1979,n1991);
and (n1979,n583,n1980);
wire s0n1980,s1n1980,notn1980;
or (n1980,s0n1980,s1n1980);
not(notn1980,n566);
and (s0n1980,notn1980,n1981);
and (s1n1980,n566,n1983);
wire s0n1981,s1n1981,notn1981;
or (n1981,s0n1981,s1n1981);
not(notn1981,n13);
and (s0n1981,notn1981,1'b0);
and (s1n1981,n13,n1982);
or (n1983,1'b0,n1984,n1986,n1988,n1990);
and (n1984,n1985,n547);
and (n1986,n1987,n558);
and (n1988,n1989,n562);
and (n1990,n1982,n564);
and (n1991,n754,n1961);
xor (n1992,n1956,n1957);
xor (n1993,n1953,n1958);
or (n1994,n1995,n2010);
and (n1995,n1996,n2009);
xor (n1996,n1997,n2000);
and (n1997,n1998,n1999);
wire s0n1998,s1n1998,notn1998;
or (n1998,s0n1998,s1n1998);
not(notn1998,n690);
and (s0n1998,notn1998,1'b0);
and (s1n1998,n690,n1932);
and (n1999,n761,n1961);
or (n2000,n2001,n2008);
and (n2001,n2002,n2007);
xor (n2002,n2003,n2006);
and (n2003,n2004,n2005);
and (n2004,n761,n1980);
wire s0n2005,s1n2005,notn2005;
or (n2005,s0n2005,s1n2005);
not(notn2005,n690);
and (s0n2005,notn2005,1'b0);
and (s1n2005,n690,n1961);
xor (n2006,n1998,n1999);
and (n2007,n754,n1980);
and (n2008,n2003,n2006);
xor (n2009,n1978,n1992);
and (n2010,n1997,n2000);
and (n2011,n1977,n1993);
and (n2012,n1951,n1973);
and (n2013,n1925,n1947);
and (n2014,n1899,n1921);
and (n2015,n1873,n1895);
and (n2016,n2017,n2018);
and (n2017,n1817,n977);
or (n2018,n2019,n2023,n2082);
and (n2019,n2020,n2022);
and (n2020,n2021,n977);
xor (n2021,n1833,n1870);
and (n2022,n1817,n1025);
and (n2023,n2022,n2024);
or (n2024,n2025,n2029,n2081);
and (n2025,n2026,n2028);
and (n2026,n2027,n977);
xor (n2027,n1872,n1896);
and (n2028,n2021,n1025);
and (n2029,n2028,n2030);
or (n2030,n2031,n2035,n2080);
and (n2031,n2032,n2034);
and (n2032,n2033,n977);
xor (n2033,n1898,n1922);
and (n2034,n2027,n1025);
and (n2035,n2034,n2036);
or (n2036,n2037,n2041,n2079);
and (n2037,n2038,n2040);
and (n2038,n2039,n977);
xor (n2039,n1924,n1948);
and (n2040,n2033,n1025);
and (n2041,n2040,n2042);
or (n2042,n2043,n2047,n2078);
and (n2043,n2044,n2046);
and (n2044,n2045,n977);
xor (n2045,n1950,n1974);
and (n2046,n2039,n1025);
and (n2047,n2046,n2048);
or (n2048,n2049,n2053,n2077);
and (n2049,n2050,n2052);
and (n2050,n2051,n977);
xor (n2051,n1976,n1994);
and (n2052,n2045,n1025);
and (n2053,n2052,n2054);
or (n2054,n2055,n2059,n2076);
and (n2055,n2056,n2058);
and (n2056,n2057,n977);
xor (n2057,n1996,n2009);
and (n2058,n2051,n1025);
and (n2059,n2058,n2060);
or (n2060,n2061,n2065,n2067);
and (n2061,n2062,n2064);
and (n2062,n2063,n977);
xor (n2063,n2002,n2007);
and (n2064,n2057,n1025);
and (n2065,n2064,n2066);
or (n2066,n2067,n2071,n2072);
and (n2067,n2068,n2070);
and (n2068,n2069,n977);
xor (n2069,n2004,n2005);
and (n2070,n2063,n1025);
and (n2071,n2070,n2072);
and (n2072,n2073,n2075);
wire s0n2073,s1n2073,notn2073;
or (n2073,s0n2073,s1n2073);
not(notn2073,n977);
and (s0n2073,notn2073,1'b0);
and (s1n2073,n977,n2074);
wire s0n2074,s1n2074,notn2074;
or (n2074,s0n2074,s1n2074);
not(notn2074,n690);
and (s0n2074,notn2074,1'b0);
and (s1n2074,n690,n1980);
and (n2075,n2069,n1025);
and (n2076,n2056,n2060);
and (n2077,n2050,n2054);
and (n2078,n2044,n2048);
and (n2079,n2038,n2042);
and (n2080,n2032,n2036);
and (n2081,n2026,n2030);
and (n2082,n2020,n2024);
and (n2083,n2016,n2084);
or (n2084,n2085,n2088,n2149);
and (n2085,n2086,n2087);
and (n2086,n2021,n928);
xor (n2087,n2017,n2018);
and (n2088,n2087,n2089);
or (n2089,n2090,n2094,n2148);
and (n2090,n2091,n2092);
and (n2091,n2027,n928);
xor (n2092,n2093,n2024);
xor (n2093,n2020,n2022);
and (n2094,n2092,n2095);
or (n2095,n2096,n2100,n2147);
and (n2096,n2097,n2098);
and (n2097,n2033,n928);
xor (n2098,n2099,n2030);
xor (n2099,n2026,n2028);
and (n2100,n2098,n2101);
or (n2101,n2102,n2106,n2146);
and (n2102,n2103,n2104);
and (n2103,n2039,n928);
xor (n2104,n2105,n2036);
xor (n2105,n2032,n2034);
and (n2106,n2104,n2107);
or (n2107,n2108,n2112,n2145);
and (n2108,n2109,n2110);
and (n2109,n2045,n928);
xor (n2110,n2111,n2042);
xor (n2111,n2038,n2040);
and (n2112,n2110,n2113);
or (n2113,n2114,n2118,n2144);
and (n2114,n2115,n2116);
and (n2115,n2051,n928);
xor (n2116,n2117,n2048);
xor (n2117,n2044,n2046);
and (n2118,n2116,n2119);
or (n2119,n2120,n2124,n2143);
and (n2120,n2121,n2122);
and (n2121,n2057,n928);
xor (n2122,n2123,n2054);
xor (n2123,n2050,n2052);
and (n2124,n2122,n2125);
or (n2125,n2126,n2130,n2142);
and (n2126,n2127,n2128);
and (n2127,n2063,n928);
xor (n2128,n2129,n2060);
xor (n2129,n2056,n2058);
and (n2130,n2128,n2131);
or (n2131,n2132,n2136,n2141);
and (n2132,n2133,n2134);
and (n2133,n2069,n928);
xor (n2134,n2135,n2066);
xor (n2135,n2062,n2064);
and (n2136,n2134,n2137);
and (n2137,n2138,n2139);
wire s0n2138,s1n2138,notn2138;
or (n2138,s0n2138,s1n2138);
not(notn2138,n928);
and (s0n2138,notn2138,1'b0);
and (s1n2138,n928,n2074);
xor (n2139,n2140,n2072);
xor (n2140,n2068,n2070);
and (n2141,n2133,n2137);
and (n2142,n2127,n2131);
and (n2143,n2121,n2125);
and (n2144,n2115,n2119);
and (n2145,n2109,n2113);
and (n2146,n2103,n2107);
and (n2147,n2097,n2101);
and (n2148,n2091,n2095);
and (n2149,n2086,n2089);
and (n2150,n1816,n2084);
or (n2151,n2152,n2405,n2472);
and (n2152,n2153,n2331);
wire s0n2153,s1n2153,notn2153;
or (n2153,s0n2153,s1n2153);
not(notn2153,n928);
and (s0n2153,notn2153,1'b0);
and (s1n2153,n928,n2154);
or (n2154,n2155,n2284,n2330);
and (n2155,n2156,n2168);
wire s0n2156,s1n2156,notn2156;
or (n2156,s0n2156,s1n2156);
not(notn2156,n585);
and (s0n2156,notn2156,1'b0);
and (s1n2156,n585,n2157);
wire s0n2157,s1n2157,notn2157;
or (n2157,s0n2157,s1n2157);
not(notn2157,n566);
and (s0n2157,notn2157,n2158);
and (s1n2157,n566,n2160);
wire s0n2158,s1n2158,notn2158;
or (n2158,s0n2158,s1n2158);
not(notn2158,n13);
and (s0n2158,notn2158,1'b0);
and (s1n2158,n13,n2159);
or (n2160,1'b0,n2161,n2163,n2165,n2167);
and (n2161,n2162,n547);
and (n2163,n2164,n558);
and (n2165,n2166,n562);
and (n2167,n2159,n564);
and (n2168,n2169,n2170);
wire s0n2169,s1n2169,notn2169;
or (n2169,s0n2169,s1n2169);
not(notn2169,n642);
and (s0n2169,notn2169,1'b0);
and (s1n2169,n642,n2157);
or (n2170,n2171,n2185,n2283);
and (n2171,n2172,n2184);
wire s0n2172,s1n2172,notn2172;
or (n2172,s0n2172,s1n2172);
not(notn2172,n642);
and (s0n2172,notn2172,1'b0);
and (s1n2172,n642,n2173);
wire s0n2173,s1n2173,notn2173;
or (n2173,s0n2173,s1n2173);
not(notn2173,n566);
and (s0n2173,notn2173,n2174);
and (s1n2173,n566,n2176);
wire s0n2174,s1n2174,notn2174;
or (n2174,s0n2174,s1n2174);
not(notn2174,n13);
and (s0n2174,notn2174,1'b0);
and (s1n2174,n13,n2175);
or (n2176,1'b0,n2177,n2179,n2181,n2183);
and (n2177,n2178,n547);
and (n2179,n2180,n558);
and (n2181,n2182,n562);
and (n2183,n2175,n564);
wire s0n2184,s1n2184,notn2184;
or (n2184,s0n2184,s1n2184);
not(notn2184,n690);
and (s0n2184,notn2184,1'b0);
and (s1n2184,n690,n2157);
and (n2185,n2184,n2186);
or (n2186,n2187,n2201,n2282);
and (n2187,n2188,n2200);
wire s0n2188,s1n2188,notn2188;
or (n2188,s0n2188,s1n2188);
not(notn2188,n642);
and (s0n2188,notn2188,1'b0);
and (s1n2188,n642,n2189);
wire s0n2189,s1n2189,notn2189;
or (n2189,s0n2189,s1n2189);
not(notn2189,n566);
and (s0n2189,notn2189,n2190);
and (s1n2189,n566,n2192);
wire s0n2190,s1n2190,notn2190;
or (n2190,s0n2190,s1n2190);
not(notn2190,n13);
and (s0n2190,notn2190,1'b0);
and (s1n2190,n13,n2191);
or (n2192,1'b0,n2193,n2195,n2197,n2199);
and (n2193,n2194,n547);
and (n2195,n2196,n558);
and (n2197,n2198,n562);
and (n2199,n2191,n564);
wire s0n2200,s1n2200,notn2200;
or (n2200,s0n2200,s1n2200);
not(notn2200,n690);
and (s0n2200,notn2200,1'b0);
and (s1n2200,n690,n2173);
and (n2201,n2200,n2202);
or (n2202,n2203,n2217,n2281);
and (n2203,n2204,n2216);
wire s0n2204,s1n2204,notn2204;
or (n2204,s0n2204,s1n2204);
not(notn2204,n642);
and (s0n2204,notn2204,1'b0);
and (s1n2204,n642,n2205);
wire s0n2205,s1n2205,notn2205;
or (n2205,s0n2205,s1n2205);
not(notn2205,n566);
and (s0n2205,notn2205,n2206);
and (s1n2205,n566,n2208);
wire s0n2206,s1n2206,notn2206;
or (n2206,s0n2206,s1n2206);
not(notn2206,n13);
and (s0n2206,notn2206,1'b0);
and (s1n2206,n13,n2207);
or (n2208,1'b0,n2209,n2211,n2213,n2215);
and (n2209,n2210,n547);
and (n2211,n2212,n558);
and (n2213,n2214,n562);
and (n2215,n2207,n564);
wire s0n2216,s1n2216,notn2216;
or (n2216,s0n2216,s1n2216);
not(notn2216,n690);
and (s0n2216,notn2216,1'b0);
and (s1n2216,n690,n2189);
and (n2217,n2216,n2218);
or (n2218,n2219,n2233,n2280);
and (n2219,n2220,n2232);
wire s0n2220,s1n2220,notn2220;
or (n2220,s0n2220,s1n2220);
not(notn2220,n642);
and (s0n2220,notn2220,1'b0);
and (s1n2220,n642,n2221);
wire s0n2221,s1n2221,notn2221;
or (n2221,s0n2221,s1n2221);
not(notn2221,n566);
and (s0n2221,notn2221,n2222);
and (s1n2221,n566,n2224);
wire s0n2222,s1n2222,notn2222;
or (n2222,s0n2222,s1n2222);
not(notn2222,n13);
and (s0n2222,notn2222,1'b0);
and (s1n2222,n13,n2223);
or (n2224,1'b0,n2225,n2227,n2229,n2231);
and (n2225,n2226,n547);
and (n2227,n2228,n558);
and (n2229,n2230,n562);
and (n2231,n2223,n564);
wire s0n2232,s1n2232,notn2232;
or (n2232,s0n2232,s1n2232);
not(notn2232,n690);
and (s0n2232,notn2232,1'b0);
and (s1n2232,n690,n2205);
and (n2233,n2232,n2234);
or (n2234,n2235,n2249,n2251);
and (n2235,n2236,n2248);
wire s0n2236,s1n2236,notn2236;
or (n2236,s0n2236,s1n2236);
not(notn2236,n642);
and (s0n2236,notn2236,1'b0);
and (s1n2236,n642,n2237);
wire s0n2237,s1n2237,notn2237;
or (n2237,s0n2237,s1n2237);
not(notn2237,n566);
and (s0n2237,notn2237,n2238);
and (s1n2237,n566,n2240);
wire s0n2238,s1n2238,notn2238;
or (n2238,s0n2238,s1n2238);
not(notn2238,n13);
and (s0n2238,notn2238,1'b0);
and (s1n2238,n13,n2239);
or (n2240,1'b0,n2241,n2243,n2245,n2247);
and (n2241,n2242,n547);
and (n2243,n2244,n558);
and (n2245,n2246,n562);
and (n2247,n2239,n564);
wire s0n2248,s1n2248,notn2248;
or (n2248,s0n2248,s1n2248);
not(notn2248,n690);
and (s0n2248,notn2248,1'b0);
and (s1n2248,n690,n2221);
and (n2249,n2248,n2250);
or (n2250,n2251,n2265,n2266);
and (n2251,n2252,n2264);
wire s0n2252,s1n2252,notn2252;
or (n2252,s0n2252,s1n2252);
not(notn2252,n642);
and (s0n2252,notn2252,1'b0);
and (s1n2252,n642,n2253);
wire s0n2253,s1n2253,notn2253;
or (n2253,s0n2253,s1n2253);
not(notn2253,n566);
and (s0n2253,notn2253,n2254);
and (s1n2253,n566,n2256);
wire s0n2254,s1n2254,notn2254;
or (n2254,s0n2254,s1n2254);
not(notn2254,n13);
and (s0n2254,notn2254,1'b0);
and (s1n2254,n13,n2255);
or (n2256,1'b0,n2257,n2259,n2261,n2263);
and (n2257,n2258,n547);
and (n2259,n2260,n558);
and (n2261,n2262,n562);
and (n2263,n2255,n564);
wire s0n2264,s1n2264,notn2264;
or (n2264,s0n2264,s1n2264);
not(notn2264,n690);
and (s0n2264,notn2264,1'b0);
and (s1n2264,n690,n2237);
and (n2265,n2264,n2266);
and (n2266,n2267,n2279);
wire s0n2267,s1n2267,notn2267;
or (n2267,s0n2267,s1n2267);
not(notn2267,n642);
and (s0n2267,notn2267,1'b0);
and (s1n2267,n642,n2268);
wire s0n2268,s1n2268,notn2268;
or (n2268,s0n2268,s1n2268);
not(notn2268,n566);
and (s0n2268,notn2268,n2269);
and (s1n2268,n566,n2271);
wire s0n2269,s1n2269,notn2269;
or (n2269,s0n2269,s1n2269);
not(notn2269,n13);
and (s0n2269,notn2269,1'b0);
and (s1n2269,n13,n2270);
or (n2271,1'b0,n2272,n2274,n2276,n2278);
and (n2272,n2273,n547);
and (n2274,n2275,n558);
and (n2276,n2277,n562);
and (n2278,n2270,n564);
wire s0n2279,s1n2279,notn2279;
or (n2279,s0n2279,s1n2279);
not(notn2279,n690);
and (s0n2279,notn2279,1'b0);
and (s1n2279,n690,n2253);
and (n2280,n2220,n2234);
and (n2281,n2204,n2218);
and (n2282,n2188,n2202);
and (n2283,n2172,n2186);
and (n2284,n2168,n2285);
or (n2285,n2286,n2289,n2329);
and (n2286,n2287,n2288);
wire s0n2287,s1n2287,notn2287;
or (n2287,s0n2287,s1n2287);
not(notn2287,n585);
and (s0n2287,notn2287,1'b0);
and (s1n2287,n585,n2173);
xor (n2288,n2169,n2170);
and (n2289,n2288,n2290);
or (n2290,n2291,n2295,n2328);
and (n2291,n2292,n2293);
wire s0n2292,s1n2292,notn2292;
or (n2292,s0n2292,s1n2292);
not(notn2292,n585);
and (s0n2292,notn2292,1'b0);
and (s1n2292,n585,n2189);
xor (n2293,n2294,n2186);
xor (n2294,n2172,n2184);
and (n2295,n2293,n2296);
or (n2296,n2297,n2301,n2327);
and (n2297,n2298,n2299);
wire s0n2298,s1n2298,notn2298;
or (n2298,s0n2298,s1n2298);
not(notn2298,n585);
and (s0n2298,notn2298,1'b0);
and (s1n2298,n585,n2205);
xor (n2299,n2300,n2202);
xor (n2300,n2188,n2200);
and (n2301,n2299,n2302);
or (n2302,n2303,n2307,n2326);
and (n2303,n2304,n2305);
wire s0n2304,s1n2304,notn2304;
or (n2304,s0n2304,s1n2304);
not(notn2304,n585);
and (s0n2304,notn2304,1'b0);
and (s1n2304,n585,n2221);
xor (n2305,n2306,n2218);
xor (n2306,n2204,n2216);
and (n2307,n2305,n2308);
or (n2308,n2309,n2313,n2325);
and (n2309,n2310,n2311);
wire s0n2310,s1n2310,notn2310;
or (n2310,s0n2310,s1n2310);
not(notn2310,n585);
and (s0n2310,notn2310,1'b0);
and (s1n2310,n585,n2237);
xor (n2311,n2312,n2234);
xor (n2312,n2220,n2232);
and (n2313,n2311,n2314);
or (n2314,n2315,n2319,n2324);
and (n2315,n2316,n2317);
wire s0n2316,s1n2316,notn2316;
or (n2316,s0n2316,s1n2316);
not(notn2316,n585);
and (s0n2316,notn2316,1'b0);
and (s1n2316,n585,n2253);
xor (n2317,n2318,n2250);
xor (n2318,n2236,n2248);
and (n2319,n2317,n2320);
and (n2320,n2321,n2322);
wire s0n2321,s1n2321,notn2321;
or (n2321,s0n2321,s1n2321);
not(notn2321,n585);
and (s0n2321,notn2321,1'b0);
and (s1n2321,n585,n2268);
xor (n2322,n2323,n2266);
xor (n2323,n2252,n2264);
and (n2324,n2316,n2320);
and (n2325,n2310,n2314);
and (n2326,n2304,n2308);
and (n2327,n2298,n2302);
and (n2328,n2292,n2296);
and (n2329,n2287,n2290);
and (n2330,n2156,n2285);
and (n2331,n2332,n2333);
wire s0n2332,s1n2332,notn2332;
or (n2332,s0n2332,s1n2332);
not(notn2332,n977);
and (s0n2332,notn2332,1'b0);
and (s1n2332,n977,n2154);
or (n2333,n2334,n2339,n2404);
and (n2334,n2335,n2338);
wire s0n2335,s1n2335,notn2335;
or (n2335,s0n2335,s1n2335);
not(notn2335,n977);
and (s0n2335,notn2335,1'b0);
and (s1n2335,n977,n2336);
xor (n2336,n2337,n2285);
xor (n2337,n2156,n2168);
wire s0n2338,s1n2338,notn2338;
or (n2338,s0n2338,s1n2338);
not(notn2338,n1025);
and (s0n2338,notn2338,1'b0);
and (s1n2338,n1025,n2154);
and (n2339,n2338,n2340);
or (n2340,n2341,n2346,n2403);
and (n2341,n2342,n2345);
wire s0n2342,s1n2342,notn2342;
or (n2342,s0n2342,s1n2342);
not(notn2342,n977);
and (s0n2342,notn2342,1'b0);
and (s1n2342,n977,n2343);
xor (n2343,n2344,n2290);
xor (n2344,n2287,n2288);
wire s0n2345,s1n2345,notn2345;
or (n2345,s0n2345,s1n2345);
not(notn2345,n1025);
and (s0n2345,notn2345,1'b0);
and (s1n2345,n1025,n2336);
and (n2346,n2345,n2347);
or (n2347,n2348,n2353,n2402);
and (n2348,n2349,n2352);
wire s0n2349,s1n2349,notn2349;
or (n2349,s0n2349,s1n2349);
not(notn2349,n977);
and (s0n2349,notn2349,1'b0);
and (s1n2349,n977,n2350);
xor (n2350,n2351,n2296);
xor (n2351,n2292,n2293);
wire s0n2352,s1n2352,notn2352;
or (n2352,s0n2352,s1n2352);
not(notn2352,n1025);
and (s0n2352,notn2352,1'b0);
and (s1n2352,n1025,n2343);
and (n2353,n2352,n2354);
or (n2354,n2355,n2360,n2401);
and (n2355,n2356,n2359);
wire s0n2356,s1n2356,notn2356;
or (n2356,s0n2356,s1n2356);
not(notn2356,n977);
and (s0n2356,notn2356,1'b0);
and (s1n2356,n977,n2357);
xor (n2357,n2358,n2302);
xor (n2358,n2298,n2299);
wire s0n2359,s1n2359,notn2359;
or (n2359,s0n2359,s1n2359);
not(notn2359,n1025);
and (s0n2359,notn2359,1'b0);
and (s1n2359,n1025,n2350);
and (n2360,n2359,n2361);
or (n2361,n2362,n2367,n2400);
and (n2362,n2363,n2366);
wire s0n2363,s1n2363,notn2363;
or (n2363,s0n2363,s1n2363);
not(notn2363,n977);
and (s0n2363,notn2363,1'b0);
and (s1n2363,n977,n2364);
xor (n2364,n2365,n2308);
xor (n2365,n2304,n2305);
wire s0n2366,s1n2366,notn2366;
or (n2366,s0n2366,s1n2366);
not(notn2366,n1025);
and (s0n2366,notn2366,1'b0);
and (s1n2366,n1025,n2357);
and (n2367,n2366,n2368);
or (n2368,n2369,n2374,n2399);
and (n2369,n2370,n2373);
wire s0n2370,s1n2370,notn2370;
or (n2370,s0n2370,s1n2370);
not(notn2370,n977);
and (s0n2370,notn2370,1'b0);
and (s1n2370,n977,n2371);
xor (n2371,n2372,n2314);
xor (n2372,n2310,n2311);
wire s0n2373,s1n2373,notn2373;
or (n2373,s0n2373,s1n2373);
not(notn2373,n1025);
and (s0n2373,notn2373,1'b0);
and (s1n2373,n1025,n2364);
and (n2374,n2373,n2375);
or (n2375,n2376,n2381,n2398);
and (n2376,n2377,n2380);
wire s0n2377,s1n2377,notn2377;
or (n2377,s0n2377,s1n2377);
not(notn2377,n977);
and (s0n2377,notn2377,1'b0);
and (s1n2377,n977,n2378);
xor (n2378,n2379,n2320);
xor (n2379,n2316,n2317);
wire s0n2380,s1n2380,notn2380;
or (n2380,s0n2380,s1n2380);
not(notn2380,n1025);
and (s0n2380,notn2380,1'b0);
and (s1n2380,n1025,n2371);
and (n2381,n2380,n2382);
or (n2382,n2383,n2387,n2389);
and (n2383,n2384,n2386);
wire s0n2384,s1n2384,notn2384;
or (n2384,s0n2384,s1n2384);
not(notn2384,n977);
and (s0n2384,notn2384,1'b0);
and (s1n2384,n977,n2385);
xor (n2385,n2321,n2322);
wire s0n2386,s1n2386,notn2386;
or (n2386,s0n2386,s1n2386);
not(notn2386,n1025);
and (s0n2386,notn2386,1'b0);
and (s1n2386,n1025,n2378);
and (n2387,n2386,n2388);
or (n2388,n2389,n2393,n2394);
and (n2389,n2390,n2392);
wire s0n2390,s1n2390,notn2390;
or (n2390,s0n2390,s1n2390);
not(notn2390,n977);
and (s0n2390,notn2390,1'b0);
and (s1n2390,n977,n2391);
xor (n2391,n2267,n2279);
wire s0n2392,s1n2392,notn2392;
or (n2392,s0n2392,s1n2392);
not(notn2392,n1025);
and (s0n2392,notn2392,1'b0);
and (s1n2392,n1025,n2385);
and (n2393,n2392,n2394);
and (n2394,n2395,n2397);
wire s0n2395,s1n2395,notn2395;
or (n2395,s0n2395,s1n2395);
not(notn2395,n977);
and (s0n2395,notn2395,1'b0);
and (s1n2395,n977,n2396);
wire s0n2396,s1n2396,notn2396;
or (n2396,s0n2396,s1n2396);
not(notn2396,n690);
and (s0n2396,notn2396,1'b0);
and (s1n2396,n690,n2268);
wire s0n2397,s1n2397,notn2397;
or (n2397,s0n2397,s1n2397);
not(notn2397,n1025);
and (s0n2397,notn2397,1'b0);
and (s1n2397,n1025,n2391);
and (n2398,n2377,n2382);
and (n2399,n2370,n2375);
and (n2400,n2363,n2368);
and (n2401,n2356,n2361);
and (n2402,n2349,n2354);
and (n2403,n2342,n2347);
and (n2404,n2335,n2340);
and (n2405,n2331,n2406);
or (n2406,n2407,n2410,n2471);
and (n2407,n2408,n2409);
wire s0n2408,s1n2408,notn2408;
or (n2408,s0n2408,s1n2408);
not(notn2408,n928);
and (s0n2408,notn2408,1'b0);
and (s1n2408,n928,n2336);
xor (n2409,n2332,n2333);
and (n2410,n2409,n2411);
or (n2411,n2412,n2416,n2470);
and (n2412,n2413,n2414);
wire s0n2413,s1n2413,notn2413;
or (n2413,s0n2413,s1n2413);
not(notn2413,n928);
and (s0n2413,notn2413,1'b0);
and (s1n2413,n928,n2343);
xor (n2414,n2415,n2340);
xor (n2415,n2335,n2338);
and (n2416,n2414,n2417);
or (n2417,n2418,n2422,n2469);
and (n2418,n2419,n2420);
wire s0n2419,s1n2419,notn2419;
or (n2419,s0n2419,s1n2419);
not(notn2419,n928);
and (s0n2419,notn2419,1'b0);
and (s1n2419,n928,n2350);
xor (n2420,n2421,n2347);
xor (n2421,n2342,n2345);
and (n2422,n2420,n2423);
or (n2423,n2424,n2428,n2468);
and (n2424,n2425,n2426);
wire s0n2425,s1n2425,notn2425;
or (n2425,s0n2425,s1n2425);
not(notn2425,n928);
and (s0n2425,notn2425,1'b0);
and (s1n2425,n928,n2357);
xor (n2426,n2427,n2354);
xor (n2427,n2349,n2352);
and (n2428,n2426,n2429);
or (n2429,n2430,n2434,n2467);
and (n2430,n2431,n2432);
wire s0n2431,s1n2431,notn2431;
or (n2431,s0n2431,s1n2431);
not(notn2431,n928);
and (s0n2431,notn2431,1'b0);
and (s1n2431,n928,n2364);
xor (n2432,n2433,n2361);
xor (n2433,n2356,n2359);
and (n2434,n2432,n2435);
or (n2435,n2436,n2440,n2466);
and (n2436,n2437,n2438);
wire s0n2437,s1n2437,notn2437;
or (n2437,s0n2437,s1n2437);
not(notn2437,n928);
and (s0n2437,notn2437,1'b0);
and (s1n2437,n928,n2371);
xor (n2438,n2439,n2368);
xor (n2439,n2363,n2366);
and (n2440,n2438,n2441);
or (n2441,n2442,n2446,n2465);
and (n2442,n2443,n2444);
wire s0n2443,s1n2443,notn2443;
or (n2443,s0n2443,s1n2443);
not(notn2443,n928);
and (s0n2443,notn2443,1'b0);
and (s1n2443,n928,n2378);
xor (n2444,n2445,n2375);
xor (n2445,n2370,n2373);
and (n2446,n2444,n2447);
or (n2447,n2448,n2452,n2464);
and (n2448,n2449,n2450);
wire s0n2449,s1n2449,notn2449;
or (n2449,s0n2449,s1n2449);
not(notn2449,n928);
and (s0n2449,notn2449,1'b0);
and (s1n2449,n928,n2385);
xor (n2450,n2451,n2382);
xor (n2451,n2377,n2380);
and (n2452,n2450,n2453);
or (n2453,n2454,n2458,n2463);
and (n2454,n2455,n2456);
wire s0n2455,s1n2455,notn2455;
or (n2455,s0n2455,s1n2455);
not(notn2455,n928);
and (s0n2455,notn2455,1'b0);
and (s1n2455,n928,n2391);
xor (n2456,n2457,n2388);
xor (n2457,n2384,n2386);
and (n2458,n2456,n2459);
and (n2459,n2460,n2461);
wire s0n2460,s1n2460,notn2460;
or (n2460,s0n2460,s1n2460);
not(notn2460,n928);
and (s0n2460,notn2460,1'b0);
and (s1n2460,n928,n2396);
xor (n2461,n2462,n2394);
xor (n2462,n2390,n2392);
and (n2463,n2455,n2459);
and (n2464,n2449,n2453);
and (n2465,n2443,n2447);
and (n2466,n2437,n2441);
and (n2467,n2431,n2435);
and (n2468,n2425,n2429);
and (n2469,n2419,n2423);
and (n2470,n2413,n2417);
and (n2471,n2408,n2411);
and (n2472,n2153,n2406);
or (n2473,n2474,n2479,n2567);
and (n2474,n2475,n2477);
xor (n2475,n2476,n2084);
xor (n2476,n1816,n2016);
xor (n2477,n2478,n2406);
xor (n2478,n2153,n2331);
and (n2479,n2477,n2480);
or (n2480,n2481,n2486,n2566);
and (n2481,n2482,n2484);
xor (n2482,n2483,n2089);
xor (n2483,n2086,n2087);
xor (n2484,n2485,n2411);
xor (n2485,n2408,n2409);
and (n2486,n2484,n2487);
or (n2487,n2488,n2493,n2565);
and (n2488,n2489,n2491);
xor (n2489,n2490,n2095);
xor (n2490,n2091,n2092);
xor (n2491,n2492,n2417);
xor (n2492,n2413,n2414);
and (n2493,n2491,n2494);
or (n2494,n2495,n2500,n2564);
and (n2495,n2496,n2498);
xor (n2496,n2497,n2101);
xor (n2497,n2097,n2098);
xor (n2498,n2499,n2423);
xor (n2499,n2419,n2420);
and (n2500,n2498,n2501);
or (n2501,n2502,n2507,n2563);
and (n2502,n2503,n2505);
xor (n2503,n2504,n2107);
xor (n2504,n2103,n2104);
xor (n2505,n2506,n2429);
xor (n2506,n2425,n2426);
and (n2507,n2505,n2508);
or (n2508,n2509,n2514,n2562);
and (n2509,n2510,n2512);
xor (n2510,n2511,n2113);
xor (n2511,n2109,n2110);
xor (n2512,n2513,n2435);
xor (n2513,n2431,n2432);
and (n2514,n2512,n2515);
or (n2515,n2516,n2521,n2561);
and (n2516,n2517,n2519);
xor (n2517,n2518,n2119);
xor (n2518,n2115,n2116);
xor (n2519,n2520,n2441);
xor (n2520,n2437,n2438);
and (n2521,n2519,n2522);
or (n2522,n2523,n2528,n2560);
and (n2523,n2524,n2526);
xor (n2524,n2525,n2125);
xor (n2525,n2121,n2122);
xor (n2526,n2527,n2447);
xor (n2527,n2443,n2444);
and (n2528,n2526,n2529);
or (n2529,n2530,n2535,n2559);
and (n2530,n2531,n2533);
xor (n2531,n2532,n2131);
xor (n2532,n2127,n2128);
xor (n2533,n2534,n2453);
xor (n2534,n2449,n2450);
and (n2535,n2533,n2536);
or (n2536,n2537,n2542,n2558);
and (n2537,n2538,n2540);
xor (n2538,n2539,n2137);
xor (n2539,n2133,n2134);
xor (n2540,n2541,n2459);
xor (n2541,n2455,n2456);
and (n2542,n2540,n2543);
or (n2543,n2544,n2547,n2557);
and (n2544,n2545,n2546);
xor (n2545,n2138,n2139);
xor (n2546,n2460,n2461);
and (n2547,n2546,n2548);
or (n2548,n2549,n2552,n2556);
and (n2549,n2550,n2551);
xor (n2550,n2073,n2075);
xor (n2551,n2395,n2397);
and (n2552,n2551,n2553);
and (n2553,n2554,n2555);
wire s0n2554,s1n2554,notn2554;
or (n2554,s0n2554,s1n2554);
not(notn2554,n1025);
and (s0n2554,notn2554,1'b0);
and (s1n2554,n1025,n2074);
wire s0n2555,s1n2555,notn2555;
or (n2555,s0n2555,s1n2555);
not(notn2555,n1025);
and (s0n2555,notn2555,1'b0);
and (s1n2555,n1025,n2396);
and (n2556,n2550,n2553);
and (n2557,n2545,n2548);
and (n2558,n2538,n2543);
and (n2559,n2531,n2536);
and (n2560,n2524,n2529);
and (n2561,n2517,n2522);
and (n2562,n2510,n2515);
and (n2563,n2503,n2508);
and (n2564,n2496,n2501);
and (n2565,n2489,n2494);
and (n2566,n2482,n2487);
and (n2567,n2475,n2480);
or (n2568,n2569,n2574,n2666);
and (n2569,n2570,n2572);
xor (n2570,n2571,n1724);
xor (n2571,n1719,n1721);
xor (n2572,n2573,n2480);
xor (n2573,n2475,n2477);
and (n2574,n2572,n2575);
or (n2575,n2576,n2581,n2665);
and (n2576,n2577,n2579);
xor (n2577,n2578,n1731);
xor (n2578,n1726,n1728);
xor (n2579,n2580,n2487);
xor (n2580,n2482,n2484);
and (n2581,n2579,n2582);
or (n2582,n2583,n2588,n2664);
and (n2583,n2584,n2586);
xor (n2584,n2585,n1738);
xor (n2585,n1733,n1735);
xor (n2586,n2587,n2494);
xor (n2587,n2489,n2491);
and (n2588,n2586,n2589);
or (n2589,n2590,n2595,n2663);
and (n2590,n2591,n2593);
xor (n2591,n2592,n1745);
xor (n2592,n1740,n1742);
xor (n2593,n2594,n2501);
xor (n2594,n2496,n2498);
and (n2595,n2593,n2596);
or (n2596,n2597,n2602,n2662);
and (n2597,n2598,n2600);
xor (n2598,n2599,n1752);
xor (n2599,n1747,n1749);
xor (n2600,n2601,n2508);
xor (n2601,n2503,n2505);
and (n2602,n2600,n2603);
or (n2603,n2604,n2609,n2661);
and (n2604,n2605,n2607);
xor (n2605,n2606,n1759);
xor (n2606,n1754,n1756);
xor (n2607,n2608,n2515);
xor (n2608,n2510,n2512);
and (n2609,n2607,n2610);
or (n2610,n2611,n2616,n2660);
and (n2611,n2612,n2614);
xor (n2612,n2613,n1766);
xor (n2613,n1761,n1763);
xor (n2614,n2615,n2522);
xor (n2615,n2517,n2519);
and (n2616,n2614,n2617);
or (n2617,n2618,n2623,n2659);
and (n2618,n2619,n2621);
xor (n2619,n2620,n1773);
xor (n2620,n1768,n1770);
xor (n2621,n2622,n2529);
xor (n2622,n2524,n2526);
and (n2623,n2621,n2624);
or (n2624,n2625,n2630,n2658);
and (n2625,n2626,n2628);
xor (n2626,n2627,n1780);
xor (n2627,n1775,n1777);
xor (n2628,n2629,n2536);
xor (n2629,n2531,n2533);
and (n2630,n2628,n2631);
or (n2631,n2632,n2637,n2657);
and (n2632,n2633,n2635);
xor (n2633,n2634,n1787);
xor (n2634,n1782,n1784);
xor (n2635,n2636,n2543);
xor (n2636,n2538,n2540);
and (n2637,n2635,n2638);
or (n2638,n2639,n2644,n2656);
and (n2639,n2640,n2642);
xor (n2640,n2641,n1792);
xor (n2641,n1789,n1790);
xor (n2642,n2643,n2548);
xor (n2643,n2545,n2546);
and (n2644,n2642,n2645);
or (n2645,n2646,n2651,n2655);
and (n2646,n2647,n2649);
xor (n2647,n2648,n1797);
xor (n2648,n1794,n1795);
xor (n2649,n2650,n2553);
xor (n2650,n2550,n2551);
and (n2651,n2649,n2652);
and (n2652,n2653,n2654);
xor (n2653,n1798,n1799);
xor (n2654,n2554,n2555);
and (n2655,n2647,n2652);
and (n2656,n2640,n2645);
and (n2657,n2633,n2638);
and (n2658,n2626,n2631);
and (n2659,n2619,n2624);
and (n2660,n2612,n2617);
and (n2661,n2605,n2610);
and (n2662,n2598,n2603);
and (n2663,n2591,n2596);
and (n2664,n2584,n2589);
and (n2665,n2577,n2582);
and (n2666,n2570,n2575);
and (n2667,n2668,n2670);
xor (n2668,n2669,n2575);
xor (n2669,n2570,n2572);
and (n2670,n2671,n2673);
xor (n2671,n2672,n2582);
xor (n2672,n2577,n2579);
and (n2673,n2674,n2676);
xor (n2674,n2675,n2589);
xor (n2675,n2584,n2586);
and (n2676,n2677,n2679);
xor (n2677,n2678,n2596);
xor (n2678,n2591,n2593);
and (n2679,n2680,n2682);
xor (n2680,n2681,n2603);
xor (n2681,n2598,n2600);
and (n2682,n2683,n2685);
xor (n2683,n2684,n2610);
xor (n2684,n2605,n2607);
and (n2685,n2686,n2688);
xor (n2686,n2687,n2617);
xor (n2687,n2612,n2614);
xor (n2688,n2689,n2624);
xor (n2689,n2619,n2621);
nand (n2690,n2691,n3517);
or (n2691,n2692,n3054);
not (n2692,n2693);
nand (n2693,n2694,n3053);
or (n2694,n2695,n2941);
not (n2695,n2696);
nand (n2696,n2697,n2903);
not (n2697,n2698);
or (n2698,n2699,n2902);
and (n2699,n2700,n2807);
xor (n2700,n2701,n2799);
or (n2701,n2702,n2798);
and (n2702,n2703,n2747);
xor (n2703,n2704,n2706);
xor (n2704,n2705,n1207);
xor (n2705,n1080,n2086);
xor (n2706,n2707,n2332);
xor (n2707,n2708,n2745);
or (n2708,n2709,n2744);
and (n2709,n2710,n2413);
xor (n2710,n2711,n1643);
and (n2711,n2712,n1651);
xor (n2712,n1650,n2713);
xor (n2713,n2714,n2724);
xor (n2714,n2715,n2721);
xor (n2715,n2716,n2720);
xor (n2716,n2717,n2719);
nor (n2717,n2718,n1024);
not (n2718,n2156);
and (n2719,n1292,n1025);
and (n2720,n2719,n1308);
and (n2721,n2717,n2722);
not (n2722,n2723);
not (n2723,n2172);
or (n2724,n2725,n2743);
and (n2725,n2726,n2735);
xor (n2726,n2727,n2728);
nor (n2727,n1503,n1024);
and (n2728,n2729,n1025);
nand (n2729,n2730,n2734);
or (n2730,n2731,n2732);
not (n2731,n2169);
not (n2732,n2733);
not (n2733,n2287);
or (n2734,n2733,n2169);
and (n2735,n2736,n1025);
or (n2736,n2737,n2741);
nor (n2737,n2738,n2723);
and (n2738,n2739,n2740);
not (n2739,n2292);
not (n2740,n2184);
nor (n2741,n2742,n2718);
not (n2742,n2216);
and (n2743,n2727,n2728);
and (n2744,n2711,n1643);
xor (n2745,n2746,n1636);
xor (n2746,n1483,n1635);
or (n2747,n2748,n2797);
and (n2748,n2749,n2755);
xor (n2749,n2750,n2754);
or (n2750,n2751,n2753);
and (n2751,n2752,n1222);
xor (n2752,n2097,n2026);
and (n2753,n2097,n2026);
xor (n2754,n2710,n2413);
and (n2755,n2756,n1089);
xor (n2756,n1221,n2757);
or (n2757,n2758,n2796);
and (n2758,n2759,n2781);
xor (n2759,n2425,n2760);
and (n2760,n2761,n2775);
or (n2761,n2762,n2774);
and (n2762,n2763,n2773);
xor (n2763,n2764,n2772);
and (n2764,n2765,n1025);
nand (n2765,n2766,n2768,n2771);
or (n2766,n2767,n2739);
not (n2767,n2248);
or (n2768,n2769,n2770);
not (n2769,n2298);
not (n2770,n2220);
not (n2771,n2203);
and (n2772,n1527,n1025);
nor (n2773,n1524,n1024);
and (n2774,n2764,n2772);
and (n2775,n2776,n1025);
nor (n2776,n2777,n2779);
and (n2777,n2778,n2722);
xor (n2778,n2739,n2740);
and (n2779,n2780,n2723);
not (n2780,n2778);
or (n2781,n2782,n2795);
and (n2782,n2783,n2431);
xor (n2783,n1667,n2784);
xor (n2784,n2785,n2794);
xor (n2785,n2786,n2787);
and (n2786,n1514,n1025);
and (n2787,n2788,n1025);
nand (n2788,n2789,n2793);
or (n2789,n2790,n2769);
and (n2790,n2791,n2792);
not (n2791,n2188);
not (n2792,n2200);
not (n2793,n2187);
and (n2794,n1509,n1025);
and (n2795,n1667,n2784);
and (n2796,n2425,n2760);
and (n2797,n2750,n2754);
and (n2798,n2704,n2706);
xor (n2799,n2800,n2805);
xor (n2800,n2801,n2804);
or (n2801,n2802,n2803);
and (n2802,n2707,n2332);
and (n2803,n2708,n2745);
xor (n2804,n1477,n1075);
xor (n2805,n2806,n1077);
xor (n2806,n1816,n2153);
or (n2807,n2808,n2901);
and (n2808,n2809,n2857);
xor (n2809,n2810,n2847);
or (n2810,n2811,n2846);
and (n2811,n2812,n2838);
xor (n2812,n2813,n2828);
or (n2813,n2814,n2827);
and (n2814,n2815,n1142);
xor (n2815,n2028,n2816);
xor (n2816,n2817,n2419);
xor (n2817,n1491,n2818);
or (n2818,n2819,n2826);
and (n2819,n2820,n2823);
xor (n2820,n2821,n2822);
xor (n2821,n2726,n2735);
and (n2822,n1494,n1025);
or (n2823,n2824,n2825);
and (n2824,n2785,n2794);
and (n2825,n2786,n2787);
and (n2826,n2821,n2822);
and (n2827,n2028,n2816);
xor (n2828,n2829,n2020);
xor (n2829,n1486,n2830);
xor (n2830,n2831,n1642);
xor (n2831,n2832,n2835);
or (n2832,n2833,n2834);
and (n2833,n2714,n2724);
and (n2834,n2715,n2721);
or (n2835,n2836,n2837);
and (n2836,n2716,n2720);
and (n2837,n2717,n2719);
xor (n2838,n2839,n1214);
xor (n2839,n2840,n2091);
or (n2840,n2841,n2845);
and (n2841,n2842,n2342);
xor (n2842,n2843,n2844);
xor (n2843,n2712,n1651);
and (n2844,n1657,n1579);
and (n2845,n2843,n2844);
and (n2846,n2813,n2828);
xor (n2847,n2848,n2852);
xor (n2848,n2849,n2017);
or (n2849,n2850,n2851);
and (n2850,n2829,n2020);
and (n2851,n1486,n2830);
and (n2852,n2853,n2335);
xor (n2853,n1213,n2854);
or (n2854,n2855,n2856);
and (n2855,n2817,n2419);
and (n2856,n1491,n2818);
or (n2857,n2858,n2900);
and (n2858,n2859,n2898);
xor (n2859,n2860,n2861);
xor (n2860,n2853,n2335);
or (n2861,n2862,n2897);
and (n2862,n2863,n2892);
xor (n2863,n2864,n2865);
xor (n2864,n2842,n2342);
or (n2865,n2866,n2891);
and (n2866,n2867,n2349);
xor (n2867,n2868,n2890);
or (n2868,n2869,n2889);
and (n2869,n2870,n2356);
xor (n2870,n1585,n2871);
or (n2871,n2872,n2888);
and (n2872,n2873,n1675);
xor (n2873,n2874,n2886);
or (n2874,n2875,n2876);
and (n2875,n1538,n1025);
and (n2876,n2877,n1025);
nand (n2877,n2878,n2879);
not (n2878,n2219);
nand (n2879,n2880,n2884);
or (n2880,n2881,n2882);
not (n2881,n2770);
not (n2882,n2883);
not (n2883,n2232);
not (n2884,n2885);
not (n2885,n2310);
nor (n2886,n1024,n2887);
xor (n2887,n2300,n2769);
and (n2888,n2874,n2886);
and (n2889,n1585,n2871);
xor (n2890,n2820,n2823);
and (n2891,n2868,n2890);
or (n2892,n2893,n2896);
and (n2893,n2894,n2103);
xor (n2894,n1229,n2895);
xor (n2895,n1657,n1579);
and (n2896,n1229,n2895);
and (n2897,n2864,n2865);
xor (n2898,n2899,n1084);
xor (n2899,n1085,n2022);
and (n2900,n2860,n2861);
and (n2901,n2810,n2847);
and (n2902,n2701,n2799);
or (n2903,n2904,n2698);
nor (n2904,n2905,n2918);
not (n2905,n2906);
nor (n2906,n2907,n2915);
not (n2907,n2908);
nor (n2908,n2909,n2910);
and (n2909,n2806,n1077);
not (n2910,n2911);
nor (n2911,n2912,n2913);
and (n2912,n1477,n1075);
not (n2913,n2914);
xnor (n2914,n6,n1289);
or (n2915,n2916,n2917);
and (n2916,n2800,n2805);
and (n2917,n2801,n2804);
and (n2918,n2919,n2930);
xor (n2919,n2920,n2929);
xor (n2920,n2921,n2926);
xor (n2921,n2922,n2925);
and (n2922,n2923,n2408);
xor (n2923,n1206,n2924);
and (n2924,n2832,n2835);
and (n2925,n2746,n1636);
or (n2926,n2927,n2928);
and (n2927,n2705,n1207);
and (n2928,n1080,n2086);
and (n2929,n2848,n2852);
or (n2930,n2931,n2940);
and (n2931,n2932,n2937);
xor (n2932,n2933,n2934);
xor (n2933,n2923,n2408);
or (n2934,n2935,n2936);
and (n2935,n2839,n1214);
and (n2936,n2840,n2091);
or (n2937,n2938,n2939);
and (n2938,n2899,n1084);
and (n2939,n1085,n2022);
and (n2940,n2933,n2934);
not (n2941,n2942);
or (n2942,n2943,n3052);
and (n2943,n2944,n3051);
xor (n2944,n2945,n3050);
or (n2945,n2946,n3049);
and (n2946,n2947,n2950);
xor (n2947,n2948,n2949);
xor (n2948,n2703,n2747);
xor (n2949,n2932,n2937);
or (n2950,n2951,n3048);
and (n2951,n2952,n2977);
xor (n2952,n2953,n2954);
xor (n2953,n2749,n2755);
or (n2954,n2955,n2976);
and (n2955,n2956,n2963);
xor (n2956,n2957,n2962);
or (n2957,n2958,n2961);
and (n2958,n2959,n2034);
xor (n2959,n1230,n2960);
xor (n2960,n2759,n2781);
and (n2961,n1230,n2960);
xor (n2962,n2756,n1089);
or (n2963,n2964,n2975);
and (n2964,n2965,n1146);
xor (n2965,n2032,n2966);
or (n2966,n2967,n2974);
and (n2967,n2968,n1237);
xor (n2968,n2969,n2971);
xor (n2969,n2970,n1666);
xor (n2970,n2761,n2775);
and (n2971,n2972,n2437);
xor (n2972,n2973,n1674);
xor (n2973,n2763,n2773);
and (n2974,n2969,n2971);
and (n2975,n2032,n2966);
and (n2976,n2957,n2962);
or (n2977,n2978,n3047);
and (n2978,n2979,n3046);
xor (n2979,n2980,n3045);
or (n2980,n2981,n3044);
and (n2981,n2982,n1150);
xor (n2982,n2983,n3020);
or (n2983,n2984,n3019);
and (n2984,n2985,n1238);
xor (n2985,n2986,n2987);
xor (n2986,n2870,n2356);
and (n2987,n2988,n3018);
xor (n2988,n2989,n3016);
or (n2989,n2990,n3015);
and (n2990,n2991,n2443);
xor (n2991,n2992,n3000);
and (n2992,n2993,n2996);
xor (n2993,n2994,n1690);
and (n2994,n2995,n1025);
xnor (n2995,n2885,n2312);
and (n2996,n2997,n2998);
and (n2997,n2555,n2884);
nor (n2998,n2999,n1557);
not (n2999,n1799);
or (n3000,n3001,n3014);
and (n3001,n3002,n3013);
xor (n3002,n3003,n3012);
and (n3003,n3004,n1025);
not (n3004,n3005);
nor (n3005,n3006,n3007);
and (n3006,n2884,n2252);
and (n3007,n3008,n3011);
nand (n3008,n3009,n3010);
not (n3009,n2316);
not (n3010,n2236);
not (n3011,n2767);
and (n3012,n1550,n1025);
and (n3013,n1556,n1025);
and (n3014,n3003,n3012);
and (n3015,n2992,n3000);
and (n3016,n3017,n1598);
xor (n3017,n2370,n1682);
xor (n3018,n2972,n2437);
and (n3019,n2986,n2987);
or (n3020,n3021,n3043);
and (n3021,n3022,n2109);
xor (n3022,n3023,n3024);
xor (n3023,n2783,n2431);
or (n3024,n3025,n3042);
and (n3025,n3026,n2363);
xor (n3026,n1592,n3027);
or (n3027,n3028,n3041);
and (n3028,n3029,n1683);
xor (n3029,n3030,n3040);
and (n3030,n3031,n1025);
not (n3031,n3032);
nor (n3032,n3033,n3039);
and (n3033,n3034,n3037);
not (n3034,n3035);
xor (n3035,n2742,n3036);
not (n3036,n2304);
not (n3037,n3038);
not (n3038,n2204);
and (n3039,n3035,n3038);
and (n3040,n1544,n1025);
and (n3041,n3030,n3040);
and (n3042,n1592,n3027);
and (n3043,n3023,n3024);
and (n3044,n2983,n3020);
xor (n3045,n2752,n1222);
xor (n3046,n2815,n1142);
and (n3047,n2980,n3045);
and (n3048,n2953,n2954);
and (n3049,n2948,n2949);
xor (n3050,n2919,n2930);
xor (n3051,n2700,n2807);
and (n3052,n2945,n3050);
or (n3053,n2942,n2696);
not (n3054,n3055);
or (n3055,n3056,n3516);
and (n3056,n3057,n3117);
xor (n3057,n3058,n3059);
xor (n3058,n2944,n3051);
or (n3059,n3060,n3116);
and (n3060,n3061,n3115);
xor (n3061,n3062,n3114);
or (n3062,n3063,n3113);
and (n3063,n3064,n3067);
xor (n3064,n3065,n3066);
xor (n3065,n2859,n2898);
xor (n3066,n2812,n2838);
or (n3067,n3068,n3112);
and (n3068,n3069,n3102);
xor (n3069,n3070,n3101);
or (n3070,n3071,n3100);
and (n3071,n3072,n3075);
xor (n3072,n3073,n3074);
xor (n3073,n2894,n2103);
xor (n3074,n2867,n2349);
or (n3075,n3076,n3099);
and (n3076,n3077,n2040);
xor (n3077,n3078,n3081);
and (n3078,n3079,n2115);
xor (n3079,n1245,n3080);
xor (n3080,n2873,n1675);
or (n3081,n3082,n3098);
and (n3082,n3083,n1246);
xor (n3083,n3084,n3085);
xor (n3084,n3026,n2363);
or (n3085,n3086,n3097);
and (n3086,n3087,n3093);
xor (n3087,n3088,n3089);
xor (n3088,n3029,n1683);
nand (n3089,n3090,n2874);
or (n3090,n3091,n3092);
not (n3091,n2876);
not (n3092,n2875);
or (n3093,n3094,n3096);
and (n3094,n3095,n1604);
xor (n3095,n1691,n2449);
and (n3096,n1691,n2449);
and (n3097,n3088,n3089);
and (n3098,n3084,n3085);
and (n3099,n3078,n3081);
and (n3100,n3073,n3074);
xor (n3101,n2863,n2892);
or (n3102,n3103,n3111);
and (n3103,n3104,n3110);
xor (n3104,n3105,n3106);
xor (n3105,n2959,n2034);
or (n3106,n3107,n3109);
and (n3107,n3108,n1157);
xor (n3108,n1154,n2038);
and (n3109,n1154,n2038);
xor (n3110,n2965,n1146);
and (n3111,n3105,n3106);
and (n3112,n3070,n3101);
and (n3113,n3065,n3066);
xor (n3114,n2809,n2857);
xor (n3115,n2947,n2950);
and (n3116,n3062,n3114);
or (n3117,n3118,n3515);
and (n3118,n3119,n3190);
xor (n3119,n3120,n3121);
xor (n3120,n3061,n3115);
or (n3121,n3122,n3189);
and (n3122,n3123,n3188);
xor (n3123,n3124,n3187);
or (n3124,n3125,n3186);
and (n3125,n3126,n3185);
xor (n3126,n3127,n3128);
xor (n3127,n2956,n2963);
or (n3128,n3129,n3184);
and (n3129,n3130,n3161);
xor (n3130,n3131,n3132);
xor (n3131,n2982,n1150);
or (n3132,n3133,n3160);
and (n3133,n3134,n3137);
xor (n3134,n3135,n3136);
xor (n3135,n2968,n1237);
xor (n3136,n3022,n2109);
or (n3137,n3138,n3159);
and (n3138,n3139,n2044);
xor (n3139,n3140,n1161);
and (n3140,n3141,n3158);
and (n3141,n3142,n3147);
or (n3142,n3143,n3146);
and (n3143,n3144,n2384);
xor (n3144,n1699,n3145);
xor (n3145,n2997,n2998);
and (n3146,n1699,n3145);
and (n3147,n3148,n3157);
xor (n3148,n3149,n1269);
and (n3149,n3150,n1025);
nand (n3150,n3151,n3156);
or (n3151,n3010,n3152);
nand (n3152,n3153,n3155);
or (n3153,n3154,n2767);
not (n3154,n3009);
nand (n3155,n3154,n2767);
nand (n3156,n3152,n3010);
and (n3157,n1562,n1025);
xor (n3158,n2991,n2443);
and (n3159,n3140,n1161);
and (n3160,n3135,n3136);
or (n3161,n3162,n3183);
and (n3162,n3163,n3182);
xor (n3163,n3164,n3181);
or (n3164,n3165,n3180);
and (n3165,n3166,n1164);
xor (n3166,n3167,n3179);
or (n3167,n3168,n3178);
and (n3168,n3169,n1254);
xor (n3169,n3170,n3171);
xor (n3170,n3017,n1598);
or (n3171,n3172,n3177);
and (n3172,n3173,n2377);
xor (n3173,n3174,n3175);
xor (n3174,n3002,n3013);
and (n3175,n2455,n3176);
and (n3176,n2460,n2138);
and (n3177,n3174,n3175);
and (n3178,n3170,n3171);
xor (n3179,n2988,n3018);
and (n3180,n3167,n3179);
xor (n3181,n2985,n1238);
xor (n3182,n3108,n1157);
and (n3183,n3164,n3181);
and (n3184,n3131,n3132);
xor (n3185,n2979,n3046);
and (n3186,n3127,n3128);
xor (n3187,n2952,n2977);
xor (n3188,n3064,n3067);
and (n3189,n3124,n3187);
or (n3190,n3191,n3514);
and (n3191,n3192,n3283);
xor (n3192,n3193,n3194);
xor (n3193,n3123,n3188);
or (n3194,n3195,n3282);
and (n3195,n3196,n3281);
xor (n3196,n3197,n3198);
xor (n3197,n3069,n3102);
or (n3198,n3199,n3280);
and (n3199,n3200,n3279);
xor (n3200,n3201,n3202);
xor (n3201,n3072,n3075);
or (n3202,n3203,n3278);
and (n3203,n3204,n3220);
xor (n3204,n3205,n3219);
or (n3205,n3206,n3218);
and (n3206,n3207,n3209);
xor (n3207,n2046,n3208);
xor (n3208,n3079,n2115);
or (n3209,n3210,n3217);
and (n3210,n3211,n1168);
xor (n3211,n3212,n2121);
or (n3212,n3213,n3216);
and (n3213,n3214,n1262);
xor (n3214,n2127,n3215);
xor (n3215,n2993,n2996);
and (n3216,n2127,n3215);
and (n3217,n3212,n2121);
and (n3218,n2046,n3208);
xor (n3219,n3077,n2040);
or (n3220,n3221,n3277);
and (n3221,n3222,n3276);
xor (n3222,n3223,n3224);
xor (n3223,n3083,n1246);
or (n3224,n3225,n3275);
and (n3225,n3226,n2052);
xor (n3226,n2050,n3227);
or (n3227,n3228,n3274);
and (n3228,n3229,n3252);
xor (n3229,n3230,n3231);
xor (n3230,n3095,n1604);
or (n3231,n3232,n3251);
and (n3232,n3233,n1610);
xor (n3233,n3234,n3241);
or (n3234,n3235,n3240);
and (n3235,n3236,n3238);
xor (n3236,n3237,n2390);
xor (n3237,n2460,n2138);
and (n3238,n3239,n1025);
not (n3239,n1568);
and (n3240,n3237,n2390);
or (n3241,n3242,n3250);
and (n3242,n3243,n3246);
xor (n3243,n3244,n3245);
and (n3244,n1388,n1025);
and (n3245,n2252,n1025);
and (n3246,n3247,n1025);
xor (n3247,n3248,n3249);
not (n3248,n2264);
not (n3249,n2321);
and (n3250,n3244,n3245);
and (n3251,n3234,n3241);
or (n3252,n3253,n3273);
and (n3253,n3254,n2133);
xor (n3254,n3255,n3271);
or (n3255,n3256,n3270);
and (n3256,n3257,n1275);
xor (n3257,n3258,n3265);
or (n3258,n3259,n3264);
and (n3259,n3260,n3262);
xor (n3260,n3261,n2395);
nor (n3261,n1554,n1024);
nor (n3262,n3263,n1024);
not (n3263,n2279);
and (n3264,n3261,n2395);
and (n3265,n3266,n3268);
nor (n3266,n3267,n1024);
not (n3267,n1404);
nor (n3268,n3269,n1024);
not (n3269,n2267);
and (n3270,n3258,n3265);
xor (n3271,n3272,n1698);
xor (n3272,n2455,n3176);
and (n3273,n3255,n3271);
and (n3274,n3230,n3231);
and (n3275,n2050,n3227);
xor (n3276,n3139,n2044);
and (n3277,n3223,n3224);
and (n3278,n3205,n3219);
xor (n3279,n3104,n3110);
and (n3280,n3201,n3202);
xor (n3281,n3126,n3185);
and (n3282,n3197,n3198);
or (n3283,n3284,n3513);
and (n3284,n3285,n3337);
xor (n3285,n3286,n3336);
or (n3286,n3287,n3335);
and (n3287,n3288,n3334);
xor (n3288,n3289,n3333);
or (n3289,n3290,n3332);
and (n3290,n3291,n3331);
xor (n3291,n3292,n3330);
or (n3292,n3293,n3329);
and (n3293,n3294,n3328);
xor (n3294,n3295,n3322);
or (n3295,n3296,n3321);
and (n3296,n3297,n3316);
xor (n3297,n3298,n3300);
xor (n3298,n3299,n1253);
xor (n3299,n3141,n3158);
or (n3300,n3301,n3315);
and (n3301,n3302,n1175);
xor (n3302,n3303,n3313);
or (n3303,n3304,n3312);
and (n3304,n3305,n3311);
xor (n3305,n1270,n3306);
or (n3306,n3307,n3310);
and (n3307,n3308,n1704);
xor (n3308,n3309,n1616);
xor (n3309,n3243,n3246);
and (n3310,n3309,n1616);
xor (n3311,n3144,n2384);
and (n3312,n1270,n3306);
xor (n3313,n3314,n1261);
xor (n3314,n3142,n3147);
and (n3315,n3303,n3313);
or (n3316,n3317,n3320);
and (n3317,n3318,n1177);
xor (n3318,n2056,n3319);
xor (n3319,n3173,n2377);
and (n3320,n2056,n3319);
and (n3321,n3298,n3300);
or (n3322,n3323,n3327);
and (n3323,n3324,n1171);
xor (n3324,n3325,n3326);
xor (n3325,n3087,n3093);
xor (n3326,n3169,n1254);
and (n3327,n3325,n3326);
xor (n3328,n3166,n1164);
and (n3329,n3295,n3322);
xor (n3330,n3134,n3137);
xor (n3331,n3163,n3182);
and (n3332,n3292,n3330);
xor (n3333,n3130,n3161);
xor (n3334,n3200,n3279);
and (n3335,n3289,n3333);
xor (n3336,n3196,n3281);
or (n3337,n3338,n3512);
and (n3338,n3339,n3404);
xor (n3339,n3340,n3403);
or (n3340,n3341,n3402);
and (n3341,n3342,n3401);
xor (n3342,n3343,n3344);
xor (n3343,n3204,n3220);
or (n3344,n3345,n3400);
and (n3345,n3346,n3399);
xor (n3346,n3347,n3348);
xor (n3347,n3207,n3209);
or (n3348,n3349,n3398);
and (n3349,n3350,n3362);
xor (n3350,n3351,n3352);
xor (n3351,n3211,n1168);
or (n3352,n3353,n3361);
and (n3353,n3354,n2058);
xor (n3354,n3355,n3356);
xor (n3355,n3214,n1262);
or (n3356,n3357,n3360);
and (n3357,n3358,n1181);
xor (n3358,n2062,n3359);
xor (n3359,n3148,n3157);
and (n3360,n2062,n3359);
and (n3361,n3355,n3356);
or (n3362,n3363,n3397);
and (n3363,n3364,n3382);
xor (n3364,n3365,n3366);
xor (n3365,n3229,n3252);
or (n3366,n3367,n3381);
and (n3367,n3368,n2064);
xor (n3368,n3369,n3380);
or (n3369,n3370,n3379);
and (n3370,n3371,n1187);
xor (n3371,n3372,n3373);
xor (n3372,n3236,n3238);
or (n3373,n3374,n3378);
and (n3374,n3375,n3377);
xor (n3375,n3376,n2073);
and (n3376,n1799,n2554);
xor (n3377,n3266,n3268);
and (n3378,n3376,n2073);
and (n3379,n3372,n3373);
xor (n3380,n3233,n1610);
and (n3381,n3369,n3380);
or (n3382,n3383,n3396);
and (n3383,n3384,n1183);
xor (n3384,n3385,n3386);
xor (n3385,n3254,n2133);
or (n3386,n3387,n3395);
and (n3387,n3388,n2068);
xor (n3388,n3389,n3390);
xor (n3389,n3308,n1704);
or (n3390,n3391,n3394);
and (n3391,n3392,n1621);
xor (n3392,n1192,n3393);
xor (n3393,n3260,n3262);
and (n3394,n1192,n3393);
and (n3395,n3389,n3390);
and (n3396,n3385,n3386);
and (n3397,n3365,n3366);
and (n3398,n3351,n3352);
xor (n3399,n3222,n3276);
and (n3400,n3347,n3348);
xor (n3401,n3291,n3331);
and (n3402,n3343,n3344);
xor (n3403,n3288,n3334);
nand (n3404,n3405,n3511);
or (n3405,n3406,n3421);
nor (n3406,n3407,n3408);
xor (n3407,n3342,n3401);
or (n3408,n3409,n3420);
and (n3409,n3410,n3419);
xor (n3410,n3411,n3412);
xor (n3411,n3294,n3328);
or (n3412,n3413,n3418);
and (n3413,n3414,n3417);
xor (n3414,n3415,n3416);
xor (n3415,n3226,n2052);
xor (n3416,n3324,n1171);
xor (n3417,n3297,n3316);
and (n3418,n3415,n3416);
xor (n3419,n3346,n3399);
and (n3420,n3411,n3412);
and (n3421,n3422,n3510);
nand (n3422,n3423,n3438);
or (n3423,n3424,n3425);
xor (n3424,n3410,n3419);
or (n3425,n3426,n3437);
and (n3426,n3427,n3436);
xor (n3427,n3428,n3435);
or (n3428,n3429,n3434);
and (n3429,n3430,n3433);
xor (n3430,n3431,n3432);
xor (n3431,n3318,n1177);
xor (n3432,n3302,n1175);
xor (n3433,n3354,n2058);
and (n3434,n3431,n3432);
xor (n3435,n3350,n3362);
xor (n3436,n3414,n3417);
and (n3437,n3428,n3435);
nand (n3438,n3439,n3503);
nand (n3439,n3440,n3475,n3478);
or (n3440,n3441,n3474);
or (n3441,n3442,n3473);
and (n3442,n3443,n3472);
xor (n3443,n3444,n3461);
or (n3444,n3445,n3460);
and (n3445,n3446,n3459);
xor (n3446,n3447,n3448);
xor (n3447,n3368,n2064);
or (n3448,n3449,n3458);
and (n3449,n3450,n3457);
xor (n3450,n3451,n3452);
xor (n3451,n3371,n1187);
or (n3452,n3453,n3456);
and (n3453,n3454,n2075);
xor (n3454,n3455,n1194);
xor (n3455,n3375,n3377);
and (n3456,n3455,n1194);
xor (n3457,n3388,n2068);
and (n3458,n3451,n3452);
xor (n3459,n3384,n1183);
and (n3460,n3447,n3448);
or (n3461,n3462,n3471);
and (n3462,n3463,n3470);
xor (n3463,n3464,n3469);
or (n3464,n3465,n3468);
and (n3465,n3466,n1189);
xor (n3466,n2070,n3467);
xor (n3467,n3257,n1275);
and (n3468,n2070,n3467);
xor (n3469,n3305,n3311);
xor (n3470,n3358,n1181);
and (n3471,n3464,n3469);
xor (n3472,n3364,n3382);
and (n3473,n3444,n3461);
xor (n3474,n3427,n3436);
or (n3475,n3476,n3477);
xor (n3476,n3443,n3472);
xor (n3477,n3430,n3433);
nand (n3478,n3479,n3499);
or (n3479,n3480,n3483);
nor (n3480,n3481,n3482);
xor (n3481,n3446,n3459);
xor (n3482,n3463,n3470);
nand (n3483,n3484,n3487,n3490);
or (n3484,n3485,n3486);
xor (n3485,n3466,n1189);
xor (n3486,n3450,n3457);
or (n3487,n3488,n3489);
xor (n3488,n3392,n1621);
xor (n3489,n3454,n2075);
nand (n3490,n3491,n3494);
or (n3491,n3492,n3493);
not (n3492,n3488);
not (n3493,n3489);
nor (n3494,n3495,n3498);
and (n3495,n3496,n3497);
xor (n3496,n1799,n2554);
or (n3497,n1798,n2555);
and (n3498,n1798,n2555);
nor (n3499,n3500,n3502);
and (n3500,n3501,n3485,n3486);
not (n3501,n3480);
and (n3502,n3481,n3482);
nor (n3503,n3504,n3508);
and (n3504,n3474,n3505);
nand (n3505,n3506,n3507);
not (n3506,n3441);
nand (n3507,n3476,n3477);
and (n3508,n3509,n3441);
not (n3509,n3507);
nand (n3510,n3424,n3425);
nand (n3511,n3407,n3408);
and (n3512,n3340,n3403);
and (n3513,n3286,n3336);
and (n3514,n3193,n3194);
and (n3515,n3120,n3121);
and (n3516,n3058,n3059);
or (n3517,n3055,n2693);
endmodule
