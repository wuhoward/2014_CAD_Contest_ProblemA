module top (out,n4,n5,n24,n25,n31,n33,n40,n54,n55
        ,n61,n65,n71,n80,n81,n89,n95,n106,n112,n116
        ,n134,n140,n144,n158,n166,n174,n180,n188,n209,n216
        ,n218,n223,n227,n247,n281,n1065);
output out;
input n4;
input n5;
input n24;
input n25;
input n31;
input n33;
input n40;
input n54;
input n55;
input n61;
input n65;
input n71;
input n80;
input n81;
input n89;
input n95;
input n106;
input n112;
input n116;
input n134;
input n140;
input n144;
input n158;
input n166;
input n174;
input n180;
input n188;
input n209;
input n216;
input n218;
input n223;
input n227;
input n247;
input n281;
input n1065;
wire n0;
wire n1;
wire n2;
wire n3;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n217;
wire n219;
wire n220;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
xor (out,n0,n1067);
or (n0,n1,n1064);
and (n1,n2,n6);
nor (n2,n3,n5);
not (n3,n4);
nand (n6,n7,n1063);
or (n7,n8,n490);
not (n8,n9);
nand (n9,n10,n489);
not (n10,n11);
nor (n11,n12,n397);
xor (n12,n13,n349);
xor (n13,n14,n191);
xor (n14,n15,n151);
xor (n15,n16,n99);
or (n16,n17,n98);
and (n17,n18,n74);
xor (n18,n19,n48);
nand (n19,n20,n36);
or (n20,n21,n28);
nor (n21,n22,n26);
and (n22,n23,n25);
not (n23,n24);
and (n26,n24,n27);
not (n27,n25);
not (n28,n29);
nand (n29,n30,n34);
or (n30,n31,n32);
not (n32,n33);
or (n34,n35,n33);
not (n35,n31);
nand (n36,n37,n43);
not (n37,n38);
nor (n38,n39,n41);
and (n39,n40,n35);
and (n41,n42,n31);
not (n42,n40);
not (n43,n44);
nand (n44,n21,n45);
nand (n45,n46,n47);
or (n46,n24,n35);
nand (n47,n35,n24);
nand (n48,n49,n68);
or (n49,n50,n63);
nand (n50,n51,n58);
nor (n51,n52,n56);
and (n52,n53,n55);
not (n53,n54);
and (n56,n54,n57);
not (n57,n55);
nand (n58,n59,n62);
nand (n59,n60,n55);
not (n60,n61);
nand (n62,n61,n57);
nor (n63,n64,n66);
and (n64,n65,n60);
and (n66,n61,n67);
not (n67,n65);
or (n68,n69,n51);
nor (n69,n70,n72);
and (n70,n71,n60);
and (n72,n61,n73);
not (n73,n71);
nand (n74,n75,n92);
or (n75,n76,n87);
nand (n76,n77,n84);
or (n77,n78,n82);
and (n78,n79,n81);
not (n79,n80);
and (n82,n80,n83);
not (n83,n81);
nor (n84,n85,n86);
and (n85,n61,n79);
and (n86,n60,n80);
nor (n87,n88,n90);
and (n88,n89,n83);
and (n90,n81,n91);
not (n91,n89);
or (n92,n93,n84);
nor (n93,n94,n96);
and (n94,n95,n83);
and (n96,n81,n97);
not (n97,n95);
and (n98,n19,n48);
xor (n99,n100,n129);
xor (n100,n101,n123);
nand (n101,n102,n119);
or (n102,n103,n114);
nand (n103,n104,n109);
nor (n104,n105,n107);
and (n105,n35,n106);
and (n107,n31,n108);
not (n108,n106);
nand (n109,n110,n113);
or (n110,n106,n111);
not (n111,n112);
nand (n113,n111,n106);
nor (n114,n115,n117);
and (n115,n111,n116);
and (n117,n112,n118);
not (n118,n116);
or (n119,n104,n120);
nor (n120,n121,n122);
and (n121,n111,n40);
and (n122,n112,n42);
nand (n123,n124,n125);
or (n124,n76,n93);
or (n125,n126,n84);
nor (n126,n127,n128);
and (n127,n65,n83);
and (n128,n81,n67);
nand (n129,n130,n147);
or (n130,n131,n142);
nand (n131,n132,n137);
nor (n132,n133,n135);
and (n133,n83,n134);
and (n135,n81,n136);
not (n136,n134);
nand (n137,n138,n141);
or (n138,n139,n134);
not (n139,n140);
nand (n141,n139,n134);
nor (n142,n143,n145);
and (n143,n144,n139);
and (n145,n140,n146);
not (n146,n144);
or (n147,n148,n132);
nor (n148,n149,n150);
and (n149,n89,n139);
and (n150,n140,n91);
xor (n151,n152,n183);
xor (n152,n153,n161);
nand (n153,n154,n155);
or (n154,n28,n44);
or (n155,n21,n156);
nor (n156,n157,n159);
and (n157,n35,n158);
and (n159,n31,n160);
not (n160,n158);
nand (n161,n162,n177);
or (n162,n163,n172);
nand (n163,n164,n169);
nor (n164,n165,n167);
and (n165,n111,n166);
and (n167,n112,n168);
not (n168,n166);
nand (n169,n170,n171);
or (n170,n53,n166);
nand (n171,n53,n166);
nor (n172,n173,n175);
and (n173,n53,n174);
and (n175,n54,n176);
not (n176,n174);
or (n177,n164,n178);
nor (n178,n179,n181);
and (n179,n53,n180);
and (n181,n54,n182);
not (n182,n180);
nand (n183,n184,n185);
or (n184,n50,n69);
or (n185,n51,n186);
nor (n186,n187,n189);
and (n187,n188,n60);
and (n189,n61,n190);
not (n190,n188);
or (n191,n192,n348);
and (n192,n193,n320);
xor (n193,n194,n261);
or (n194,n195,n260);
and (n195,n196,n230);
xor (n196,n197,n204);
nand (n197,n198,n203);
or (n198,n76,n199);
not (n199,n200);
nand (n200,n201,n202);
or (n201,n146,n81);
or (n202,n83,n144);
or (n203,n87,n84);
xor (n204,n205,n212);
nor (n205,n206,n139);
nor (n206,n207,n210);
and (n207,n208,n83);
nand (n208,n209,n134);
and (n210,n211,n136);
not (n211,n209);
nand (n212,n213,n224);
or (n213,n214,n221);
nor (n214,n215,n219);
and (n215,n216,n217);
not (n217,n218);
and (n219,n220,n218);
not (n220,n216);
nand (n221,n222,n218);
not (n222,n223);
or (n224,n225,n222);
nor (n225,n226,n228);
and (n226,n217,n227);
and (n228,n218,n229);
not (n229,n227);
or (n230,n231,n259);
and (n231,n232,n240);
xor (n232,n233,n234);
nor (n233,n132,n211);
nand (n234,n235,n239);
or (n235,n236,n221);
nor (n236,n237,n238);
and (n237,n218,n160);
nor (n238,n218,n160);
or (n239,n214,n222);
nand (n240,n241,n255);
or (n241,n242,n252);
nand (n242,n243,n249);
not (n243,n244);
nand (n244,n245,n248);
or (n245,n246,n218);
not (n246,n247);
nand (n248,n246,n218);
nand (n249,n250,n251);
or (n250,n246,n25);
nand (n251,n25,n246);
nor (n252,n253,n254);
and (n253,n27,n40);
and (n254,n25,n42);
or (n255,n243,n256);
nor (n256,n257,n258);
and (n257,n27,n33);
and (n258,n25,n32);
and (n259,n233,n234);
and (n260,n197,n204);
xor (n261,n262,n294);
xor (n262,n263,n264);
and (n263,n205,n212);
or (n264,n265,n293);
and (n265,n266,n284);
xor (n266,n267,n273);
nand (n267,n268,n269);
or (n268,n242,n256);
or (n269,n243,n270);
nor (n270,n271,n272);
and (n271,n27,n158);
and (n272,n25,n160);
nand (n273,n274,n278);
or (n274,n131,n275);
nor (n275,n276,n277);
and (n276,n211,n140);
and (n277,n209,n139);
or (n278,n279,n132);
nor (n279,n280,n282);
and (n280,n281,n139);
and (n282,n283,n140);
not (n283,n281);
nand (n284,n285,n289);
or (n285,n103,n286);
nor (n286,n287,n288);
and (n287,n111,n174);
and (n288,n112,n176);
or (n289,n104,n290);
nor (n290,n291,n292);
and (n291,n111,n180);
and (n292,n112,n182);
and (n293,n267,n273);
or (n294,n295,n319);
and (n295,n296,n313);
xor (n296,n297,n307);
nand (n297,n298,n303);
or (n298,n164,n299);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n190,n53);
and (n302,n188,n54);
or (n303,n163,n304);
nor (n304,n305,n306);
and (n305,n53,n71);
and (n306,n54,n73);
nand (n307,n308,n312);
or (n308,n44,n309);
nor (n309,n310,n311);
and (n310,n35,n116);
and (n311,n31,n118);
or (n312,n21,n38);
nand (n313,n314,n318);
or (n314,n50,n315);
nor (n315,n316,n317);
and (n316,n60,n95);
and (n317,n61,n97);
or (n318,n51,n63);
and (n319,n297,n307);
or (n320,n321,n347);
and (n321,n322,n346);
xor (n322,n323,n345);
or (n323,n324,n344);
and (n324,n325,n338);
xor (n325,n326,n332);
nand (n326,n327,n331);
or (n327,n103,n328);
nor (n328,n329,n330);
and (n329,n188,n111);
and (n330,n112,n190);
or (n331,n286,n104);
nand (n332,n333,n337);
or (n333,n163,n334);
nor (n334,n335,n336);
and (n335,n53,n65);
and (n336,n54,n67);
or (n337,n304,n164);
nand (n338,n339,n343);
or (n339,n44,n340);
nor (n340,n341,n342);
and (n341,n35,n180);
and (n342,n31,n182);
or (n343,n21,n309);
and (n344,n326,n332);
xor (n345,n296,n313);
xor (n346,n266,n284);
and (n347,n323,n345);
and (n348,n194,n261);
xor (n349,n350,n389);
xor (n350,n351,n354);
or (n351,n352,n353);
and (n352,n262,n294);
and (n353,n263,n264);
xor (n354,n355,n376);
xor (n355,n356,n366);
not (n356,n357);
nand (n357,n358,n362);
or (n358,n242,n359);
nor (n359,n360,n361);
and (n360,n27,n216);
and (n361,n25,n220);
or (n362,n243,n363);
nor (n363,n364,n365);
and (n364,n27,n227);
and (n365,n25,n229);
nand (n366,n367,n372);
not (n367,n368);
nand (n368,n369,n371);
or (n369,n370,n223);
not (n370,n221);
not (n371,n225);
not (n372,n373);
nand (n373,n374,n375);
or (n374,n242,n270);
or (n375,n243,n359);
or (n376,n377,n388);
and (n377,n378,n385);
xor (n378,n379,n382);
nand (n379,n380,n381);
or (n380,n131,n279);
or (n381,n142,n132);
nand (n382,n383,n384);
or (n383,n103,n290);
or (n384,n104,n114);
nand (n385,n386,n387);
or (n386,n163,n299);
or (n387,n172,n164);
and (n388,n379,n382);
or (n389,n390,n396);
and (n390,n391,n395);
xor (n391,n392,n393);
xor (n392,n18,n74);
nand (n393,n394,n366);
or (n394,n367,n372);
xor (n395,n378,n385);
and (n396,n392,n393);
or (n397,n398,n488);
and (n398,n399,n487);
xor (n399,n400,n401);
xor (n400,n391,n395);
or (n401,n402,n486);
and (n402,n403,n435);
xor (n403,n404,n434);
or (n404,n405,n433);
and (n405,n406,n421);
xor (n406,n407,n413);
nand (n407,n408,n412);
or (n408,n50,n409);
nor (n409,n410,n411);
and (n410,n89,n60);
and (n411,n61,n91);
or (n412,n51,n315);
nand (n413,n414,n415);
or (n414,n84,n199);
nand (n415,n416,n420);
not (n416,n417);
nor (n417,n418,n419);
and (n418,n83,n281);
and (n419,n283,n81);
not (n420,n76);
and (n421,n422,n427);
nor (n422,n423,n83);
nor (n423,n424,n426);
and (n424,n425,n60);
nand (n425,n80,n209);
and (n426,n211,n79);
nand (n427,n428,n432);
or (n428,n429,n221);
nor (n429,n430,n431);
and (n430,n217,n33);
and (n431,n218,n32);
or (n432,n236,n222);
and (n433,n407,n413);
xor (n434,n196,n230);
or (n435,n436,n485);
and (n436,n437,n484);
xor (n437,n438,n462);
or (n438,n439,n461);
and (n439,n440,n454);
xor (n440,n441,n447);
nand (n441,n442,n446);
or (n442,n242,n443);
nor (n443,n444,n445);
and (n444,n116,n27);
and (n445,n118,n25);
or (n446,n243,n252);
nand (n447,n448,n453);
or (n448,n449,n103);
not (n449,n450);
nand (n450,n451,n452);
or (n451,n112,n73);
or (n452,n111,n71);
or (n453,n328,n104);
nand (n454,n455,n460);
or (n455,n163,n456);
not (n456,n457);
nor (n457,n458,n459);
and (n458,n97,n53);
and (n459,n95,n54);
or (n460,n334,n164);
and (n461,n441,n447);
or (n462,n463,n483);
and (n463,n464,n477);
xor (n464,n465,n471);
nand (n465,n466,n470);
or (n466,n44,n467);
nor (n467,n468,n469);
and (n468,n35,n174);
and (n469,n31,n176);
or (n470,n21,n340);
nand (n471,n472,n476);
or (n472,n50,n473);
nor (n473,n474,n475);
and (n474,n144,n60);
and (n475,n61,n146);
or (n476,n409,n51);
nand (n477,n478,n482);
or (n478,n76,n479);
nor (n479,n480,n481);
and (n480,n211,n81);
and (n481,n209,n83);
or (n482,n417,n84);
and (n483,n465,n471);
xor (n484,n232,n240);
and (n485,n438,n462);
and (n486,n404,n434);
xor (n487,n193,n320);
and (n488,n400,n401);
nand (n489,n12,n397);
not (n490,n491);
nand (n491,n492,n1062);
or (n492,n493,n1057);
not (n493,n494);
or (n494,n495,n1056);
and (n495,n496,n619);
xor (n496,n497,n612);
or (n497,n498,n611);
and (n498,n499,n555);
xor (n499,n500,n501);
xor (n500,n437,n484);
xor (n501,n502,n505);
xor (n502,n503,n504);
xor (n503,n325,n338);
xor (n504,n406,n421);
or (n505,n506,n554);
and (n506,n507,n530);
xor (n507,n508,n509);
xor (n508,n422,n427);
or (n509,n510,n529);
and (n510,n511,n522);
xor (n511,n512,n514);
and (n512,n513,n209);
not (n513,n84);
nand (n514,n515,n520);
or (n515,n516,n242);
not (n516,n517);
nand (n517,n518,n519);
or (n518,n25,n182);
or (n519,n27,n180);
nand (n520,n521,n244);
not (n521,n443);
nand (n522,n523,n528);
or (n523,n103,n524);
not (n524,n525);
nand (n525,n526,n527);
or (n526,n112,n67);
or (n527,n111,n65);
or (n528,n104,n449);
and (n529,n512,n514);
or (n530,n531,n553);
and (n531,n532,n547);
xor (n532,n533,n541);
nand (n533,n534,n539);
or (n534,n535,n163);
not (n535,n536);
nand (n536,n537,n538);
or (n537,n54,n91);
or (n538,n53,n89);
nand (n539,n457,n540);
not (n540,n164);
nand (n541,n542,n543);
or (n542,n222,n429);
or (n543,n544,n221);
nor (n544,n545,n546);
and (n545,n217,n40);
and (n546,n218,n42);
nand (n547,n548,n552);
or (n548,n549,n50);
nor (n549,n550,n551);
and (n550,n281,n60);
and (n551,n61,n283);
or (n552,n473,n51);
and (n553,n533,n541);
and (n554,n508,n509);
or (n555,n556,n610);
and (n556,n557,n560);
xor (n557,n558,n559);
xor (n558,n464,n477);
xor (n559,n440,n454);
or (n560,n561,n609);
and (n561,n562,n583);
xor (n562,n563,n569);
nand (n563,n564,n568);
or (n564,n44,n565);
nor (n565,n566,n567);
and (n566,n35,n188);
and (n567,n31,n190);
or (n568,n21,n467);
nor (n569,n570,n577);
not (n570,n571);
nand (n571,n572,n576);
or (n572,n573,n242);
nor (n573,n574,n575);
and (n574,n174,n27);
and (n575,n176,n25);
nand (n576,n244,n517);
nand (n577,n578,n61);
nand (n578,n579,n580);
or (n579,n209,n55);
nand (n580,n581,n53);
not (n581,n582);
and (n582,n209,n55);
or (n583,n584,n608);
and (n584,n585,n601);
xor (n585,n586,n594);
nand (n586,n587,n588);
or (n587,n104,n524);
nand (n588,n589,n593);
not (n589,n590);
nor (n590,n591,n592);
and (n591,n97,n112);
and (n592,n95,n111);
not (n593,n103);
nand (n594,n595,n600);
or (n595,n596,n163);
not (n596,n597);
nor (n597,n598,n599);
and (n598,n53,n146);
and (n599,n54,n144);
nand (n600,n540,n536);
nand (n601,n602,n607);
or (n602,n603,n221);
not (n603,n604);
or (n604,n605,n606);
and (n605,n118,n218);
and (n606,n116,n217);
or (n607,n544,n222);
and (n608,n586,n594);
and (n609,n563,n569);
and (n610,n558,n559);
and (n611,n500,n501);
xor (n612,n613,n618);
xor (n613,n614,n615);
xor (n614,n322,n346);
or (n615,n616,n617);
and (n616,n502,n505);
and (n617,n503,n504);
xor (n618,n403,n435);
or (n619,n620,n1055);
and (n620,n621,n655);
xor (n621,n622,n654);
or (n622,n623,n653);
and (n623,n624,n652);
xor (n624,n625,n626);
xor (n625,n507,n530);
or (n626,n627,n651);
and (n627,n628,n631);
xor (n628,n629,n630);
xor (n629,n532,n547);
xor (n630,n511,n522);
or (n631,n632,n650);
and (n632,n633,n646);
xor (n633,n634,n640);
nand (n634,n635,n639);
or (n635,n50,n636);
nor (n636,n637,n638);
and (n637,n211,n61);
and (n638,n209,n60);
or (n639,n549,n51);
nand (n640,n641,n645);
or (n641,n44,n642);
nor (n642,n643,n644);
and (n643,n35,n71);
and (n644,n31,n73);
or (n645,n21,n565);
nand (n646,n647,n649);
or (n647,n648,n570);
not (n648,n577);
or (n649,n571,n577);
and (n650,n634,n640);
and (n651,n629,n630);
xor (n652,n557,n560);
and (n653,n625,n626);
xor (n654,n499,n555);
nand (n655,n656,n1051);
or (n656,n657,n1029);
nor (n657,n658,n1028);
and (n658,n659,n1009);
or (n659,n660,n1008);
and (n660,n661,n804);
xor (n661,n662,n773);
or (n662,n663,n772);
and (n663,n664,n734);
xor (n664,n665,n695);
xor (n665,n666,n685);
xor (n666,n667,n676);
nand (n667,n668,n672);
or (n668,n103,n669);
nor (n669,n670,n671);
and (n670,n144,n111);
and (n671,n146,n112);
or (n672,n673,n104);
nor (n673,n674,n675);
and (n674,n111,n89);
and (n675,n112,n91);
nand (n676,n677,n681);
or (n677,n163,n678);
nor (n678,n679,n680);
and (n679,n211,n54);
and (n680,n209,n53);
or (n681,n682,n164);
nor (n682,n683,n684);
and (n683,n281,n53);
and (n684,n283,n54);
nand (n685,n686,n691);
or (n686,n221,n687);
not (n687,n688);
nor (n688,n689,n690);
and (n689,n174,n218);
and (n690,n176,n217);
or (n691,n692,n222);
nor (n692,n693,n694);
and (n693,n180,n217);
and (n694,n182,n218);
or (n695,n696,n733);
and (n696,n697,n716);
xor (n697,n698,n707);
nand (n698,n699,n703);
or (n699,n242,n700);
nor (n700,n701,n702);
and (n701,n27,n65);
and (n702,n25,n67);
or (n703,n243,n704);
nor (n704,n705,n706);
and (n705,n73,n25);
and (n706,n71,n27);
nand (n707,n708,n712);
or (n708,n44,n709);
nor (n709,n710,n711);
and (n710,n89,n35);
and (n711,n31,n91);
or (n712,n21,n713);
nor (n713,n714,n715);
and (n714,n35,n95);
and (n715,n31,n97);
and (n716,n717,n723);
nor (n717,n718,n111);
nor (n718,n719,n722);
and (n719,n720,n35);
not (n720,n721);
and (n721,n209,n106);
and (n722,n211,n108);
nand (n723,n724,n729);
or (n724,n725,n221);
not (n725,n726);
nor (n726,n727,n728);
and (n727,n73,n217);
and (n728,n71,n218);
or (n729,n730,n222);
nor (n730,n731,n732);
and (n731,n188,n217);
and (n732,n190,n218);
and (n733,n698,n707);
xor (n734,n735,n757);
xor (n735,n736,n742);
nand (n736,n737,n738);
or (n737,n44,n713);
or (n738,n21,n739);
nor (n739,n740,n741);
and (n740,n35,n65);
and (n741,n31,n67);
xor (n742,n743,n748);
nor (n743,n744,n53);
nor (n744,n745,n747);
and (n745,n746,n111);
nand (n746,n209,n166);
and (n747,n211,n168);
nand (n748,n749,n754);
or (n749,n243,n750);
not (n750,n751);
nand (n751,n752,n753);
or (n752,n25,n190);
or (n753,n27,n188);
nand (n754,n755,n756);
not (n755,n704);
not (n756,n242);
or (n757,n758,n771);
and (n758,n759,n764);
xor (n759,n760,n761);
nor (n760,n164,n211);
nand (n761,n762,n763);
or (n762,n222,n687);
or (n763,n730,n221);
nand (n764,n765,n766);
or (n765,n104,n669);
nand (n766,n767,n593);
not (n767,n768);
or (n768,n769,n770);
and (n769,n283,n111);
and (n770,n281,n112);
and (n771,n760,n761);
and (n772,n665,n695);
xor (n773,n774,n789);
xor (n774,n775,n786);
xor (n775,n776,n783);
xor (n776,n777,n780);
nand (n777,n778,n779);
or (n778,n164,n596);
or (n779,n163,n682);
nand (n780,n781,n782);
or (n781,n692,n221);
nand (n782,n604,n223);
nand (n783,n784,n785);
or (n784,n44,n739);
or (n785,n21,n642);
or (n786,n787,n788);
and (n787,n735,n757);
and (n788,n736,n742);
xor (n789,n790,n795);
xor (n790,n791,n792);
and (n791,n743,n748);
or (n792,n793,n794);
and (n793,n666,n685);
and (n794,n667,n676);
xor (n795,n796,n801);
xor (n796,n797,n798);
nor (n797,n51,n211);
nand (n798,n799,n800);
or (n799,n750,n242);
or (n800,n243,n573);
nand (n801,n802,n803);
or (n802,n103,n673);
or (n803,n104,n590);
nand (n804,n805,n1004,n1007);
nand (n805,n806,n861,n997);
not (n806,n807);
nor (n807,n808,n835);
xor (n808,n809,n834);
xor (n809,n810,n833);
or (n810,n811,n832);
and (n811,n812,n826);
xor (n812,n813,n819);
nand (n813,n814,n818);
or (n814,n103,n815);
nor (n815,n816,n817);
and (n816,n211,n112);
and (n817,n209,n111);
or (n818,n768,n104);
nand (n819,n820,n825);
or (n820,n821,n242);
not (n821,n822);
nor (n822,n823,n824);
and (n823,n95,n25);
and (n824,n97,n27);
or (n825,n243,n700);
nand (n826,n827,n831);
or (n827,n44,n828);
nor (n828,n829,n830);
and (n829,n144,n35);
and (n830,n31,n146);
or (n831,n21,n709);
and (n832,n813,n819);
xor (n833,n759,n764);
xor (n834,n697,n716);
or (n835,n836,n860);
and (n836,n837,n859);
xor (n837,n838,n839);
xor (n838,n717,n723);
or (n839,n840,n858);
and (n840,n841,n851);
xor (n841,n842,n844);
and (n842,n843,n209);
not (n843,n104);
nand (n844,n845,n850);
or (n845,n221,n846);
not (n846,n847);
nor (n847,n848,n849);
and (n848,n67,n217);
and (n849,n65,n218);
nand (n850,n726,n223);
nand (n851,n852,n857);
or (n852,n853,n242);
not (n853,n854);
nor (n854,n855,n856);
and (n855,n91,n27);
and (n856,n89,n25);
nand (n857,n822,n244);
and (n858,n842,n844);
xor (n859,n812,n826);
and (n860,n838,n839);
or (n861,n862,n996);
and (n862,n863,n889);
xor (n863,n864,n888);
or (n864,n865,n887);
and (n865,n866,n886);
xor (n866,n867,n873);
nand (n867,n868,n872);
or (n868,n44,n869);
nor (n869,n870,n871);
and (n870,n35,n281);
and (n871,n31,n283);
or (n872,n828,n21);
and (n873,n874,n880);
and (n874,n875,n31);
nand (n875,n876,n877);
or (n876,n209,n24);
nand (n877,n878,n27);
not (n878,n879);
and (n879,n209,n24);
nand (n880,n881,n882);
or (n881,n222,n846);
or (n882,n883,n221);
nor (n883,n884,n885);
and (n884,n217,n95);
and (n885,n218,n97);
xor (n886,n841,n851);
and (n887,n867,n873);
xor (n888,n837,n859);
nand (n889,n890,n995);
or (n890,n891,n990);
nor (n891,n892,n989);
and (n892,n893,n968);
nand (n893,n894,n966);
or (n894,n895,n949);
not (n895,n896);
or (n896,n897,n948);
and (n897,n898,n927);
xor (n898,n899,n908);
nand (n899,n900,n904);
or (n900,n242,n901);
nor (n901,n902,n903);
and (n902,n25,n211);
and (n903,n209,n27);
or (n904,n243,n905);
nor (n905,n906,n907);
and (n906,n283,n25);
and (n907,n281,n27);
nand (n908,n909,n926);
or (n909,n910,n916);
not (n910,n911);
nand (n911,n912,n25);
nand (n912,n913,n915);
or (n913,n914,n218);
and (n914,n209,n247);
nand (n915,n211,n246);
not (n916,n917);
nand (n917,n918,n922);
or (n918,n919,n221);
or (n919,n920,n921);
and (n920,n144,n218);
and (n921,n146,n217);
or (n922,n923,n222);
nor (n923,n924,n925);
and (n924,n91,n218);
and (n925,n89,n217);
or (n926,n917,n911);
or (n927,n928,n947);
and (n928,n929,n937);
xor (n929,n930,n931);
nor (n930,n243,n211);
nand (n931,n932,n936);
or (n932,n933,n221);
nor (n933,n934,n935);
and (n934,n283,n218);
and (n935,n281,n217);
or (n936,n919,n222);
nor (n937,n938,n945);
nor (n938,n939,n941);
and (n939,n940,n223);
not (n940,n933);
and (n941,n942,n370);
nand (n942,n943,n944);
or (n943,n211,n218);
nand (n944,n218,n211);
or (n945,n946,n217);
and (n946,n209,n223);
and (n947,n930,n931);
and (n948,n899,n908);
not (n949,n950);
nand (n950,n951,n965);
not (n951,n952);
xor (n952,n953,n962);
xor (n953,n954,n956);
and (n954,n955,n209);
not (n955,n21);
nand (n956,n957,n958);
or (n957,n905,n242);
nand (n958,n959,n244);
nor (n959,n960,n961);
and (n960,n146,n27);
and (n961,n144,n25);
nand (n962,n963,n964);
or (n963,n923,n221);
or (n964,n883,n222);
nand (n965,n910,n917);
nand (n966,n967,n952);
not (n967,n965);
nand (n968,n969,n985);
not (n969,n970);
xor (n970,n971,n984);
xor (n971,n972,n976);
nand (n972,n973,n975);
or (n973,n974,n242);
not (n974,n959);
nand (n975,n854,n244);
nand (n976,n977,n982);
or (n977,n978,n44);
not (n978,n979);
nand (n979,n980,n981);
or (n980,n209,n35);
or (n981,n211,n31);
nand (n982,n983,n955);
not (n983,n869);
xor (n984,n874,n880);
not (n985,n986);
or (n986,n987,n988);
and (n987,n953,n962);
and (n988,n954,n956);
nor (n989,n969,n985);
nor (n990,n991,n992);
xor (n991,n866,n886);
or (n992,n993,n994);
and (n993,n971,n984);
and (n994,n972,n976);
nand (n995,n991,n992);
and (n996,n864,n888);
nand (n997,n998,n1002);
not (n998,n999);
or (n999,n1000,n1001);
and (n1000,n809,n834);
and (n1001,n810,n833);
not (n1002,n1003);
xor (n1003,n664,n734);
nand (n1004,n1005,n997);
not (n1005,n1006);
nand (n1006,n808,n835);
nand (n1007,n1003,n999);
and (n1008,n662,n773);
or (n1009,n1010,n1025);
xor (n1010,n1011,n1022);
xor (n1011,n1012,n1013);
xor (n1012,n633,n646);
xor (n1013,n1014,n1021);
xor (n1014,n1015,n1018);
or (n1015,n1016,n1017);
and (n1016,n796,n801);
and (n1017,n797,n798);
or (n1018,n1019,n1020);
and (n1019,n776,n783);
and (n1020,n777,n780);
xor (n1021,n585,n601);
or (n1022,n1023,n1024);
and (n1023,n790,n795);
and (n1024,n791,n792);
or (n1025,n1026,n1027);
and (n1026,n774,n789);
and (n1027,n775,n786);
and (n1028,n1010,n1025);
nand (n1029,n1030,n1044);
not (n1030,n1031);
and (n1031,n1032,n1040);
not (n1032,n1033);
xor (n1033,n1034,n1039);
xor (n1034,n1035,n1036);
xor (n1035,n562,n583);
or (n1036,n1037,n1038);
and (n1037,n1014,n1021);
and (n1038,n1015,n1018);
xor (n1039,n628,n631);
not (n1040,n1041);
or (n1041,n1042,n1043);
and (n1042,n1011,n1022);
and (n1043,n1012,n1013);
nand (n1044,n1045,n1047);
not (n1045,n1046);
xor (n1046,n624,n652);
not (n1047,n1048);
or (n1048,n1049,n1050);
and (n1049,n1034,n1039);
and (n1050,n1035,n1036);
nor (n1051,n1052,n1054);
and (n1052,n1044,n1053);
nor (n1053,n1032,n1040);
nor (n1054,n1045,n1047);
and (n1055,n622,n654);
and (n1056,n497,n612);
nor (n1057,n1058,n1061);
or (n1058,n1059,n1060);
and (n1059,n613,n618);
and (n1060,n614,n615);
xor (n1061,n399,n487);
nand (n1062,n1061,n1058);
or (n1063,n491,n9);
and (n1064,n1065,n1066);
not (n1066,n2);
or (n1067,n1068,n1064);
and (n1068,n1069,n2);
xor (n1069,n1070,n1861);
xor (n1070,n1071,n1862);
xor (n1071,n1072,n1856);
xor (n1072,n1073,n1853);
xor (n1073,n1074,n1852);
xor (n1074,n1075,n1837);
xor (n1075,n1076,n1836);
xor (n1076,n1077,n1815);
xor (n1077,n1078,n1814);
xor (n1078,n1079,n1787);
xor (n1079,n1080,n1786);
xor (n1080,n1081,n1753);
xor (n1081,n1082,n1752);
xor (n1082,n1083,n1714);
xor (n1083,n1084,n1713);
xor (n1084,n1085,n1671);
xor (n1085,n1086,n1670);
xor (n1086,n1087,n1619);
xor (n1087,n1088,n1618);
xor (n1088,n1089,n1562);
xor (n1089,n1090,n1561);
xor (n1090,n1091,n1499);
xor (n1091,n1092,n1498);
xor (n1092,n1093,n1429);
xor (n1093,n1094,n1428);
xor (n1094,n1095,n1354);
xor (n1095,n1096,n1353);
xor (n1096,n1097,n1275);
xor (n1097,n1098,n1274);
xor (n1098,n1099,n1106);
xor (n1099,n1100,n1105);
xor (n1100,n1101,n1104);
xor (n1101,n1102,n1103);
and (n1102,n227,n223);
and (n1103,n227,n218);
and (n1104,n1102,n1103);
and (n1105,n227,n247);
or (n1106,n1107,n1192);
and (n1107,n1108,n1191);
xor (n1108,n1101,n1109);
or (n1109,n1110,n1112);
and (n1110,n1102,n1111);
and (n1111,n216,n218);
and (n1112,n1113,n1114);
xor (n1113,n1102,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
and (n1116,n216,n223);
and (n1117,n158,n218);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
and (n1122,n158,n223);
and (n1123,n33,n218);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
and (n1128,n33,n223);
and (n1129,n40,n218);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
and (n1134,n40,n223);
and (n1135,n116,n218);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n116,n223);
and (n1141,n180,n218);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1147);
and (n1145,n1146,n689);
and (n1146,n180,n223);
and (n1147,n1148,n1149);
xor (n1148,n1146,n689);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
and (n1151,n174,n223);
and (n1152,n188,n218);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1158);
and (n1156,n1157,n728);
and (n1157,n188,n223);
and (n1158,n1159,n1160);
xor (n1159,n1157,n728);
or (n1160,n1161,n1163);
and (n1161,n1162,n849);
and (n1162,n71,n223);
and (n1163,n1164,n1165);
xor (n1164,n1162,n849);
or (n1165,n1166,n1169);
and (n1166,n1167,n1168);
and (n1167,n65,n223);
and (n1168,n95,n218);
and (n1169,n1170,n1171);
xor (n1170,n1167,n1168);
or (n1171,n1172,n1175);
and (n1172,n1173,n1174);
and (n1173,n95,n223);
and (n1174,n89,n218);
and (n1175,n1176,n1177);
xor (n1176,n1173,n1174);
or (n1177,n1178,n1180);
and (n1178,n1179,n920);
and (n1179,n89,n223);
and (n1180,n1181,n1182);
xor (n1181,n1179,n920);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
and (n1184,n144,n223);
and (n1185,n281,n218);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
and (n1188,n1189,n1190);
and (n1189,n281,n223);
and (n1190,n209,n218);
and (n1191,n216,n247);
and (n1192,n1193,n1194);
xor (n1193,n1108,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1113,n1114);
and (n1197,n158,n247);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1119,n1120);
and (n1203,n33,n247);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1125,n1126);
and (n1209,n40,n247);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1131,n1132);
and (n1215,n116,n247);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1137,n1138);
and (n1221,n180,n247);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1143,n1144);
and (n1227,n174,n247);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1148,n1149);
and (n1233,n188,n247);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1154,n1155);
and (n1239,n71,n247);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1246);
and (n1243,n1244,n1245);
xor (n1244,n1159,n1160);
and (n1245,n65,n247);
and (n1246,n1247,n1248);
xor (n1247,n1244,n1245);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1164,n1165);
and (n1251,n95,n247);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1170,n1171);
and (n1257,n89,n247);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1176,n1177);
and (n1263,n144,n247);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
or (n1266,n1267,n1270);
and (n1267,n1268,n1269);
xor (n1268,n1181,n1182);
and (n1269,n281,n247);
and (n1270,n1271,n1272);
xor (n1271,n1268,n1269);
and (n1272,n1273,n914);
xor (n1273,n1187,n1188);
and (n1274,n216,n25);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1193,n1194);
and (n1278,n158,n25);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1199,n1200);
and (n1284,n33,n25);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1205,n1206);
and (n1290,n40,n25);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1211,n1212);
and (n1296,n116,n25);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1217,n1218);
and (n1302,n180,n25);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1223,n1224);
and (n1308,n174,n25);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1229,n1230);
and (n1314,n188,n25);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1235,n1236);
and (n1320,n71,n25);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1241,n1242);
and (n1326,n65,n25);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1332);
and (n1330,n1331,n823);
xor (n1331,n1247,n1248);
and (n1332,n1333,n1334);
xor (n1333,n1331,n823);
or (n1334,n1335,n1337);
and (n1335,n1336,n856);
xor (n1336,n1253,n1254);
and (n1337,n1338,n1339);
xor (n1338,n1336,n856);
or (n1339,n1340,n1342);
and (n1340,n1341,n961);
xor (n1341,n1259,n1260);
and (n1342,n1343,n1344);
xor (n1343,n1341,n961);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1265,n1266);
and (n1347,n281,n25);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
and (n1350,n1351,n1352);
xor (n1351,n1271,n1272);
and (n1352,n209,n25);
and (n1353,n158,n24);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1280,n1281);
and (n1357,n33,n24);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1286,n1287);
and (n1363,n40,n24);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1292,n1293);
and (n1369,n116,n24);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1298,n1299);
and (n1375,n180,n24);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1304,n1305);
and (n1381,n174,n24);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1310,n1311);
and (n1387,n188,n24);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1316,n1317);
and (n1393,n71,n24);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1322,n1323);
and (n1399,n65,n24);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1328,n1329);
and (n1405,n95,n24);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1333,n1334);
and (n1411,n89,n24);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1338,n1339);
and (n1417,n144,n24);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1343,n1344);
and (n1423,n281,n24);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
and (n1426,n1427,n879);
xor (n1427,n1349,n1350);
and (n1428,n33,n31);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1359,n1360);
and (n1432,n40,n31);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1365,n1366);
and (n1438,n116,n31);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1371,n1372);
and (n1444,n180,n31);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1377,n1378);
and (n1450,n174,n31);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1383,n1384);
and (n1456,n188,n31);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
or (n1459,n1460,n1463);
and (n1460,n1461,n1462);
xor (n1461,n1389,n1390);
and (n1462,n71,n31);
and (n1463,n1464,n1465);
xor (n1464,n1461,n1462);
or (n1465,n1466,n1469);
and (n1466,n1467,n1468);
xor (n1467,n1395,n1396);
and (n1468,n65,n31);
and (n1469,n1470,n1471);
xor (n1470,n1467,n1468);
or (n1471,n1472,n1475);
and (n1472,n1473,n1474);
xor (n1473,n1401,n1402);
and (n1474,n95,n31);
and (n1475,n1476,n1477);
xor (n1476,n1473,n1474);
or (n1477,n1478,n1481);
and (n1478,n1479,n1480);
xor (n1479,n1407,n1408);
and (n1480,n89,n31);
and (n1481,n1482,n1483);
xor (n1482,n1479,n1480);
or (n1483,n1484,n1487);
and (n1484,n1485,n1486);
xor (n1485,n1413,n1414);
and (n1486,n144,n31);
and (n1487,n1488,n1489);
xor (n1488,n1485,n1486);
or (n1489,n1490,n1493);
and (n1490,n1491,n1492);
xor (n1491,n1419,n1420);
and (n1492,n281,n31);
and (n1493,n1494,n1495);
xor (n1494,n1491,n1492);
and (n1495,n1496,n1497);
xor (n1496,n1425,n1426);
and (n1497,n209,n31);
and (n1498,n40,n106);
or (n1499,n1500,n1503);
and (n1500,n1501,n1502);
xor (n1501,n1434,n1435);
and (n1502,n116,n106);
and (n1503,n1504,n1505);
xor (n1504,n1501,n1502);
or (n1505,n1506,n1509);
and (n1506,n1507,n1508);
xor (n1507,n1440,n1441);
and (n1508,n180,n106);
and (n1509,n1510,n1511);
xor (n1510,n1507,n1508);
or (n1511,n1512,n1515);
and (n1512,n1513,n1514);
xor (n1513,n1446,n1447);
and (n1514,n174,n106);
and (n1515,n1516,n1517);
xor (n1516,n1513,n1514);
or (n1517,n1518,n1521);
and (n1518,n1519,n1520);
xor (n1519,n1452,n1453);
and (n1520,n188,n106);
and (n1521,n1522,n1523);
xor (n1522,n1519,n1520);
or (n1523,n1524,n1527);
and (n1524,n1525,n1526);
xor (n1525,n1458,n1459);
and (n1526,n71,n106);
and (n1527,n1528,n1529);
xor (n1528,n1525,n1526);
or (n1529,n1530,n1533);
and (n1530,n1531,n1532);
xor (n1531,n1464,n1465);
and (n1532,n65,n106);
and (n1533,n1534,n1535);
xor (n1534,n1531,n1532);
or (n1535,n1536,n1539);
and (n1536,n1537,n1538);
xor (n1537,n1470,n1471);
and (n1538,n95,n106);
and (n1539,n1540,n1541);
xor (n1540,n1537,n1538);
or (n1541,n1542,n1545);
and (n1542,n1543,n1544);
xor (n1543,n1476,n1477);
and (n1544,n89,n106);
and (n1545,n1546,n1547);
xor (n1546,n1543,n1544);
or (n1547,n1548,n1551);
and (n1548,n1549,n1550);
xor (n1549,n1482,n1483);
and (n1550,n144,n106);
and (n1551,n1552,n1553);
xor (n1552,n1549,n1550);
or (n1553,n1554,n1557);
and (n1554,n1555,n1556);
xor (n1555,n1488,n1489);
and (n1556,n281,n106);
and (n1557,n1558,n1559);
xor (n1558,n1555,n1556);
and (n1559,n1560,n721);
xor (n1560,n1494,n1495);
and (n1561,n116,n112);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
xor (n1564,n1504,n1505);
and (n1565,n180,n112);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
or (n1568,n1569,n1572);
and (n1569,n1570,n1571);
xor (n1570,n1510,n1511);
and (n1571,n174,n112);
and (n1572,n1573,n1574);
xor (n1573,n1570,n1571);
or (n1574,n1575,n1578);
and (n1575,n1576,n1577);
xor (n1576,n1516,n1517);
and (n1577,n188,n112);
and (n1578,n1579,n1580);
xor (n1579,n1576,n1577);
or (n1580,n1581,n1584);
and (n1581,n1582,n1583);
xor (n1582,n1522,n1523);
and (n1583,n71,n112);
and (n1584,n1585,n1586);
xor (n1585,n1582,n1583);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
xor (n1588,n1528,n1529);
and (n1589,n65,n112);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1534,n1535);
and (n1595,n95,n112);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1540,n1541);
and (n1601,n89,n112);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
xor (n1606,n1546,n1547);
and (n1607,n144,n112);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1613);
and (n1611,n1612,n770);
xor (n1612,n1552,n1553);
and (n1613,n1614,n1615);
xor (n1614,n1612,n770);
and (n1615,n1616,n1617);
xor (n1616,n1558,n1559);
and (n1617,n209,n112);
and (n1618,n180,n166);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1567,n1568);
and (n1622,n174,n166);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1573,n1574);
and (n1628,n188,n166);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1579,n1580);
and (n1634,n71,n166);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1585,n1586);
and (n1640,n65,n166);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1591,n1592);
and (n1646,n95,n166);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1597,n1598);
and (n1652,n89,n166);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1603,n1604);
and (n1658,n144,n166);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1609,n1610);
and (n1664,n281,n166);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
and (n1667,n1668,n1669);
xor (n1668,n1614,n1615);
not (n1669,n746);
and (n1670,n174,n54);
or (n1671,n1672,n1674);
and (n1672,n1673,n302);
xor (n1673,n1624,n1625);
and (n1674,n1675,n1676);
xor (n1675,n1673,n302);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1630,n1631);
and (n1679,n71,n54);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1636,n1637);
and (n1685,n65,n54);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1691);
and (n1689,n1690,n459);
xor (n1690,n1642,n1643);
and (n1691,n1692,n1693);
xor (n1692,n1690,n459);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1648,n1649);
and (n1696,n89,n54);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1702);
and (n1700,n1701,n599);
xor (n1701,n1654,n1655);
and (n1702,n1703,n1704);
xor (n1703,n1701,n599);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1660,n1661);
and (n1707,n281,n54);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
and (n1710,n1711,n1712);
xor (n1711,n1666,n1667);
and (n1712,n209,n54);
and (n1713,n188,n55);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
xor (n1716,n1675,n1676);
and (n1717,n71,n55);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
xor (n1722,n1681,n1682);
and (n1723,n65,n55);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
xor (n1728,n1687,n1688);
and (n1729,n95,n55);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1736);
and (n1733,n1734,n1735);
xor (n1734,n1692,n1693);
and (n1735,n89,n55);
and (n1736,n1737,n1738);
xor (n1737,n1734,n1735);
or (n1738,n1739,n1742);
and (n1739,n1740,n1741);
xor (n1740,n1698,n1699);
and (n1741,n144,n55);
and (n1742,n1743,n1744);
xor (n1743,n1740,n1741);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1703,n1704);
and (n1747,n281,n55);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
and (n1750,n1751,n582);
xor (n1751,n1709,n1710);
and (n1752,n71,n61);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1719,n1720);
and (n1756,n65,n61);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1725,n1726);
and (n1762,n95,n61);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1731,n1732);
and (n1768,n89,n61);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1737,n1738);
and (n1774,n144,n61);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1743,n1744);
and (n1780,n281,n61);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
and (n1783,n1784,n1785);
xor (n1784,n1749,n1750);
and (n1785,n209,n61);
and (n1786,n65,n80);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1758,n1759);
and (n1790,n95,n80);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1764,n1765);
and (n1796,n89,n80);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1770,n1771);
and (n1802,n144,n80);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1776,n1777);
and (n1808,n281,n80);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
and (n1811,n1812,n1813);
xor (n1812,n1782,n1783);
not (n1813,n425);
and (n1814,n95,n81);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1792,n1793);
and (n1818,n89,n81);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1825);
and (n1822,n1823,n1824);
xor (n1823,n1798,n1799);
and (n1824,n144,n81);
and (n1825,n1826,n1827);
xor (n1826,n1823,n1824);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1804,n1805);
and (n1830,n281,n81);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
and (n1833,n1834,n1835);
xor (n1834,n1810,n1811);
and (n1835,n209,n81);
and (n1836,n89,n134);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
xor (n1839,n1820,n1821);
and (n1840,n144,n134);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
or (n1843,n1844,n1847);
and (n1844,n1845,n1846);
xor (n1845,n1826,n1827);
and (n1846,n281,n134);
and (n1847,n1848,n1849);
xor (n1848,n1845,n1846);
and (n1849,n1850,n1851);
xor (n1850,n1832,n1833);
not (n1851,n208);
and (n1852,n144,n140);
or (n1853,n1854,n1857);
and (n1854,n1855,n1856);
xor (n1855,n1842,n1843);
and (n1856,n281,n140);
and (n1857,n1858,n1859);
xor (n1858,n1855,n1856);
and (n1859,n1860,n1861);
xor (n1860,n1848,n1849);
and (n1861,n209,n140);
and (n1862,n1863,n1861);
xor (n1863,n1858,n1859);
endmodule
