module top (out,n16,n17,n22,n29,n34,n38,n42,n71,n72
        ,n86,n115,n121,n130,n136,n142,n154,n160,n171,n172
        ,n178,n186,n207,n215,n220,n249,n270,n329,n351,n352
        ,n381,n770,n803,n864,n943);
output out;
input n16;
input n17;
input n22;
input n29;
input n34;
input n38;
input n42;
input n71;
input n72;
input n86;
input n115;
input n121;
input n130;
input n136;
input n142;
input n154;
input n160;
input n171;
input n172;
input n178;
input n186;
input n207;
input n215;
input n220;
input n249;
input n270;
input n329;
input n351;
input n352;
input n381;
input n770;
input n803;
input n864;
input n943;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
xor (out,n0,n1949);
nor (n0,n1,n1946);
and (n1,n2,n48);
nor (n2,n3,n47);
and (n3,n4,n45);
not (n4,n5);
or (n5,n6,n44);
and (n6,n7,n39);
xor (n7,n8,n24);
nand (n8,n9,n22);
or (n9,n10,n13);
not (n10,n11);
nand (n11,n12,n19);
not (n12,n13);
nand (n13,n14,n18);
or (n14,n15,n17);
not (n15,n16);
nand (n18,n15,n17);
nand (n19,n20,n23);
or (n20,n17,n21);
not (n21,n22);
nand (n23,n21,n17);
nand (n24,n25,n35);
or (n25,n26,n33);
not (n26,n27);
nor (n27,n28,n30);
not (n28,n29);
nand (n30,n31,n32);
or (n31,n21,n29);
nand (n32,n29,n21);
not (n33,n34);
or (n35,n36,n37);
not (n36,n30);
not (n37,n38);
not (n39,n40);
nor (n40,n41,n43);
and (n41,n27,n42);
and (n43,n30,n34);
and (n44,n8,n24);
not (n45,n46);
nand (n46,n27,n38);
and (n47,n5,n46);
nand (n48,n49,n1945);
or (n49,n50,n92);
not (n50,n51);
or (n51,n52,n91);
or (n52,n53,n90);
and (n53,n54,n61);
xor (n54,n55,n40);
nand (n55,n56,n60);
or (n56,n11,n57);
nor (n57,n58,n59);
and (n58,n21,n38);
and (n59,n22,n37);
or (n60,n12,n21);
or (n61,n62,n89);
and (n62,n63,n83);
xor (n63,n64,n77);
nand (n64,n65,n16);
or (n65,n66,n76);
not (n66,n67);
nand (n67,n68,n75);
nor (n68,n69,n73);
and (n69,n70,n72);
not (n70,n71);
and (n73,n71,n74);
not (n74,n72);
xor (n75,n70,n15);
not (n76,n68);
nand (n77,n78,n82);
or (n78,n11,n79);
nor (n79,n80,n81);
and (n80,n21,n34);
and (n81,n22,n33);
or (n82,n12,n57);
nand (n83,n84,n87);
or (n84,n26,n85);
not (n85,n86);
or (n87,n36,n88);
not (n88,n42);
and (n89,n64,n77);
and (n90,n55,n40);
xor (n91,n7,n39);
not (n92,n93);
nand (n93,n94,n1918);
or (n94,n95,n694);
not (n95,n96);
nor (n96,n97,n617);
nand (n97,n98,n579);
and (n98,n99,n535);
nor (n99,n100,n484);
nor (n100,n101,n431);
or (n101,n102,n430);
and (n102,n103,n335);
xor (n103,n104,n242);
xor (n104,n105,n224);
xor (n105,n106,n163);
or (n106,n107,n162);
and (n107,n108,n149);
xor (n108,n109,n124);
nand (n109,n110,n117);
or (n110,n111,n67);
not (n111,n112);
nand (n112,n113,n116);
or (n113,n114,n16);
not (n114,n115);
or (n116,n115,n15);
nand (n117,n118,n76);
not (n118,n119);
nor (n119,n120,n122);
and (n120,n121,n15);
and (n122,n16,n123);
not (n123,n121);
nand (n124,n125,n144);
or (n125,n126,n132);
not (n126,n127);
nor (n127,n128,n131);
and (n128,n85,n129);
not (n129,n130);
and (n131,n86,n130);
not (n132,n133);
nor (n133,n134,n139);
nor (n134,n135,n137);
and (n135,n136,n129);
and (n137,n130,n138);
not (n138,n136);
nand (n139,n140,n143);
or (n140,n141,n136);
not (n141,n142);
nand (n143,n136,n141);
or (n144,n145,n146);
not (n145,n139);
nor (n146,n147,n148);
and (n147,n88,n130);
and (n148,n42,n129);
nand (n149,n150,n155);
or (n150,n11,n151);
not (n151,n152);
xnor (n152,n153,n22);
not (n153,n154);
or (n155,n12,n156);
not (n156,n157);
nor (n157,n158,n161);
and (n158,n159,n21);
not (n159,n160);
and (n161,n160,n22);
and (n162,n109,n124);
or (n163,n164,n223);
and (n164,n165,n200);
xor (n165,n166,n181);
nand (n166,n167,n178);
or (n167,n168,n174);
nand (n168,n169,n173);
or (n169,n170,n172);
not (n170,n171);
nand (n173,n172,n170);
nor (n174,n168,n175);
nor (n175,n176,n179);
and (n176,n177,n178);
not (n177,n172);
and (n179,n172,n180);
not (n180,n178);
nand (n181,n182,n196);
or (n182,n183,n192);
nand (n183,n184,n188);
nand (n184,n185,n187);
or (n185,n186,n141);
nand (n187,n141,n186);
not (n188,n189);
nand (n189,n190,n191);
or (n190,n180,n186);
nand (n191,n186,n180);
not (n192,n193);
nor (n193,n194,n195);
and (n194,n33,n141);
and (n195,n34,n142);
or (n196,n188,n197);
nor (n197,n198,n199);
and (n198,n141,n38);
and (n199,n142,n37);
nand (n200,n201,n217);
or (n201,n202,n212);
nand (n202,n203,n209);
not (n203,n204);
nand (n204,n205,n208);
or (n205,n206,n130);
not (n206,n207);
nand (n208,n130,n206);
nand (n209,n210,n211);
nand (n210,n206,n72);
nand (n211,n207,n74);
nor (n212,n213,n216);
and (n213,n214,n72);
not (n214,n215);
and (n216,n215,n74);
or (n217,n203,n218);
nor (n218,n219,n221);
and (n219,n74,n220);
and (n221,n72,n222);
not (n222,n220);
and (n223,n166,n181);
xor (n224,n225,n239);
xor (n225,n226,n232);
nand (n226,n227,n228);
or (n227,n67,n119);
or (n228,n229,n68);
nor (n229,n230,n231);
and (n230,n215,n15);
and (n231,n16,n214);
nand (n232,n233,n238);
or (n233,n234,n12);
not (n234,n235);
nor (n235,n236,n237);
and (n236,n114,n21);
and (n237,n115,n22);
nand (n238,n10,n157);
nand (n239,n240,n241);
or (n240,n183,n197);
or (n241,n188,n141);
xor (n242,n243,n306);
xor (n243,n244,n264);
xor (n244,n245,n257);
xor (n245,n246,n251);
nand (n246,n247,n250);
or (n247,n26,n248);
not (n248,n249);
or (n250,n36,n153);
nand (n251,n252,n253);
or (n252,n218,n202);
or (n253,n203,n254);
nor (n254,n255,n256);
and (n255,n74,n86);
and (n256,n72,n85);
not (n257,n258);
nand (n258,n259,n260);
or (n259,n132,n146);
or (n260,n145,n261);
nor (n261,n262,n263);
and (n262,n33,n130);
and (n263,n34,n129);
or (n264,n265,n305);
and (n265,n266,n280);
xor (n266,n267,n272);
nand (n267,n268,n271);
or (n268,n26,n269);
not (n269,n270);
or (n271,n36,n248);
nand (n272,n273,n279);
or (n273,n274,n278);
not (n274,n275);
nor (n275,n276,n277);
and (n276,n38,n178);
and (n277,n37,n180);
not (n278,n174);
nand (n279,n168,n178);
or (n280,n281,n304);
and (n281,n282,n297);
xor (n282,n283,n290);
nand (n283,n284,n289);
or (n284,n285,n183);
not (n285,n286);
nor (n286,n287,n288);
and (n287,n42,n142);
and (n288,n88,n141);
nand (n289,n189,n193);
nand (n290,n291,n296);
or (n291,n292,n202);
not (n292,n293);
nor (n293,n294,n295);
and (n294,n123,n74);
and (n295,n121,n72);
or (n296,n203,n212);
nand (n297,n298,n299);
or (n298,n111,n68);
nand (n299,n300,n66);
not (n300,n301);
nor (n301,n302,n303);
and (n302,n15,n160);
and (n303,n159,n16);
and (n304,n283,n290);
and (n305,n267,n272);
or (n306,n307,n334);
and (n307,n308,n333);
xor (n308,n309,n332);
or (n309,n310,n331);
and (n310,n311,n326);
xor (n311,n312,n319);
nand (n312,n313,n318);
or (n313,n314,n132);
not (n314,n315);
nor (n315,n316,n317);
and (n316,n222,n129);
and (n317,n220,n130);
nand (n318,n139,n127);
nand (n319,n320,n325);
or (n320,n321,n11);
not (n321,n322);
nand (n322,n323,n324);
or (n323,n22,n248);
or (n324,n21,n249);
nand (n325,n13,n152);
nand (n326,n327,n330);
or (n327,n328,n26);
not (n328,n329);
nand (n330,n30,n270);
and (n331,n312,n319);
xor (n332,n108,n149);
xor (n333,n165,n200);
and (n334,n309,n332);
or (n335,n336,n429);
and (n336,n337,n399);
xor (n337,n338,n339);
xor (n338,n266,n280);
or (n339,n340,n398);
and (n340,n341,n375);
xor (n341,n342,n343);
not (n342,n272);
or (n343,n344,n374);
and (n344,n345,n367);
xor (n345,n346,n360);
nand (n346,n347,n171);
or (n347,n348,n354);
nand (n348,n349,n353);
or (n349,n350,n352);
not (n350,n351);
nand (n353,n350,n352);
not (n354,n355);
nand (n355,n356,n357);
not (n356,n348);
nand (n357,n358,n359);
or (n358,n171,n350);
nand (n359,n350,n171);
nand (n360,n361,n366);
or (n361,n362,n278);
not (n362,n363);
nand (n363,n364,n365);
or (n364,n34,n180);
nand (n365,n180,n34);
nand (n366,n275,n168);
nand (n367,n368,n373);
or (n368,n369,n132);
not (n369,n370);
nand (n370,n371,n372);
or (n371,n130,n214);
or (n372,n129,n215);
nand (n373,n139,n315);
and (n374,n346,n360);
or (n375,n376,n397);
and (n376,n377,n390);
xor (n377,n378,n383);
nand (n378,n379,n382);
or (n379,n380,n26);
not (n380,n381);
nand (n382,n30,n329);
nand (n383,n384,n389);
or (n384,n385,n202);
not (n385,n386);
nor (n386,n387,n388);
and (n387,n114,n74);
and (n388,n115,n72);
nand (n389,n204,n293);
nand (n390,n391,n396);
or (n391,n183,n392);
not (n392,n393);
nor (n393,n394,n395);
and (n394,n85,n141);
and (n395,n86,n142);
or (n396,n188,n285);
and (n397,n378,n383);
and (n398,n342,n343);
or (n399,n400,n428);
and (n400,n401,n404);
xor (n401,n402,n403);
xor (n402,n311,n326);
xor (n403,n282,n297);
or (n404,n405,n427);
and (n405,n406,n420);
xor (n406,n407,n413);
nand (n407,n408,n412);
or (n408,n409,n67);
nor (n409,n410,n411);
and (n410,n16,n153);
and (n411,n15,n154);
nand (n412,n300,n76);
nand (n413,n414,n419);
or (n414,n415,n11);
not (n415,n416);
nor (n416,n417,n418);
and (n417,n269,n21);
and (n418,n270,n22);
nand (n419,n13,n322);
not (n420,n421);
nor (n421,n422,n426);
and (n422,n354,n423);
nor (n423,n424,n425);
and (n424,n37,n170);
and (n425,n38,n171);
nor (n426,n356,n170);
and (n427,n407,n413);
and (n428,n402,n403);
and (n429,n338,n339);
and (n430,n104,n242);
xor (n431,n432,n481);
xor (n432,n433,n436);
or (n433,n434,n435);
and (n434,n105,n224);
and (n435,n106,n163);
xor (n436,n437,n459);
xor (n437,n438,n456);
xor (n438,n439,n450);
xor (n439,n440,n443);
nand (n440,n441,n142);
or (n441,n442,n189);
not (n442,n183);
nand (n443,n444,n445);
or (n444,n261,n132);
nand (n445,n446,n139);
not (n446,n447);
nor (n447,n448,n449);
and (n448,n129,n38);
and (n449,n130,n37);
nand (n450,n451,n452);
or (n451,n229,n67);
or (n452,n68,n453);
nor (n453,n454,n455);
and (n454,n15,n220);
and (n455,n16,n222);
or (n456,n457,n458);
and (n457,n245,n257);
and (n458,n246,n251);
xor (n459,n460,n464);
xor (n460,n258,n461);
or (n461,n462,n463);
and (n462,n225,n239);
and (n463,n226,n232);
xor (n464,n465,n478);
xor (n465,n466,n472);
nand (n466,n467,n468);
or (n467,n234,n11);
nand (n468,n13,n469);
nor (n469,n470,n471);
and (n470,n123,n21);
and (n471,n121,n22);
nand (n472,n473,n474);
or (n473,n254,n202);
or (n474,n203,n475);
nor (n475,n476,n477);
and (n476,n88,n72);
and (n477,n42,n74);
nand (n478,n479,n480);
or (n479,n153,n26);
or (n480,n36,n159);
or (n481,n482,n483);
and (n482,n243,n306);
and (n483,n244,n264);
nor (n484,n485,n532);
xor (n485,n486,n529);
xor (n486,n487,n490);
or (n487,n488,n489);
and (n488,n460,n464);
and (n489,n258,n461);
xor (n490,n491,n510);
xor (n491,n492,n495);
or (n492,n493,n494);
and (n493,n439,n450);
and (n494,n440,n443);
xor (n495,n496,n507);
xor (n496,n497,n504);
nand (n497,n498,n500);
or (n498,n11,n499);
not (n499,n469);
or (n500,n12,n501);
nor (n501,n502,n503);
and (n502,n21,n215);
and (n503,n22,n214);
nand (n504,n505,n506);
or (n505,n159,n26);
nand (n506,n30,n115);
nand (n507,n508,n509);
or (n508,n132,n447);
or (n509,n145,n129);
xor (n510,n511,n526);
xor (n511,n512,n518);
nand (n512,n513,n514);
or (n513,n67,n453);
or (n514,n68,n515);
nor (n515,n516,n517);
and (n516,n15,n86);
and (n517,n16,n85);
not (n518,n519);
nand (n519,n520,n525);
or (n520,n521,n203);
not (n521,n522);
nand (n522,n523,n524);
or (n523,n72,n33);
or (n524,n74,n34);
or (n525,n202,n475);
or (n526,n527,n528);
and (n527,n465,n478);
and (n528,n466,n472);
or (n529,n530,n531);
and (n530,n437,n459);
and (n531,n438,n456);
or (n532,n533,n534);
and (n533,n432,n481);
and (n534,n433,n436);
or (n535,n536,n576);
xor (n536,n537,n573);
xor (n537,n538,n541);
or (n538,n539,n540);
and (n539,n511,n526);
and (n540,n512,n518);
xor (n541,n542,n562);
xor (n542,n543,n546);
or (n543,n544,n545);
and (n544,n496,n507);
and (n545,n497,n504);
xor (n546,n547,n556);
xor (n547,n548,n550);
nand (n548,n549,n130);
or (n549,n139,n133);
nand (n550,n551,n552);
or (n551,n202,n521);
or (n552,n203,n553);
nor (n553,n554,n555);
and (n554,n74,n38);
and (n555,n72,n37);
nand (n556,n557,n558);
or (n557,n11,n501);
or (n558,n12,n559);
nor (n559,n560,n561);
and (n560,n21,n220);
and (n561,n22,n222);
xor (n562,n563,n519);
xor (n563,n564,n567);
nand (n564,n565,n566);
or (n565,n26,n114);
or (n566,n36,n123);
nand (n567,n568,n569);
or (n568,n67,n515);
or (n569,n68,n570);
nor (n570,n571,n572);
and (n571,n15,n42);
and (n572,n16,n88);
or (n573,n574,n575);
and (n574,n491,n510);
and (n575,n492,n495);
or (n576,n577,n578);
and (n577,n486,n529);
and (n578,n487,n490);
or (n579,n580,n583);
or (n580,n581,n582);
and (n581,n537,n573);
and (n582,n538,n541);
xor (n583,n584,n614);
xor (n584,n585,n588);
or (n585,n586,n587);
and (n586,n563,n519);
and (n587,n564,n567);
xor (n588,n589,n597);
xor (n589,n590,n594);
not (n590,n591);
nand (n591,n592,n593);
or (n592,n202,n553);
or (n593,n203,n74);
or (n594,n595,n596);
and (n595,n547,n556);
and (n596,n548,n550);
xor (n597,n598,n608);
xor (n598,n599,n602);
nand (n599,n600,n601);
or (n600,n123,n26);
nand (n601,n30,n215);
nand (n602,n603,n604);
or (n603,n67,n570);
or (n604,n68,n605);
nor (n605,n606,n607);
and (n606,n15,n34);
and (n607,n16,n33);
nand (n608,n609,n610);
or (n609,n11,n559);
or (n610,n12,n611);
nor (n611,n612,n613);
and (n612,n21,n86);
and (n613,n22,n85);
or (n614,n615,n616);
and (n615,n542,n562);
and (n616,n543,n546);
nand (n617,n618,n647,n689);
not (n618,n619);
nor (n619,n620,n646);
or (n620,n621,n645);
and (n621,n622,n632);
xor (n622,n623,n631);
not (n623,n624);
nor (n624,n625,n630);
and (n625,n66,n626);
not (n626,n627);
nor (n627,n628,n629);
and (n628,n15,n38);
and (n629,n16,n37);
and (n630,n76,n16);
xor (n631,n63,n83);
or (n632,n633,n644);
and (n633,n634,n624);
xor (n634,n635,n641);
nand (n635,n636,n640);
or (n636,n11,n637);
nor (n637,n638,n639);
and (n638,n21,n42);
and (n639,n22,n88);
or (n640,n12,n79);
nand (n641,n642,n643);
or (n642,n26,n222);
or (n643,n36,n85);
and (n644,n635,n641);
and (n645,n623,n631);
xor (n646,n54,n61);
nor (n647,n648,n676);
nor (n648,n649,n652);
or (n649,n650,n651);
and (n650,n584,n614);
and (n651,n585,n588);
xor (n652,n653,n673);
xor (n653,n654,n665);
xor (n654,n655,n662);
xor (n655,n656,n659);
nand (n656,n657,n72);
or (n657,n658,n204);
not (n658,n202);
nand (n659,n660,n661);
or (n660,n67,n605);
or (n661,n68,n627);
nand (n662,n663,n664);
or (n663,n26,n214);
or (n664,n36,n222);
xor (n665,n666,n670);
xor (n666,n667,n591);
nand (n667,n668,n669);
or (n668,n11,n611);
or (n669,n12,n637);
or (n670,n671,n672);
and (n671,n598,n608);
and (n672,n599,n602);
or (n673,n674,n675);
and (n674,n589,n597);
and (n675,n590,n594);
nor (n676,n677,n680);
or (n677,n678,n679);
and (n678,n653,n673);
and (n679,n654,n665);
xor (n680,n681,n686);
xor (n681,n682,n685);
or (n682,n683,n684);
and (n683,n655,n662);
and (n684,n656,n659);
xor (n685,n634,n624);
or (n686,n687,n688);
and (n687,n666,n670);
and (n688,n667,n591);
or (n689,n690,n693);
or (n690,n691,n692);
and (n691,n681,n686);
and (n692,n682,n685);
xor (n693,n622,n632);
not (n694,n695);
nand (n695,n696,n1399);
nor (n696,n697,n1385);
and (n697,n698,n1060);
and (n698,n699,n1043);
nor (n699,n700,n955);
nor (n700,n701,n875);
xor (n701,n702,n783);
xor (n702,n703,n730);
or (n703,n704,n729);
and (n704,n705,n708);
xor (n705,n706,n707);
xor (n706,n377,n390);
xor (n707,n406,n420);
or (n708,n709,n728);
and (n709,n710,n718);
xor (n710,n711,n421);
nand (n711,n712,n717);
or (n712,n713,n11);
not (n713,n714);
nor (n714,n715,n716);
and (n715,n328,n21);
and (n716,n329,n22);
nand (n717,n13,n416);
nand (n718,n719,n352);
nor (n719,n720,n724);
and (n720,n442,n721);
nor (n721,n722,n723);
and (n722,n214,n141);
and (n723,n215,n142);
and (n724,n189,n725);
nor (n725,n726,n727);
and (n726,n222,n141);
and (n727,n220,n142);
and (n728,n711,n421);
and (n729,n706,n707);
xor (n730,n731,n782);
xor (n731,n732,n733);
xor (n732,n341,n375);
or (n733,n734,n781);
and (n734,n735,n780);
xor (n735,n736,n757);
or (n736,n737,n756);
and (n737,n738,n750);
xor (n738,n739,n746);
nand (n739,n740,n745);
or (n740,n741,n202);
not (n741,n742);
nand (n742,n743,n744);
or (n743,n160,n74);
nand (n744,n74,n160);
nand (n745,n386,n204);
nand (n746,n747,n749);
or (n747,n748,n183);
not (n748,n725);
nand (n749,n189,n393);
nand (n750,n751,n755);
or (n751,n67,n752);
nor (n752,n753,n754);
and (n753,n249,n15);
and (n754,n16,n248);
or (n755,n409,n68);
and (n756,n739,n746);
or (n757,n758,n779);
and (n758,n759,n772);
xor (n759,n760,n767);
nand (n760,n761,n766);
or (n761,n762,n278);
not (n762,n763);
nor (n763,n764,n765);
and (n764,n88,n180);
and (n765,n42,n178);
nand (n766,n363,n168);
nand (n767,n768,n771);
or (n768,n769,n26);
not (n769,n770);
nand (n771,n30,n381);
nand (n772,n773,n778);
or (n773,n774,n132);
not (n774,n775);
nor (n775,n776,n777);
and (n776,n123,n129);
and (n777,n121,n130);
nand (n778,n139,n370);
and (n779,n760,n767);
xor (n780,n345,n367);
and (n781,n736,n757);
xor (n782,n401,n404);
or (n783,n784,n874);
and (n784,n785,n839);
xor (n785,n786,n787);
xor (n786,n735,n780);
or (n787,n788,n838);
and (n788,n789,n837);
xor (n789,n790,n814);
or (n790,n791,n813);
and (n791,n792,n805);
xor (n792,n793,n800);
nand (n793,n794,n799);
or (n794,n795,n11);
not (n795,n796);
nor (n796,n797,n798);
and (n797,n380,n21);
and (n798,n381,n22);
nand (n799,n714,n13);
nand (n800,n801,n804);
or (n801,n802,n26);
not (n802,n803);
nand (n804,n30,n770);
nand (n805,n806,n808);
or (n806,n807,n356);
not (n807,n423);
or (n808,n355,n809);
not (n809,n810);
or (n810,n811,n812);
and (n811,n33,n171);
and (n812,n34,n170);
and (n813,n793,n800);
or (n814,n815,n836);
and (n815,n816,n830);
xor (n816,n817,n824);
nand (n817,n818,n823);
or (n818,n819,n132);
not (n819,n820);
nor (n820,n821,n822);
and (n821,n114,n129);
and (n822,n115,n130);
nand (n823,n139,n775);
nand (n824,n825,n829);
or (n825,n826,n278);
nor (n826,n827,n828);
and (n827,n85,n178);
and (n828,n86,n180);
nand (n829,n763,n168);
nand (n830,n831,n835);
or (n831,n202,n832);
nor (n832,n833,n834);
and (n833,n74,n154);
and (n834,n72,n153);
or (n835,n203,n741);
and (n836,n817,n824);
xor (n837,n738,n750);
and (n838,n790,n814);
or (n839,n840,n873);
and (n840,n841,n844);
xor (n841,n842,n843);
xor (n842,n759,n772);
xor (n843,n710,n718);
and (n844,n845,n867);
or (n845,n846,n866);
and (n846,n847,n861);
xor (n847,n848,n854);
nand (n848,n849,n853);
or (n849,n850,n183);
nor (n850,n851,n852);
and (n851,n123,n142);
and (n852,n121,n141);
nand (n853,n721,n189);
nand (n854,n855,n860);
or (n855,n856,n11);
not (n856,n857);
nand (n857,n858,n859);
or (n858,n22,n769);
or (n859,n21,n770);
nand (n860,n13,n796);
nand (n861,n862,n865);
or (n862,n863,n26);
not (n863,n864);
nand (n865,n30,n803);
and (n866,n848,n854);
nand (n867,n868,n872);
or (n868,n67,n869);
nor (n869,n870,n871);
and (n870,n15,n270);
and (n871,n16,n269);
or (n872,n68,n752);
and (n873,n842,n843);
and (n874,n786,n787);
or (n875,n876,n954);
and (n876,n877,n880);
xor (n877,n878,n879);
xor (n878,n705,n708);
xor (n879,n785,n839);
or (n880,n881,n953);
and (n881,n882,n917);
xor (n882,n883,n884);
xor (n883,n789,n837);
or (n884,n885,n916);
and (n885,n886,n914);
xor (n886,n887,n913);
or (n887,n888,n912);
and (n888,n889,n904);
xor (n889,n890,n897);
nand (n890,n891,n896);
or (n891,n892,n355);
not (n892,n893);
nor (n893,n894,n895);
and (n894,n88,n170);
and (n895,n42,n171);
nand (n896,n348,n810);
nand (n897,n898,n903);
or (n898,n899,n132);
not (n899,n900);
nand (n900,n901,n902);
or (n901,n130,n159);
or (n902,n129,n160);
nand (n903,n139,n820);
nand (n904,n905,n910);
or (n905,n278,n906);
not (n906,n907);
nor (n907,n908,n909);
and (n908,n180,n222);
and (n909,n220,n178);
or (n910,n826,n911);
not (n911,n168);
and (n912,n890,n897);
xor (n913,n816,n830);
nand (n914,n915,n718);
or (n915,n352,n719);
and (n916,n887,n913);
or (n917,n918,n952);
and (n918,n919,n951);
xor (n919,n920,n921);
xor (n920,n792,n805);
or (n921,n922,n950);
and (n922,n923,n939);
xor (n923,n924,n932);
nand (n924,n925,n930);
or (n925,n926,n202);
not (n926,n927);
nor (n927,n928,n929);
and (n928,n248,n74);
and (n929,n249,n72);
nand (n930,n931,n204);
not (n931,n832);
nand (n932,n933,n938);
or (n933,n934,n67);
not (n934,n935);
nand (n935,n936,n937);
or (n936,n16,n328);
or (n937,n15,n329);
or (n938,n68,n869);
nand (n939,n940,n949);
or (n940,n941,n944);
nand (n941,n942,n352);
not (n942,n943);
not (n944,n945);
nor (n945,n946,n948);
and (n946,n37,n947);
not (n947,n352);
and (n948,n38,n352);
or (n949,n947,n942);
and (n950,n924,n932);
xor (n951,n845,n867);
and (n952,n920,n921);
and (n953,n883,n884);
and (n954,n878,n879);
nor (n955,n956,n957);
xor (n956,n877,n880);
or (n957,n958,n1042);
and (n958,n959,n1041);
xor (n959,n960,n961);
xor (n960,n841,n844);
or (n961,n962,n1040);
and (n962,n963,n1039);
xor (n963,n964,n1032);
or (n964,n965,n1031);
and (n965,n966,n1008);
xor (n966,n967,n985);
or (n967,n968,n984);
and (n968,n969,n977);
xor (n969,n970,n971);
and (n970,n30,n864);
nand (n971,n972,n973);
or (n972,n942,n944);
or (n973,n974,n941);
nor (n974,n975,n976);
and (n975,n947,n34);
and (n976,n352,n33);
nand (n977,n978,n983);
or (n978,n355,n979);
not (n979,n980);
nor (n980,n981,n982);
and (n981,n85,n170);
and (n982,n86,n171);
nand (n983,n348,n893);
and (n984,n970,n971);
or (n985,n986,n1007);
and (n986,n987,n1001);
xor (n987,n988,n995);
nand (n988,n989,n994);
or (n989,n990,n278);
not (n990,n991);
nand (n991,n992,n993);
or (n992,n178,n214);
or (n993,n180,n215);
nand (n994,n907,n168);
nand (n995,n996,n1000);
or (n996,n997,n202);
nor (n997,n998,n999);
and (n998,n269,n72);
and (n999,n270,n74);
nand (n1000,n927,n204);
nand (n1001,n1002,n1003);
or (n1002,n934,n68);
or (n1003,n67,n1004);
nor (n1004,n1005,n1006);
and (n1005,n381,n15);
and (n1006,n16,n380);
and (n1007,n988,n995);
or (n1008,n1009,n1030);
and (n1009,n1010,n1024);
xor (n1010,n1011,n1018);
nand (n1011,n1012,n1017);
or (n1012,n1013,n11);
not (n1013,n1014);
nand (n1014,n1015,n1016);
or (n1015,n22,n802);
or (n1016,n21,n803);
nand (n1017,n857,n13);
nand (n1018,n1019,n1023);
or (n1019,n183,n1020);
nor (n1020,n1021,n1022);
and (n1021,n114,n142);
and (n1022,n115,n141);
or (n1023,n188,n850);
nand (n1024,n1025,n1029);
or (n1025,n132,n1026);
nor (n1026,n1027,n1028);
and (n1027,n153,n130);
and (n1028,n154,n129);
or (n1029,n145,n899);
and (n1030,n1011,n1018);
and (n1031,n967,n985);
or (n1032,n1033,n1038);
and (n1033,n1034,n1037);
xor (n1034,n1035,n1036);
xor (n1035,n847,n861);
xor (n1036,n889,n904);
xor (n1037,n923,n939);
and (n1038,n1035,n1036);
xor (n1039,n886,n914);
and (n1040,n964,n1032);
xor (n1041,n882,n917);
and (n1042,n960,n961);
nor (n1043,n1044,n1055);
nor (n1044,n1045,n1052);
xor (n1045,n1046,n1049);
xor (n1046,n1047,n1048);
xor (n1047,n308,n333);
xor (n1048,n337,n399);
or (n1049,n1050,n1051);
and (n1050,n731,n782);
and (n1051,n732,n733);
or (n1052,n1053,n1054);
and (n1053,n702,n783);
and (n1054,n703,n730);
nor (n1055,n1056,n1057);
xor (n1056,n103,n335);
or (n1057,n1058,n1059);
and (n1058,n1046,n1049);
and (n1059,n1047,n1048);
nand (n1060,n1061,n1379);
or (n1061,n1062,n1361);
not (n1062,n1063);
nor (n1063,n1064,n1360);
and (n1064,n1065,n1301);
nand (n1065,n1066,n1209);
xor (n1066,n1067,n1196);
xor (n1067,n1068,n1069);
xor (n1068,n1034,n1037);
or (n1069,n1070,n1195);
and (n1070,n1071,n1166);
xor (n1071,n1072,n1119);
or (n1072,n1073,n1118);
and (n1073,n1074,n1094);
xor (n1074,n1075,n1081);
nand (n1075,n1076,n1080);
or (n1076,n67,n1077);
nor (n1077,n1078,n1079);
and (n1078,n15,n770);
and (n1079,n16,n769);
or (n1080,n68,n1004);
xor (n1081,n1082,n1088);
nor (n1082,n1083,n21);
nor (n1083,n1084,n1086);
and (n1084,n1085,n15);
nand (n1085,n864,n17);
and (n1086,n863,n1087);
not (n1087,n17);
nand (n1088,n1089,n1093);
or (n1089,n1090,n941);
nor (n1090,n1091,n1092);
and (n1091,n88,n352);
and (n1092,n42,n947);
or (n1093,n974,n942);
or (n1094,n1095,n1117);
and (n1095,n1096,n1106);
xor (n1096,n1097,n1098);
nor (n1097,n12,n863);
nand (n1098,n1099,n1104);
or (n1099,n941,n1100);
not (n1100,n1101);
nor (n1101,n1102,n1103);
and (n1102,n85,n947);
and (n1103,n86,n352);
nand (n1104,n1105,n943);
not (n1105,n1090);
nand (n1106,n1107,n1112);
or (n1107,n355,n1108);
not (n1108,n1109);
nand (n1109,n1110,n1111);
or (n1110,n171,n214);
or (n1111,n170,n215);
or (n1112,n356,n1113);
not (n1113,n1114);
nand (n1114,n1115,n1116);
or (n1115,n171,n222);
or (n1116,n170,n220);
and (n1117,n1097,n1098);
and (n1118,n1075,n1081);
xor (n1119,n1120,n1143);
xor (n1120,n1121,n1122);
and (n1121,n1082,n1088);
or (n1122,n1123,n1142);
and (n1123,n1124,n1135);
xor (n1124,n1125,n1128);
nand (n1125,n1126,n1127);
or (n1126,n1113,n355);
nand (n1127,n348,n980);
nand (n1128,n1129,n1134);
or (n1129,n1130,n11);
not (n1130,n1131);
nand (n1131,n1132,n1133);
or (n1132,n21,n864);
or (n1133,n22,n863);
nand (n1134,n1014,n13);
nand (n1135,n1136,n1141);
or (n1136,n183,n1137);
not (n1137,n1138);
nor (n1138,n1139,n1140);
and (n1139,n159,n141);
and (n1140,n160,n142);
or (n1141,n188,n1020);
and (n1142,n1125,n1128);
or (n1143,n1144,n1165);
and (n1144,n1145,n1159);
xor (n1145,n1146,n1153);
nand (n1146,n1147,n1152);
or (n1147,n1148,n132);
not (n1148,n1149);
nor (n1149,n1150,n1151);
and (n1150,n248,n129);
and (n1151,n249,n130);
or (n1152,n1026,n145);
nand (n1153,n1154,n1158);
or (n1154,n1155,n278);
nor (n1155,n1156,n1157);
and (n1156,n180,n121);
and (n1157,n178,n123);
nand (n1158,n168,n991);
nand (n1159,n1160,n1164);
or (n1160,n202,n1161);
nor (n1161,n1162,n1163);
and (n1162,n74,n329);
and (n1163,n72,n328);
or (n1164,n203,n997);
and (n1165,n1146,n1153);
or (n1166,n1167,n1194);
and (n1167,n1168,n1193);
xor (n1168,n1169,n1192);
or (n1169,n1170,n1191);
and (n1170,n1171,n1185);
xor (n1171,n1172,n1179);
nand (n1172,n1173,n1178);
or (n1173,n1174,n183);
not (n1174,n1175);
nand (n1175,n1176,n1177);
or (n1176,n142,n153);
or (n1177,n141,n154);
nand (n1178,n189,n1138);
nand (n1179,n1180,n1184);
or (n1180,n132,n1181);
nor (n1181,n1182,n1183);
and (n1182,n129,n270);
and (n1183,n130,n269);
nand (n1184,n139,n1149);
nand (n1185,n1186,n1190);
or (n1186,n278,n1187);
nor (n1187,n1188,n1189);
and (n1188,n180,n115);
and (n1189,n178,n114);
or (n1190,n1155,n911);
and (n1191,n1172,n1179);
xor (n1192,n1145,n1159);
xor (n1193,n1124,n1135);
and (n1194,n1169,n1192);
and (n1195,n1072,n1119);
xor (n1196,n1197,n1202);
xor (n1197,n1198,n1201);
or (n1198,n1199,n1200);
and (n1199,n1120,n1143);
and (n1200,n1121,n1122);
xor (n1201,n966,n1008);
or (n1202,n1203,n1208);
and (n1203,n1204,n1207);
xor (n1204,n1205,n1206);
xor (n1205,n987,n1001);
xor (n1206,n969,n977);
xor (n1207,n1010,n1024);
and (n1208,n1205,n1206);
or (n1209,n1210,n1300);
and (n1210,n1211,n1299);
xor (n1211,n1212,n1213);
xor (n1212,n1204,n1207);
or (n1213,n1214,n1298);
and (n1214,n1215,n1246);
xor (n1215,n1216,n1245);
or (n1216,n1217,n1244);
and (n1217,n1218,n1232);
xor (n1218,n1219,n1226);
nand (n1219,n1220,n1224);
or (n1220,n1221,n202);
nor (n1221,n1222,n1223);
and (n1222,n380,n72);
and (n1223,n381,n74);
nand (n1224,n1225,n204);
not (n1225,n1161);
nand (n1226,n1227,n1231);
or (n1227,n1228,n67);
nor (n1228,n1229,n1230);
and (n1229,n15,n803);
and (n1230,n16,n802);
or (n1231,n68,n1077);
and (n1232,n1233,n1238);
nor (n1233,n1234,n15);
nor (n1234,n1235,n1237);
and (n1235,n1236,n74);
nand (n1236,n864,n71);
and (n1237,n863,n70);
nand (n1238,n1239,n1240);
or (n1239,n942,n1100);
or (n1240,n1241,n941);
nor (n1241,n1242,n1243);
and (n1242,n222,n352);
and (n1243,n220,n947);
and (n1244,n1219,n1226);
xor (n1245,n1074,n1094);
or (n1246,n1247,n1297);
and (n1247,n1248,n1296);
xor (n1248,n1249,n1274);
or (n1249,n1250,n1273);
and (n1250,n1251,n1266);
xor (n1251,n1252,n1259);
nand (n1252,n1253,n1258);
or (n1253,n1254,n355);
not (n1254,n1255);
nor (n1255,n1256,n1257);
and (n1256,n123,n170);
and (n1257,n121,n171);
nand (n1258,n1109,n348);
nand (n1259,n1260,n1265);
or (n1260,n1261,n183);
not (n1261,n1262);
nand (n1262,n1263,n1264);
or (n1263,n142,n248);
or (n1264,n141,n249);
nand (n1265,n189,n1175);
nand (n1266,n1267,n1272);
or (n1267,n132,n1268);
not (n1268,n1269);
nand (n1269,n1270,n1271);
or (n1270,n130,n328);
or (n1271,n129,n329);
or (n1272,n145,n1181);
and (n1273,n1252,n1259);
or (n1274,n1275,n1295);
and (n1275,n1276,n1289);
xor (n1276,n1277,n1283);
nand (n1277,n1278,n1282);
or (n1278,n278,n1279);
nor (n1279,n1280,n1281);
and (n1280,n180,n160);
and (n1281,n178,n159);
or (n1282,n1187,n911);
nand (n1283,n1284,n1288);
or (n1284,n202,n1285);
nor (n1285,n1286,n1287);
and (n1286,n74,n770);
and (n1287,n72,n769);
or (n1288,n1221,n203);
nand (n1289,n1290,n1294);
or (n1290,n67,n1291);
nor (n1291,n1292,n1293);
and (n1292,n863,n16);
and (n1293,n864,n15);
or (n1294,n1228,n68);
and (n1295,n1277,n1283);
xor (n1296,n1096,n1106);
and (n1297,n1249,n1274);
and (n1298,n1216,n1245);
xor (n1299,n1071,n1166);
and (n1300,n1212,n1213);
nand (n1301,n1302,n1303);
xor (n1302,n1211,n1299);
or (n1303,n1304,n1359);
and (n1304,n1305,n1358);
xor (n1305,n1306,n1307);
xor (n1306,n1168,n1193);
or (n1307,n1308,n1357);
and (n1308,n1309,n1312);
xor (n1309,n1310,n1311);
xor (n1310,n1171,n1185);
xor (n1311,n1218,n1232);
or (n1312,n1313,n1356);
and (n1313,n1314,n1334);
xor (n1314,n1315,n1316);
xor (n1315,n1233,n1238);
or (n1316,n1317,n1333);
and (n1317,n1318,n1327);
xor (n1318,n1319,n1320);
and (n1319,n76,n864);
nand (n1320,n1321,n1326);
or (n1321,n1322,n355);
not (n1322,n1323);
nand (n1323,n1324,n1325);
or (n1324,n171,n114);
or (n1325,n170,n115);
nand (n1326,n348,n1255);
nand (n1327,n1328,n1329);
or (n1328,n1261,n188);
or (n1329,n183,n1330);
nor (n1330,n1331,n1332);
and (n1331,n269,n142);
and (n1332,n270,n141);
and (n1333,n1319,n1320);
or (n1334,n1335,n1355);
and (n1335,n1336,n1349);
xor (n1336,n1337,n1343);
nand (n1337,n1338,n1342);
or (n1338,n1339,n132);
nor (n1339,n1340,n1341);
and (n1340,n380,n130);
and (n1341,n381,n129);
nand (n1342,n1269,n139);
nand (n1343,n1344,n1348);
or (n1344,n1345,n941);
nor (n1345,n1346,n1347);
and (n1346,n947,n215);
and (n1347,n352,n214);
or (n1348,n1241,n942);
nand (n1349,n1350,n1354);
or (n1350,n1351,n202);
nor (n1351,n1352,n1353);
and (n1352,n74,n803);
and (n1353,n72,n802);
or (n1354,n1285,n203);
and (n1355,n1337,n1343);
and (n1356,n1315,n1316);
and (n1357,n1310,n1311);
xor (n1358,n1215,n1246);
and (n1359,n1306,n1307);
nor (n1360,n1066,n1209);
not (n1361,n1362);
nor (n1362,n1363,n1374);
nor (n1363,n1364,n1365);
xor (n1364,n959,n1041);
or (n1365,n1366,n1373);
and (n1366,n1367,n1372);
xor (n1367,n1368,n1369);
xor (n1368,n919,n951);
or (n1369,n1370,n1371);
and (n1370,n1197,n1202);
and (n1371,n1198,n1201);
xor (n1372,n963,n1039);
and (n1373,n1368,n1369);
nor (n1374,n1375,n1376);
xor (n1375,n1367,n1372);
or (n1376,n1377,n1378);
and (n1377,n1067,n1196);
and (n1378,n1068,n1069);
nor (n1379,n1380,n1384);
and (n1380,n1381,n1382);
not (n1381,n1363);
not (n1382,n1383);
nand (n1383,n1375,n1376);
and (n1384,n1364,n1365);
nand (n1385,n1386,n1393);
or (n1386,n1387,n1388);
not (n1387,n1043);
not (n1388,n1389);
nor (n1389,n1390,n700);
and (n1390,n1391,n1392);
nand (n1391,n875,n701);
nand (n1392,n956,n957);
nor (n1393,n1394,n1398);
and (n1394,n1395,n1396);
not (n1395,n1055);
not (n1396,n1397);
nand (n1397,n1045,n1052);
and (n1398,n1056,n1057);
nand (n1399,n698,n1400,n1403);
and (n1400,n1362,n1401);
nor (n1401,n1360,n1402);
nor (n1402,n1302,n1303);
nand (n1403,n1404,n1905);
or (n1404,n1405,n1841);
not (n1405,n1406);
nand (n1406,n1407,n1830,n1840);
nand (n1407,n1408,n1586,n1690);
nand (n1408,n1409,n1550);
not (n1409,n1410);
xor (n1410,n1411,n1509);
xor (n1411,n1412,n1447);
xor (n1412,n1413,n1429);
xor (n1413,n1414,n1420);
nand (n1414,n1415,n1419);
or (n1415,n202,n1416);
nor (n1416,n1417,n1418);
and (n1417,n863,n72);
and (n1418,n74,n864);
or (n1419,n203,n1351);
nand (n1420,n1421,n1425);
or (n1421,n278,n1422);
nor (n1422,n1423,n1424);
and (n1423,n180,n249);
and (n1424,n178,n248);
or (n1425,n1426,n911);
nor (n1426,n1427,n1428);
and (n1427,n180,n154);
and (n1428,n178,n153);
nand (n1429,n1430,n1446);
or (n1430,n1431,n1438);
not (n1431,n1432);
nand (n1432,n1433,n72);
nand (n1433,n1434,n1435);
or (n1434,n864,n207);
nand (n1435,n1436,n129);
not (n1436,n1437);
and (n1437,n864,n207);
not (n1438,n1439);
nand (n1439,n1440,n1445);
or (n1440,n1441,n355);
not (n1441,n1442);
nand (n1442,n1443,n1444);
or (n1443,n171,n159);
or (n1444,n170,n160);
nand (n1445,n348,n1323);
or (n1446,n1439,n1432);
xor (n1447,n1448,n1498);
xor (n1448,n1449,n1470);
or (n1449,n1450,n1469);
and (n1450,n1451,n1459);
xor (n1451,n1452,n1453);
and (n1452,n204,n864);
nand (n1453,n1454,n1458);
or (n1454,n1455,n355);
nor (n1455,n1456,n1457);
and (n1456,n153,n171);
and (n1457,n154,n170);
nand (n1458,n348,n1442);
nand (n1459,n1460,n1465);
or (n1460,n183,n1461);
not (n1461,n1462);
nor (n1462,n1463,n1464);
and (n1463,n380,n141);
and (n1464,n381,n142);
or (n1465,n188,n1466);
nor (n1466,n1467,n1468);
and (n1467,n329,n141);
and (n1468,n328,n142);
and (n1469,n1452,n1453);
or (n1470,n1471,n1497);
and (n1471,n1472,n1491);
xor (n1472,n1473,n1482);
nand (n1473,n1474,n1478);
or (n1474,n132,n1475);
nor (n1475,n1476,n1477);
and (n1476,n802,n130);
and (n1477,n803,n129);
or (n1478,n145,n1479);
nor (n1479,n1480,n1481);
and (n1480,n770,n129);
and (n1481,n769,n130);
nand (n1482,n1483,n1487);
or (n1483,n1484,n941);
nor (n1484,n1485,n1486);
and (n1485,n947,n115);
and (n1486,n352,n114);
or (n1487,n1488,n942);
nor (n1488,n1489,n1490);
and (n1489,n947,n121);
and (n1490,n352,n123);
nand (n1491,n1492,n1496);
or (n1492,n278,n1493);
nor (n1493,n1494,n1495);
and (n1494,n180,n270);
and (n1495,n178,n269);
or (n1496,n1422,n911);
and (n1497,n1473,n1482);
xor (n1498,n1499,n1506);
xor (n1499,n1500,n1503);
nand (n1500,n1501,n1502);
or (n1501,n183,n1466);
or (n1502,n1330,n188);
nand (n1503,n1504,n1505);
or (n1504,n132,n1479);
or (n1505,n145,n1339);
nand (n1506,n1507,n1508);
or (n1507,n1488,n941);
or (n1508,n1345,n942);
or (n1509,n1510,n1549);
and (n1510,n1511,n1548);
xor (n1511,n1512,n1525);
and (n1512,n1513,n1519);
and (n1513,n1514,n130);
nand (n1514,n1515,n1516);
or (n1515,n864,n136);
nand (n1516,n1517,n141);
not (n1517,n1518);
and (n1518,n864,n136);
nand (n1519,n1520,n1524);
or (n1520,n355,n1521);
nor (n1521,n1522,n1523);
and (n1522,n170,n249);
and (n1523,n171,n248);
or (n1524,n356,n1455);
or (n1525,n1526,n1547);
and (n1526,n1527,n1541);
xor (n1527,n1528,n1535);
nand (n1528,n1529,n1534);
or (n1529,n1530,n183);
not (n1530,n1531);
nor (n1531,n1532,n1533);
and (n1532,n770,n142);
and (n1533,n769,n141);
nand (n1534,n189,n1462);
nand (n1535,n1536,n1540);
or (n1536,n132,n1537);
nor (n1537,n1538,n1539);
and (n1538,n130,n863);
and (n1539,n129,n864);
or (n1540,n145,n1475);
nand (n1541,n1542,n1546);
or (n1542,n941,n1543);
nor (n1543,n1544,n1545);
and (n1544,n947,n160);
and (n1545,n352,n159);
or (n1546,n1484,n942);
and (n1547,n1528,n1535);
xor (n1548,n1451,n1459);
and (n1549,n1512,n1525);
not (n1550,n1551);
or (n1551,n1552,n1585);
and (n1552,n1553,n1584);
xor (n1553,n1554,n1555);
xor (n1554,n1472,n1491);
or (n1555,n1556,n1583);
and (n1556,n1557,n1565);
xor (n1557,n1558,n1564);
nand (n1558,n1559,n1563);
or (n1559,n278,n1560);
nor (n1560,n1561,n1562);
and (n1561,n180,n329);
and (n1562,n178,n328);
or (n1563,n1493,n911);
xor (n1564,n1513,n1519);
or (n1565,n1566,n1582);
and (n1566,n1567,n1575);
xor (n1567,n1568,n1569);
and (n1568,n139,n864);
nand (n1569,n1570,n1574);
or (n1570,n1571,n941);
nor (n1571,n1572,n1573);
and (n1572,n947,n154);
and (n1573,n352,n153);
or (n1574,n1543,n942);
nand (n1575,n1576,n1581);
or (n1576,n183,n1577);
not (n1577,n1578);
nand (n1578,n1579,n1580);
or (n1579,n142,n802);
or (n1580,n141,n803);
or (n1581,n188,n1530);
and (n1582,n1568,n1569);
and (n1583,n1558,n1564);
xor (n1584,n1511,n1548);
and (n1585,n1554,n1555);
nor (n1586,n1587,n1627);
not (n1587,n1588);
or (n1588,n1589,n1590);
xor (n1589,n1553,n1584);
or (n1590,n1591,n1626);
and (n1591,n1592,n1625);
xor (n1592,n1593,n1594);
xor (n1593,n1527,n1541);
or (n1594,n1595,n1624);
and (n1595,n1596,n1609);
xor (n1596,n1597,n1603);
nand (n1597,n1598,n1602);
or (n1598,n355,n1599);
nor (n1599,n1600,n1601);
and (n1600,n170,n270);
and (n1601,n171,n269);
or (n1602,n356,n1521);
nand (n1603,n1604,n1608);
or (n1604,n278,n1605);
nor (n1605,n1606,n1607);
and (n1606,n180,n381);
and (n1607,n178,n380);
or (n1608,n1560,n911);
and (n1609,n1610,n1617);
nor (n1610,n1611,n141);
nor (n1611,n1612,n1615);
and (n1612,n1613,n180);
not (n1613,n1614);
and (n1614,n864,n186);
and (n1615,n863,n1616);
not (n1616,n186);
nand (n1617,n1618,n1623);
or (n1618,n941,n1619);
not (n1619,n1620);
nor (n1620,n1621,n1622);
and (n1621,n249,n352);
and (n1622,n248,n947);
or (n1623,n1571,n942);
and (n1624,n1597,n1603);
xor (n1625,n1557,n1565);
and (n1626,n1593,n1594);
nand (n1627,n1628,n1684);
not (n1628,n1629);
nor (n1629,n1630,n1659);
xor (n1630,n1631,n1658);
xor (n1631,n1632,n1657);
or (n1632,n1633,n1656);
and (n1633,n1634,n1650);
xor (n1634,n1635,n1642);
nand (n1635,n1636,n1641);
or (n1636,n1637,n183);
not (n1637,n1638);
nand (n1638,n1639,n1640);
or (n1639,n141,n864);
or (n1640,n142,n863);
nand (n1641,n189,n1578);
nand (n1642,n1643,n1648);
or (n1643,n1644,n355);
not (n1644,n1645);
nand (n1645,n1646,n1647);
or (n1646,n171,n328);
or (n1647,n170,n329);
nand (n1648,n1649,n348);
not (n1649,n1599);
nand (n1650,n1651,n1655);
or (n1651,n278,n1652);
nor (n1652,n1653,n1654);
and (n1653,n180,n770);
and (n1654,n178,n769);
or (n1655,n1605,n911);
and (n1656,n1635,n1642);
xor (n1657,n1567,n1575);
xor (n1658,n1596,n1609);
or (n1659,n1660,n1683);
and (n1660,n1661,n1682);
xor (n1661,n1662,n1663);
xor (n1662,n1610,n1617);
or (n1663,n1664,n1681);
and (n1664,n1665,n1674);
xor (n1665,n1666,n1667);
and (n1666,n189,n864);
nand (n1667,n1668,n1669);
or (n1668,n942,n1619);
or (n1669,n1670,n941);
not (n1670,n1671);
nand (n1671,n1672,n1673);
or (n1672,n270,n947);
nand (n1673,n947,n270);
nand (n1674,n1675,n1680);
or (n1675,n1676,n355);
not (n1676,n1677);
nand (n1677,n1678,n1679);
or (n1678,n171,n380);
or (n1679,n170,n381);
nand (n1680,n348,n1645);
and (n1681,n1666,n1667);
xor (n1682,n1634,n1650);
and (n1683,n1662,n1663);
not (n1684,n1685);
nor (n1685,n1686,n1687);
xor (n1686,n1592,n1625);
or (n1687,n1688,n1689);
and (n1688,n1631,n1658);
and (n1689,n1632,n1657);
or (n1690,n1691,n1829);
and (n1691,n1692,n1719);
xor (n1692,n1693,n1718);
or (n1693,n1694,n1717);
and (n1694,n1695,n1716);
xor (n1695,n1696,n1702);
nand (n1696,n1697,n1701);
or (n1697,n278,n1698);
nor (n1698,n1699,n1700);
and (n1699,n180,n803);
and (n1700,n178,n802);
or (n1701,n1652,n911);
nor (n1702,n1703,n1711);
not (n1703,n1704);
nand (n1704,n1705,n1710);
or (n1705,n941,n1706);
not (n1706,n1707);
nor (n1707,n1708,n1709);
and (n1708,n329,n352);
and (n1709,n328,n947);
nand (n1710,n1671,n943);
nand (n1711,n1712,n178);
nand (n1712,n1713,n1715);
or (n1713,n1714,n171);
and (n1714,n864,n172);
or (n1715,n864,n172);
xor (n1716,n1665,n1674);
and (n1717,n1696,n1702);
xor (n1718,n1661,n1682);
or (n1719,n1720,n1828);
and (n1720,n1721,n1745);
xor (n1721,n1722,n1744);
or (n1722,n1723,n1743);
and (n1723,n1724,n1739);
xor (n1724,n1725,n1732);
nand (n1725,n1726,n1731);
or (n1726,n1727,n355);
not (n1727,n1728);
nor (n1728,n1729,n1730);
and (n1729,n769,n170);
and (n1730,n770,n171);
nand (n1731,n348,n1677);
nand (n1732,n1733,n1738);
or (n1733,n1734,n278);
not (n1734,n1735);
nand (n1735,n1736,n1737);
or (n1736,n180,n864);
or (n1737,n863,n178);
or (n1738,n1698,n911);
nand (n1739,n1740,n1742);
or (n1740,n1741,n1703);
not (n1741,n1711);
or (n1742,n1704,n1711);
and (n1743,n1725,n1732);
xor (n1744,n1695,n1716);
or (n1745,n1746,n1827);
and (n1746,n1747,n1768);
xor (n1747,n1748,n1767);
or (n1748,n1749,n1766);
and (n1749,n1750,n1759);
xor (n1750,n1751,n1752);
and (n1751,n168,n864);
nand (n1752,n1753,n1758);
or (n1753,n1754,n355);
not (n1754,n1755);
nor (n1755,n1756,n1757);
and (n1756,n802,n170);
and (n1757,n803,n171);
nand (n1758,n348,n1728);
nand (n1759,n1760,n1761);
or (n1760,n942,n1706);
or (n1761,n941,n1762);
not (n1762,n1763);
nor (n1763,n1764,n1765);
and (n1764,n380,n947);
and (n1765,n381,n352);
and (n1766,n1751,n1752);
xor (n1767,n1724,n1739);
nand (n1768,n1769,n1826);
or (n1769,n1770,n1786);
nor (n1770,n1771,n1772);
xor (n1771,n1750,n1759);
and (n1772,n1773,n1780);
nand (n1773,n1774,n1775);
nand (n1774,n1763,n943);
nand (n1775,n1776,n1779);
nor (n1776,n1777,n1778);
and (n1777,n769,n947);
and (n1778,n770,n352);
not (n1779,n941);
not (n1780,n1781);
nand (n1781,n1782,n171);
nand (n1782,n1783,n1785);
or (n1783,n1784,n352);
and (n1784,n864,n351);
or (n1785,n864,n351);
nor (n1786,n1787,n1825);
and (n1787,n1788,n1799);
nand (n1788,n1789,n1793);
nor (n1789,n1790,n1792);
and (n1790,n1791,n1780);
not (n1791,n1773);
and (n1792,n1773,n1781);
nor (n1793,n1794,n1795);
and (n1794,n348,n1755);
and (n1795,n354,n1796);
nand (n1796,n1797,n1798);
or (n1797,n170,n864);
or (n1798,n863,n171);
nand (n1799,n1800,n1823);
or (n1800,n1801,n1815);
not (n1801,n1802);
and (n1802,n1803,n1813);
nand (n1803,n1804,n1809);
or (n1804,n942,n1805);
not (n1805,n1806);
nor (n1806,n1807,n1808);
and (n1807,n802,n947);
and (n1808,n803,n352);
nand (n1809,n1810,n1779);
nand (n1810,n1811,n1812);
or (n1811,n947,n864);
or (n1812,n352,n863);
nor (n1813,n1814,n947);
and (n1814,n864,n943);
not (n1815,n1816);
nand (n1816,n1817,n1822);
not (n1817,n1818);
nand (n1818,n1819,n1821);
or (n1819,n942,n1820);
not (n1820,n1776);
nand (n1821,n1806,n1779);
nand (n1822,n348,n864);
nand (n1823,n1824,n1818);
not (n1824,n1822);
nor (n1825,n1789,n1793);
nand (n1826,n1771,n1772);
and (n1827,n1748,n1767);
and (n1828,n1722,n1744);
and (n1829,n1693,n1718);
nand (n1830,n1831,n1408);
or (n1831,n1832,n1834);
not (n1832,n1833);
nand (n1833,n1589,n1590);
not (n1834,n1835);
nand (n1835,n1588,n1836);
nand (n1836,n1837,n1839);
or (n1837,n1685,n1838);
nand (n1838,n1630,n1659);
nand (n1839,n1686,n1687);
nand (n1840,n1410,n1551);
not (n1841,n1842);
nor (n1842,n1843,n1868);
nor (n1843,n1844,n1845);
xor (n1844,n1305,n1358);
or (n1845,n1846,n1867);
and (n1846,n1847,n1850);
xor (n1847,n1848,n1849);
xor (n1848,n1248,n1296);
xor (n1849,n1309,n1312);
or (n1850,n1851,n1866);
and (n1851,n1852,n1855);
xor (n1852,n1853,n1854);
xor (n1853,n1276,n1289);
xor (n1854,n1251,n1266);
or (n1855,n1856,n1865);
and (n1856,n1857,n1862);
xor (n1857,n1858,n1861);
nand (n1858,n1859,n1860);
or (n1859,n278,n1426);
or (n1860,n1279,n911);
and (n1861,n1439,n1431);
or (n1862,n1863,n1864);
and (n1863,n1499,n1506);
and (n1864,n1500,n1503);
and (n1865,n1858,n1861);
and (n1866,n1853,n1854);
and (n1867,n1848,n1849);
nand (n1868,n1869,n1898);
nor (n1869,n1870,n1893);
nor (n1870,n1871,n1884);
xor (n1871,n1872,n1883);
xor (n1872,n1873,n1874);
xor (n1873,n1314,n1334);
or (n1874,n1875,n1882);
and (n1875,n1876,n1879);
xor (n1876,n1877,n1878);
xor (n1877,n1336,n1349);
xor (n1878,n1318,n1327);
or (n1879,n1880,n1881);
and (n1880,n1413,n1429);
and (n1881,n1414,n1420);
and (n1882,n1877,n1878);
xor (n1883,n1852,n1855);
or (n1884,n1885,n1892);
and (n1885,n1886,n1891);
xor (n1886,n1887,n1888);
xor (n1887,n1857,n1862);
or (n1888,n1889,n1890);
and (n1889,n1448,n1498);
and (n1890,n1449,n1470);
xor (n1891,n1876,n1879);
and (n1892,n1887,n1888);
nor (n1893,n1894,n1897);
or (n1894,n1895,n1896);
and (n1895,n1411,n1509);
and (n1896,n1412,n1447);
xor (n1897,n1886,n1891);
nand (n1898,n1899,n1901);
not (n1899,n1900);
xor (n1900,n1847,n1850);
not (n1901,n1902);
or (n1902,n1903,n1904);
and (n1903,n1872,n1883);
and (n1904,n1873,n1874);
nor (n1905,n1906,n1917);
and (n1906,n1907,n1908);
not (n1907,n1843);
nand (n1908,n1909,n1916);
or (n1909,n1910,n1911);
not (n1910,n1898);
not (n1911,n1912);
nand (n1912,n1913,n1915);
or (n1913,n1870,n1914);
nand (n1914,n1894,n1897);
nand (n1915,n1871,n1884);
nand (n1916,n1900,n1902);
and (n1917,n1844,n1845);
nor (n1918,n1919,n1935);
and (n1919,n1920,n1934);
nand (n1920,n1921,n1933);
or (n1921,n1922,n1923);
not (n1922,n579);
not (n1923,n1924);
nand (n1924,n1925,n1932);
or (n1925,n1926,n1927);
not (n1926,n535);
not (n1927,n1928);
nand (n1928,n1929,n1931);
or (n1929,n1930,n484);
nand (n1930,n101,n431);
nand (n1931,n485,n532);
nand (n1932,n576,n536);
nand (n1933,n580,n583);
not (n1934,n617);
nand (n1935,n1936,n1944);
or (n1936,n1937,n619);
and (n1937,n1938,n1943);
nand (n1938,n1939,n689);
nand (n1939,n1940,n1942);
or (n1940,n1941,n676);
nand (n1941,n649,n652);
nand (n1942,n677,n680);
nand (n1943,n690,n693);
nand (n1944,n620,n646);
nand (n1945,n52,n91);
and (n1946,n1947,n1948);
not (n1947,n2);
not (n1948,n48);
or (n1949,n1950,n3376);
and (n1950,n1951,n3375);
or (n1951,n1952,n3286);
and (n1952,n1953,n3285);
or (n1953,n1954,n3190);
and (n1954,n1955,n3189);
or (n1955,n1956,n3094);
and (n1956,n1957,n3093);
or (n1957,n1958,n2998);
and (n1958,n1959,n2997);
or (n1959,n1960,n2905);
and (n1960,n1961,n2904);
or (n1961,n1962,n2810);
and (n1962,n1963,n2809);
or (n1963,n1964,n2719);
and (n1964,n1965,n2718);
or (n1965,n1966,n2624);
and (n1966,n1967,n2623);
or (n1967,n1968,n2536);
and (n1968,n1969,n2535);
or (n1969,n1970,n2441);
and (n1970,n1971,n2440);
or (n1971,n1972,n2347);
and (n1972,n1973,n276);
or (n1973,n1974,n2253);
and (n1974,n1975,n2252);
or (n1975,n1976,n2162);
and (n1976,n1977,n425);
or (n1977,n1978,n2068);
and (n1978,n1979,n2067);
and (n1979,n948,n1980);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
and (n1982,n38,n943);
and (n1983,n34,n352);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
and (n1988,n34,n943);
and (n1989,n42,n352);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1995);
and (n1993,n1994,n1103);
and (n1994,n42,n943);
and (n1995,n1996,n1997);
xor (n1996,n1994,n1103);
or (n1997,n1998,n2001);
and (n1998,n1999,n2000);
and (n1999,n86,n943);
and (n2000,n220,n352);
and (n2001,n2002,n2003);
xor (n2002,n1999,n2000);
or (n2003,n2004,n2007);
and (n2004,n2005,n2006);
and (n2005,n220,n943);
and (n2006,n215,n352);
and (n2007,n2008,n2009);
xor (n2008,n2005,n2006);
or (n2009,n2010,n2013);
and (n2010,n2011,n2012);
and (n2011,n215,n943);
and (n2012,n121,n352);
and (n2013,n2014,n2015);
xor (n2014,n2011,n2012);
or (n2015,n2016,n2019);
and (n2016,n2017,n2018);
and (n2017,n121,n943);
and (n2018,n115,n352);
and (n2019,n2020,n2021);
xor (n2020,n2017,n2018);
or (n2021,n2022,n2025);
and (n2022,n2023,n2024);
and (n2023,n115,n943);
and (n2024,n160,n352);
and (n2025,n2026,n2027);
xor (n2026,n2023,n2024);
or (n2027,n2028,n2031);
and (n2028,n2029,n2030);
and (n2029,n160,n943);
and (n2030,n154,n352);
and (n2031,n2032,n2033);
xor (n2032,n2029,n2030);
or (n2033,n2034,n2036);
and (n2034,n2035,n1621);
and (n2035,n154,n943);
and (n2036,n2037,n2038);
xor (n2037,n2035,n1621);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
and (n2040,n249,n943);
and (n2041,n270,n352);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
or (n2044,n2045,n2047);
and (n2045,n2046,n1708);
and (n2046,n270,n943);
and (n2047,n2048,n2049);
xor (n2048,n2046,n1708);
or (n2049,n2050,n2052);
and (n2050,n2051,n1765);
and (n2051,n329,n943);
and (n2052,n2053,n2054);
xor (n2053,n2051,n1765);
or (n2054,n2055,n2057);
and (n2055,n2056,n1778);
and (n2056,n381,n943);
and (n2057,n2058,n2059);
xor (n2058,n2056,n1778);
or (n2059,n2060,n2062);
and (n2060,n2061,n1808);
and (n2061,n770,n943);
and (n2062,n2063,n2064);
xor (n2063,n2061,n1808);
and (n2064,n2065,n2066);
and (n2065,n803,n943);
and (n2066,n864,n352);
and (n2067,n38,n351);
and (n2068,n2069,n2070);
xor (n2069,n1979,n2067);
or (n2070,n2071,n2074);
and (n2071,n2072,n2073);
xor (n2072,n948,n1980);
and (n2073,n34,n351);
and (n2074,n2075,n2076);
xor (n2075,n2072,n2073);
or (n2076,n2077,n2080);
and (n2077,n2078,n2079);
xor (n2078,n1985,n1986);
and (n2079,n42,n351);
and (n2080,n2081,n2082);
xor (n2081,n2078,n2079);
or (n2082,n2083,n2086);
and (n2083,n2084,n2085);
xor (n2084,n1991,n1992);
and (n2085,n86,n351);
and (n2086,n2087,n2088);
xor (n2087,n2084,n2085);
or (n2088,n2089,n2092);
and (n2089,n2090,n2091);
xor (n2090,n1996,n1997);
and (n2091,n220,n351);
and (n2092,n2093,n2094);
xor (n2093,n2090,n2091);
or (n2094,n2095,n2098);
and (n2095,n2096,n2097);
xor (n2096,n2002,n2003);
and (n2097,n215,n351);
and (n2098,n2099,n2100);
xor (n2099,n2096,n2097);
or (n2100,n2101,n2104);
and (n2101,n2102,n2103);
xor (n2102,n2008,n2009);
and (n2103,n121,n351);
and (n2104,n2105,n2106);
xor (n2105,n2102,n2103);
or (n2106,n2107,n2110);
and (n2107,n2108,n2109);
xor (n2108,n2014,n2015);
and (n2109,n115,n351);
and (n2110,n2111,n2112);
xor (n2111,n2108,n2109);
or (n2112,n2113,n2116);
and (n2113,n2114,n2115);
xor (n2114,n2020,n2021);
and (n2115,n160,n351);
and (n2116,n2117,n2118);
xor (n2117,n2114,n2115);
or (n2118,n2119,n2122);
and (n2119,n2120,n2121);
xor (n2120,n2026,n2027);
and (n2121,n154,n351);
and (n2122,n2123,n2124);
xor (n2123,n2120,n2121);
or (n2124,n2125,n2128);
and (n2125,n2126,n2127);
xor (n2126,n2032,n2033);
and (n2127,n249,n351);
and (n2128,n2129,n2130);
xor (n2129,n2126,n2127);
or (n2130,n2131,n2134);
and (n2131,n2132,n2133);
xor (n2132,n2037,n2038);
and (n2133,n270,n351);
and (n2134,n2135,n2136);
xor (n2135,n2132,n2133);
or (n2136,n2137,n2140);
and (n2137,n2138,n2139);
xor (n2138,n2043,n2044);
and (n2139,n329,n351);
and (n2140,n2141,n2142);
xor (n2141,n2138,n2139);
or (n2142,n2143,n2146);
and (n2143,n2144,n2145);
xor (n2144,n2048,n2049);
and (n2145,n381,n351);
and (n2146,n2147,n2148);
xor (n2147,n2144,n2145);
or (n2148,n2149,n2152);
and (n2149,n2150,n2151);
xor (n2150,n2053,n2054);
and (n2151,n770,n351);
and (n2152,n2153,n2154);
xor (n2153,n2150,n2151);
or (n2154,n2155,n2158);
and (n2155,n2156,n2157);
xor (n2156,n2058,n2059);
and (n2157,n803,n351);
and (n2158,n2159,n2160);
xor (n2159,n2156,n2157);
and (n2160,n2161,n1784);
xor (n2161,n2063,n2064);
and (n2162,n2163,n2164);
xor (n2163,n1977,n425);
or (n2164,n2165,n2168);
and (n2165,n2166,n2167);
xor (n2166,n2069,n2070);
and (n2167,n34,n171);
and (n2168,n2169,n2170);
xor (n2169,n2166,n2167);
or (n2170,n2171,n2173);
and (n2171,n2172,n895);
xor (n2172,n2075,n2076);
and (n2173,n2174,n2175);
xor (n2174,n2172,n895);
or (n2175,n2176,n2178);
and (n2176,n2177,n982);
xor (n2177,n2081,n2082);
and (n2178,n2179,n2180);
xor (n2179,n2177,n982);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2087,n2088);
and (n2183,n220,n171);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2093,n2094);
and (n2189,n215,n171);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2195);
and (n2193,n2194,n1257);
xor (n2194,n2099,n2100);
and (n2195,n2196,n2197);
xor (n2196,n2194,n1257);
or (n2197,n2198,n2201);
and (n2198,n2199,n2200);
xor (n2199,n2105,n2106);
and (n2200,n115,n171);
and (n2201,n2202,n2203);
xor (n2202,n2199,n2200);
or (n2203,n2204,n2207);
and (n2204,n2205,n2206);
xor (n2205,n2111,n2112);
and (n2206,n160,n171);
and (n2207,n2208,n2209);
xor (n2208,n2205,n2206);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2117,n2118);
and (n2212,n154,n171);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
or (n2215,n2216,n2219);
and (n2216,n2217,n2218);
xor (n2217,n2123,n2124);
and (n2218,n249,n171);
and (n2219,n2220,n2221);
xor (n2220,n2217,n2218);
or (n2221,n2222,n2225);
and (n2222,n2223,n2224);
xor (n2223,n2129,n2130);
and (n2224,n270,n171);
and (n2225,n2226,n2227);
xor (n2226,n2223,n2224);
or (n2227,n2228,n2231);
and (n2228,n2229,n2230);
xor (n2229,n2135,n2136);
and (n2230,n329,n171);
and (n2231,n2232,n2233);
xor (n2232,n2229,n2230);
or (n2233,n2234,n2237);
and (n2234,n2235,n2236);
xor (n2235,n2141,n2142);
and (n2236,n381,n171);
and (n2237,n2238,n2239);
xor (n2238,n2235,n2236);
or (n2239,n2240,n2242);
and (n2240,n2241,n1730);
xor (n2241,n2147,n2148);
and (n2242,n2243,n2244);
xor (n2243,n2241,n1730);
or (n2244,n2245,n2247);
and (n2245,n2246,n1757);
xor (n2246,n2153,n2154);
and (n2247,n2248,n2249);
xor (n2248,n2246,n1757);
and (n2249,n2250,n2251);
xor (n2250,n2159,n2160);
and (n2251,n864,n171);
and (n2252,n38,n172);
and (n2253,n2254,n2255);
xor (n2254,n1975,n2252);
or (n2255,n2256,n2259);
and (n2256,n2257,n2258);
xor (n2257,n2163,n2164);
and (n2258,n34,n172);
and (n2259,n2260,n2261);
xor (n2260,n2257,n2258);
or (n2261,n2262,n2265);
and (n2262,n2263,n2264);
xor (n2263,n2169,n2170);
and (n2264,n42,n172);
and (n2265,n2266,n2267);
xor (n2266,n2263,n2264);
or (n2267,n2268,n2271);
and (n2268,n2269,n2270);
xor (n2269,n2174,n2175);
and (n2270,n86,n172);
and (n2271,n2272,n2273);
xor (n2272,n2269,n2270);
or (n2273,n2274,n2277);
and (n2274,n2275,n2276);
xor (n2275,n2179,n2180);
and (n2276,n220,n172);
and (n2277,n2278,n2279);
xor (n2278,n2275,n2276);
or (n2279,n2280,n2283);
and (n2280,n2281,n2282);
xor (n2281,n2185,n2186);
and (n2282,n215,n172);
and (n2283,n2284,n2285);
xor (n2284,n2281,n2282);
or (n2285,n2286,n2289);
and (n2286,n2287,n2288);
xor (n2287,n2191,n2192);
and (n2288,n121,n172);
and (n2289,n2290,n2291);
xor (n2290,n2287,n2288);
or (n2291,n2292,n2295);
and (n2292,n2293,n2294);
xor (n2293,n2196,n2197);
and (n2294,n115,n172);
and (n2295,n2296,n2297);
xor (n2296,n2293,n2294);
or (n2297,n2298,n2301);
and (n2298,n2299,n2300);
xor (n2299,n2202,n2203);
and (n2300,n160,n172);
and (n2301,n2302,n2303);
xor (n2302,n2299,n2300);
or (n2303,n2304,n2307);
and (n2304,n2305,n2306);
xor (n2305,n2208,n2209);
and (n2306,n154,n172);
and (n2307,n2308,n2309);
xor (n2308,n2305,n2306);
or (n2309,n2310,n2313);
and (n2310,n2311,n2312);
xor (n2311,n2214,n2215);
and (n2312,n249,n172);
and (n2313,n2314,n2315);
xor (n2314,n2311,n2312);
or (n2315,n2316,n2319);
and (n2316,n2317,n2318);
xor (n2317,n2220,n2221);
and (n2318,n270,n172);
and (n2319,n2320,n2321);
xor (n2320,n2317,n2318);
or (n2321,n2322,n2325);
and (n2322,n2323,n2324);
xor (n2323,n2226,n2227);
and (n2324,n329,n172);
and (n2325,n2326,n2327);
xor (n2326,n2323,n2324);
or (n2327,n2328,n2331);
and (n2328,n2329,n2330);
xor (n2329,n2232,n2233);
and (n2330,n381,n172);
and (n2331,n2332,n2333);
xor (n2332,n2329,n2330);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2238,n2239);
and (n2336,n770,n172);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
or (n2339,n2340,n2343);
and (n2340,n2341,n2342);
xor (n2341,n2243,n2244);
and (n2342,n803,n172);
and (n2343,n2344,n2345);
xor (n2344,n2341,n2342);
and (n2345,n2346,n1714);
xor (n2346,n2248,n2249);
and (n2347,n2348,n2349);
xor (n2348,n1973,n276);
or (n2349,n2350,n2353);
and (n2350,n2351,n2352);
xor (n2351,n2254,n2255);
and (n2352,n34,n178);
and (n2353,n2354,n2355);
xor (n2354,n2351,n2352);
or (n2355,n2356,n2358);
and (n2356,n2357,n765);
xor (n2357,n2260,n2261);
and (n2358,n2359,n2360);
xor (n2359,n2357,n765);
or (n2360,n2361,n2364);
and (n2361,n2362,n2363);
xor (n2362,n2266,n2267);
and (n2363,n86,n178);
and (n2364,n2365,n2366);
xor (n2365,n2362,n2363);
or (n2366,n2367,n2369);
and (n2367,n2368,n909);
xor (n2368,n2272,n2273);
and (n2369,n2370,n2371);
xor (n2370,n2368,n909);
or (n2371,n2372,n2375);
and (n2372,n2373,n2374);
xor (n2373,n2278,n2279);
and (n2374,n215,n178);
and (n2375,n2376,n2377);
xor (n2376,n2373,n2374);
or (n2377,n2378,n2381);
and (n2378,n2379,n2380);
xor (n2379,n2284,n2285);
and (n2380,n121,n178);
and (n2381,n2382,n2383);
xor (n2382,n2379,n2380);
or (n2383,n2384,n2387);
and (n2384,n2385,n2386);
xor (n2385,n2290,n2291);
and (n2386,n115,n178);
and (n2387,n2388,n2389);
xor (n2388,n2385,n2386);
or (n2389,n2390,n2393);
and (n2390,n2391,n2392);
xor (n2391,n2296,n2297);
and (n2392,n160,n178);
and (n2393,n2394,n2395);
xor (n2394,n2391,n2392);
or (n2395,n2396,n2399);
and (n2396,n2397,n2398);
xor (n2397,n2302,n2303);
and (n2398,n154,n178);
and (n2399,n2400,n2401);
xor (n2400,n2397,n2398);
or (n2401,n2402,n2405);
and (n2402,n2403,n2404);
xor (n2403,n2308,n2309);
and (n2404,n249,n178);
and (n2405,n2406,n2407);
xor (n2406,n2403,n2404);
or (n2407,n2408,n2411);
and (n2408,n2409,n2410);
xor (n2409,n2314,n2315);
and (n2410,n270,n178);
and (n2411,n2412,n2413);
xor (n2412,n2409,n2410);
or (n2413,n2414,n2417);
and (n2414,n2415,n2416);
xor (n2415,n2320,n2321);
and (n2416,n329,n178);
and (n2417,n2418,n2419);
xor (n2418,n2415,n2416);
or (n2419,n2420,n2423);
and (n2420,n2421,n2422);
xor (n2421,n2326,n2327);
and (n2422,n381,n178);
and (n2423,n2424,n2425);
xor (n2424,n2421,n2422);
or (n2425,n2426,n2429);
and (n2426,n2427,n2428);
xor (n2427,n2332,n2333);
and (n2428,n770,n178);
and (n2429,n2430,n2431);
xor (n2430,n2427,n2428);
or (n2431,n2432,n2435);
and (n2432,n2433,n2434);
xor (n2433,n2338,n2339);
and (n2434,n803,n178);
and (n2435,n2436,n2437);
xor (n2436,n2433,n2434);
and (n2437,n2438,n2439);
xor (n2438,n2344,n2345);
and (n2439,n864,n178);
and (n2440,n38,n186);
and (n2441,n2442,n2443);
xor (n2442,n1971,n2440);
or (n2443,n2444,n2447);
and (n2444,n2445,n2446);
xor (n2445,n2348,n2349);
and (n2446,n34,n186);
and (n2447,n2448,n2449);
xor (n2448,n2445,n2446);
or (n2449,n2450,n2453);
and (n2450,n2451,n2452);
xor (n2451,n2354,n2355);
and (n2452,n42,n186);
and (n2453,n2454,n2455);
xor (n2454,n2451,n2452);
or (n2455,n2456,n2459);
and (n2456,n2457,n2458);
xor (n2457,n2359,n2360);
and (n2458,n86,n186);
and (n2459,n2460,n2461);
xor (n2460,n2457,n2458);
or (n2461,n2462,n2465);
and (n2462,n2463,n2464);
xor (n2463,n2365,n2366);
and (n2464,n220,n186);
and (n2465,n2466,n2467);
xor (n2466,n2463,n2464);
or (n2467,n2468,n2471);
and (n2468,n2469,n2470);
xor (n2469,n2370,n2371);
and (n2470,n215,n186);
and (n2471,n2472,n2473);
xor (n2472,n2469,n2470);
or (n2473,n2474,n2477);
and (n2474,n2475,n2476);
xor (n2475,n2376,n2377);
and (n2476,n121,n186);
and (n2477,n2478,n2479);
xor (n2478,n2475,n2476);
or (n2479,n2480,n2483);
and (n2480,n2481,n2482);
xor (n2481,n2382,n2383);
and (n2482,n115,n186);
and (n2483,n2484,n2485);
xor (n2484,n2481,n2482);
or (n2485,n2486,n2489);
and (n2486,n2487,n2488);
xor (n2487,n2388,n2389);
and (n2488,n160,n186);
and (n2489,n2490,n2491);
xor (n2490,n2487,n2488);
or (n2491,n2492,n2495);
and (n2492,n2493,n2494);
xor (n2493,n2394,n2395);
and (n2494,n154,n186);
and (n2495,n2496,n2497);
xor (n2496,n2493,n2494);
or (n2497,n2498,n2501);
and (n2498,n2499,n2500);
xor (n2499,n2400,n2401);
and (n2500,n249,n186);
and (n2501,n2502,n2503);
xor (n2502,n2499,n2500);
or (n2503,n2504,n2507);
and (n2504,n2505,n2506);
xor (n2505,n2406,n2407);
and (n2506,n270,n186);
and (n2507,n2508,n2509);
xor (n2508,n2505,n2506);
or (n2509,n2510,n2513);
and (n2510,n2511,n2512);
xor (n2511,n2412,n2413);
and (n2512,n329,n186);
and (n2513,n2514,n2515);
xor (n2514,n2511,n2512);
or (n2515,n2516,n2519);
and (n2516,n2517,n2518);
xor (n2517,n2418,n2419);
and (n2518,n381,n186);
and (n2519,n2520,n2521);
xor (n2520,n2517,n2518);
or (n2521,n2522,n2525);
and (n2522,n2523,n2524);
xor (n2523,n2424,n2425);
and (n2524,n770,n186);
and (n2525,n2526,n2527);
xor (n2526,n2523,n2524);
or (n2527,n2528,n2531);
and (n2528,n2529,n2530);
xor (n2529,n2430,n2431);
and (n2530,n803,n186);
and (n2531,n2532,n2533);
xor (n2532,n2529,n2530);
and (n2533,n2534,n1614);
xor (n2534,n2436,n2437);
and (n2535,n38,n142);
and (n2536,n2537,n2538);
xor (n2537,n1969,n2535);
or (n2538,n2539,n2541);
and (n2539,n2540,n195);
xor (n2540,n2442,n2443);
and (n2541,n2542,n2543);
xor (n2542,n2540,n195);
or (n2543,n2544,n2546);
and (n2544,n2545,n287);
xor (n2545,n2448,n2449);
and (n2546,n2547,n2548);
xor (n2547,n2545,n287);
or (n2548,n2549,n2551);
and (n2549,n2550,n395);
xor (n2550,n2454,n2455);
and (n2551,n2552,n2553);
xor (n2552,n2550,n395);
or (n2553,n2554,n2556);
and (n2554,n2555,n727);
xor (n2555,n2460,n2461);
and (n2556,n2557,n2558);
xor (n2557,n2555,n727);
or (n2558,n2559,n2561);
and (n2559,n2560,n723);
xor (n2560,n2466,n2467);
and (n2561,n2562,n2563);
xor (n2562,n2560,n723);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2472,n2473);
and (n2566,n121,n142);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2478,n2479);
and (n2572,n115,n142);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
or (n2575,n2576,n2578);
and (n2576,n2577,n1140);
xor (n2577,n2484,n2485);
and (n2578,n2579,n2580);
xor (n2579,n2577,n1140);
or (n2580,n2581,n2584);
and (n2581,n2582,n2583);
xor (n2582,n2490,n2491);
and (n2583,n154,n142);
and (n2584,n2585,n2586);
xor (n2585,n2582,n2583);
or (n2586,n2587,n2590);
and (n2587,n2588,n2589);
xor (n2588,n2496,n2497);
and (n2589,n249,n142);
and (n2590,n2591,n2592);
xor (n2591,n2588,n2589);
or (n2592,n2593,n2596);
and (n2593,n2594,n2595);
xor (n2594,n2502,n2503);
and (n2595,n270,n142);
and (n2596,n2597,n2598);
xor (n2597,n2594,n2595);
or (n2598,n2599,n2602);
and (n2599,n2600,n2601);
xor (n2600,n2508,n2509);
and (n2601,n329,n142);
and (n2602,n2603,n2604);
xor (n2603,n2600,n2601);
or (n2604,n2605,n2607);
and (n2605,n2606,n1464);
xor (n2606,n2514,n2515);
and (n2607,n2608,n2609);
xor (n2608,n2606,n1464);
or (n2609,n2610,n2612);
and (n2610,n2611,n1532);
xor (n2611,n2520,n2521);
and (n2612,n2613,n2614);
xor (n2613,n2611,n1532);
or (n2614,n2615,n2618);
and (n2615,n2616,n2617);
xor (n2616,n2526,n2527);
and (n2617,n803,n142);
and (n2618,n2619,n2620);
xor (n2619,n2616,n2617);
and (n2620,n2621,n2622);
xor (n2621,n2532,n2533);
and (n2622,n864,n142);
and (n2623,n38,n136);
and (n2624,n2625,n2626);
xor (n2625,n1967,n2623);
or (n2626,n2627,n2630);
and (n2627,n2628,n2629);
xor (n2628,n2537,n2538);
and (n2629,n34,n136);
and (n2630,n2631,n2632);
xor (n2631,n2628,n2629);
or (n2632,n2633,n2636);
and (n2633,n2634,n2635);
xor (n2634,n2542,n2543);
and (n2635,n42,n136);
and (n2636,n2637,n2638);
xor (n2637,n2634,n2635);
or (n2638,n2639,n2642);
and (n2639,n2640,n2641);
xor (n2640,n2547,n2548);
and (n2641,n86,n136);
and (n2642,n2643,n2644);
xor (n2643,n2640,n2641);
or (n2644,n2645,n2648);
and (n2645,n2646,n2647);
xor (n2646,n2552,n2553);
and (n2647,n220,n136);
and (n2648,n2649,n2650);
xor (n2649,n2646,n2647);
or (n2650,n2651,n2654);
and (n2651,n2652,n2653);
xor (n2652,n2557,n2558);
and (n2653,n215,n136);
and (n2654,n2655,n2656);
xor (n2655,n2652,n2653);
or (n2656,n2657,n2660);
and (n2657,n2658,n2659);
xor (n2658,n2562,n2563);
and (n2659,n121,n136);
and (n2660,n2661,n2662);
xor (n2661,n2658,n2659);
or (n2662,n2663,n2666);
and (n2663,n2664,n2665);
xor (n2664,n2568,n2569);
and (n2665,n115,n136);
and (n2666,n2667,n2668);
xor (n2667,n2664,n2665);
or (n2668,n2669,n2672);
and (n2669,n2670,n2671);
xor (n2670,n2574,n2575);
and (n2671,n160,n136);
and (n2672,n2673,n2674);
xor (n2673,n2670,n2671);
or (n2674,n2675,n2678);
and (n2675,n2676,n2677);
xor (n2676,n2579,n2580);
and (n2677,n154,n136);
and (n2678,n2679,n2680);
xor (n2679,n2676,n2677);
or (n2680,n2681,n2684);
and (n2681,n2682,n2683);
xor (n2682,n2585,n2586);
and (n2683,n249,n136);
and (n2684,n2685,n2686);
xor (n2685,n2682,n2683);
or (n2686,n2687,n2690);
and (n2687,n2688,n2689);
xor (n2688,n2591,n2592);
and (n2689,n270,n136);
and (n2690,n2691,n2692);
xor (n2691,n2688,n2689);
or (n2692,n2693,n2696);
and (n2693,n2694,n2695);
xor (n2694,n2597,n2598);
and (n2695,n329,n136);
and (n2696,n2697,n2698);
xor (n2697,n2694,n2695);
or (n2698,n2699,n2702);
and (n2699,n2700,n2701);
xor (n2700,n2603,n2604);
and (n2701,n381,n136);
and (n2702,n2703,n2704);
xor (n2703,n2700,n2701);
or (n2704,n2705,n2708);
and (n2705,n2706,n2707);
xor (n2706,n2608,n2609);
and (n2707,n770,n136);
and (n2708,n2709,n2710);
xor (n2709,n2706,n2707);
or (n2710,n2711,n2714);
and (n2711,n2712,n2713);
xor (n2712,n2613,n2614);
and (n2713,n803,n136);
and (n2714,n2715,n2716);
xor (n2715,n2712,n2713);
and (n2716,n2717,n1518);
xor (n2717,n2619,n2620);
and (n2718,n38,n130);
and (n2719,n2720,n2721);
xor (n2720,n1965,n2718);
or (n2721,n2722,n2725);
and (n2722,n2723,n2724);
xor (n2723,n2625,n2626);
and (n2724,n34,n130);
and (n2725,n2726,n2727);
xor (n2726,n2723,n2724);
or (n2727,n2728,n2731);
and (n2728,n2729,n2730);
xor (n2729,n2631,n2632);
and (n2730,n42,n130);
and (n2731,n2732,n2733);
xor (n2732,n2729,n2730);
or (n2733,n2734,n2736);
and (n2734,n2735,n131);
xor (n2735,n2637,n2638);
and (n2736,n2737,n2738);
xor (n2737,n2735,n131);
or (n2738,n2739,n2741);
and (n2739,n2740,n317);
xor (n2740,n2643,n2644);
and (n2741,n2742,n2743);
xor (n2742,n2740,n317);
or (n2743,n2744,n2747);
and (n2744,n2745,n2746);
xor (n2745,n2649,n2650);
and (n2746,n215,n130);
and (n2747,n2748,n2749);
xor (n2748,n2745,n2746);
or (n2749,n2750,n2752);
and (n2750,n2751,n777);
xor (n2751,n2655,n2656);
and (n2752,n2753,n2754);
xor (n2753,n2751,n777);
or (n2754,n2755,n2757);
and (n2755,n2756,n822);
xor (n2756,n2661,n2662);
and (n2757,n2758,n2759);
xor (n2758,n2756,n822);
or (n2759,n2760,n2763);
and (n2760,n2761,n2762);
xor (n2761,n2667,n2668);
and (n2762,n160,n130);
and (n2763,n2764,n2765);
xor (n2764,n2761,n2762);
or (n2765,n2766,n2769);
and (n2766,n2767,n2768);
xor (n2767,n2673,n2674);
and (n2768,n154,n130);
and (n2769,n2770,n2771);
xor (n2770,n2767,n2768);
or (n2771,n2772,n2774);
and (n2772,n2773,n1151);
xor (n2773,n2679,n2680);
and (n2774,n2775,n2776);
xor (n2775,n2773,n1151);
or (n2776,n2777,n2780);
and (n2777,n2778,n2779);
xor (n2778,n2685,n2686);
and (n2779,n270,n130);
and (n2780,n2781,n2782);
xor (n2781,n2778,n2779);
or (n2782,n2783,n2786);
and (n2783,n2784,n2785);
xor (n2784,n2691,n2692);
and (n2785,n329,n130);
and (n2786,n2787,n2788);
xor (n2787,n2784,n2785);
or (n2788,n2789,n2792);
and (n2789,n2790,n2791);
xor (n2790,n2697,n2698);
and (n2791,n381,n130);
and (n2792,n2793,n2794);
xor (n2793,n2790,n2791);
or (n2794,n2795,n2798);
and (n2795,n2796,n2797);
xor (n2796,n2703,n2704);
and (n2797,n770,n130);
and (n2798,n2799,n2800);
xor (n2799,n2796,n2797);
or (n2800,n2801,n2804);
and (n2801,n2802,n2803);
xor (n2802,n2709,n2710);
and (n2803,n803,n130);
and (n2804,n2805,n2806);
xor (n2805,n2802,n2803);
and (n2806,n2807,n2808);
xor (n2807,n2715,n2716);
and (n2808,n864,n130);
and (n2809,n38,n207);
and (n2810,n2811,n2812);
xor (n2811,n1963,n2809);
or (n2812,n2813,n2816);
and (n2813,n2814,n2815);
xor (n2814,n2720,n2721);
and (n2815,n34,n207);
and (n2816,n2817,n2818);
xor (n2817,n2814,n2815);
or (n2818,n2819,n2822);
and (n2819,n2820,n2821);
xor (n2820,n2726,n2727);
and (n2821,n42,n207);
and (n2822,n2823,n2824);
xor (n2823,n2820,n2821);
or (n2824,n2825,n2828);
and (n2825,n2826,n2827);
xor (n2826,n2732,n2733);
and (n2827,n86,n207);
and (n2828,n2829,n2830);
xor (n2829,n2826,n2827);
or (n2830,n2831,n2834);
and (n2831,n2832,n2833);
xor (n2832,n2737,n2738);
and (n2833,n220,n207);
and (n2834,n2835,n2836);
xor (n2835,n2832,n2833);
or (n2836,n2837,n2840);
and (n2837,n2838,n2839);
xor (n2838,n2742,n2743);
and (n2839,n215,n207);
and (n2840,n2841,n2842);
xor (n2841,n2838,n2839);
or (n2842,n2843,n2846);
and (n2843,n2844,n2845);
xor (n2844,n2748,n2749);
and (n2845,n121,n207);
and (n2846,n2847,n2848);
xor (n2847,n2844,n2845);
or (n2848,n2849,n2852);
and (n2849,n2850,n2851);
xor (n2850,n2753,n2754);
and (n2851,n115,n207);
and (n2852,n2853,n2854);
xor (n2853,n2850,n2851);
or (n2854,n2855,n2858);
and (n2855,n2856,n2857);
xor (n2856,n2758,n2759);
and (n2857,n160,n207);
and (n2858,n2859,n2860);
xor (n2859,n2856,n2857);
or (n2860,n2861,n2864);
and (n2861,n2862,n2863);
xor (n2862,n2764,n2765);
and (n2863,n154,n207);
and (n2864,n2865,n2866);
xor (n2865,n2862,n2863);
or (n2866,n2867,n2870);
and (n2867,n2868,n2869);
xor (n2868,n2770,n2771);
and (n2869,n249,n207);
and (n2870,n2871,n2872);
xor (n2871,n2868,n2869);
or (n2872,n2873,n2876);
and (n2873,n2874,n2875);
xor (n2874,n2775,n2776);
and (n2875,n270,n207);
and (n2876,n2877,n2878);
xor (n2877,n2874,n2875);
or (n2878,n2879,n2882);
and (n2879,n2880,n2881);
xor (n2880,n2781,n2782);
and (n2881,n329,n207);
and (n2882,n2883,n2884);
xor (n2883,n2880,n2881);
or (n2884,n2885,n2888);
and (n2885,n2886,n2887);
xor (n2886,n2787,n2788);
and (n2887,n381,n207);
and (n2888,n2889,n2890);
xor (n2889,n2886,n2887);
or (n2890,n2891,n2894);
and (n2891,n2892,n2893);
xor (n2892,n2793,n2794);
and (n2893,n770,n207);
and (n2894,n2895,n2896);
xor (n2895,n2892,n2893);
or (n2896,n2897,n2900);
and (n2897,n2898,n2899);
xor (n2898,n2799,n2800);
and (n2899,n803,n207);
and (n2900,n2901,n2902);
xor (n2901,n2898,n2899);
and (n2902,n2903,n1437);
xor (n2903,n2805,n2806);
and (n2904,n38,n72);
and (n2905,n2906,n2907);
xor (n2906,n1961,n2904);
or (n2907,n2908,n2911);
and (n2908,n2909,n2910);
xor (n2909,n2811,n2812);
and (n2910,n34,n72);
and (n2911,n2912,n2913);
xor (n2912,n2909,n2910);
or (n2913,n2914,n2917);
and (n2914,n2915,n2916);
xor (n2915,n2817,n2818);
and (n2916,n42,n72);
and (n2917,n2918,n2919);
xor (n2918,n2915,n2916);
or (n2919,n2920,n2923);
and (n2920,n2921,n2922);
xor (n2921,n2823,n2824);
and (n2922,n86,n72);
and (n2923,n2924,n2925);
xor (n2924,n2921,n2922);
or (n2925,n2926,n2929);
and (n2926,n2927,n2928);
xor (n2927,n2829,n2830);
and (n2928,n220,n72);
and (n2929,n2930,n2931);
xor (n2930,n2927,n2928);
or (n2931,n2932,n2935);
and (n2932,n2933,n2934);
xor (n2933,n2835,n2836);
and (n2934,n215,n72);
and (n2935,n2936,n2937);
xor (n2936,n2933,n2934);
or (n2937,n2938,n2940);
and (n2938,n2939,n295);
xor (n2939,n2841,n2842);
and (n2940,n2941,n2942);
xor (n2941,n2939,n295);
or (n2942,n2943,n2945);
and (n2943,n2944,n388);
xor (n2944,n2847,n2848);
and (n2945,n2946,n2947);
xor (n2946,n2944,n388);
or (n2947,n2948,n2951);
and (n2948,n2949,n2950);
xor (n2949,n2853,n2854);
and (n2950,n160,n72);
and (n2951,n2952,n2953);
xor (n2952,n2949,n2950);
or (n2953,n2954,n2957);
and (n2954,n2955,n2956);
xor (n2955,n2859,n2860);
and (n2956,n154,n72);
and (n2957,n2958,n2959);
xor (n2958,n2955,n2956);
or (n2959,n2960,n2962);
and (n2960,n2961,n929);
xor (n2961,n2865,n2866);
and (n2962,n2963,n2964);
xor (n2963,n2961,n929);
or (n2964,n2965,n2968);
and (n2965,n2966,n2967);
xor (n2966,n2871,n2872);
and (n2967,n270,n72);
and (n2968,n2969,n2970);
xor (n2969,n2966,n2967);
or (n2970,n2971,n2974);
and (n2971,n2972,n2973);
xor (n2972,n2877,n2878);
and (n2973,n329,n72);
and (n2974,n2975,n2976);
xor (n2975,n2972,n2973);
or (n2976,n2977,n2980);
and (n2977,n2978,n2979);
xor (n2978,n2883,n2884);
and (n2979,n381,n72);
and (n2980,n2981,n2982);
xor (n2981,n2978,n2979);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
xor (n2984,n2889,n2890);
and (n2985,n770,n72);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
or (n2988,n2989,n2992);
and (n2989,n2990,n2991);
xor (n2990,n2895,n2896);
and (n2991,n803,n72);
and (n2992,n2993,n2994);
xor (n2993,n2990,n2991);
and (n2994,n2995,n2996);
xor (n2995,n2901,n2902);
and (n2996,n864,n72);
and (n2997,n38,n71);
and (n2998,n2999,n3000);
xor (n2999,n1959,n2997);
or (n3000,n3001,n3004);
and (n3001,n3002,n3003);
xor (n3002,n2906,n2907);
and (n3003,n34,n71);
and (n3004,n3005,n3006);
xor (n3005,n3002,n3003);
or (n3006,n3007,n3010);
and (n3007,n3008,n3009);
xor (n3008,n2912,n2913);
and (n3009,n42,n71);
and (n3010,n3011,n3012);
xor (n3011,n3008,n3009);
or (n3012,n3013,n3016);
and (n3013,n3014,n3015);
xor (n3014,n2918,n2919);
and (n3015,n86,n71);
and (n3016,n3017,n3018);
xor (n3017,n3014,n3015);
or (n3018,n3019,n3022);
and (n3019,n3020,n3021);
xor (n3020,n2924,n2925);
and (n3021,n220,n71);
and (n3022,n3023,n3024);
xor (n3023,n3020,n3021);
or (n3024,n3025,n3028);
and (n3025,n3026,n3027);
xor (n3026,n2930,n2931);
and (n3027,n215,n71);
and (n3028,n3029,n3030);
xor (n3029,n3026,n3027);
or (n3030,n3031,n3034);
and (n3031,n3032,n3033);
xor (n3032,n2936,n2937);
and (n3033,n121,n71);
and (n3034,n3035,n3036);
xor (n3035,n3032,n3033);
or (n3036,n3037,n3040);
and (n3037,n3038,n3039);
xor (n3038,n2941,n2942);
and (n3039,n115,n71);
and (n3040,n3041,n3042);
xor (n3041,n3038,n3039);
or (n3042,n3043,n3046);
and (n3043,n3044,n3045);
xor (n3044,n2946,n2947);
and (n3045,n160,n71);
and (n3046,n3047,n3048);
xor (n3047,n3044,n3045);
or (n3048,n3049,n3052);
and (n3049,n3050,n3051);
xor (n3050,n2952,n2953);
and (n3051,n154,n71);
and (n3052,n3053,n3054);
xor (n3053,n3050,n3051);
or (n3054,n3055,n3058);
and (n3055,n3056,n3057);
xor (n3056,n2958,n2959);
and (n3057,n249,n71);
and (n3058,n3059,n3060);
xor (n3059,n3056,n3057);
or (n3060,n3061,n3064);
and (n3061,n3062,n3063);
xor (n3062,n2963,n2964);
and (n3063,n270,n71);
and (n3064,n3065,n3066);
xor (n3065,n3062,n3063);
or (n3066,n3067,n3070);
and (n3067,n3068,n3069);
xor (n3068,n2969,n2970);
and (n3069,n329,n71);
and (n3070,n3071,n3072);
xor (n3071,n3068,n3069);
or (n3072,n3073,n3076);
and (n3073,n3074,n3075);
xor (n3074,n2975,n2976);
and (n3075,n381,n71);
and (n3076,n3077,n3078);
xor (n3077,n3074,n3075);
or (n3078,n3079,n3082);
and (n3079,n3080,n3081);
xor (n3080,n2981,n2982);
and (n3081,n770,n71);
and (n3082,n3083,n3084);
xor (n3083,n3080,n3081);
or (n3084,n3085,n3088);
and (n3085,n3086,n3087);
xor (n3086,n2987,n2988);
and (n3087,n803,n71);
and (n3088,n3089,n3090);
xor (n3089,n3086,n3087);
and (n3090,n3091,n3092);
xor (n3091,n2993,n2994);
not (n3092,n1236);
and (n3093,n38,n16);
and (n3094,n3095,n3096);
xor (n3095,n1957,n3093);
or (n3096,n3097,n3100);
and (n3097,n3098,n3099);
xor (n3098,n2999,n3000);
and (n3099,n34,n16);
and (n3100,n3101,n3102);
xor (n3101,n3098,n3099);
or (n3102,n3103,n3106);
and (n3103,n3104,n3105);
xor (n3104,n3005,n3006);
and (n3105,n42,n16);
and (n3106,n3107,n3108);
xor (n3107,n3104,n3105);
or (n3108,n3109,n3112);
and (n3109,n3110,n3111);
xor (n3110,n3011,n3012);
and (n3111,n86,n16);
and (n3112,n3113,n3114);
xor (n3113,n3110,n3111);
or (n3114,n3115,n3118);
and (n3115,n3116,n3117);
xor (n3116,n3017,n3018);
and (n3117,n220,n16);
and (n3118,n3119,n3120);
xor (n3119,n3116,n3117);
or (n3120,n3121,n3124);
and (n3121,n3122,n3123);
xor (n3122,n3023,n3024);
and (n3123,n215,n16);
and (n3124,n3125,n3126);
xor (n3125,n3122,n3123);
or (n3126,n3127,n3130);
and (n3127,n3128,n3129);
xor (n3128,n3029,n3030);
and (n3129,n121,n16);
and (n3130,n3131,n3132);
xor (n3131,n3128,n3129);
or (n3132,n3133,n3136);
and (n3133,n3134,n3135);
xor (n3134,n3035,n3036);
and (n3135,n115,n16);
and (n3136,n3137,n3138);
xor (n3137,n3134,n3135);
or (n3138,n3139,n3142);
and (n3139,n3140,n3141);
xor (n3140,n3041,n3042);
and (n3141,n160,n16);
and (n3142,n3143,n3144);
xor (n3143,n3140,n3141);
or (n3144,n3145,n3148);
and (n3145,n3146,n3147);
xor (n3146,n3047,n3048);
and (n3147,n154,n16);
and (n3148,n3149,n3150);
xor (n3149,n3146,n3147);
or (n3150,n3151,n3154);
and (n3151,n3152,n3153);
xor (n3152,n3053,n3054);
and (n3153,n249,n16);
and (n3154,n3155,n3156);
xor (n3155,n3152,n3153);
or (n3156,n3157,n3160);
and (n3157,n3158,n3159);
xor (n3158,n3059,n3060);
and (n3159,n270,n16);
and (n3160,n3161,n3162);
xor (n3161,n3158,n3159);
or (n3162,n3163,n3166);
and (n3163,n3164,n3165);
xor (n3164,n3065,n3066);
and (n3165,n329,n16);
and (n3166,n3167,n3168);
xor (n3167,n3164,n3165);
or (n3168,n3169,n3172);
and (n3169,n3170,n3171);
xor (n3170,n3071,n3072);
and (n3171,n381,n16);
and (n3172,n3173,n3174);
xor (n3173,n3170,n3171);
or (n3174,n3175,n3178);
and (n3175,n3176,n3177);
xor (n3176,n3077,n3078);
and (n3177,n770,n16);
and (n3178,n3179,n3180);
xor (n3179,n3176,n3177);
or (n3180,n3181,n3184);
and (n3181,n3182,n3183);
xor (n3182,n3083,n3084);
and (n3183,n803,n16);
and (n3184,n3185,n3186);
xor (n3185,n3182,n3183);
and (n3186,n3187,n3188);
xor (n3187,n3089,n3090);
and (n3188,n864,n16);
and (n3189,n38,n17);
and (n3190,n3191,n3192);
xor (n3191,n1955,n3189);
or (n3192,n3193,n3196);
and (n3193,n3194,n3195);
xor (n3194,n3095,n3096);
and (n3195,n34,n17);
and (n3196,n3197,n3198);
xor (n3197,n3194,n3195);
or (n3198,n3199,n3202);
and (n3199,n3200,n3201);
xor (n3200,n3101,n3102);
and (n3201,n42,n17);
and (n3202,n3203,n3204);
xor (n3203,n3200,n3201);
or (n3204,n3205,n3208);
and (n3205,n3206,n3207);
xor (n3206,n3107,n3108);
and (n3207,n86,n17);
and (n3208,n3209,n3210);
xor (n3209,n3206,n3207);
or (n3210,n3211,n3214);
and (n3211,n3212,n3213);
xor (n3212,n3113,n3114);
and (n3213,n220,n17);
and (n3214,n3215,n3216);
xor (n3215,n3212,n3213);
or (n3216,n3217,n3220);
and (n3217,n3218,n3219);
xor (n3218,n3119,n3120);
and (n3219,n215,n17);
and (n3220,n3221,n3222);
xor (n3221,n3218,n3219);
or (n3222,n3223,n3226);
and (n3223,n3224,n3225);
xor (n3224,n3125,n3126);
and (n3225,n121,n17);
and (n3226,n3227,n3228);
xor (n3227,n3224,n3225);
or (n3228,n3229,n3232);
and (n3229,n3230,n3231);
xor (n3230,n3131,n3132);
and (n3231,n115,n17);
and (n3232,n3233,n3234);
xor (n3233,n3230,n3231);
or (n3234,n3235,n3238);
and (n3235,n3236,n3237);
xor (n3236,n3137,n3138);
and (n3237,n160,n17);
and (n3238,n3239,n3240);
xor (n3239,n3236,n3237);
or (n3240,n3241,n3244);
and (n3241,n3242,n3243);
xor (n3242,n3143,n3144);
and (n3243,n154,n17);
and (n3244,n3245,n3246);
xor (n3245,n3242,n3243);
or (n3246,n3247,n3250);
and (n3247,n3248,n3249);
xor (n3248,n3149,n3150);
and (n3249,n249,n17);
and (n3250,n3251,n3252);
xor (n3251,n3248,n3249);
or (n3252,n3253,n3256);
and (n3253,n3254,n3255);
xor (n3254,n3155,n3156);
and (n3255,n270,n17);
and (n3256,n3257,n3258);
xor (n3257,n3254,n3255);
or (n3258,n3259,n3262);
and (n3259,n3260,n3261);
xor (n3260,n3161,n3162);
and (n3261,n329,n17);
and (n3262,n3263,n3264);
xor (n3263,n3260,n3261);
or (n3264,n3265,n3268);
and (n3265,n3266,n3267);
xor (n3266,n3167,n3168);
and (n3267,n381,n17);
and (n3268,n3269,n3270);
xor (n3269,n3266,n3267);
or (n3270,n3271,n3274);
and (n3271,n3272,n3273);
xor (n3272,n3173,n3174);
and (n3273,n770,n17);
and (n3274,n3275,n3276);
xor (n3275,n3272,n3273);
or (n3276,n3277,n3280);
and (n3277,n3278,n3279);
xor (n3278,n3179,n3180);
and (n3279,n803,n17);
and (n3280,n3281,n3282);
xor (n3281,n3278,n3279);
and (n3282,n3283,n3284);
xor (n3283,n3185,n3186);
not (n3284,n1085);
and (n3285,n38,n22);
and (n3286,n3287,n3288);
xor (n3287,n1953,n3285);
or (n3288,n3289,n3292);
and (n3289,n3290,n3291);
xor (n3290,n3191,n3192);
and (n3291,n34,n22);
and (n3292,n3293,n3294);
xor (n3293,n3290,n3291);
or (n3294,n3295,n3298);
and (n3295,n3296,n3297);
xor (n3296,n3197,n3198);
and (n3297,n42,n22);
and (n3298,n3299,n3300);
xor (n3299,n3296,n3297);
or (n3300,n3301,n3304);
and (n3301,n3302,n3303);
xor (n3302,n3203,n3204);
and (n3303,n86,n22);
and (n3304,n3305,n3306);
xor (n3305,n3302,n3303);
or (n3306,n3307,n3310);
and (n3307,n3308,n3309);
xor (n3308,n3209,n3210);
and (n3309,n220,n22);
and (n3310,n3311,n3312);
xor (n3311,n3308,n3309);
or (n3312,n3313,n3316);
and (n3313,n3314,n3315);
xor (n3314,n3215,n3216);
and (n3315,n215,n22);
and (n3316,n3317,n3318);
xor (n3317,n3314,n3315);
or (n3318,n3319,n3321);
and (n3319,n3320,n471);
xor (n3320,n3221,n3222);
and (n3321,n3322,n3323);
xor (n3322,n3320,n471);
or (n3323,n3324,n3326);
and (n3324,n3325,n237);
xor (n3325,n3227,n3228);
and (n3326,n3327,n3328);
xor (n3327,n3325,n237);
or (n3328,n3329,n3331);
and (n3329,n3330,n161);
xor (n3330,n3233,n3234);
and (n3331,n3332,n3333);
xor (n3332,n3330,n161);
or (n3333,n3334,n3337);
and (n3334,n3335,n3336);
xor (n3335,n3239,n3240);
and (n3336,n154,n22);
and (n3337,n3338,n3339);
xor (n3338,n3335,n3336);
or (n3339,n3340,n3343);
and (n3340,n3341,n3342);
xor (n3341,n3245,n3246);
and (n3342,n249,n22);
and (n3343,n3344,n3345);
xor (n3344,n3341,n3342);
or (n3345,n3346,n3348);
and (n3346,n3347,n418);
xor (n3347,n3251,n3252);
and (n3348,n3349,n3350);
xor (n3349,n3347,n418);
or (n3350,n3351,n3353);
and (n3351,n3352,n716);
xor (n3352,n3257,n3258);
and (n3353,n3354,n3355);
xor (n3354,n3352,n716);
or (n3355,n3356,n3358);
and (n3356,n3357,n798);
xor (n3357,n3263,n3264);
and (n3358,n3359,n3360);
xor (n3359,n3357,n798);
or (n3360,n3361,n3364);
and (n3361,n3362,n3363);
xor (n3362,n3269,n3270);
and (n3363,n770,n22);
and (n3364,n3365,n3366);
xor (n3365,n3362,n3363);
or (n3366,n3367,n3370);
and (n3367,n3368,n3369);
xor (n3368,n3275,n3276);
and (n3369,n803,n22);
and (n3370,n3371,n3372);
xor (n3371,n3368,n3369);
and (n3372,n3373,n3374);
xor (n3373,n3281,n3282);
and (n3374,n864,n22);
and (n3375,n38,n29);
and (n3376,n3377,n3378);
xor (n3377,n1951,n3375);
or (n3378,n3379,n3382);
and (n3379,n3380,n3381);
xor (n3380,n3287,n3288);
and (n3381,n34,n29);
and (n3382,n3383,n3384);
xor (n3383,n3380,n3381);
or (n3384,n3385,n3388);
and (n3385,n3386,n3387);
xor (n3386,n3293,n3294);
and (n3387,n42,n29);
and (n3388,n3389,n3390);
xor (n3389,n3386,n3387);
or (n3390,n3391,n3394);
and (n3391,n3392,n3393);
xor (n3392,n3299,n3300);
and (n3393,n86,n29);
and (n3394,n3395,n3396);
xor (n3395,n3392,n3393);
or (n3396,n3397,n3400);
and (n3397,n3398,n3399);
xor (n3398,n3305,n3306);
and (n3399,n220,n29);
and (n3400,n3401,n3402);
xor (n3401,n3398,n3399);
or (n3402,n3403,n3406);
and (n3403,n3404,n3405);
xor (n3404,n3311,n3312);
and (n3405,n215,n29);
and (n3406,n3407,n3408);
xor (n3407,n3404,n3405);
or (n3408,n3409,n3412);
and (n3409,n3410,n3411);
xor (n3410,n3317,n3318);
and (n3411,n121,n29);
and (n3412,n3413,n3414);
xor (n3413,n3410,n3411);
or (n3414,n3415,n3418);
and (n3415,n3416,n3417);
xor (n3416,n3322,n3323);
and (n3417,n115,n29);
and (n3418,n3419,n3420);
xor (n3419,n3416,n3417);
or (n3420,n3421,n3424);
and (n3421,n3422,n3423);
xor (n3422,n3327,n3328);
and (n3423,n160,n29);
and (n3424,n3425,n3426);
xor (n3425,n3422,n3423);
or (n3426,n3427,n3430);
and (n3427,n3428,n3429);
xor (n3428,n3332,n3333);
and (n3429,n154,n29);
and (n3430,n3431,n3432);
xor (n3431,n3428,n3429);
or (n3432,n3433,n3436);
and (n3433,n3434,n3435);
xor (n3434,n3338,n3339);
and (n3435,n249,n29);
and (n3436,n3437,n3438);
xor (n3437,n3434,n3435);
or (n3438,n3439,n3442);
and (n3439,n3440,n3441);
xor (n3440,n3344,n3345);
and (n3441,n270,n29);
and (n3442,n3443,n3444);
xor (n3443,n3440,n3441);
or (n3444,n3445,n3448);
and (n3445,n3446,n3447);
xor (n3446,n3349,n3350);
and (n3447,n329,n29);
and (n3448,n3449,n3450);
xor (n3449,n3446,n3447);
or (n3450,n3451,n3454);
and (n3451,n3452,n3453);
xor (n3452,n3354,n3355);
and (n3453,n381,n29);
and (n3454,n3455,n3456);
xor (n3455,n3452,n3453);
or (n3456,n3457,n3460);
and (n3457,n3458,n3459);
xor (n3458,n3359,n3360);
and (n3459,n770,n29);
and (n3460,n3461,n3462);
xor (n3461,n3458,n3459);
or (n3462,n3463,n3466);
and (n3463,n3464,n3465);
xor (n3464,n3365,n3366);
and (n3465,n803,n29);
and (n3466,n3467,n3468);
xor (n3467,n3464,n3465);
and (n3468,n3469,n3470);
xor (n3469,n3371,n3372);
and (n3470,n864,n29);
endmodule
