module top (out,n16,n17,n22,n27,n33,n42,n43,n49,n53
        ,n59,n77,n84,n85,n95,n118,n120,n125,n135,n152
        ,n161,n170,n174,n181,n209);
output out;
input n16;
input n17;
input n22;
input n27;
input n33;
input n42;
input n43;
input n49;
input n53;
input n59;
input n77;
input n84;
input n85;
input n95;
input n118;
input n120;
input n125;
input n135;
input n152;
input n161;
input n170;
input n174;
input n181;
input n209;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
xor (out,n0,n538);
nand (n0,n1,n537);
or (n1,n2,n290);
not (n2,n3);
nand (n3,n4,n289);
nand (n4,n5,n253);
not (n5,n6);
xor (n6,n7,n211);
xor (n7,n8,n98);
xor (n8,n9,n62);
xor (n9,n10,n36);
nand (n10,n11,n30);
or (n11,n12,n24);
nand (n12,n13,n20);
nor (n13,n14,n18);
and (n14,n15,n17);
not (n15,n16);
and (n18,n16,n19);
not (n19,n17);
nand (n20,n21,n23);
or (n21,n19,n22);
nand (n23,n19,n22);
nor (n24,n25,n28);
and (n25,n26,n27);
not (n26,n22);
and (n28,n29,n22);
not (n29,n27);
or (n30,n13,n31);
nor (n31,n32,n34);
and (n32,n33,n26);
and (n34,n35,n22);
not (n35,n33);
nand (n36,n37,n56);
or (n37,n38,n51);
nand (n38,n39,n46);
nor (n39,n40,n44);
and (n40,n41,n43);
not (n41,n42);
and (n44,n42,n45);
not (n45,n43);
nand (n46,n47,n50);
or (n47,n43,n48);
not (n48,n49);
nand (n50,n48,n43);
nor (n51,n52,n54);
and (n52,n48,n53);
and (n54,n49,n55);
not (n55,n53);
or (n56,n39,n57);
nor (n57,n58,n60);
and (n58,n48,n59);
and (n60,n49,n61);
not (n61,n59);
nand (n62,n63,n97);
or (n63,n64,n70);
not (n64,n65);
nand (n65,n66,n22);
nand (n66,n67,n68);
or (n67,n16,n17);
nand (n68,n69,n29);
or (n69,n19,n15);
not (n70,n71);
nand (n71,n72,n91);
or (n72,n73,n79);
not (n73,n74);
nor (n74,n75,n78);
and (n75,n76,n41);
not (n76,n77);
and (n78,n42,n77);
not (n79,n80);
nor (n80,n81,n87);
nand (n81,n82,n86);
or (n82,n83,n85);
not (n83,n84);
nand (n86,n83,n85);
nor (n87,n88,n89);
and (n88,n41,n85);
and (n89,n42,n90);
not (n90,n85);
nand (n91,n81,n92);
nand (n92,n93,n96);
or (n93,n42,n94);
not (n94,n95);
or (n96,n41,n95);
or (n97,n71,n65);
xor (n98,n99,n186);
xor (n99,n100,n138);
or (n100,n101,n137);
and (n101,n102,n112);
xor (n102,n103,n105);
and (n103,n104,n27);
not (n104,n13);
nand (n105,n106,n111);
or (n106,n107,n79);
not (n107,n108);
nand (n108,n109,n110);
or (n109,n42,n61);
or (n110,n41,n59);
nand (n111,n81,n74);
nand (n112,n113,n131);
or (n113,n114,n122);
not (n114,n115);
nor (n115,n116,n121);
and (n116,n117,n119);
not (n117,n118);
not (n119,n120);
and (n121,n120,n118);
nand (n122,n123,n127);
nand (n123,n124,n126);
or (n124,n125,n119);
nand (n126,n119,n125);
not (n127,n128);
nand (n128,n129,n130);
or (n129,n48,n125);
nand (n130,n48,n125);
nand (n131,n128,n132);
nand (n132,n133,n136);
or (n133,n120,n134);
not (n134,n135);
or (n136,n119,n135);
and (n137,n103,n105);
or (n138,n139,n185);
and (n139,n140,n177);
xor (n140,n141,n163);
nand (n141,n142,n157);
or (n142,n143,n147);
not (n143,n144);
nand (n144,n145,n146);
or (n145,n16,n35);
or (n146,n15,n33);
not (n147,n148);
and (n148,n149,n154);
not (n149,n150);
nand (n150,n151,n153);
or (n151,n152,n119);
nand (n153,n152,n119);
nand (n154,n155,n156);
or (n155,n152,n15);
nand (n156,n15,n152);
nand (n157,n150,n158);
nand (n158,n159,n162);
or (n159,n16,n160);
not (n160,n161);
or (n162,n15,n161);
nand (n163,n164,n171);
or (n164,n165,n168);
nor (n165,n166,n167);
and (n166,n83,n95);
and (n167,n84,n94);
nand (n168,n84,n169);
not (n169,n170);
or (n171,n172,n169);
nor (n172,n173,n175);
and (n173,n83,n174);
and (n175,n84,n176);
not (n176,n174);
nand (n177,n178,n184);
or (n178,n38,n179);
nor (n179,n180,n182);
and (n180,n48,n181);
and (n182,n49,n183);
not (n183,n181);
or (n184,n51,n39);
and (n185,n141,n163);
xor (n186,n187,n203);
xor (n187,n188,n196);
nand (n188,n189,n191);
or (n189,n190,n122);
not (n190,n132);
nand (n191,n192,n128);
not (n192,n193);
nor (n193,n194,n195);
and (n194,n119,n181);
and (n195,n120,n183);
nand (n196,n197,n199);
or (n197,n198,n147);
not (n198,n158);
or (n199,n149,n200);
nor (n200,n201,n202);
and (n201,n15,n118);
and (n202,n16,n117);
nand (n203,n204,n205);
or (n204,n172,n168);
or (n205,n206,n169);
nor (n206,n207,n210);
and (n207,n208,n84);
not (n208,n209);
and (n210,n209,n83);
or (n211,n212,n252);
and (n212,n213,n251);
xor (n213,n214,n229);
and (n214,n215,n221);
and (n215,n216,n16);
nand (n216,n217,n218);
or (n217,n120,n152);
nand (n218,n219,n29);
or (n219,n220,n119);
not (n220,n152);
nand (n221,n222,n224);
or (n222,n223,n107);
not (n223,n81);
nand (n224,n225,n80);
not (n225,n226);
nor (n226,n227,n228);
and (n227,n41,n53);
and (n228,n42,n55);
or (n229,n230,n250);
and (n230,n231,n244);
xor (n231,n232,n238);
nand (n232,n233,n237);
or (n233,n122,n234);
nor (n234,n235,n236);
and (n235,n160,n120);
and (n236,n161,n119);
nand (n237,n115,n128);
nand (n238,n239,n240);
or (n239,n149,n143);
nand (n240,n148,n241);
nand (n241,n242,n243);
or (n242,n16,n29);
or (n243,n15,n27);
nand (n244,n245,n249);
or (n245,n168,n246);
nor (n246,n247,n248);
and (n247,n83,n77);
and (n248,n84,n76);
or (n249,n165,n169);
and (n250,n232,n238);
xor (n251,n102,n112);
and (n252,n214,n229);
not (n253,n254);
or (n254,n255,n288);
and (n255,n256,n287);
xor (n256,n257,n258);
xor (n257,n140,n177);
or (n258,n259,n286);
and (n259,n260,n268);
xor (n260,n261,n267);
nand (n261,n262,n266);
or (n262,n38,n263);
nor (n263,n264,n265);
and (n264,n135,n48);
and (n265,n49,n134);
or (n266,n179,n39);
xor (n267,n215,n221);
or (n268,n269,n285);
and (n269,n270,n278);
xor (n270,n271,n272);
and (n271,n150,n27);
nand (n272,n273,n277);
or (n273,n274,n168);
nor (n274,n275,n276);
and (n275,n61,n84);
and (n276,n59,n83);
or (n277,n246,n169);
nand (n278,n279,n284);
or (n279,n122,n280);
not (n280,n281);
nor (n281,n282,n283);
and (n282,n35,n119);
and (n283,n120,n33);
or (n284,n127,n234);
and (n285,n271,n272);
and (n286,n261,n267);
xor (n287,n213,n251);
and (n288,n257,n258);
nand (n289,n6,n254);
not (n290,n291);
nand (n291,n292,n536);
or (n292,n293,n528);
nor (n293,n294,n524);
and (n294,n295,n491);
or (n295,n296,n490);
and (n296,n297,n384);
xor (n297,n298,n346);
or (n298,n299,n345);
and (n299,n300,n325);
xor (n300,n301,n310);
nand (n301,n302,n306);
or (n302,n38,n303);
nor (n303,n304,n305);
and (n304,n48,n33);
and (n305,n49,n35);
or (n306,n39,n307);
nor (n307,n308,n309);
and (n308,n48,n161);
and (n309,n49,n160);
and (n310,n311,n316);
and (n311,n312,n49);
nand (n312,n313,n314);
or (n313,n42,n43);
nand (n314,n315,n29);
or (n315,n45,n41);
nand (n316,n317,n321);
or (n317,n318,n168);
nor (n318,n319,n320);
and (n319,n83,n135);
and (n320,n84,n134);
or (n321,n322,n169);
nor (n322,n323,n324);
and (n323,n83,n181);
and (n324,n84,n183);
xor (n325,n326,n335);
xor (n326,n327,n328);
and (n327,n128,n27);
nand (n328,n329,n334);
or (n329,n169,n330);
not (n330,n331);
nor (n331,n332,n333);
and (n332,n84,n53);
and (n333,n55,n83);
or (n334,n168,n322);
nand (n335,n336,n341);
or (n336,n337,n79);
not (n337,n338);
nor (n338,n339,n340);
and (n339,n42,n118);
and (n340,n117,n41);
nand (n341,n81,n342);
nand (n342,n343,n344);
or (n343,n42,n134);
or (n344,n41,n135);
and (n345,n301,n310);
xor (n346,n347,n361);
xor (n347,n348,n358);
xor (n348,n349,n355);
nor (n349,n350,n119);
nor (n350,n351,n353);
and (n351,n352,n29);
nand (n352,n49,n125);
and (n353,n48,n354);
not (n354,n125);
nand (n355,n356,n357);
or (n356,n168,n330);
or (n357,n274,n169);
or (n358,n359,n360);
and (n359,n326,n335);
and (n360,n327,n328);
xor (n361,n362,n378);
xor (n362,n363,n370);
nand (n363,n364,n369);
or (n364,n365,n122);
not (n365,n366);
nand (n366,n367,n368);
or (n367,n120,n29);
or (n368,n119,n27);
nand (n369,n281,n128);
nand (n370,n371,n373);
or (n371,n372,n79);
not (n372,n342);
nand (n373,n374,n81);
not (n374,n375);
nor (n375,n376,n377);
and (n376,n183,n42);
and (n377,n181,n41);
nand (n378,n379,n380);
or (n379,n38,n307);
or (n380,n39,n381);
nor (n381,n382,n383);
and (n382,n118,n48);
and (n383,n49,n117);
or (n384,n385,n489);
and (n385,n386,n407);
xor (n386,n387,n406);
or (n387,n388,n405);
and (n388,n389,n404);
xor (n389,n390,n397);
nand (n390,n391,n396);
or (n391,n392,n79);
not (n392,n393);
nor (n393,n394,n395);
and (n394,n160,n41);
and (n395,n42,n161);
nand (n396,n81,n338);
nand (n397,n398,n403);
or (n398,n399,n38);
not (n399,n400);
nand (n400,n401,n402);
or (n401,n29,n49);
or (n402,n48,n27);
or (n403,n39,n303);
xor (n404,n311,n316);
and (n405,n390,n397);
xor (n406,n300,n325);
or (n407,n408,n488);
and (n408,n409,n429);
xor (n409,n410,n428);
or (n410,n411,n427);
and (n411,n412,n420);
xor (n412,n413,n414);
nor (n413,n39,n29);
nand (n414,n415,n419);
or (n415,n416,n79);
nor (n416,n417,n418);
and (n417,n33,n41);
and (n418,n35,n42);
nand (n419,n393,n81);
nand (n420,n421,n426);
or (n421,n168,n422);
not (n422,n423);
nand (n423,n424,n425);
or (n424,n118,n83);
nand (n425,n83,n118);
or (n426,n318,n169);
and (n427,n413,n414);
xor (n428,n389,n404);
or (n429,n430,n487);
and (n430,n431,n486);
xor (n431,n432,n447);
nor (n432,n433,n441);
not (n433,n434);
nand (n434,n435,n440);
or (n435,n168,n436);
not (n436,n437);
nand (n437,n438,n439);
or (n438,n161,n83);
nand (n439,n83,n161);
nand (n440,n423,n170);
nand (n441,n442,n42);
nand (n442,n443,n446);
nand (n443,n444,n29);
not (n444,n445);
and (n445,n84,n85);
or (n446,n85,n84);
nand (n447,n448,n485);
nand (n448,n449,n462);
or (n449,n450,n457);
not (n450,n451);
nor (n451,n452,n456);
and (n452,n80,n453);
nand (n453,n454,n455);
or (n454,n42,n29);
or (n455,n41,n27);
nor (n456,n223,n416);
not (n457,n458);
nor (n458,n459,n460);
and (n459,n441,n434);
and (n460,n461,n433);
not (n461,n441);
nand (n462,n463,n484);
or (n463,n464,n474);
nor (n464,n465,n467);
not (n465,n466);
nand (n466,n81,n27);
nand (n467,n468,n469);
or (n468,n169,n436);
nand (n469,n470,n473);
nand (n470,n471,n472);
or (n471,n35,n84);
nand (n472,n84,n35);
not (n473,n168);
nand (n474,n475,n482);
nand (n475,n476,n480);
or (n476,n477,n168);
nor (n477,n478,n479);
and (n478,n29,n84);
and (n479,n27,n83);
or (n480,n481,n169);
not (n481,n470);
nor (n482,n483,n83);
and (n483,n27,n170);
nand (n484,n465,n467);
or (n485,n458,n451);
xor (n486,n412,n420);
and (n487,n432,n447);
and (n488,n410,n428);
and (n489,n387,n406);
and (n490,n298,n346);
not (n491,n492);
nand (n492,n493,n519);
not (n493,n494);
nor (n494,n495,n510);
xor (n495,n496,n509);
xor (n496,n497,n498);
xor (n497,n231,n244);
or (n498,n499,n508);
and (n499,n500,n507);
xor (n500,n501,n504);
nand (n501,n502,n503);
or (n502,n79,n375);
or (n503,n223,n226);
nand (n504,n505,n506);
or (n505,n38,n381);
or (n506,n39,n263);
and (n507,n349,n355);
and (n508,n501,n504);
xor (n509,n260,n268);
or (n510,n511,n518);
and (n511,n512,n517);
xor (n512,n513,n516);
or (n513,n514,n515);
and (n514,n362,n378);
and (n515,n363,n370);
xor (n516,n270,n278);
xor (n517,n500,n507);
and (n518,n513,n516);
or (n519,n520,n521);
xor (n520,n512,n517);
or (n521,n522,n523);
and (n522,n347,n361);
and (n523,n348,n358);
nand (n524,n525,n527);
or (n525,n494,n526);
nand (n526,n520,n521);
nand (n527,n495,n510);
not (n528,n529);
nand (n529,n530,n532);
not (n530,n531);
xor (n531,n256,n287);
not (n532,n533);
or (n533,n534,n535);
and (n534,n496,n509);
and (n535,n497,n498);
nand (n536,n531,n533);
or (n537,n291,n3);
xor (n538,n539,n864);
xor (n539,n540,n861);
xor (n540,n541,n860);
xor (n541,n542,n851);
xor (n542,n543,n850);
xor (n543,n544,n835);
xor (n544,n545,n78);
xor (n545,n546,n814);
xor (n546,n547,n813);
xor (n547,n548,n787);
xor (n548,n549,n786);
xor (n549,n550,n753);
xor (n550,n551,n752);
xor (n551,n552,n713);
xor (n552,n553,n712);
xor (n553,n554,n669);
xor (n554,n555,n668);
xor (n555,n556,n618);
xor (n556,n557,n617);
xor (n557,n558,n561);
xor (n558,n559,n560);
and (n559,n22,n27);
and (n560,n17,n33);
or (n561,n562,n565);
and (n562,n563,n564);
and (n563,n17,n27);
and (n564,n16,n33);
and (n565,n566,n567);
xor (n566,n563,n564);
or (n567,n568,n571);
and (n568,n569,n570);
and (n569,n16,n27);
and (n570,n152,n33);
and (n571,n572,n573);
xor (n572,n569,n570);
or (n573,n574,n576);
and (n574,n575,n283);
and (n575,n152,n27);
and (n576,n577,n578);
xor (n577,n575,n283);
or (n578,n579,n582);
and (n579,n580,n581);
and (n580,n120,n27);
and (n581,n125,n33);
and (n582,n583,n584);
xor (n583,n580,n581);
or (n584,n585,n588);
and (n585,n586,n587);
and (n586,n125,n27);
and (n587,n49,n33);
and (n588,n589,n590);
xor (n589,n586,n587);
or (n590,n591,n594);
and (n591,n592,n593);
and (n592,n49,n27);
and (n593,n43,n33);
and (n594,n595,n596);
xor (n595,n592,n593);
or (n596,n597,n600);
and (n597,n598,n599);
and (n598,n43,n27);
and (n599,n42,n33);
and (n600,n601,n602);
xor (n601,n598,n599);
or (n602,n603,n606);
and (n603,n604,n605);
and (n604,n42,n27);
and (n605,n85,n33);
and (n606,n607,n608);
xor (n607,n604,n605);
or (n608,n609,n612);
and (n609,n610,n611);
and (n610,n85,n27);
and (n611,n84,n33);
and (n612,n613,n614);
xor (n613,n610,n611);
and (n614,n615,n616);
and (n615,n84,n27);
and (n616,n170,n33);
and (n617,n16,n161);
or (n618,n619,n622);
and (n619,n620,n621);
xor (n620,n566,n567);
and (n621,n152,n161);
and (n622,n623,n624);
xor (n623,n620,n621);
or (n624,n625,n628);
and (n625,n626,n627);
xor (n626,n572,n573);
and (n627,n120,n161);
and (n628,n629,n630);
xor (n629,n626,n627);
or (n630,n631,n634);
and (n631,n632,n633);
xor (n632,n577,n578);
and (n633,n125,n161);
and (n634,n635,n636);
xor (n635,n632,n633);
or (n636,n637,n640);
and (n637,n638,n639);
xor (n638,n583,n584);
and (n639,n49,n161);
and (n640,n641,n642);
xor (n641,n638,n639);
or (n642,n643,n646);
and (n643,n644,n645);
xor (n644,n589,n590);
and (n645,n43,n161);
and (n646,n647,n648);
xor (n647,n644,n645);
or (n648,n649,n651);
and (n649,n650,n395);
xor (n650,n595,n596);
and (n651,n652,n653);
xor (n652,n650,n395);
or (n653,n654,n657);
and (n654,n655,n656);
xor (n655,n601,n602);
and (n656,n85,n161);
and (n657,n658,n659);
xor (n658,n655,n656);
or (n659,n660,n663);
and (n660,n661,n662);
xor (n661,n607,n608);
and (n662,n84,n161);
and (n663,n664,n665);
xor (n664,n661,n662);
and (n665,n666,n667);
xor (n666,n613,n614);
and (n667,n170,n161);
and (n668,n152,n118);
or (n669,n670,n672);
and (n670,n671,n121);
xor (n671,n623,n624);
and (n672,n673,n674);
xor (n673,n671,n121);
or (n674,n675,n678);
and (n675,n676,n677);
xor (n676,n629,n630);
and (n677,n125,n118);
and (n678,n679,n680);
xor (n679,n676,n677);
or (n680,n681,n684);
and (n681,n682,n683);
xor (n682,n635,n636);
and (n683,n49,n118);
and (n684,n685,n686);
xor (n685,n682,n683);
or (n686,n687,n690);
and (n687,n688,n689);
xor (n688,n641,n642);
and (n689,n43,n118);
and (n690,n691,n692);
xor (n691,n688,n689);
or (n692,n693,n695);
and (n693,n694,n339);
xor (n694,n647,n648);
and (n695,n696,n697);
xor (n696,n694,n339);
or (n697,n698,n701);
and (n698,n699,n700);
xor (n699,n652,n653);
and (n700,n85,n118);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n658,n659);
and (n706,n84,n118);
and (n707,n708,n709);
xor (n708,n705,n706);
and (n709,n710,n711);
xor (n710,n664,n665);
and (n711,n170,n118);
and (n712,n120,n135);
or (n713,n714,n717);
and (n714,n715,n716);
xor (n715,n673,n674);
and (n716,n125,n135);
and (n717,n718,n719);
xor (n718,n715,n716);
or (n719,n720,n723);
and (n720,n721,n722);
xor (n721,n679,n680);
and (n722,n49,n135);
and (n723,n724,n725);
xor (n724,n721,n722);
or (n725,n726,n729);
and (n726,n727,n728);
xor (n727,n685,n686);
and (n728,n43,n135);
and (n729,n730,n731);
xor (n730,n727,n728);
or (n731,n732,n735);
and (n732,n733,n734);
xor (n733,n691,n692);
and (n734,n42,n135);
and (n735,n736,n737);
xor (n736,n733,n734);
or (n737,n738,n741);
and (n738,n739,n740);
xor (n739,n696,n697);
and (n740,n85,n135);
and (n741,n742,n743);
xor (n742,n739,n740);
or (n743,n744,n747);
and (n744,n745,n746);
xor (n745,n702,n703);
and (n746,n84,n135);
and (n747,n748,n749);
xor (n748,n745,n746);
and (n749,n750,n751);
xor (n750,n708,n709);
and (n751,n170,n135);
and (n752,n125,n181);
or (n753,n754,n757);
and (n754,n755,n756);
xor (n755,n718,n719);
and (n756,n49,n181);
and (n757,n758,n759);
xor (n758,n755,n756);
or (n759,n760,n763);
and (n760,n761,n762);
xor (n761,n724,n725);
and (n762,n43,n181);
and (n763,n764,n765);
xor (n764,n761,n762);
or (n765,n766,n769);
and (n766,n767,n768);
xor (n767,n730,n731);
and (n768,n42,n181);
and (n769,n770,n771);
xor (n770,n767,n768);
or (n771,n772,n775);
and (n772,n773,n774);
xor (n773,n736,n737);
and (n774,n85,n181);
and (n775,n776,n777);
xor (n776,n773,n774);
or (n777,n778,n781);
and (n778,n779,n780);
xor (n779,n742,n743);
and (n780,n84,n181);
and (n781,n782,n783);
xor (n782,n779,n780);
and (n783,n784,n785);
xor (n784,n748,n749);
and (n785,n170,n181);
and (n786,n49,n53);
or (n787,n788,n791);
and (n788,n789,n790);
xor (n789,n758,n759);
and (n790,n43,n53);
and (n791,n792,n793);
xor (n792,n789,n790);
or (n793,n794,n797);
and (n794,n795,n796);
xor (n795,n764,n765);
and (n796,n42,n53);
and (n797,n798,n799);
xor (n798,n795,n796);
or (n799,n800,n803);
and (n800,n801,n802);
xor (n801,n770,n771);
and (n802,n85,n53);
and (n803,n804,n805);
xor (n804,n801,n802);
or (n805,n806,n808);
and (n806,n807,n332);
xor (n807,n776,n777);
and (n808,n809,n810);
xor (n809,n807,n332);
and (n810,n811,n812);
xor (n811,n782,n783);
and (n812,n170,n53);
and (n813,n43,n59);
or (n814,n815,n818);
and (n815,n816,n817);
xor (n816,n792,n793);
and (n817,n42,n59);
and (n818,n819,n820);
xor (n819,n816,n817);
or (n820,n821,n824);
and (n821,n822,n823);
xor (n822,n798,n799);
and (n823,n85,n59);
and (n824,n825,n826);
xor (n825,n822,n823);
or (n826,n827,n830);
and (n827,n828,n829);
xor (n828,n804,n805);
and (n829,n84,n59);
and (n830,n831,n832);
xor (n831,n828,n829);
and (n832,n833,n834);
xor (n833,n809,n810);
and (n834,n170,n59);
or (n835,n836,n839);
and (n836,n837,n838);
xor (n837,n819,n820);
and (n838,n85,n77);
and (n839,n840,n841);
xor (n840,n837,n838);
or (n841,n842,n845);
and (n842,n843,n844);
xor (n843,n825,n826);
and (n844,n84,n77);
and (n845,n846,n847);
xor (n846,n843,n844);
and (n847,n848,n849);
xor (n848,n831,n832);
and (n849,n170,n77);
and (n850,n85,n95);
or (n851,n852,n855);
and (n852,n853,n854);
xor (n853,n840,n841);
and (n854,n84,n95);
and (n855,n856,n857);
xor (n856,n853,n854);
and (n857,n858,n859);
xor (n858,n846,n847);
and (n859,n170,n95);
and (n860,n84,n174);
and (n861,n862,n863);
xor (n862,n856,n857);
and (n863,n170,n174);
and (n864,n170,n209);
endmodule
