module top (out,n22,n23,n29,n33,n39,n49,n54,n58,n64
        ,n73,n75,n80,n84,n90,n102,n107,n111,n117,n125
        ,n131,n135,n141,n150,n151,n157,n161,n167,n178,n180
        ,n185,n192,n200,n208,n214,n222,n230,n236,n301,n306
        ,n310,n335,n342,n348,n356,n448,n474,n493,n495,n625
        ,n826,n832,n839,n847,n858,n859,n864,n887,n897,n898
        ,n952,n983,n1002,n1030,n1037);
output out;
input n22;
input n23;
input n29;
input n33;
input n39;
input n49;
input n54;
input n58;
input n64;
input n73;
input n75;
input n80;
input n84;
input n90;
input n102;
input n107;
input n111;
input n117;
input n125;
input n131;
input n135;
input n141;
input n150;
input n151;
input n157;
input n161;
input n167;
input n178;
input n180;
input n185;
input n192;
input n200;
input n208;
input n214;
input n222;
input n230;
input n236;
input n301;
input n306;
input n310;
input n335;
input n342;
input n348;
input n356;
input n448;
input n474;
input n493;
input n495;
input n625;
input n826;
input n832;
input n839;
input n847;
input n858;
input n859;
input n864;
input n887;
input n897;
input n898;
input n952;
input n983;
input n1002;
input n1030;
input n1037;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n302;
wire n303;
wire n304;
wire n305;
wire n307;
wire n308;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n494;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n860;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
xor (out,n0,n5163);
nand (n0,n1,n5162);
or (n1,n2,n761);
not (n2,n3);
and (n3,n4,n760);
not (n4,n5);
nor (n5,n6,n659);
or (n6,n7,n658);
and (n7,n8,n588);
xor (n8,n9,n317);
xor (n9,n10,n255);
xor (n10,n11,n240);
or (n11,n12,n239);
and (n12,n13,n170);
xor (n13,n14,n93);
xor (n14,n15,n67);
xor (n15,n16,n42);
nand (n16,n17,n36);
or (n17,n18,n31);
nand (n18,n19,n26);
nor (n19,n20,n24);
and (n20,n21,n23);
not (n21,n22);
and (n24,n22,n25);
not (n25,n23);
nand (n26,n27,n30);
or (n27,n23,n28);
not (n28,n29);
nand (n30,n28,n23);
nor (n31,n32,n34);
and (n32,n28,n33);
and (n34,n29,n35);
not (n35,n33);
or (n36,n19,n37);
nor (n37,n38,n40);
and (n38,n28,n39);
and (n40,n29,n41);
not (n41,n39);
nand (n42,n43,n61);
or (n43,n44,n56);
nand (n44,n45,n51);
not (n45,n46);
nand (n46,n47,n50);
or (n47,n29,n48);
not (n48,n49);
nand (n50,n29,n48);
nand (n51,n52,n55);
or (n52,n49,n53);
not (n53,n54);
nand (n55,n53,n49);
nor (n56,n57,n59);
and (n57,n53,n58);
and (n59,n54,n60);
not (n60,n58);
or (n61,n45,n62);
nor (n62,n63,n65);
and (n63,n53,n64);
and (n65,n54,n66);
not (n66,n64);
nand (n67,n68,n87);
or (n68,n69,n82);
nand (n69,n70,n77);
not (n70,n71);
nand (n71,n72,n76);
or (n72,n73,n74);
not (n74,n75);
nand (n76,n73,n74);
nand (n77,n78,n81);
or (n78,n73,n79);
not (n79,n80);
nand (n81,n79,n73);
nor (n82,n83,n85);
and (n83,n79,n84);
and (n85,n80,n86);
not (n86,n84);
or (n87,n70,n88);
nor (n88,n89,n91);
and (n89,n79,n90);
and (n91,n80,n92);
not (n92,n90);
xor (n93,n94,n144);
xor (n94,n95,n120);
nand (n95,n96,n114);
or (n96,n97,n109);
not (n97,n98);
and (n98,n99,n104);
nor (n99,n100,n103);
and (n100,n54,n101);
not (n101,n102);
and (n103,n53,n102);
nor (n104,n105,n108);
and (n105,n101,n106);
not (n106,n107);
and (n108,n102,n107);
nor (n109,n110,n112);
and (n110,n106,n111);
and (n112,n107,n113);
not (n113,n111);
or (n114,n99,n115);
nor (n115,n116,n118);
and (n116,n106,n117);
and (n118,n107,n119);
not (n119,n117);
nand (n120,n121,n138);
or (n121,n122,n133);
nand (n122,n123,n128);
nor (n123,n124,n126);
and (n124,n106,n125);
and (n126,n107,n127);
not (n127,n125);
nor (n128,n129,n132);
and (n129,n130,n127);
not (n130,n131);
and (n132,n131,n125);
nor (n133,n134,n136);
and (n134,n130,n135);
and (n136,n137,n131);
not (n137,n135);
or (n138,n123,n139);
nor (n139,n140,n142);
and (n140,n130,n141);
and (n142,n143,n131);
not (n143,n141);
nand (n144,n145,n164);
or (n145,n146,n159);
nand (n146,n147,n154);
nor (n147,n148,n152);
and (n148,n149,n151);
not (n149,n150);
and (n152,n150,n153);
not (n153,n151);
nand (n154,n155,n158);
or (n155,n151,n156);
not (n156,n157);
nand (n158,n156,n151);
nor (n159,n160,n162);
and (n160,n156,n161);
and (n162,n157,n163);
not (n163,n161);
or (n164,n147,n165);
nor (n165,n166,n168);
and (n166,n156,n167);
and (n168,n157,n169);
not (n169,n167);
xor (n170,n171,n217);
xor (n171,n172,n195);
nand (n172,n173,n189);
or (n173,n174,n182);
nor (n174,n175,n182);
not (n175,n176);
nand (n176,n177,n181);
or (n177,n178,n179);
not (n179,n180);
nand (n181,n179,n178);
not (n182,n183);
nor (n183,n184,n187);
and (n184,n185,n186);
not (n186,n178);
and (n187,n188,n178);
not (n188,n185);
not (n189,n190);
nor (n190,n191,n193);
and (n191,n179,n192);
and (n193,n180,n194);
not (n194,n192);
nand (n195,n196,n211);
or (n196,n197,n206);
nand (n197,n198,n203);
nor (n198,n199,n201);
and (n199,n179,n200);
and (n201,n180,n202);
not (n202,n200);
nand (n203,n204,n205);
or (n204,n200,n149);
nand (n205,n149,n200);
nor (n206,n207,n209);
and (n207,n149,n208);
and (n209,n150,n210);
not (n210,n208);
or (n211,n198,n212);
nor (n212,n213,n215);
and (n213,n149,n214);
and (n215,n150,n216);
not (n216,n214);
nand (n217,n218,n233);
or (n218,n219,n228);
nand (n219,n220,n225);
nor (n220,n221,n223);
and (n221,n156,n222);
and (n223,n157,n224);
not (n224,n222);
nand (n225,n226,n227);
or (n226,n222,n74);
nand (n227,n74,n222);
nor (n228,n229,n231);
and (n229,n74,n230);
and (n231,n75,n232);
not (n232,n230);
or (n233,n220,n234);
nor (n234,n235,n237);
and (n235,n74,n236);
and (n237,n75,n238);
not (n238,n236);
and (n239,n14,n93);
xor (n240,n241,n252);
xor (n241,n242,n249);
not (n242,n243);
nand (n243,n244,n245);
or (n244,n197,n212);
or (n245,n198,n246);
nor (n246,n247,n248);
and (n247,n149,n192);
and (n248,n150,n194);
or (n249,n250,n251);
and (n250,n171,n217);
and (n251,n172,n195);
or (n252,n253,n254);
and (n253,n15,n67);
and (n254,n16,n42);
xor (n255,n256,n280);
xor (n256,n257,n260);
or (n257,n258,n259);
and (n258,n94,n144);
and (n259,n95,n120);
xor (n260,n261,n274);
xor (n261,n262,n268);
nand (n262,n263,n264);
or (n263,n69,n88);
or (n264,n70,n265);
nor (n265,n266,n267);
and (n266,n79,n230);
and (n267,n80,n232);
nand (n268,n269,n270);
or (n269,n44,n62);
or (n270,n45,n271);
nor (n271,n272,n273);
and (n272,n53,n33);
and (n273,n54,n35);
nand (n274,n275,n279);
or (n275,n276,n99);
nor (n276,n277,n278);
and (n277,n106,n58);
and (n278,n60,n107);
or (n279,n97,n115);
xor (n280,n281,n294);
xor (n281,n282,n288);
nand (n282,n283,n284);
or (n283,n146,n165);
or (n284,n147,n285);
nor (n285,n286,n287);
and (n286,n156,n208);
and (n287,n157,n210);
nand (n288,n289,n290);
or (n289,n122,n139);
or (n290,n123,n291);
nor (n291,n292,n293);
and (n292,n130,n111);
and (n293,n131,n113);
nand (n294,n295,n313);
or (n295,n296,n308);
nand (n296,n297,n303);
not (n297,n298);
nor (n298,n299,n302);
and (n299,n79,n300);
not (n300,n301);
and (n302,n80,n301);
nand (n303,n304,n307);
or (n304,n301,n305);
not (n305,n306);
nand (n307,n301,n305);
nor (n308,n309,n311);
and (n309,n305,n310);
and (n311,n306,n312);
not (n312,n310);
or (n313,n297,n314);
nor (n314,n315,n316);
and (n315,n305,n84);
and (n316,n306,n86);
xor (n317,n318,n575);
xor (n318,n319,n454);
xor (n319,n320,n381);
xor (n320,n321,n359);
xor (n321,n322,n351);
xor (n322,n323,n329);
nand (n323,n324,n325);
or (n324,n219,n234);
or (n325,n220,n326);
nor (n326,n327,n328);
and (n327,n74,n161);
and (n328,n75,n163);
nand (n329,n330,n345);
or (n330,n331,n340);
nand (n331,n332,n337);
or (n332,n333,n336);
and (n333,n334,n305);
not (n334,n335);
and (n336,n335,n306);
nand (n337,n338,n339);
or (n338,n335,n21);
nand (n339,n21,n335);
nor (n340,n341,n343);
and (n341,n21,n342);
and (n343,n22,n344);
not (n344,n342);
or (n345,n332,n346);
nor (n346,n347,n349);
and (n347,n21,n348);
and (n349,n22,n350);
not (n350,n348);
nand (n351,n352,n353);
or (n352,n18,n37);
or (n353,n19,n354);
nor (n354,n355,n357);
and (n355,n28,n356);
and (n357,n29,n358);
not (n358,n356);
or (n359,n360,n380);
and (n360,n361,n374);
xor (n361,n362,n368);
nand (n362,n363,n367);
or (n363,n296,n364);
nor (n364,n365,n366);
and (n365,n305,n348);
and (n366,n306,n350);
or (n367,n297,n308);
nand (n368,n369,n373);
or (n369,n331,n370);
nor (n370,n371,n372);
and (n371,n21,n356);
and (n372,n22,n358);
or (n373,n332,n340);
nand (n374,n375,n379);
or (n375,n197,n376);
nor (n376,n377,n378);
and (n377,n149,n167);
and (n378,n150,n169);
or (n379,n198,n206);
and (n380,n362,n368);
or (n381,n382,n453);
and (n382,n383,n429);
xor (n383,n384,n407);
or (n384,n385,n406);
and (n385,n386,n400);
xor (n386,n387,n394);
nand (n387,n388,n393);
or (n388,n389,n390);
not (n389,n174);
nor (n390,n391,n392);
and (n391,n179,n214);
and (n392,n180,n216);
or (n393,n183,n190);
nand (n394,n395,n399);
or (n395,n146,n396);
nor (n396,n397,n398);
and (n397,n156,n236);
and (n398,n157,n238);
or (n399,n147,n159);
nand (n400,n401,n405);
or (n401,n296,n402);
nor (n402,n403,n404);
and (n403,n305,n342);
and (n404,n306,n344);
or (n405,n297,n364);
and (n406,n387,n394);
or (n407,n408,n428);
and (n408,n409,n422);
xor (n409,n410,n416);
nand (n410,n411,n415);
or (n411,n219,n412);
nor (n412,n413,n414);
and (n413,n74,n90);
and (n414,n75,n92);
or (n415,n220,n228);
nand (n416,n417,n421);
or (n417,n18,n418);
nor (n418,n419,n420);
and (n419,n28,n64);
and (n420,n29,n66);
or (n421,n19,n31);
nand (n422,n423,n424);
or (n423,n56,n45);
or (n424,n44,n425);
nor (n425,n426,n427);
and (n426,n53,n117);
and (n427,n54,n119);
and (n428,n410,n416);
or (n429,n430,n452);
and (n430,n431,n444);
xor (n431,n432,n438);
nand (n432,n433,n437);
or (n433,n69,n434);
nor (n434,n435,n436);
and (n435,n79,n310);
and (n436,n80,n312);
or (n437,n70,n82);
nand (n438,n439,n443);
or (n439,n97,n440);
nor (n440,n441,n442);
and (n441,n106,n141);
and (n442,n143,n107);
or (n443,n99,n109);
nand (n444,n445,n451);
or (n445,n122,n446);
nor (n446,n447,n449);
and (n447,n448,n130);
and (n449,n450,n131);
not (n450,n448);
or (n451,n123,n133);
and (n452,n432,n438);
and (n453,n384,n407);
or (n454,n455,n574);
and (n455,n456,n544);
xor (n456,n457,n458);
xor (n457,n361,n374);
or (n458,n459,n543);
and (n459,n460,n518);
xor (n460,n461,n485);
or (n461,n462,n484);
and (n462,n463,n478);
xor (n463,n464,n470);
nand (n464,n465,n469);
or (n465,n69,n466);
nor (n466,n467,n468);
and (n467,n79,n348);
and (n468,n80,n350);
or (n469,n70,n434);
nand (n470,n471,n477);
or (n471,n122,n472);
nor (n472,n473,n475);
and (n473,n474,n130);
and (n475,n476,n131);
not (n476,n474);
or (n477,n446,n123);
nand (n478,n479,n483);
or (n479,n480,n296);
nor (n480,n481,n482);
and (n481,n305,n356);
and (n482,n306,n358);
or (n483,n297,n402);
and (n484,n464,n470);
or (n485,n486,n517);
and (n486,n487,n511);
xor (n487,n488,n505);
nand (n488,n489,n501);
or (n489,n490,n491);
nor (n490,n491,n497);
nand (n491,n492,n496);
or (n492,n493,n494);
not (n494,n495);
nand (n496,n493,n494);
nor (n497,n498,n499);
and (n498,n188,n493);
and (n499,n185,n500);
not (n500,n493);
not (n501,n502);
nor (n502,n503,n504);
and (n503,n188,n192);
and (n504,n185,n194);
nand (n505,n506,n510);
or (n506,n389,n507);
nor (n507,n508,n509);
and (n508,n179,n208);
and (n509,n180,n210);
or (n510,n183,n390);
nand (n511,n512,n516);
or (n512,n146,n513);
nor (n513,n514,n515);
and (n514,n156,n230);
and (n515,n157,n232);
or (n516,n147,n396);
and (n517,n488,n505);
or (n518,n519,n542);
and (n519,n520,n536);
xor (n520,n521,n530);
nand (n521,n522,n526);
or (n522,n331,n523);
nor (n523,n524,n525);
and (n524,n21,n33);
and (n525,n22,n35);
or (n526,n332,n527);
nor (n527,n528,n529);
and (n528,n21,n39);
and (n529,n22,n41);
nand (n530,n531,n535);
or (n531,n18,n532);
nor (n532,n533,n534);
and (n533,n28,n58);
and (n534,n29,n60);
or (n535,n19,n418);
nand (n536,n537,n541);
or (n537,n538,n219);
nor (n538,n539,n540);
and (n539,n74,n84);
and (n540,n75,n86);
or (n541,n220,n412);
and (n542,n521,n530);
and (n543,n461,n485);
or (n544,n545,n573);
and (n545,n546,n551);
xor (n546,n547,n550);
nand (n547,n548,n549);
or (n548,n331,n527);
or (n549,n332,n370);
not (n550,n374);
or (n551,n552,n572);
and (n552,n553,n566);
xor (n553,n554,n560);
nand (n554,n555,n559);
or (n555,n44,n556);
nor (n556,n557,n558);
and (n557,n53,n111);
and (n558,n54,n113);
or (n559,n45,n425);
nand (n560,n561,n565);
or (n561,n97,n562);
nor (n562,n563,n564);
and (n563,n106,n135);
and (n564,n137,n107);
or (n565,n99,n440);
nand (n566,n567,n571);
or (n567,n197,n568);
nor (n568,n569,n570);
and (n569,n149,n161);
and (n570,n150,n163);
or (n571,n198,n376);
and (n572,n554,n560);
and (n573,n547,n550);
and (n574,n457,n458);
or (n575,n576,n587);
and (n576,n577,n586);
xor (n577,n578,n579);
xor (n578,n383,n429);
or (n579,n580,n585);
and (n580,n581,n584);
xor (n581,n582,n583);
xor (n582,n386,n400);
xor (n583,n431,n444);
xor (n584,n409,n422);
and (n585,n582,n583);
xor (n586,n13,n170);
and (n587,n578,n579);
or (n588,n589,n657);
and (n589,n590,n656);
xor (n590,n591,n592);
xor (n591,n456,n544);
or (n592,n593,n655);
and (n593,n594,n654);
xor (n594,n595,n653);
or (n595,n596,n652);
and (n596,n597,n630);
xor (n597,n598,n604);
nand (n598,n599,n603);
or (n599,n389,n600);
nor (n600,n601,n602);
and (n601,n179,n167);
and (n602,n180,n169);
or (n603,n183,n507);
or (n604,n605,n629);
and (n605,n606,n621);
xor (n606,n607,n615);
nand (n607,n608,n613);
or (n608,n609,n610);
not (n609,n490);
nor (n610,n611,n612);
and (n611,n188,n214);
and (n612,n185,n216);
or (n613,n614,n502);
not (n614,n491);
nand (n615,n616,n620);
or (n616,n197,n617);
nor (n617,n618,n619);
and (n618,n149,n236);
and (n619,n150,n238);
or (n620,n198,n568);
nand (n621,n622,n628);
or (n622,n122,n623);
nor (n623,n624,n626);
and (n624,n625,n130);
and (n626,n627,n131);
not (n627,n625);
or (n628,n123,n472);
and (n629,n607,n615);
or (n630,n631,n651);
and (n631,n632,n645);
xor (n632,n633,n639);
nand (n633,n634,n638);
or (n634,n146,n635);
nor (n635,n636,n637);
and (n636,n156,n90);
and (n637,n157,n92);
or (n638,n147,n513);
nand (n639,n640,n644);
or (n640,n331,n641);
nor (n641,n642,n643);
and (n642,n21,n64);
and (n643,n22,n66);
or (n644,n332,n523);
nand (n645,n646,n650);
or (n646,n18,n647);
nor (n647,n648,n649);
and (n648,n28,n117);
and (n649,n29,n119);
or (n650,n19,n532);
and (n651,n633,n639);
and (n652,n598,n604);
xor (n653,n546,n551);
xor (n654,n460,n518);
and (n655,n595,n653);
xor (n656,n577,n586);
and (n657,n591,n592);
and (n658,n9,n317);
xor (n659,n660,n757);
xor (n660,n661,n697);
xor (n661,n662,n669);
xor (n662,n663,n666);
or (n663,n664,n665);
and (n664,n241,n252);
and (n665,n242,n249);
or (n666,n667,n668);
and (n667,n256,n280);
and (n668,n257,n260);
xor (n669,n670,n677);
xor (n670,n671,n674);
or (n671,n672,n673);
and (n672,n281,n294);
and (n673,n282,n288);
or (n674,n675,n676);
and (n675,n322,n351);
and (n676,n323,n329);
xor (n677,n678,n691);
xor (n678,n679,n685);
nand (n679,n680,n681);
or (n680,n122,n291);
or (n681,n123,n682);
nor (n682,n683,n684);
and (n683,n130,n117);
and (n684,n131,n119);
nand (n685,n686,n687);
or (n686,n219,n326);
or (n687,n220,n688);
nor (n688,n689,n690);
and (n689,n74,n167);
and (n690,n75,n169);
nand (n691,n692,n693);
or (n692,n331,n346);
or (n693,n332,n694);
nor (n694,n695,n696);
and (n695,n21,n310);
and (n696,n22,n312);
xor (n697,n698,n754);
xor (n698,n699,n751);
xor (n699,n700,n740);
xor (n700,n701,n720);
xor (n701,n702,n714);
xor (n702,n703,n708);
nand (n703,n704,n707);
or (n704,n705,n706);
not (n705,n197);
not (n706,n198);
not (n707,n246);
nand (n708,n709,n710);
or (n709,n146,n285);
or (n710,n147,n711);
nor (n711,n712,n713);
and (n712,n156,n214);
and (n713,n157,n216);
nand (n714,n715,n716);
or (n715,n69,n265);
or (n716,n70,n717);
nor (n717,n718,n719);
and (n718,n79,n236);
and (n719,n80,n238);
xor (n720,n721,n734);
xor (n721,n722,n728);
nand (n722,n723,n724);
or (n723,n44,n271);
or (n724,n45,n725);
nor (n725,n726,n727);
and (n726,n53,n39);
and (n727,n54,n41);
nand (n728,n729,n730);
or (n729,n97,n276);
or (n730,n99,n731);
nor (n731,n732,n733);
and (n732,n106,n64);
and (n733,n107,n66);
nand (n734,n735,n736);
or (n735,n296,n314);
or (n736,n297,n737);
nor (n737,n738,n739);
and (n738,n305,n90);
and (n739,n306,n92);
xor (n740,n741,n748);
xor (n741,n742,n243);
nand (n742,n743,n744);
or (n743,n18,n354);
or (n744,n19,n745);
nor (n745,n746,n747);
and (n746,n28,n342);
and (n747,n29,n344);
or (n748,n749,n750);
and (n749,n261,n274);
and (n750,n262,n268);
or (n751,n752,n753);
and (n752,n320,n381);
and (n753,n321,n359);
or (n754,n755,n756);
and (n755,n10,n255);
and (n756,n11,n240);
or (n757,n758,n759);
and (n758,n318,n575);
and (n759,n319,n454);
nand (n760,n6,n659);
not (n761,n762);
nor (n762,n763,n5119);
nor (n763,n764,n3863);
nor (n764,n765,n3851);
nand (n765,n766,n2659);
or (n766,n767,n1976);
not (n767,n768);
nand (n768,n769,n1975);
or (n769,n770,n1604);
nor (n770,n771,n1466);
xor (n771,n772,n1408);
xor (n772,n773,n1086);
xor (n773,n774,n1005);
xor (n774,n775,n913);
or (n775,n776,n912);
and (n776,n777,n849);
xor (n777,n778,n810);
xor (n778,n779,n800);
xor (n779,n780,n791);
nand (n780,n781,n786);
or (n781,n782,n146);
not (n782,n783);
nor (n783,n784,n785);
and (n784,n137,n156);
and (n785,n135,n157);
nand (n786,n787,n790);
nor (n787,n788,n789);
and (n788,n143,n156);
and (n789,n141,n157);
not (n790,n147);
nand (n791,n792,n796);
or (n792,n793,n219);
nor (n793,n794,n795);
and (n794,n476,n75);
and (n795,n474,n74);
or (n796,n220,n797);
nor (n797,n798,n799);
and (n798,n450,n75);
and (n799,n448,n74);
nand (n800,n801,n806);
or (n801,n802,n614);
not (n802,n803);
nor (n803,n804,n805);
and (n804,n39,n185);
and (n805,n41,n188);
or (n806,n609,n807);
nor (n807,n808,n809);
and (n808,n188,n33);
and (n809,n185,n35);
xor (n810,n811,n835);
xor (n811,n812,n822);
nand (n812,n813,n817);
or (n813,n389,n814);
nor (n814,n815,n816);
and (n815,n179,n58);
and (n816,n180,n60);
or (n817,n183,n818);
not (n818,n819);
nor (n819,n820,n821);
and (n820,n64,n180);
and (n821,n66,n179);
nand (n822,n823,n829);
or (n823,n331,n824);
nor (n824,n825,n827);
and (n825,n21,n826);
and (n827,n22,n828);
not (n828,n826);
or (n829,n332,n830);
nor (n830,n831,n833);
and (n831,n21,n832);
and (n833,n834,n22);
not (n834,n832);
nand (n835,n836,n842);
or (n836,n18,n837);
nor (n837,n838,n840);
and (n838,n28,n839);
and (n840,n29,n841);
not (n841,n839);
or (n842,n19,n843);
not (n843,n844);
nand (n844,n845,n848);
or (n845,n29,n846);
not (n846,n847);
or (n848,n28,n847);
xor (n849,n850,n883);
xor (n850,n851,n874);
nand (n851,n852,n869);
or (n852,n853,n866);
not (n853,n854);
nor (n854,n855,n861);
nand (n855,n856,n860);
or (n856,n857,n859);
not (n857,n858);
nand (n860,n859,n857);
nor (n861,n862,n865);
and (n862,n863,n858);
not (n863,n864);
and (n865,n864,n857);
nor (n866,n867,n868);
and (n867,n863,n348);
and (n868,n864,n350);
or (n869,n870,n871);
not (n870,n855);
nor (n871,n872,n873);
and (n872,n863,n310);
and (n873,n864,n312);
nand (n874,n875,n879);
or (n875,n197,n876);
nor (n876,n877,n878);
and (n877,n149,n111);
and (n878,n150,n113);
or (n879,n198,n880);
nor (n880,n881,n882);
and (n881,n149,n117);
and (n882,n150,n119);
and (n883,n884,n891);
and (n884,n885,n29);
nand (n885,n886,n888);
or (n886,n887,n23);
nand (n888,n889,n21);
not (n889,n890);
and (n890,n887,n23);
nand (n891,n892,n908);
or (n892,n893,n905);
nand (n893,n894,n901);
nor (n894,n895,n899);
and (n895,n896,n898);
not (n896,n897);
and (n899,n897,n900);
not (n900,n898);
nand (n901,n902,n904);
or (n902,n898,n903);
not (n903,n859);
nand (n904,n903,n898);
nor (n905,n906,n907);
and (n906,n903,n310);
and (n907,n859,n312);
or (n908,n894,n909);
nor (n909,n910,n911);
and (n910,n903,n84);
and (n911,n859,n86);
and (n912,n778,n810);
xor (n913,n914,n977);
xor (n914,n915,n941);
xor (n915,n916,n931);
xor (n916,n917,n924);
nand (n917,n918,n919);
or (n918,n843,n18);
nand (n919,n920,n923);
nor (n920,n921,n922);
and (n921,n28,n828);
and (n922,n29,n826);
not (n923,n19);
nand (n924,n925,n926);
or (n925,n871,n853);
nand (n926,n927,n855);
not (n927,n928);
nor (n928,n929,n930);
and (n929,n86,n864);
and (n930,n84,n863);
nand (n931,n932,n937);
or (n932,n44,n933);
nor (n933,n934,n936);
and (n934,n935,n54);
not (n935,n887);
and (n936,n887,n53);
or (n937,n938,n45);
nor (n938,n939,n940);
and (n939,n53,n839);
and (n940,n841,n54);
xor (n941,n942,n971);
xor (n942,n943,n964);
nand (n943,n944,n958);
or (n944,n945,n949);
not (n945,n946);
nor (n946,n947,n948);
and (n947,n342,n495);
and (n948,n344,n494);
nand (n949,n950,n955);
nor (n950,n951,n953);
and (n951,n863,n952);
and (n953,n864,n954);
not (n954,n952);
nand (n955,n956,n957);
or (n956,n952,n494);
nand (n957,n494,n952);
nand (n958,n959,n963);
not (n959,n960);
nor (n960,n961,n962);
and (n961,n350,n495);
and (n962,n348,n494);
not (n963,n950);
nand (n964,n965,n967);
or (n965,n966,n146);
not (n966,n787);
nand (n967,n790,n968);
nand (n968,n969,n970);
or (n969,n157,n113);
or (n970,n156,n111);
nand (n971,n972,n973);
or (n972,n219,n797);
or (n973,n220,n974);
nor (n974,n975,n976);
and (n975,n74,n135);
and (n976,n75,n137);
xor (n977,n978,n997);
xor (n978,n979,n991);
nand (n979,n980,n987);
or (n980,n981,n984);
nand (n981,n897,n982);
not (n982,n983);
nor (n984,n985,n986);
and (n985,n238,n897);
and (n986,n236,n896);
or (n987,n988,n982);
nor (n988,n989,n990);
and (n989,n896,n161);
and (n990,n897,n163);
nand (n991,n992,n993);
or (n992,n818,n389);
nand (n993,n182,n994);
nand (n994,n995,n996);
or (n995,n180,n35);
or (n996,n179,n33);
nand (n997,n998,n999);
or (n998,n331,n830);
or (n999,n332,n1000);
nor (n1000,n1001,n1003);
and (n1001,n21,n1002);
and (n1003,n22,n1004);
not (n1004,n1002);
xor (n1005,n1006,n1042);
xor (n1006,n1007,n1039);
xor (n1007,n1008,n1026);
xor (n1008,n1009,n1016);
nand (n1009,n1010,n1011);
or (n1010,n802,n609);
nand (n1011,n1012,n491);
not (n1012,n1013);
nor (n1013,n1014,n1015);
and (n1014,n188,n356);
and (n1015,n185,n358);
nand (n1016,n1017,n1022);
or (n1017,n1018,n69);
not (n1018,n1019);
nor (n1019,n1020,n1021);
and (n1020,n627,n79);
and (n1021,n625,n80);
nand (n1022,n71,n1023);
nand (n1023,n1024,n1025);
or (n1024,n80,n476);
or (n1025,n79,n474);
nand (n1026,n1027,n1033);
or (n1027,n296,n1028);
nor (n1028,n1029,n1031);
and (n1029,n305,n1030);
and (n1031,n306,n1032);
not (n1032,n1030);
or (n1033,n297,n1034);
nor (n1034,n1035,n1038);
and (n1035,n1036,n306);
not (n1036,n1037);
and (n1038,n1037,n305);
or (n1039,n1040,n1041);
and (n1040,n850,n883);
and (n1041,n851,n874);
xor (n1042,n1043,n1072);
xor (n1043,n1044,n1050);
nand (n1044,n1045,n1046);
or (n1045,n197,n880);
or (n1046,n198,n1047);
nor (n1047,n1048,n1049);
and (n1048,n149,n58);
and (n1049,n150,n60);
nand (n1050,n1051,n1071);
or (n1051,n1052,n1059);
not (n1052,n1053);
nand (n1053,n1054,n54);
nand (n1054,n1055,n1056);
or (n1055,n887,n49);
nand (n1056,n1057,n28);
not (n1057,n1058);
and (n1058,n887,n49);
not (n1059,n1060);
nand (n1060,n1061,n1066);
or (n1061,n1062,n893);
not (n1062,n1063);
nand (n1063,n1064,n1065);
or (n1064,n859,n92);
or (n1065,n903,n90);
nand (n1066,n1067,n1068);
not (n1067,n894);
nor (n1068,n1069,n1070);
and (n1069,n230,n859);
and (n1070,n232,n903);
nand (n1071,n1059,n1052);
or (n1072,n1073,n1085);
and (n1073,n1074,n1079);
xor (n1074,n1075,n1076);
nor (n1075,n45,n935);
nand (n1076,n1077,n1078);
or (n1077,n909,n893);
nand (n1078,n1067,n1063);
nand (n1079,n1080,n1084);
or (n1080,n949,n1081);
nor (n1081,n1082,n1083);
and (n1082,n494,n356);
and (n1083,n495,n358);
or (n1084,n950,n945);
and (n1085,n1075,n1076);
or (n1086,n1087,n1407);
and (n1087,n1088,n1346);
xor (n1088,n1089,n1283);
or (n1089,n1090,n1282);
and (n1090,n1091,n1225);
xor (n1091,n1092,n1156);
or (n1092,n1093,n1155);
and (n1093,n1094,n1121);
xor (n1094,n1095,n1104);
nand (n1095,n1096,n1100);
or (n1096,n197,n1097);
nor (n1097,n1098,n1099);
and (n1098,n149,n135);
and (n1099,n150,n137);
or (n1100,n198,n1101);
nor (n1101,n1102,n1103);
and (n1102,n149,n141);
and (n1103,n150,n143);
and (n1104,n1105,n1111);
and (n1105,n1106,n22);
nand (n1106,n1107,n1108);
or (n1107,n887,n335);
nand (n1108,n1109,n305);
not (n1109,n1110);
and (n1110,n887,n335);
nand (n1111,n1112,n1117);
or (n1112,n1113,n893);
not (n1113,n1114);
nor (n1114,n1115,n1116);
and (n1115,n342,n859);
and (n1116,n344,n903);
nand (n1117,n1067,n1118);
nand (n1118,n1119,n1120);
or (n1119,n859,n350);
or (n1120,n903,n348);
or (n1121,n1122,n1154);
and (n1122,n1123,n1144);
xor (n1123,n1124,n1134);
nand (n1124,n1125,n1129);
or (n1125,n1126,n609);
nor (n1126,n1127,n1128);
and (n1127,n188,n117);
and (n1128,n185,n119);
nand (n1129,n1130,n491);
not (n1130,n1131);
nor (n1131,n1132,n1133);
and (n1132,n188,n58);
and (n1133,n185,n60);
nand (n1134,n1135,n1140);
or (n1135,n69,n1136);
not (n1136,n1137);
nor (n1137,n1138,n1139);
and (n1138,n834,n79);
and (n1139,n832,n80);
or (n1140,n70,n1141);
nor (n1141,n1142,n1143);
and (n1142,n79,n1002);
and (n1143,n80,n1004);
nand (n1144,n1145,n1149);
or (n1145,n296,n1146);
nor (n1146,n1147,n1148);
and (n1147,n847,n305);
and (n1148,n846,n306);
or (n1149,n297,n1150);
not (n1150,n1151);
nand (n1151,n1152,n1153);
or (n1152,n306,n828);
or (n1153,n305,n826);
and (n1154,n1124,n1134);
and (n1155,n1095,n1104);
xor (n1156,n1157,n1211);
xor (n1157,n1158,n1191);
or (n1158,n1159,n1190);
and (n1159,n1160,n1181);
xor (n1160,n1161,n1172);
nand (n1161,n1162,n1167);
or (n1162,n1163,n853);
not (n1163,n1164);
nor (n1164,n1165,n1166);
and (n1165,n356,n864);
and (n1166,n358,n863);
nand (n1167,n1168,n855);
not (n1168,n1169);
nor (n1169,n1170,n1171);
and (n1170,n863,n342);
and (n1171,n864,n344);
nand (n1172,n1173,n1177);
or (n1173,n1174,n331);
nor (n1174,n1175,n1176);
and (n1175,n21,n839);
and (n1176,n22,n841);
or (n1177,n332,n1178);
nor (n1178,n1179,n1180);
and (n1179,n21,n847);
and (n1180,n22,n846);
nand (n1181,n1182,n1186);
or (n1182,n389,n1183);
nor (n1183,n1184,n1185);
and (n1184,n179,n111);
and (n1185,n180,n113);
or (n1186,n183,n1187);
nor (n1187,n1188,n1189);
and (n1188,n179,n117);
and (n1189,n180,n119);
and (n1190,n1161,n1172);
or (n1191,n1192,n1210);
and (n1192,n1193,n1200);
xor (n1193,n1194,n1195);
nor (n1194,n19,n935);
nand (n1195,n1196,n1198);
or (n1196,n1197,n893);
not (n1197,n1118);
nand (n1198,n1199,n1067);
not (n1199,n905);
nand (n1200,n1201,n1205);
or (n1201,n949,n1202);
nor (n1202,n1203,n1204);
and (n1203,n35,n495);
and (n1204,n33,n494);
or (n1205,n950,n1206);
not (n1206,n1207);
nand (n1207,n1208,n1209);
or (n1208,n495,n41);
or (n1209,n494,n39);
and (n1210,n1194,n1195);
xor (n1211,n1212,n1222);
xor (n1212,n1213,n1219);
nand (n1213,n1214,n1218);
or (n1214,n18,n1215);
nor (n1215,n1216,n1217);
and (n1216,n935,n29);
and (n1217,n887,n28);
or (n1218,n837,n19);
nand (n1219,n1220,n1221);
or (n1220,n853,n1169);
or (n1221,n870,n866);
nand (n1222,n1223,n1224);
or (n1223,n197,n1101);
or (n1224,n198,n876);
or (n1225,n1226,n1281);
and (n1226,n1227,n1255);
xor (n1227,n1228,n1254);
xor (n1228,n1229,n1244);
xor (n1229,n1230,n1237);
nand (n1230,n1231,n1232);
or (n1231,n1141,n69);
nand (n1232,n1233,n71);
not (n1233,n1234);
nor (n1234,n1235,n1236);
and (n1235,n1032,n80);
and (n1236,n1030,n79);
nand (n1237,n1238,n1239);
or (n1238,n1150,n296);
nand (n1239,n1240,n298);
not (n1240,n1241);
nor (n1241,n1242,n1243);
and (n1242,n305,n832);
and (n1243,n306,n834);
nand (n1244,n1245,n1250);
or (n1245,n1246,n981);
not (n1246,n1247);
nor (n1247,n1248,n1249);
and (n1248,n84,n897);
and (n1249,n86,n896);
or (n1250,n1251,n982);
nor (n1251,n1252,n1253);
and (n1252,n896,n90);
and (n1253,n897,n92);
xor (n1254,n1193,n1200);
xor (n1255,n1256,n1275);
xor (n1256,n1257,n1266);
nand (n1257,n1258,n1262);
or (n1258,n146,n1259);
nor (n1259,n1260,n1261);
and (n1260,n476,n157);
and (n1261,n474,n156);
or (n1262,n147,n1263);
nor (n1263,n1264,n1265);
and (n1264,n450,n157);
and (n1265,n448,n156);
nand (n1266,n1267,n1271);
or (n1267,n219,n1268);
nor (n1268,n1269,n1270);
and (n1269,n74,n1037);
and (n1270,n75,n1036);
or (n1271,n220,n1272);
nor (n1272,n1273,n1274);
and (n1273,n74,n625);
and (n1274,n75,n627);
nand (n1275,n1276,n1277);
or (n1276,n609,n1131);
or (n1277,n614,n1278);
nor (n1278,n1279,n1280);
and (n1279,n188,n64);
and (n1280,n185,n66);
and (n1281,n1228,n1254);
and (n1282,n1092,n1156);
xor (n1283,n1284,n1299);
xor (n1284,n1285,n1296);
or (n1285,n1286,n1295);
and (n1286,n1287,n1292);
xor (n1287,n1288,n1289);
xor (n1288,n884,n891);
or (n1289,n1290,n1291);
and (n1290,n1256,n1275);
and (n1291,n1257,n1266);
or (n1292,n1293,n1294);
and (n1293,n1229,n1244);
and (n1294,n1230,n1237);
and (n1295,n1288,n1289);
or (n1296,n1297,n1298);
and (n1297,n1157,n1211);
and (n1298,n1158,n1191);
or (n1299,n1300,n1345);
and (n1300,n1301,n1331);
xor (n1301,n1302,n1314);
xor (n1302,n1303,n1311);
xor (n1303,n1304,n1308);
nand (n1304,n1305,n1306);
or (n1305,n1206,n949);
nand (n1306,n1307,n963);
not (n1307,n1081);
nand (n1308,n1309,n1310);
or (n1309,n1263,n146);
nand (n1310,n790,n783);
nand (n1311,n1312,n1313);
or (n1312,n219,n1272);
or (n1313,n220,n793);
xor (n1314,n1315,n1325);
xor (n1315,n1316,n1319);
nand (n1316,n1317,n1318);
or (n1317,n609,n1278);
or (n1318,n614,n807);
nand (n1319,n1320,n1321);
or (n1320,n69,n1234);
or (n1321,n70,n1322);
nor (n1322,n1323,n1324);
and (n1323,n1036,n80);
and (n1324,n1037,n79);
nand (n1325,n1326,n1327);
or (n1326,n296,n1241);
or (n1327,n297,n1328);
nor (n1328,n1329,n1330);
and (n1329,n1004,n306);
and (n1330,n1002,n305);
xor (n1331,n1332,n1342);
xor (n1332,n1333,n1339);
nand (n1333,n1334,n1335);
or (n1334,n981,n1251);
or (n1335,n1336,n982);
nor (n1336,n1337,n1338);
and (n1337,n896,n230);
and (n1338,n897,n232);
nand (n1339,n1340,n1341);
or (n1340,n389,n1187);
or (n1341,n183,n814);
nand (n1342,n1343,n1344);
or (n1343,n331,n1178);
or (n1344,n332,n824);
and (n1345,n1302,n1314);
or (n1346,n1347,n1406);
and (n1347,n1348,n1405);
xor (n1348,n1349,n1404);
or (n1349,n1350,n1403);
and (n1350,n1351,n1402);
xor (n1351,n1352,n1377);
or (n1352,n1353,n1376);
and (n1353,n1354,n1369);
xor (n1354,n1355,n1362);
nand (n1355,n1356,n1357);
or (n1356,n982,n1246);
nand (n1357,n1358,n1361);
nand (n1358,n1359,n1360);
or (n1359,n312,n897);
nand (n1360,n897,n312);
not (n1361,n981);
nand (n1362,n1363,n1368);
or (n1363,n1364,n853);
not (n1364,n1365);
nor (n1365,n1366,n1367);
and (n1366,n39,n864);
and (n1367,n41,n863);
nand (n1368,n855,n1164);
nand (n1369,n1370,n1375);
or (n1370,n1371,n331);
not (n1371,n1372);
nand (n1372,n1373,n1374);
or (n1373,n887,n21);
or (n1374,n935,n22);
or (n1375,n332,n1174);
and (n1376,n1355,n1362);
or (n1377,n1378,n1401);
and (n1378,n1379,n1395);
xor (n1379,n1380,n1387);
nand (n1380,n1381,n1385);
or (n1381,n1382,n949);
nor (n1382,n1383,n1384);
and (n1383,n66,n495);
and (n1384,n64,n494);
nand (n1385,n1386,n963);
not (n1386,n1202);
nand (n1387,n1388,n1393);
or (n1388,n1389,n146);
not (n1389,n1390);
nor (n1390,n1391,n1392);
and (n1391,n625,n157);
and (n1392,n627,n156);
nand (n1393,n1394,n790);
not (n1394,n1259);
nand (n1395,n1396,n1400);
or (n1396,n219,n1397);
nor (n1397,n1398,n1399);
and (n1398,n74,n1030);
and (n1399,n75,n1032);
or (n1400,n220,n1268);
and (n1401,n1380,n1387);
xor (n1402,n1160,n1181);
and (n1403,n1352,n1377);
xor (n1404,n1287,n1292);
xor (n1405,n1301,n1331);
and (n1406,n1349,n1404);
and (n1407,n1089,n1283);
xor (n1408,n1409,n1447);
xor (n1409,n1410,n1413);
or (n1410,n1411,n1412);
and (n1411,n1284,n1299);
and (n1412,n1285,n1296);
or (n1413,n1414,n1446);
and (n1414,n1415,n1428);
xor (n1415,n1416,n1427);
xor (n1416,n1417,n1424);
xor (n1417,n1418,n1421);
or (n1418,n1419,n1420);
and (n1419,n1303,n1311);
and (n1420,n1304,n1308);
or (n1421,n1422,n1423);
and (n1422,n1315,n1325);
and (n1423,n1316,n1319);
or (n1424,n1425,n1426);
and (n1425,n1332,n1342);
and (n1426,n1333,n1339);
xor (n1427,n777,n849);
xor (n1428,n1429,n1434);
xor (n1429,n1430,n1433);
or (n1430,n1431,n1432);
and (n1431,n1212,n1222);
and (n1432,n1213,n1219);
xor (n1433,n1074,n1079);
xor (n1434,n1435,n1443);
xor (n1435,n1436,n1439);
nand (n1436,n1437,n1438);
or (n1437,n1018,n70);
or (n1438,n69,n1322);
nand (n1439,n1440,n1441);
or (n1440,n1328,n296);
nand (n1441,n1442,n298);
not (n1442,n1028);
nand (n1443,n1444,n1445);
or (n1444,n981,n1336);
or (n1445,n984,n982);
and (n1446,n1416,n1427);
xor (n1447,n1448,n1455);
xor (n1448,n1449,n1452);
or (n1449,n1450,n1451);
and (n1450,n1417,n1424);
and (n1451,n1418,n1421);
or (n1452,n1453,n1454);
and (n1453,n1429,n1434);
and (n1454,n1430,n1433);
xor (n1455,n1456,n1463);
xor (n1456,n1457,n1460);
or (n1457,n1458,n1459);
and (n1458,n779,n800);
and (n1459,n780,n791);
or (n1460,n1461,n1462);
and (n1461,n1435,n1443);
and (n1462,n1436,n1439);
or (n1463,n1464,n1465);
and (n1464,n811,n835);
and (n1465,n812,n822);
or (n1466,n1467,n1603);
and (n1467,n1468,n1602);
xor (n1468,n1469,n1470);
xor (n1469,n1415,n1428);
or (n1470,n1471,n1601);
and (n1471,n1472,n1600);
xor (n1472,n1473,n1565);
or (n1473,n1474,n1564);
and (n1474,n1475,n1563);
xor (n1475,n1476,n1494);
or (n1476,n1477,n1493);
and (n1477,n1478,n1492);
xor (n1478,n1479,n1485);
nand (n1479,n1480,n1484);
or (n1480,n389,n1481);
nor (n1481,n1482,n1483);
and (n1482,n179,n141);
and (n1483,n180,n143);
or (n1484,n183,n1183);
nand (n1485,n1486,n1490);
or (n1486,n1487,n197);
nor (n1487,n1488,n1489);
and (n1488,n149,n448);
and (n1489,n150,n450);
nand (n1490,n1491,n706);
not (n1491,n1097);
xor (n1492,n1105,n1111);
and (n1493,n1479,n1485);
or (n1494,n1495,n1562);
and (n1495,n1496,n1545);
xor (n1496,n1497,n1522);
or (n1497,n1498,n1521);
and (n1498,n1499,n1514);
xor (n1499,n1500,n1507);
nand (n1500,n1501,n1506);
or (n1501,n1502,n69);
not (n1502,n1503);
nor (n1503,n1504,n1505);
and (n1504,n828,n79);
and (n1505,n826,n80);
nand (n1506,n71,n1137);
nand (n1507,n1508,n1512);
or (n1508,n1509,n296);
nor (n1509,n1510,n1511);
and (n1510,n839,n305);
and (n1511,n841,n306);
nand (n1512,n1513,n298);
not (n1513,n1146);
nand (n1514,n1515,n1519);
or (n1515,n981,n1516);
nor (n1516,n1517,n1518);
and (n1517,n896,n348);
and (n1518,n897,n350);
or (n1519,n1520,n982);
not (n1520,n1358);
and (n1521,n1500,n1507);
or (n1522,n1523,n1544);
and (n1523,n1524,n1538);
xor (n1524,n1525,n1531);
nand (n1525,n1526,n1530);
or (n1526,n1527,n853);
nor (n1527,n1528,n1529);
and (n1528,n863,n33);
and (n1529,n864,n35);
nand (n1530,n855,n1365);
nand (n1531,n1532,n1533);
or (n1532,n183,n1481);
nand (n1533,n1534,n174);
not (n1534,n1535);
nor (n1535,n1536,n1537);
and (n1536,n137,n180);
and (n1537,n135,n179);
nand (n1538,n1539,n1543);
or (n1539,n197,n1540);
nor (n1540,n1541,n1542);
and (n1541,n149,n474);
and (n1542,n150,n476);
or (n1543,n198,n1487);
and (n1544,n1525,n1531);
or (n1545,n1546,n1561);
and (n1546,n1547,n1555);
xor (n1547,n1548,n1549);
nor (n1548,n332,n935);
nand (n1549,n1550,n1554);
or (n1550,n1551,n893);
nor (n1551,n1552,n1553);
and (n1552,n358,n859);
and (n1553,n356,n903);
nand (n1554,n1067,n1114);
nand (n1555,n1556,n1560);
or (n1556,n949,n1557);
nor (n1557,n1558,n1559);
and (n1558,n60,n495);
and (n1559,n58,n494);
or (n1560,n950,n1382);
and (n1561,n1548,n1549);
and (n1562,n1497,n1522);
xor (n1563,n1094,n1121);
and (n1564,n1476,n1494);
or (n1565,n1566,n1599);
and (n1566,n1567,n1598);
xor (n1567,n1568,n1569);
xor (n1568,n1351,n1402);
or (n1569,n1570,n1597);
and (n1570,n1571,n1596);
xor (n1571,n1572,n1595);
or (n1572,n1573,n1594);
and (n1573,n1574,n1588);
xor (n1574,n1575,n1582);
nand (n1575,n1576,n1581);
or (n1576,n1577,n146);
not (n1577,n1578);
nand (n1578,n1579,n1580);
or (n1579,n157,n1036);
or (n1580,n156,n1037);
nand (n1581,n1390,n790);
nand (n1582,n1583,n1587);
or (n1583,n1584,n219);
nor (n1584,n1585,n1586);
and (n1585,n74,n1002);
and (n1586,n75,n1004);
or (n1587,n1397,n220);
nand (n1588,n1589,n1593);
or (n1589,n609,n1590);
nor (n1590,n1591,n1592);
and (n1591,n188,n111);
and (n1592,n185,n113);
or (n1593,n614,n1126);
and (n1594,n1575,n1582);
xor (n1595,n1354,n1369);
xor (n1596,n1123,n1144);
and (n1597,n1572,n1595);
xor (n1598,n1227,n1255);
and (n1599,n1568,n1569);
xor (n1600,n1091,n1225);
and (n1601,n1473,n1565);
xor (n1602,n1088,n1346);
and (n1603,n1469,n1470);
not (n1604,n1605);
nand (n1605,n1606,n1974);
or (n1606,n1607,n1728);
not (n1607,n1608);
nand (n1608,n1609,n1611);
not (n1609,n1610);
xor (n1610,n1468,n1602);
not (n1611,n1612);
or (n1612,n1613,n1727);
and (n1613,n1614,n1726);
xor (n1614,n1615,n1616);
xor (n1615,n1348,n1405);
or (n1616,n1617,n1725);
and (n1617,n1618,n1689);
xor (n1618,n1619,n1688);
or (n1619,n1620,n1687);
and (n1620,n1621,n1624);
xor (n1621,n1622,n1623);
xor (n1622,n1379,n1395);
xor (n1623,n1478,n1492);
or (n1624,n1625,n1686);
and (n1625,n1626,n1663);
xor (n1626,n1627,n1640);
and (n1627,n1628,n1634);
and (n1628,n1629,n306);
nand (n1629,n1630,n1631);
or (n1630,n887,n301);
nand (n1631,n1632,n79);
not (n1632,n1633);
and (n1633,n887,n301);
nand (n1634,n1635,n1639);
or (n1635,n893,n1636);
nor (n1636,n1637,n1638);
and (n1637,n903,n39);
and (n1638,n859,n41);
or (n1639,n894,n1551);
or (n1640,n1641,n1662);
and (n1641,n1642,n1656);
xor (n1642,n1643,n1650);
nand (n1643,n1644,n1649);
or (n1644,n981,n1645);
not (n1645,n1646);
nor (n1646,n1647,n1648);
and (n1647,n344,n896);
and (n1648,n342,n897);
or (n1649,n1516,n982);
nand (n1650,n1651,n1655);
or (n1651,n853,n1652);
nor (n1652,n1653,n1654);
and (n1653,n863,n64);
and (n1654,n864,n66);
or (n1655,n870,n1527);
nand (n1656,n1657,n1661);
or (n1657,n389,n1658);
nor (n1658,n1659,n1660);
and (n1659,n179,n448);
and (n1660,n180,n450);
or (n1661,n183,n1535);
and (n1662,n1643,n1650);
or (n1663,n1664,n1685);
and (n1664,n1665,n1679);
xor (n1665,n1666,n1672);
nand (n1666,n1667,n1671);
or (n1667,n609,n1668);
nor (n1668,n1669,n1670);
and (n1669,n188,n141);
and (n1670,n185,n143);
or (n1671,n614,n1590);
nand (n1672,n1673,n1678);
or (n1673,n69,n1674);
not (n1674,n1675);
nand (n1675,n1676,n1677);
or (n1676,n80,n846);
or (n1677,n79,n847);
or (n1678,n70,n1502);
nand (n1679,n1680,n1684);
or (n1680,n296,n1681);
nor (n1681,n1682,n1683);
and (n1682,n935,n306);
and (n1683,n305,n887);
or (n1684,n297,n1509);
and (n1685,n1666,n1672);
and (n1686,n1627,n1640);
and (n1687,n1622,n1623);
xor (n1688,n1475,n1563);
or (n1689,n1690,n1724);
and (n1690,n1691,n1723);
xor (n1691,n1692,n1693);
xor (n1692,n1496,n1545);
or (n1693,n1694,n1722);
and (n1694,n1695,n1721);
xor (n1695,n1696,n1720);
or (n1696,n1697,n1719);
and (n1697,n1698,n1713);
xor (n1698,n1699,n1706);
nand (n1699,n1700,n1704);
or (n1700,n1701,n949);
nor (n1701,n1702,n1703);
and (n1702,n117,n494);
and (n1703,n119,n495);
nand (n1704,n1705,n963);
not (n1705,n1557);
nand (n1706,n1707,n1708);
or (n1707,n1577,n147);
nand (n1708,n1709,n1710);
not (n1709,n146);
nor (n1710,n1711,n1712);
and (n1711,n1030,n157);
and (n1712,n1032,n156);
nand (n1713,n1714,n1718);
or (n1714,n219,n1715);
nor (n1715,n1716,n1717);
and (n1716,n74,n832);
and (n1717,n75,n834);
or (n1718,n220,n1584);
and (n1719,n1699,n1706);
xor (n1720,n1524,n1538);
xor (n1721,n1574,n1588);
and (n1722,n1696,n1720);
xor (n1723,n1571,n1596);
and (n1724,n1692,n1693);
and (n1725,n1619,n1688);
xor (n1726,n1472,n1600);
and (n1727,n1615,n1616);
not (n1728,n1729);
nand (n1729,n1730,n1973);
or (n1730,n1731,n1789);
nor (n1731,n1732,n1788);
or (n1732,n1733,n1787);
and (n1733,n1734,n1737);
xor (n1734,n1735,n1736);
xor (n1735,n1567,n1598);
xor (n1736,n1618,n1689);
or (n1737,n1738,n1786);
and (n1738,n1739,n1785);
xor (n1739,n1740,n1741);
xor (n1740,n1621,n1624);
or (n1741,n1742,n1784);
and (n1742,n1743,n1746);
xor (n1743,n1744,n1745);
xor (n1744,n1499,n1514);
xor (n1745,n1547,n1555);
or (n1746,n1747,n1783);
and (n1747,n1748,n1756);
xor (n1748,n1749,n1755);
nand (n1749,n1750,n1754);
or (n1750,n197,n1751);
nor (n1751,n1752,n1753);
and (n1752,n149,n625);
and (n1753,n150,n627);
or (n1754,n198,n1540);
xor (n1755,n1628,n1634);
or (n1756,n1757,n1782);
and (n1757,n1758,n1774);
xor (n1758,n1759,n1766);
nand (n1759,n1760,n1765);
or (n1760,n1761,n146);
not (n1761,n1762);
nor (n1762,n1763,n1764);
and (n1763,n1004,n156);
and (n1764,n1002,n157);
nand (n1765,n790,n1710);
nand (n1766,n1767,n1771);
or (n1767,n1768,n219);
nor (n1768,n1769,n1770);
and (n1769,n826,n74);
and (n1770,n75,n828);
nand (n1771,n1772,n1773);
not (n1772,n1715);
not (n1773,n220);
nand (n1774,n1775,n1780);
or (n1775,n1776,n893);
not (n1776,n1777);
nand (n1777,n1778,n1779);
or (n1778,n859,n35);
or (n1779,n903,n33);
nand (n1780,n1781,n1067);
not (n1781,n1636);
and (n1782,n1759,n1766);
and (n1783,n1749,n1755);
and (n1784,n1744,n1745);
xor (n1785,n1691,n1723);
and (n1786,n1740,n1741);
and (n1787,n1735,n1736);
xor (n1788,n1614,n1726);
nand (n1789,n1790,n1791);
xor (n1790,n1734,n1737);
or (n1791,n1792,n1972);
and (n1792,n1793,n1971);
xor (n1793,n1794,n1884);
or (n1794,n1795,n1883);
and (n1795,n1796,n1846);
xor (n1796,n1797,n1845);
or (n1797,n1798,n1844);
and (n1798,n1799,n1843);
xor (n1799,n1800,n1818);
or (n1800,n1801,n1817);
and (n1801,n1802,n1810);
xor (n1802,n1803,n1804);
and (n1803,n298,n887);
nand (n1804,n1805,n1806);
or (n1805,n982,n1645);
or (n1806,n981,n1807);
nor (n1807,n1808,n1809);
and (n1808,n896,n356);
and (n1809,n897,n358);
nand (n1810,n1811,n1816);
or (n1811,n949,n1812);
not (n1812,n1813);
nor (n1813,n1814,n1815);
and (n1814,n111,n495);
and (n1815,n113,n494);
or (n1816,n950,n1701);
and (n1817,n1803,n1804);
or (n1818,n1819,n1842);
and (n1819,n1820,n1836);
xor (n1820,n1821,n1829);
nand (n1821,n1822,n1823);
or (n1822,n1674,n70);
nand (n1823,n1824,n1828);
not (n1824,n1825);
nor (n1825,n1826,n1827);
and (n1826,n841,n80);
and (n1827,n839,n79);
not (n1828,n69);
nand (n1829,n1830,n1835);
or (n1830,n1831,n609);
not (n1831,n1832);
nand (n1832,n1833,n1834);
or (n1833,n185,n137);
or (n1834,n188,n135);
or (n1835,n614,n1668);
nand (n1836,n1837,n1841);
or (n1837,n853,n1838);
nor (n1838,n1839,n1840);
and (n1839,n60,n864);
and (n1840,n58,n863);
or (n1841,n870,n1652);
and (n1842,n1821,n1829);
xor (n1843,n1642,n1656);
and (n1844,n1800,n1818);
xor (n1845,n1626,n1663);
or (n1846,n1847,n1882);
and (n1847,n1848,n1851);
xor (n1848,n1849,n1850);
xor (n1849,n1698,n1713);
xor (n1850,n1665,n1679);
or (n1851,n1852,n1881);
and (n1852,n1853,n1866);
xor (n1853,n1854,n1860);
nand (n1854,n1855,n1859);
or (n1855,n389,n1856);
nor (n1856,n1857,n1858);
and (n1857,n474,n179);
and (n1858,n180,n476);
or (n1859,n183,n1658);
nand (n1860,n1861,n1865);
or (n1861,n197,n1862);
nor (n1862,n1863,n1864);
and (n1863,n149,n1037);
and (n1864,n150,n1036);
or (n1865,n198,n1751);
and (n1866,n1867,n1874);
nor (n1867,n1868,n79);
nor (n1868,n1869,n1872);
and (n1869,n1870,n74);
not (n1870,n1871);
and (n1871,n887,n73);
and (n1872,n935,n1873);
not (n1873,n73);
nand (n1874,n1875,n1880);
or (n1875,n981,n1876);
not (n1876,n1877);
nor (n1877,n1878,n1879);
and (n1878,n41,n896);
and (n1879,n39,n897);
or (n1880,n1807,n982);
and (n1881,n1854,n1860);
and (n1882,n1849,n1850);
and (n1883,n1797,n1845);
or (n1884,n1885,n1970);
and (n1885,n1886,n1889);
xor (n1886,n1887,n1888);
xor (n1887,n1695,n1721);
xor (n1888,n1743,n1746);
or (n1889,n1890,n1969);
and (n1890,n1891,n1968);
xor (n1891,n1892,n1967);
or (n1892,n1893,n1966);
and (n1893,n1894,n1944);
xor (n1894,n1895,n1919);
or (n1895,n1896,n1918);
and (n1896,n1897,n1912);
xor (n1897,n1898,n1905);
nand (n1898,n1899,n1904);
or (n1899,n1900,n949);
not (n1900,n1901);
nor (n1901,n1902,n1903);
and (n1902,n141,n495);
and (n1903,n143,n494);
nand (n1904,n963,n1813);
nand (n1905,n1906,n1911);
or (n1906,n1907,n146);
not (n1907,n1908);
nor (n1908,n1909,n1910);
and (n1909,n834,n156);
and (n1910,n832,n157);
nand (n1911,n1762,n790);
nand (n1912,n1913,n1917);
or (n1913,n219,n1914);
nor (n1914,n1915,n1916);
and (n1915,n847,n74);
and (n1916,n75,n846);
or (n1917,n1768,n220);
and (n1918,n1898,n1905);
or (n1919,n1920,n1943);
and (n1920,n1921,n1937);
xor (n1921,n1922,n1930);
nand (n1922,n1923,n1928);
or (n1923,n1924,n853);
not (n1924,n1925);
nor (n1925,n1926,n1927);
and (n1926,n117,n864);
and (n1927,n119,n863);
nand (n1928,n1929,n855);
not (n1929,n1838);
nand (n1930,n1931,n1932);
or (n1931,n183,n1856);
nand (n1932,n1933,n174);
not (n1933,n1934);
nor (n1934,n1935,n1936);
and (n1935,n625,n179);
and (n1936,n180,n627);
nand (n1937,n1938,n1942);
or (n1938,n197,n1939);
nor (n1939,n1940,n1941);
and (n1940,n149,n1030);
and (n1941,n150,n1032);
or (n1942,n198,n1862);
and (n1943,n1922,n1930);
or (n1944,n1945,n1965);
and (n1945,n1946,n1959);
xor (n1946,n1947,n1953);
nand (n1947,n1948,n1949);
or (n1948,n1776,n894);
or (n1949,n893,n1950);
nor (n1950,n1951,n1952);
and (n1951,n903,n64);
and (n1952,n859,n66);
nand (n1953,n1954,n1958);
or (n1954,n69,n1955);
nor (n1955,n1956,n1957);
and (n1956,n935,n80);
and (n1957,n887,n79);
or (n1958,n70,n1825);
nand (n1959,n1960,n1964);
or (n1960,n609,n1961);
nor (n1961,n1962,n1963);
and (n1962,n188,n448);
and (n1963,n185,n450);
or (n1964,n614,n1831);
and (n1965,n1947,n1953);
and (n1966,n1895,n1919);
xor (n1967,n1748,n1756);
xor (n1968,n1799,n1843);
and (n1969,n1892,n1967);
and (n1970,n1887,n1888);
xor (n1971,n1739,n1785);
and (n1972,n1794,n1884);
nand (n1973,n1732,n1788);
nand (n1974,n1610,n1612);
nand (n1975,n771,n1466);
not (n1976,n1977);
nor (n1977,n1978,n2311,n2654);
nand (n1978,n1979,n2304);
nand (n1979,n1980,n2294);
not (n1980,n1981);
xor (n1981,n1982,n2138);
xor (n1982,n1983,n2056);
or (n1983,n1984,n2055);
and (n1984,n1985,n2052);
xor (n1985,n1986,n2049);
xor (n1986,n1987,n2026);
xor (n1987,n1988,n2008);
xor (n1988,n1989,n2002);
xor (n1989,n1990,n1996);
nand (n1990,n1991,n1992);
or (n1991,n853,n928);
or (n1992,n870,n1993);
nor (n1993,n1994,n1995);
and (n1994,n863,n90);
and (n1995,n864,n92);
nand (n1996,n1997,n1998);
or (n1997,n44,n938);
or (n1998,n45,n1999);
nor (n1999,n2000,n2001);
and (n2000,n53,n847);
and (n2001,n846,n54);
nand (n2002,n2003,n2004);
or (n2003,n197,n1047);
or (n2004,n198,n2005);
nor (n2005,n2006,n2007);
and (n2006,n149,n64);
and (n2007,n150,n66);
xor (n2008,n2009,n2020);
xor (n2009,n2010,n2012);
and (n2010,n2011,n887);
not (n2011,n99);
nand (n2012,n2013,n2015);
or (n2013,n2014,n893);
not (n2014,n1068);
nand (n2015,n2016,n1067);
not (n2016,n2017);
nor (n2017,n2018,n2019);
and (n2018,n238,n859);
and (n2019,n236,n903);
nand (n2020,n2021,n2022);
or (n2021,n949,n960);
or (n2022,n950,n2023);
nor (n2023,n2024,n2025);
and (n2024,n494,n310);
and (n2025,n495,n312);
xor (n2026,n2027,n2043);
xor (n2027,n2028,n2036);
nand (n2028,n2029,n2031);
or (n2029,n2030,n69);
not (n2030,n1023);
nand (n2031,n2032,n71);
not (n2032,n2033);
nor (n2033,n2034,n2035);
and (n2034,n450,n80);
and (n2035,n448,n79);
nand (n2036,n2037,n2038);
or (n2037,n1034,n296);
nand (n2038,n2039,n298);
not (n2039,n2040);
nor (n2040,n2041,n2042);
and (n2041,n627,n306);
and (n2042,n625,n305);
nand (n2043,n2044,n2045);
or (n2044,n981,n988);
or (n2045,n2046,n982);
nor (n2046,n2047,n2048);
and (n2047,n896,n167);
and (n2048,n897,n169);
or (n2049,n2050,n2051);
and (n2050,n1006,n1042);
and (n2051,n1007,n1039);
or (n2052,n2053,n2054);
and (n2053,n1448,n1455);
and (n2054,n1449,n1452);
and (n2055,n1986,n2049);
or (n2056,n2057,n2137);
and (n2057,n2058,n2134);
xor (n2058,n2059,n2090);
xor (n2059,n2060,n2087);
xor (n2060,n2061,n2084);
xor (n2061,n2062,n2077);
xor (n2062,n2063,n2071);
nand (n2063,n2064,n2066);
or (n2064,n2065,n389);
not (n2065,n994);
nand (n2066,n2067,n182);
not (n2067,n2068);
nor (n2068,n2069,n2070);
and (n2069,n179,n39);
and (n2070,n180,n41);
nand (n2071,n2072,n2073);
or (n2072,n331,n1000);
or (n2073,n332,n2074);
nor (n2074,n2075,n2076);
and (n2075,n21,n1030);
and (n2076,n22,n1032);
nand (n2077,n2078,n2080);
or (n2078,n18,n2079);
not (n2079,n920);
or (n2080,n2081,n19);
nor (n2081,n2082,n2083);
and (n2082,n28,n832);
and (n2083,n29,n834);
or (n2084,n2085,n2086);
and (n2085,n1456,n1463);
and (n2086,n1457,n1460);
or (n2087,n2088,n2089);
and (n2088,n1043,n1072);
and (n2089,n1044,n1050);
xor (n2090,n2091,n2131);
xor (n2091,n2092,n2101);
xor (n2092,n2093,n2098);
xor (n2093,n2094,n2095);
and (n2094,n1060,n1052);
or (n2095,n2096,n2097);
and (n2096,n942,n971);
and (n2097,n943,n964);
or (n2098,n2099,n2100);
and (n2099,n1008,n1026);
and (n2100,n1009,n1016);
xor (n2101,n2102,n2109);
xor (n2102,n2103,n2106);
or (n2103,n2104,n2105);
and (n2104,n916,n931);
and (n2105,n917,n924);
or (n2106,n2107,n2108);
and (n2107,n978,n997);
and (n2108,n979,n991);
xor (n2109,n2110,n2125);
xor (n2110,n2111,n2119);
nand (n2111,n2112,n2114);
or (n2112,n2113,n146);
not (n2113,n968);
nand (n2114,n2115,n790);
not (n2115,n2116);
nor (n2116,n2117,n2118);
and (n2117,n156,n117);
and (n2118,n157,n119);
nand (n2119,n2120,n2121);
or (n2120,n219,n974);
or (n2121,n220,n2122);
nor (n2122,n2123,n2124);
and (n2123,n74,n141);
and (n2124,n75,n143);
nand (n2125,n2126,n2127);
or (n2126,n609,n1013);
or (n2127,n614,n2128);
nor (n2128,n2129,n2130);
and (n2129,n188,n342);
and (n2130,n185,n344);
or (n2131,n2132,n2133);
and (n2132,n914,n977);
and (n2133,n915,n941);
or (n2134,n2135,n2136);
and (n2135,n774,n1005);
and (n2136,n775,n913);
and (n2137,n2059,n2090);
xor (n2138,n2139,n2223);
xor (n2139,n2140,n2179);
xor (n2140,n2141,n2176);
xor (n2141,n2142,n2173);
xor (n2142,n2143,n2159);
xor (n2143,n2144,n2150);
nand (n2144,n2145,n2146);
or (n2145,n44,n1999);
or (n2146,n45,n2147);
nor (n2147,n2148,n2149);
and (n2148,n53,n826);
and (n2149,n54,n828);
nand (n2150,n2151,n2155);
or (n2151,n97,n2152);
nor (n2152,n2153,n2154);
and (n2153,n935,n107);
and (n2154,n887,n106);
or (n2155,n99,n2156);
nor (n2156,n2157,n2158);
and (n2157,n839,n106);
and (n2158,n841,n107);
xor (n2159,n2160,n2166);
nor (n2160,n2161,n106);
nor (n2161,n2162,n2165);
and (n2162,n2163,n53);
not (n2163,n2164);
and (n2164,n887,n102);
and (n2165,n935,n101);
nand (n2166,n2167,n2172);
or (n2167,n982,n2168);
not (n2168,n2169);
nor (n2169,n2170,n2171);
and (n2170,n210,n896);
and (n2171,n208,n897);
or (n2172,n981,n2046);
or (n2173,n2174,n2175);
and (n2174,n2093,n2098);
and (n2175,n2094,n2095);
or (n2176,n2177,n2178);
and (n2177,n1987,n2026);
and (n2178,n1988,n2008);
xor (n2179,n2180,n2195);
xor (n2180,n2181,n2192);
xor (n2181,n2182,n2189);
xor (n2182,n2183,n2186);
or (n2183,n2184,n2185);
and (n2184,n2027,n2043);
and (n2185,n2028,n2036);
or (n2186,n2187,n2188);
and (n2187,n2009,n2020);
and (n2188,n2010,n2012);
or (n2189,n2190,n2191);
and (n2190,n2110,n2125);
and (n2191,n2111,n2119);
or (n2192,n2193,n2194);
and (n2193,n2102,n2109);
and (n2194,n2103,n2106);
xor (n2195,n2196,n2203);
xor (n2196,n2197,n2200);
or (n2197,n2198,n2199);
and (n2198,n2062,n2077);
and (n2199,n2063,n2071);
or (n2200,n2201,n2202);
and (n2201,n1989,n2002);
and (n2202,n1990,n1996);
xor (n2203,n2204,n2217);
xor (n2204,n2205,n2211);
nand (n2205,n2206,n2207);
or (n2206,n893,n2017);
or (n2207,n894,n2208);
nor (n2208,n2209,n2210);
and (n2209,n163,n859);
and (n2210,n161,n903);
nand (n2211,n2212,n2213);
or (n2212,n949,n2023);
or (n2213,n950,n2214);
nor (n2214,n2215,n2216);
and (n2215,n86,n495);
and (n2216,n84,n494);
nand (n2217,n2218,n2219);
or (n2218,n146,n2116);
or (n2219,n147,n2220);
nor (n2220,n2221,n2222);
and (n2221,n156,n58);
and (n2222,n157,n60);
xor (n2223,n2224,n2291);
xor (n2224,n2225,n2288);
xor (n2225,n2226,n2268);
xor (n2226,n2227,n2247);
xor (n2227,n2228,n2241);
xor (n2228,n2229,n2235);
nand (n2229,n2230,n2231);
or (n2230,n331,n2074);
or (n2231,n332,n2232);
nor (n2232,n2233,n2234);
and (n2233,n21,n1037);
and (n2234,n22,n1036);
nand (n2235,n2236,n2237);
or (n2236,n18,n2081);
or (n2237,n19,n2238);
nor (n2238,n2239,n2240);
and (n2239,n1004,n29);
and (n2240,n1002,n28);
nand (n2241,n2242,n2243);
or (n2242,n197,n2005);
or (n2243,n198,n2244);
nor (n2244,n2245,n2246);
and (n2245,n149,n33);
and (n2246,n150,n35);
xor (n2247,n2248,n2262);
xor (n2248,n2249,n2255);
nand (n2249,n2250,n2251);
or (n2250,n2122,n219);
or (n2251,n2252,n220);
nor (n2252,n2253,n2254);
and (n2253,n74,n111);
and (n2254,n75,n113);
nand (n2255,n2256,n2257);
or (n2256,n609,n2128);
or (n2257,n614,n2258);
not (n2258,n2259);
nand (n2259,n2260,n2261);
or (n2260,n185,n350);
or (n2261,n188,n348);
nand (n2262,n2263,n2264);
or (n2263,n69,n2033);
or (n2264,n70,n2265);
nor (n2265,n2266,n2267);
and (n2266,n79,n135);
and (n2267,n80,n137);
xor (n2268,n2269,n2282);
xor (n2269,n2270,n2276);
nand (n2270,n2271,n2272);
or (n2271,n296,n2040);
or (n2272,n297,n2273);
nor (n2273,n2274,n2275);
and (n2274,n305,n474);
and (n2275,n306,n476);
nand (n2276,n2277,n2278);
or (n2277,n853,n1993);
or (n2278,n870,n2279);
nor (n2279,n2280,n2281);
and (n2280,n230,n863);
and (n2281,n232,n864);
nand (n2282,n2283,n2284);
or (n2283,n389,n2068);
or (n2284,n183,n2285);
nor (n2285,n2286,n2287);
and (n2286,n179,n356);
and (n2287,n180,n358);
or (n2288,n2289,n2290);
and (n2289,n2060,n2087);
and (n2290,n2061,n2084);
or (n2291,n2292,n2293);
and (n2292,n2091,n2131);
and (n2293,n2092,n2101);
not (n2294,n2295);
or (n2295,n2296,n2303);
and (n2296,n2297,n2302);
xor (n2297,n2298,n2299);
xor (n2298,n1985,n2052);
or (n2299,n2300,n2301);
and (n2300,n1409,n1447);
and (n2301,n1410,n1413);
xor (n2302,n2058,n2134);
and (n2303,n2298,n2299);
nand (n2304,n2305,n2307);
not (n2305,n2306);
xor (n2306,n2297,n2302);
not (n2307,n2308);
or (n2308,n2309,n2310);
and (n2309,n772,n1408);
and (n2310,n773,n1086);
nor (n2311,n2312,n2645);
xor (n2312,n2313,n2636);
xor (n2313,n2314,n2460);
xor (n2314,n2315,n2411);
xor (n2315,n2316,n2389);
xor (n2316,n2317,n2376);
xor (n2317,n2318,n2347);
xor (n2318,n2319,n2338);
xor (n2319,n2320,n2329);
nand (n2320,n2321,n2325);
or (n2321,n69,n2322);
nor (n2322,n2323,n2324);
and (n2323,n79,n141);
and (n2324,n80,n143);
or (n2325,n70,n2326);
nor (n2326,n2327,n2328);
and (n2327,n79,n111);
and (n2328,n80,n113);
nand (n2329,n2330,n2334);
or (n2330,n296,n2331);
nor (n2331,n2332,n2333);
and (n2332,n305,n448);
and (n2333,n306,n450);
or (n2334,n297,n2335);
nor (n2335,n2336,n2337);
and (n2336,n305,n135);
and (n2337,n306,n137);
nand (n2338,n2339,n2343);
or (n2339,n853,n2340);
nor (n2340,n2341,n2342);
and (n2341,n236,n863);
and (n2342,n238,n864);
or (n2343,n870,n2344);
nor (n2344,n2345,n2346);
and (n2345,n863,n161);
and (n2346,n864,n163);
xor (n2347,n2348,n2367);
xor (n2348,n2349,n2358);
nand (n2349,n2350,n2354);
or (n2350,n389,n2351);
nor (n2351,n2352,n2353);
and (n2352,n179,n342);
and (n2353,n180,n344);
or (n2354,n183,n2355);
nor (n2355,n2356,n2357);
and (n2356,n179,n348);
and (n2357,n180,n350);
nand (n2358,n2359,n2363);
or (n2359,n331,n2360);
nor (n2360,n2361,n2362);
and (n2361,n21,n625);
and (n2362,n22,n627);
or (n2363,n332,n2364);
nor (n2364,n2365,n2366);
and (n2365,n21,n474);
and (n2366,n22,n476);
nand (n2367,n2368,n2372);
or (n2368,n18,n2369);
nor (n2369,n2370,n2371);
and (n2370,n28,n1030);
and (n2371,n29,n1032);
or (n2372,n2373,n19);
nor (n2373,n2374,n2375);
and (n2374,n28,n1037);
and (n2375,n29,n1036);
or (n2376,n2377,n2388);
and (n2377,n2378,n2385);
xor (n2378,n2379,n2382);
or (n2379,n2380,n2381);
and (n2380,n2248,n2262);
and (n2381,n2249,n2255);
or (n2382,n2383,n2384);
and (n2383,n2269,n2282);
and (n2384,n2270,n2276);
or (n2385,n2386,n2387);
and (n2386,n2228,n2241);
and (n2387,n2229,n2235);
and (n2388,n2379,n2382);
or (n2389,n2390,n2410);
and (n2390,n2391,n2407);
xor (n2391,n2392,n2404);
xor (n2392,n2393,n2401);
xor (n2393,n2394,n2400);
nand (n2394,n2395,n2396);
or (n2395,n97,n2156);
or (n2396,n99,n2397);
nor (n2397,n2398,n2399);
and (n2398,n847,n106);
and (n2399,n846,n107);
and (n2400,n2160,n2166);
or (n2401,n2402,n2403);
and (n2402,n2204,n2217);
and (n2403,n2205,n2211);
or (n2404,n2405,n2406);
and (n2405,n2182,n2189);
and (n2406,n2183,n2186);
or (n2407,n2408,n2409);
and (n2408,n2226,n2268);
and (n2409,n2227,n2247);
and (n2410,n2392,n2404);
or (n2411,n2412,n2459);
and (n2412,n2413,n2418);
xor (n2413,n2414,n2415);
xor (n2414,n2378,n2385);
or (n2415,n2416,n2417);
and (n2416,n2196,n2203);
and (n2417,n2197,n2200);
xor (n2418,n2419,n2456);
xor (n2419,n2420,n2436);
xor (n2420,n2421,n2433);
xor (n2421,n2422,n2429);
nand (n2422,n2423,n2424);
or (n2423,n2258,n609);
nand (n2424,n2425,n491);
not (n2425,n2426);
nor (n2426,n2427,n2428);
and (n2427,n188,n310);
and (n2428,n185,n312);
nand (n2429,n2430,n2431);
or (n2430,n2265,n69);
nand (n2431,n2432,n71);
not (n2432,n2322);
nand (n2433,n2434,n2435);
or (n2434,n296,n2273);
or (n2435,n297,n2331);
xor (n2436,n2437,n2450);
xor (n2437,n2438,n2444);
nand (n2438,n2439,n2440);
or (n2439,n2214,n949);
nand (n2440,n963,n2441);
nand (n2441,n2442,n2443);
or (n2442,n495,n92);
or (n2443,n494,n90);
nand (n2444,n2445,n2446);
or (n2445,n146,n2220);
or (n2446,n147,n2447);
nor (n2447,n2448,n2449);
and (n2448,n66,n157);
and (n2449,n64,n156);
nand (n2450,n2451,n2452);
or (n2451,n219,n2252);
or (n2452,n220,n2453);
nor (n2453,n2454,n2455);
and (n2454,n74,n117);
and (n2455,n75,n119);
or (n2456,n2457,n2458);
and (n2457,n2143,n2159);
and (n2458,n2144,n2150);
and (n2459,n2414,n2415);
xor (n2460,n2461,n2625);
xor (n2461,n2462,n2543);
xor (n2462,n2463,n2507);
xor (n2463,n2464,n2467);
or (n2464,n2465,n2466);
and (n2465,n2393,n2401);
and (n2466,n2394,n2400);
xor (n2467,n2468,n2486);
xor (n2468,n2469,n2472);
or (n2469,n2470,n2471);
and (n2470,n2421,n2433);
and (n2471,n2422,n2429);
or (n2472,n2473,n2485);
and (n2473,n2474,n2482);
xor (n2474,n2475,n2479);
nand (n2475,n2476,n2477);
or (n2476,n853,n2279);
nand (n2477,n2478,n855);
not (n2478,n2340);
nand (n2479,n2480,n2481);
or (n2480,n389,n2285);
or (n2481,n183,n2351);
nand (n2482,n2483,n2484);
or (n2483,n331,n2232);
or (n2484,n332,n2360);
and (n2485,n2475,n2479);
or (n2486,n2487,n2506);
and (n2487,n2488,n2500);
xor (n2488,n2489,n2492);
nand (n2489,n2490,n2491);
or (n2490,n18,n2238);
or (n2491,n2369,n19);
nand (n2492,n2493,n2498);
or (n2493,n2494,n198);
not (n2494,n2495);
nand (n2495,n2496,n2497);
or (n2496,n150,n41);
or (n2497,n149,n39);
nand (n2498,n2499,n705);
not (n2499,n2244);
nand (n2500,n2501,n2502);
or (n2501,n44,n2147);
or (n2502,n45,n2503);
nor (n2503,n2504,n2505);
and (n2504,n832,n53);
and (n2505,n54,n834);
and (n2506,n2489,n2492);
xor (n2507,n2508,n2540);
xor (n2508,n2509,n2526);
xor (n2509,n2510,n2516);
nor (n2510,n2511,n130);
nor (n2511,n2512,n2515);
and (n2512,n2513,n106);
not (n2513,n2514);
and (n2514,n887,n125);
and (n2515,n935,n127);
nand (n2516,n2517,n2522);
or (n2517,n981,n2518);
not (n2518,n2519);
nor (n2519,n2520,n2521);
and (n2520,n216,n896);
and (n2521,n214,n897);
or (n2522,n2523,n982);
nor (n2523,n2524,n2525);
and (n2524,n896,n192);
and (n2525,n897,n194);
or (n2526,n2527,n2539);
and (n2527,n2528,n2533);
xor (n2528,n2529,n2530);
nor (n2529,n123,n935);
nand (n2530,n2531,n2532);
or (n2531,n981,n2168);
nand (n2532,n2519,n983);
nand (n2533,n2534,n2535);
or (n2534,n2208,n893);
nand (n2535,n1067,n2536);
nor (n2536,n2537,n2538);
and (n2537,n167,n859);
and (n2538,n169,n903);
and (n2539,n2529,n2530);
or (n2540,n2541,n2542);
and (n2541,n2437,n2450);
and (n2542,n2438,n2444);
xor (n2543,n2544,n2555);
xor (n2544,n2545,n2552);
or (n2545,n2546,n2551);
and (n2546,n2547,n2550);
xor (n2547,n2548,n2549);
xor (n2548,n2528,n2533);
xor (n2549,n2488,n2500);
xor (n2550,n2474,n2482);
and (n2551,n2548,n2549);
or (n2552,n2553,n2554);
and (n2553,n2419,n2456);
and (n2554,n2420,n2436);
xor (n2555,n2556,n2604);
xor (n2556,n2557,n2577);
xor (n2557,n2558,n2571);
xor (n2558,n2559,n2565);
nand (n2559,n2560,n2561);
or (n2560,n2494,n197);
nand (n2561,n706,n2562);
nand (n2562,n2563,n2564);
or (n2563,n150,n358);
or (n2564,n149,n356);
nand (n2565,n2566,n2567);
or (n2566,n44,n2503);
or (n2567,n45,n2568);
nor (n2568,n2569,n2570);
and (n2569,n1002,n53);
and (n2570,n54,n1004);
nand (n2571,n2572,n2573);
or (n2572,n97,n2397);
or (n2573,n99,n2574);
nor (n2574,n2575,n2576);
and (n2575,n826,n106);
and (n2576,n107,n828);
xor (n2577,n2578,n2595);
xor (n2578,n2579,n2587);
nand (n2579,n2580,n2582);
or (n2580,n2581,n893);
not (n2581,n2536);
nand (n2582,n2583,n1067);
not (n2583,n2584);
nor (n2584,n2585,n2586);
and (n2585,n210,n859);
and (n2586,n208,n903);
nand (n2587,n2588,n2590);
or (n2588,n2589,n949);
not (n2589,n2441);
nand (n2590,n2591,n963);
not (n2591,n2592);
nor (n2592,n2593,n2594);
and (n2593,n494,n230);
and (n2594,n495,n232);
nand (n2595,n2596,n2600);
or (n2596,n122,n2597);
nor (n2597,n2598,n2599);
and (n2598,n935,n131);
and (n2599,n887,n130);
or (n2600,n2601,n123);
nor (n2601,n2602,n2603);
and (n2602,n839,n130);
and (n2603,n841,n131);
xor (n2604,n2605,n2619);
xor (n2605,n2606,n2613);
nand (n2606,n2607,n2608);
or (n2607,n2447,n146);
nand (n2608,n2609,n790);
not (n2609,n2610);
nor (n2610,n2611,n2612);
and (n2611,n156,n33);
and (n2612,n157,n35);
nand (n2613,n2614,n2615);
or (n2614,n219,n2453);
or (n2615,n220,n2616);
nor (n2616,n2617,n2618);
and (n2617,n60,n75);
and (n2618,n58,n74);
nand (n2619,n2620,n2621);
or (n2620,n609,n2426);
or (n2621,n614,n2622);
nor (n2622,n2623,n2624);
and (n2623,n188,n84);
and (n2624,n185,n86);
or (n2625,n2626,n2635);
and (n2626,n2627,n2632);
xor (n2627,n2628,n2629);
xor (n2628,n2547,n2550);
or (n2629,n2630,n2631);
and (n2630,n2180,n2195);
and (n2631,n2181,n2192);
or (n2632,n2633,n2634);
and (n2633,n2141,n2176);
and (n2634,n2142,n2173);
and (n2635,n2628,n2629);
or (n2636,n2637,n2644);
and (n2637,n2638,n2641);
xor (n2638,n2639,n2640);
xor (n2639,n2391,n2407);
xor (n2640,n2413,n2418);
or (n2641,n2642,n2643);
and (n2642,n2224,n2291);
and (n2643,n2225,n2288);
and (n2644,n2639,n2640);
or (n2645,n2646,n2653);
and (n2646,n2647,n2650);
xor (n2647,n2648,n2649);
xor (n2648,n2627,n2632);
xor (n2649,n2638,n2641);
or (n2650,n2651,n2652);
and (n2651,n2139,n2223);
and (n2652,n2140,n2179);
and (n2653,n2648,n2649);
nor (n2654,n2655,n2656);
xor (n2655,n2647,n2650);
or (n2656,n2657,n2658);
and (n2657,n1982,n2138);
and (n2658,n1983,n2056);
or (n2659,n2660,n2668);
nand (n2660,n2661,n2662,n2663,n2667);
not (n2661,n1978);
not (n2662,n2311);
nor (n2663,n2664,n770);
nand (n2664,n2665,n1608);
nor (n2665,n2666,n1731);
nor (n2666,n1790,n1791);
not (n2667,n2654);
not (n2668,n2669);
nand (n2669,n2670,n3825,n3837,n3850);
nand (n2670,n2671,n2989,n3755);
and (n2671,n2672,n2971,n2984);
nor (n2672,n2673,n2886);
nor (n2673,n2674,n2774);
xor (n2674,n2675,n2767);
xor (n2675,n2676,n2756);
or (n2676,n2677,n2755);
and (n2677,n2678,n2725);
xor (n2678,n2679,n2680);
xor (n2679,n1853,n1866);
or (n2680,n2681,n2724);
and (n2681,n2682,n2702);
xor (n2682,n2683,n2684);
xor (n2683,n1867,n1874);
or (n2684,n2685,n2701);
and (n2685,n2686,n2695);
xor (n2686,n2687,n2688);
and (n2687,n71,n887);
nand (n2688,n2689,n2694);
or (n2689,n981,n2690);
not (n2690,n2691);
nor (n2691,n2692,n2693);
and (n2692,n33,n897);
and (n2693,n35,n896);
nand (n2694,n1877,n983);
nand (n2695,n2696,n2700);
or (n2696,n949,n2697);
nor (n2697,n2698,n2699);
and (n2698,n494,n135);
and (n2699,n495,n137);
or (n2700,n950,n1900);
and (n2701,n2687,n2688);
or (n2702,n2703,n2723);
and (n2703,n2704,n2717);
xor (n2704,n2705,n2711);
nand (n2705,n2706,n2710);
or (n2706,n146,n2707);
nor (n2707,n2708,n2709);
and (n2708,n828,n157);
and (n2709,n826,n156);
or (n2710,n147,n1907);
nand (n2711,n2712,n2716);
or (n2712,n219,n2713);
nor (n2713,n2714,n2715);
and (n2714,n74,n839);
and (n2715,n75,n841);
or (n2716,n220,n1914);
nand (n2717,n2718,n2722);
or (n2718,n893,n2719);
nor (n2719,n2720,n2721);
and (n2720,n903,n58);
and (n2721,n859,n60);
or (n2722,n894,n1950);
and (n2723,n2705,n2711);
and (n2724,n2683,n2684);
or (n2725,n2726,n2754);
and (n2726,n2727,n2753);
xor (n2727,n2728,n2752);
or (n2728,n2729,n2751);
and (n2729,n2730,n2745);
xor (n2730,n2731,n2739);
nand (n2731,n2732,n2737);
or (n2732,n2733,n609);
not (n2733,n2734);
nand (n2734,n2735,n2736);
or (n2735,n185,n476);
or (n2736,n188,n474);
nand (n2737,n2738,n491);
not (n2738,n1961);
nand (n2739,n2740,n2744);
or (n2740,n2741,n853);
nor (n2741,n2742,n2743);
and (n2742,n863,n111);
and (n2743,n864,n113);
nand (n2744,n855,n1925);
nand (n2745,n2746,n2750);
or (n2746,n389,n2747);
nor (n2747,n2748,n2749);
and (n2748,n179,n1037);
and (n2749,n180,n1036);
or (n2750,n183,n1934);
and (n2751,n2731,n2739);
xor (n2752,n1921,n1937);
xor (n2753,n1897,n1912);
and (n2754,n2728,n2752);
and (n2755,n2679,n2680);
xor (n2756,n2757,n2766);
xor (n2757,n2758,n2765);
or (n2758,n2759,n2764);
and (n2759,n2760,n2763);
xor (n2760,n2761,n2762);
xor (n2761,n1802,n1810);
xor (n2762,n1758,n1774);
xor (n2763,n1820,n1836);
and (n2764,n2761,n2762);
xor (n2765,n1848,n1851);
xor (n2766,n1891,n1968);
or (n2767,n2768,n2773);
and (n2768,n2769,n2772);
xor (n2769,n2770,n2771);
xor (n2770,n1894,n1944);
xor (n2771,n2760,n2763);
xor (n2772,n2678,n2725);
and (n2773,n2770,n2771);
or (n2774,n2775,n2885);
and (n2775,n2776,n2884);
xor (n2776,n2777,n2828);
or (n2777,n2778,n2827);
and (n2778,n2779,n2826);
xor (n2779,n2780,n2781);
xor (n2780,n1946,n1959);
or (n2781,n2782,n2825);
and (n2782,n2783,n2803);
xor (n2783,n2784,n2790);
nand (n2784,n2785,n2789);
or (n2785,n197,n2786);
nor (n2786,n2787,n2788);
and (n2787,n149,n1002);
and (n2788,n150,n1004);
or (n2789,n198,n1939);
and (n2790,n2791,n2797);
nor (n2791,n2792,n74);
nor (n2792,n2793,n2796);
and (n2793,n2794,n156);
not (n2794,n2795);
and (n2795,n887,n222);
and (n2796,n935,n224);
nand (n2797,n2798,n2799);
or (n2798,n982,n2690);
or (n2799,n981,n2800);
nor (n2800,n2801,n2802);
and (n2801,n66,n897);
and (n2802,n64,n896);
or (n2803,n2804,n2824);
and (n2804,n2805,n2818);
xor (n2805,n2806,n2812);
nand (n2806,n2807,n2811);
or (n2807,n949,n2808);
nor (n2808,n2809,n2810);
and (n2809,n494,n448);
and (n2810,n495,n450);
or (n2811,n950,n2697);
nand (n2812,n2813,n2817);
or (n2813,n146,n2814);
nor (n2814,n2815,n2816);
and (n2815,n156,n847);
and (n2816,n157,n846);
or (n2817,n147,n2707);
nand (n2818,n2819,n2823);
or (n2819,n219,n2820);
nor (n2820,n2821,n2822);
and (n2821,n935,n75);
and (n2822,n74,n887);
or (n2823,n220,n2713);
and (n2824,n2806,n2812);
and (n2825,n2784,n2790);
xor (n2826,n2682,n2702);
and (n2827,n2780,n2781);
or (n2828,n2829,n2883);
and (n2829,n2830,n2860);
xor (n2830,n2831,n2859);
or (n2831,n2832,n2858);
and (n2832,n2833,n2857);
xor (n2833,n2834,n2856);
or (n2834,n2835,n2855);
and (n2835,n2836,n2849);
xor (n2836,n2837,n2843);
nand (n2837,n2838,n2842);
or (n2838,n893,n2839);
nor (n2839,n2840,n2841);
and (n2840,n903,n117);
and (n2841,n859,n119);
or (n2842,n894,n2719);
nand (n2843,n2844,n2848);
or (n2844,n609,n2845);
nor (n2845,n2846,n2847);
and (n2846,n188,n625);
and (n2847,n185,n627);
or (n2848,n614,n2733);
nand (n2849,n2850,n2854);
or (n2850,n853,n2851);
nor (n2851,n2852,n2853);
and (n2852,n863,n141);
and (n2853,n864,n143);
or (n2854,n870,n2741);
and (n2855,n2837,n2843);
xor (n2856,n2730,n2745);
xor (n2857,n2686,n2695);
and (n2858,n2834,n2856);
xor (n2859,n2727,n2753);
or (n2860,n2861,n2882);
and (n2861,n2862,n2881);
xor (n2862,n2863,n2864);
xor (n2863,n2704,n2717);
or (n2864,n2865,n2880);
and (n2865,n2866,n2879);
xor (n2866,n2867,n2873);
nand (n2867,n2868,n2872);
or (n2868,n389,n2869);
nor (n2869,n2870,n2871);
and (n2870,n179,n1030);
and (n2871,n180,n1032);
or (n2872,n183,n2747);
nand (n2873,n2874,n2878);
or (n2874,n197,n2875);
nor (n2875,n2876,n2877);
and (n2876,n149,n832);
and (n2877,n150,n834);
or (n2878,n198,n2786);
xor (n2879,n2791,n2797);
and (n2880,n2867,n2873);
xor (n2881,n2783,n2803);
and (n2882,n2863,n2864);
and (n2883,n2831,n2859);
xor (n2884,n2769,n2772);
and (n2885,n2777,n2828);
nor (n2886,n2887,n2888);
xor (n2887,n2776,n2884);
or (n2888,n2889,n2970);
and (n2889,n2890,n2969);
xor (n2890,n2891,n2892);
xor (n2891,n2779,n2826);
or (n2892,n2893,n2968);
and (n2893,n2894,n2967);
xor (n2894,n2895,n2960);
or (n2895,n2896,n2959);
and (n2896,n2897,n2937);
xor (n2897,n2898,n2915);
or (n2898,n2899,n2914);
and (n2899,n2900,n2908);
xor (n2900,n2901,n2902);
nor (n2901,n220,n935);
nand (n2902,n2903,n2907);
or (n2903,n981,n2904);
nor (n2904,n2905,n2906);
and (n2905,n896,n58);
and (n2906,n897,n60);
or (n2907,n2800,n982);
nand (n2908,n2909,n2913);
or (n2909,n893,n2910);
nor (n2910,n2911,n2912);
and (n2911,n903,n111);
and (n2912,n859,n113);
or (n2913,n894,n2839);
and (n2914,n2901,n2902);
or (n2915,n2916,n2936);
and (n2916,n2917,n2930);
xor (n2917,n2918,n2924);
nand (n2918,n2919,n2923);
or (n2919,n853,n2920);
nor (n2920,n2921,n2922);
and (n2921,n863,n135);
and (n2922,n864,n137);
or (n2923,n870,n2851);
nand (n2924,n2925,n2929);
or (n2925,n389,n2926);
nor (n2926,n2927,n2928);
and (n2927,n179,n1002);
and (n2928,n180,n1004);
or (n2929,n183,n2869);
nand (n2930,n2931,n2935);
or (n2931,n197,n2932);
nor (n2932,n2933,n2934);
and (n2933,n149,n826);
and (n2934,n150,n828);
or (n2935,n198,n2875);
and (n2936,n2918,n2924);
or (n2937,n2938,n2958);
and (n2938,n2939,n2952);
xor (n2939,n2940,n2946);
nand (n2940,n2941,n2945);
or (n2941,n146,n2942);
nor (n2942,n2943,n2944);
and (n2943,n156,n839);
and (n2944,n157,n841);
or (n2945,n147,n2814);
nand (n2946,n2947,n2951);
or (n2947,n949,n2948);
nor (n2948,n2949,n2950);
and (n2949,n494,n474);
and (n2950,n495,n476);
or (n2951,n950,n2808);
nand (n2952,n2953,n2957);
or (n2953,n609,n2954);
nor (n2954,n2955,n2956);
and (n2955,n188,n1037);
and (n2956,n185,n1036);
or (n2957,n614,n2845);
and (n2958,n2940,n2946);
and (n2959,n2898,n2915);
or (n2960,n2961,n2966);
and (n2961,n2962,n2965);
xor (n2962,n2963,n2964);
xor (n2963,n2805,n2818);
xor (n2964,n2836,n2849);
xor (n2965,n2866,n2879);
and (n2966,n2963,n2964);
xor (n2967,n2833,n2857);
and (n2968,n2895,n2960);
xor (n2969,n2830,n2860);
and (n2970,n2891,n2892);
nand (n2971,n2972,n2980);
not (n2972,n2973);
xor (n2973,n2974,n2977);
xor (n2974,n2975,n2976);
xor (n2975,n1796,n1846);
xor (n2976,n1886,n1889);
or (n2977,n2978,n2979);
and (n2978,n2757,n2766);
and (n2979,n2758,n2765);
not (n2980,n2981);
or (n2981,n2982,n2983);
and (n2982,n2675,n2767);
and (n2983,n2676,n2756);
or (n2984,n2985,n2988);
or (n2985,n2986,n2987);
and (n2986,n2974,n2977);
and (n2987,n2975,n2976);
xor (n2988,n1793,n1971);
or (n2989,n2990,n3754);
and (n2990,n2991,n3297);
xor (n2991,n2992,n3235);
or (n2992,n2993,n3234);
and (n2993,n2994,n3181);
xor (n2994,n2995,n3085);
xor (n2995,n2996,n3067);
xor (n2996,n2997,n3034);
or (n2997,n2998,n3033);
and (n2998,n2999,n3022);
xor (n2999,n3000,n3011);
nand (n3000,n3001,n3006);
or (n3001,n3002,n893);
not (n3002,n3003);
nor (n3003,n3004,n3005);
and (n3004,n448,n859);
and (n3005,n450,n903);
nand (n3006,n3007,n1067);
not (n3007,n3008);
nor (n3008,n3009,n3010);
and (n3009,n137,n859);
and (n3010,n135,n903);
nand (n3011,n3012,n3017);
or (n3012,n3013,n949);
not (n3013,n3014);
nand (n3014,n3015,n3016);
or (n3015,n495,n1032);
or (n3016,n494,n1030);
nand (n3017,n3018,n963);
not (n3018,n3019);
nor (n3019,n3020,n3021);
and (n3020,n494,n1037);
and (n3021,n495,n1036);
nand (n3022,n3023,n3028);
or (n3023,n3024,n609);
not (n3024,n3025);
nor (n3025,n3026,n3027);
and (n3026,n832,n185);
and (n3027,n834,n188);
nand (n3028,n3029,n491);
not (n3029,n3030);
nor (n3030,n3031,n3032);
and (n3031,n188,n1002);
and (n3032,n185,n1004);
and (n3033,n3000,n3011);
or (n3034,n3035,n3066);
and (n3035,n3036,n3057);
xor (n3036,n3037,n3047);
nand (n3037,n3038,n3042);
or (n3038,n3039,n853);
nor (n3039,n3040,n3041);
and (n3040,n627,n864);
and (n3041,n625,n863);
nand (n3042,n3043,n855);
not (n3043,n3044);
nor (n3044,n3045,n3046);
and (n3045,n863,n474);
and (n3046,n864,n476);
nand (n3047,n3048,n3052);
or (n3048,n3049,n389);
nor (n3049,n3050,n3051);
and (n3050,n179,n847);
and (n3051,n180,n846);
nand (n3052,n3053,n182);
not (n3053,n3054);
nor (n3054,n3055,n3056);
and (n3055,n179,n826);
and (n3056,n180,n828);
nand (n3057,n3058,n3062);
or (n3058,n197,n3059);
nor (n3059,n3060,n3061);
and (n3060,n935,n150);
and (n3061,n887,n149);
or (n3062,n198,n3063);
nor (n3063,n3064,n3065);
and (n3064,n149,n839);
and (n3065,n150,n841);
and (n3066,n3037,n3047);
xor (n3067,n3068,n3079);
xor (n3068,n3069,n3070);
nor (n3069,n147,n935);
nand (n3070,n3071,n3075);
or (n3071,n981,n3072);
nor (n3072,n3073,n3074);
and (n3073,n113,n897);
and (n3074,n111,n896);
or (n3075,n3076,n982);
nor (n3076,n3077,n3078);
and (n3077,n896,n117);
and (n3078,n897,n119);
nand (n3079,n3080,n3081);
or (n3080,n893,n3008);
or (n3081,n894,n3082);
nor (n3082,n3083,n3084);
and (n3083,n903,n141);
and (n3084,n859,n143);
xor (n3085,n3086,n3134);
xor (n3086,n3087,n3107);
xor (n3087,n3088,n3101);
xor (n3088,n3089,n3095);
nand (n3089,n3090,n3091);
or (n3090,n949,n3019);
or (n3091,n950,n3092);
nor (n3092,n3093,n3094);
and (n3093,n494,n625);
and (n3094,n495,n627);
nand (n3095,n3096,n3097);
or (n3096,n609,n3030);
or (n3097,n614,n3098);
nor (n3098,n3099,n3100);
and (n3099,n188,n1030);
and (n3100,n185,n1032);
nand (n3101,n3102,n3103);
or (n3102,n853,n3044);
or (n3103,n870,n3104);
nor (n3104,n3105,n3106);
and (n3105,n863,n448);
and (n3106,n864,n450);
xor (n3107,n3108,n3121);
xor (n3108,n3109,n3115);
nand (n3109,n3110,n3111);
or (n3110,n389,n3054);
or (n3111,n183,n3112);
nor (n3112,n3113,n3114);
and (n3113,n179,n832);
and (n3114,n180,n834);
nand (n3115,n3116,n3117);
or (n3116,n197,n3063);
or (n3117,n198,n3118);
nor (n3118,n3119,n3120);
and (n3119,n149,n847);
and (n3120,n150,n846);
and (n3121,n3122,n3128);
nor (n3122,n3123,n149);
nor (n3123,n3124,n3127);
and (n3124,n3125,n179);
not (n3125,n3126);
and (n3126,n887,n200);
and (n3127,n935,n202);
nand (n3128,n3129,n3133);
or (n3129,n981,n3130);
nor (n3130,n3131,n3132);
and (n3131,n896,n141);
and (n3132,n897,n143);
or (n3133,n3072,n982);
or (n3134,n3135,n3180);
and (n3135,n3136,n3157);
xor (n3136,n3137,n3138);
xor (n3137,n3122,n3128);
or (n3138,n3139,n3156);
and (n3139,n3140,n3149);
xor (n3140,n3141,n3142);
nor (n3141,n198,n935);
nand (n3142,n3143,n3148);
or (n3143,n3144,n893);
not (n3144,n3145);
nand (n3145,n3146,n3147);
or (n3146,n859,n476);
or (n3147,n903,n474);
nand (n3148,n1067,n3003);
nand (n3149,n3150,n3155);
or (n3150,n949,n3151);
not (n3151,n3152);
nor (n3152,n3153,n3154);
and (n3153,n1004,n494);
and (n3154,n1002,n495);
or (n3155,n950,n3013);
and (n3156,n3141,n3142);
or (n3157,n3158,n3179);
and (n3158,n3159,n3173);
xor (n3159,n3160,n3167);
nand (n3160,n3161,n3166);
or (n3161,n3162,n609);
not (n3162,n3163);
nor (n3163,n3164,n3165);
and (n3164,n828,n188);
and (n3165,n826,n185);
nand (n3166,n491,n3025);
nand (n3167,n3168,n3172);
or (n3168,n981,n3169);
nor (n3169,n3170,n3171);
and (n3170,n896,n135);
and (n3171,n897,n137);
or (n3172,n3130,n982);
nand (n3173,n3174,n3178);
or (n3174,n389,n3175);
nor (n3175,n3176,n3177);
and (n3176,n179,n839);
and (n3177,n180,n841);
or (n3178,n183,n3049);
and (n3179,n3160,n3167);
and (n3180,n3137,n3138);
or (n3181,n3182,n3233);
and (n3182,n3183,n3186);
xor (n3183,n3184,n3185);
xor (n3184,n3036,n3057);
xor (n3185,n2999,n3022);
or (n3186,n3187,n3232);
and (n3187,n3188,n3210);
xor (n3188,n3189,n3195);
nand (n3189,n3190,n3194);
or (n3190,n853,n3191);
nor (n3191,n3192,n3193);
and (n3192,n863,n1037);
and (n3193,n864,n1036);
or (n3194,n870,n3039);
nor (n3195,n3196,n3204);
not (n3196,n3197);
nand (n3197,n3198,n3203);
or (n3198,n3199,n893);
not (n3199,n3200);
nand (n3200,n3201,n3202);
or (n3201,n859,n627);
or (n3202,n903,n625);
nand (n3203,n1067,n3145);
nand (n3204,n3205,n180);
nand (n3205,n3206,n3207);
or (n3206,n887,n178);
nand (n3207,n3208,n188);
not (n3208,n3209);
and (n3209,n887,n178);
or (n3210,n3211,n3231);
and (n3211,n3212,n3225);
xor (n3212,n3213,n3219);
nand (n3213,n3214,n3215);
or (n3214,n3151,n950);
or (n3215,n949,n3216);
nor (n3216,n3217,n3218);
and (n3217,n494,n832);
and (n3218,n495,n834);
nand (n3219,n3220,n3224);
or (n3220,n609,n3221);
or (n3221,n3222,n3223);
and (n3222,n847,n185);
and (n3223,n846,n188);
nand (n3224,n491,n3163);
nand (n3225,n3226,n3230);
or (n3226,n981,n3227);
nor (n3227,n3228,n3229);
and (n3228,n896,n448);
and (n3229,n897,n450);
or (n3230,n3169,n982);
and (n3231,n3213,n3219);
and (n3232,n3189,n3195);
and (n3233,n3184,n3185);
and (n3234,n2995,n3085);
xor (n3235,n3236,n3271);
xor (n3236,n3237,n3268);
xor (n3237,n3238,n3253);
xor (n3238,n3239,n3242);
or (n3239,n3240,n3241);
and (n3240,n3088,n3101);
and (n3241,n3089,n3095);
xor (n3242,n3243,n3250);
xor (n3243,n3244,n3247);
nand (n3244,n3245,n3246);
or (n3245,n609,n3098);
or (n3246,n614,n2954);
nand (n3247,n3248,n3249);
or (n3248,n853,n3104);
or (n3249,n870,n2920);
nand (n3250,n3251,n3252);
or (n3251,n389,n3112);
or (n3252,n183,n2926);
xor (n3253,n3254,n3265);
xor (n3254,n3255,n3259);
nand (n3255,n3256,n3257);
or (n3256,n3082,n893);
nand (n3257,n3258,n1067);
not (n3258,n2910);
nand (n3259,n3260,n3264);
or (n3260,n146,n3261);
nor (n3261,n3262,n3263);
and (n3262,n935,n157);
and (n3263,n887,n156);
or (n3264,n147,n2942);
nand (n3265,n3266,n3267);
or (n3266,n949,n3092);
or (n3267,n950,n2948);
or (n3268,n3269,n3270);
and (n3269,n3086,n3134);
and (n3270,n3087,n3107);
xor (n3271,n3272,n3294);
xor (n3272,n3273,n3276);
or (n3273,n3274,n3275);
and (n3274,n3108,n3121);
and (n3275,n3109,n3115);
xor (n3276,n3277,n3291);
xor (n3277,n3278,n3281);
nand (n3278,n3279,n3280);
or (n3279,n197,n3118);
or (n3280,n198,n2932);
xor (n3281,n3282,n3288);
nor (n3282,n3283,n156);
nor (n3283,n3284,n3287);
and (n3284,n3285,n149);
not (n3285,n3286);
and (n3286,n887,n151);
and (n3287,n935,n153);
nand (n3288,n3289,n3290);
or (n3289,n981,n3076);
or (n3290,n2904,n982);
or (n3291,n3292,n3293);
and (n3292,n3068,n3079);
and (n3293,n3069,n3070);
or (n3294,n3295,n3296);
and (n3295,n2996,n3067);
and (n3296,n2997,n3034);
or (n3297,n3298,n3753);
and (n3298,n3299,n3333);
xor (n3299,n3300,n3332);
or (n3300,n3301,n3331);
and (n3301,n3302,n3330);
xor (n3302,n3303,n3304);
xor (n3303,n3136,n3157);
or (n3304,n3305,n3329);
and (n3305,n3306,n3309);
xor (n3306,n3307,n3308);
xor (n3307,n3159,n3173);
xor (n3308,n3140,n3149);
or (n3309,n3310,n3328);
and (n3310,n3311,n3324);
xor (n3311,n3312,n3318);
nand (n3312,n3313,n3317);
or (n3313,n389,n3314);
nor (n3314,n3315,n3316);
and (n3315,n935,n180);
and (n3316,n179,n887);
or (n3317,n183,n3175);
nand (n3318,n3319,n3323);
or (n3319,n853,n3320);
nor (n3320,n3321,n3322);
and (n3321,n863,n1030);
and (n3322,n864,n1032);
or (n3323,n870,n3191);
nand (n3324,n3325,n3327);
or (n3325,n3326,n3196);
not (n3326,n3204);
or (n3327,n3197,n3204);
and (n3328,n3312,n3318);
and (n3329,n3307,n3308);
xor (n3330,n3183,n3186);
and (n3331,n3303,n3304);
xor (n3332,n2994,n3181);
nand (n3333,n3334,n3747);
nand (n3334,n3335,n3730);
nand (n3335,n3336,n3729);
or (n3336,n3337,n3467);
not (n3337,n3338);
nand (n3338,n3339,n3430);
not (n3339,n3340);
xor (n3340,n3341,n3388);
xor (n3341,n3342,n3343);
xor (n3342,n3311,n3324);
xor (n3343,n3344,n3387);
xor (n3344,n3345,n3363);
or (n3345,n3346,n3362);
and (n3346,n3347,n3356);
xor (n3347,n3348,n3349);
nor (n3348,n183,n935);
nand (n3349,n3350,n3355);
or (n3350,n3351,n893);
not (n3351,n3352);
nand (n3352,n3353,n3354);
or (n3353,n859,n1036);
or (n3354,n903,n1037);
nand (n3355,n1067,n3200);
nand (n3356,n3357,n3361);
or (n3357,n949,n3358);
nor (n3358,n3359,n3360);
and (n3359,n494,n826);
and (n3360,n495,n828);
or (n3361,n950,n3216);
and (n3362,n3348,n3349);
or (n3363,n3364,n3386);
and (n3364,n3365,n3380);
xor (n3365,n3366,n3374);
nand (n3366,n3367,n3372);
or (n3367,n3368,n609);
not (n3368,n3369);
nand (n3369,n3370,n3371);
or (n3370,n185,n841);
or (n3371,n188,n839);
nand (n3372,n3373,n491);
not (n3373,n3221);
nand (n3374,n3375,n3379);
or (n3375,n981,n3376);
nor (n3376,n3377,n3378);
and (n3377,n896,n474);
and (n3378,n897,n476);
or (n3379,n3227,n982);
nand (n3380,n3381,n3385);
or (n3381,n853,n3382);
nor (n3382,n3383,n3384);
and (n3383,n863,n1002);
and (n3384,n864,n1004);
or (n3385,n870,n3320);
and (n3386,n3366,n3374);
xor (n3387,n3212,n3225);
or (n3388,n3389,n3429);
and (n3389,n3390,n3428);
xor (n3390,n3391,n3405);
and (n3391,n3392,n3398);
and (n3392,n3393,n185);
nand (n3393,n3394,n3395);
or (n3394,n887,n493);
nand (n3395,n3396,n494);
not (n3396,n3397);
and (n3397,n887,n493);
nand (n3398,n3399,n3404);
or (n3399,n3400,n893);
not (n3400,n3401);
nor (n3401,n3402,n3403);
and (n3402,n1030,n859);
and (n3403,n1032,n903);
nand (n3404,n1067,n3352);
or (n3405,n3406,n3427);
and (n3406,n3407,n3421);
xor (n3407,n3408,n3415);
nand (n3408,n3409,n3413);
or (n3409,n3410,n949);
nor (n3410,n3411,n3412);
and (n3411,n847,n494);
and (n3412,n846,n495);
nand (n3413,n3414,n963);
not (n3414,n3358);
nand (n3415,n3416,n3417);
or (n3416,n3368,n614);
nand (n3417,n490,n3418);
nand (n3418,n3419,n3420);
or (n3419,n887,n188);
or (n3420,n935,n185);
nand (n3421,n3422,n3426);
or (n3422,n981,n3423);
nor (n3423,n3424,n3425);
and (n3424,n896,n625);
and (n3425,n897,n627);
or (n3426,n3376,n982);
and (n3427,n3408,n3415);
xor (n3428,n3347,n3356);
and (n3429,n3391,n3405);
not (n3430,n3431);
or (n3431,n3432,n3466);
and (n3432,n3433,n3465);
xor (n3433,n3434,n3435);
xor (n3434,n3365,n3380);
or (n3435,n3436,n3464);
and (n3436,n3437,n3445);
xor (n3437,n3438,n3444);
nand (n3438,n3439,n3443);
or (n3439,n853,n3440);
nor (n3440,n3441,n3442);
and (n3441,n863,n832);
and (n3442,n864,n834);
or (n3443,n870,n3382);
xor (n3444,n3392,n3398);
or (n3445,n3446,n3463);
and (n3446,n3447,n3456);
xor (n3447,n3448,n3449);
and (n3448,n491,n887);
nand (n3449,n3450,n3451);
or (n3450,n3423,n982);
nand (n3451,n3452,n1361);
not (n3452,n3453);
nor (n3453,n3454,n3455);
and (n3454,n896,n1037);
and (n3455,n897,n1036);
nand (n3456,n3457,n3462);
or (n3457,n3458,n949);
not (n3458,n3459);
nor (n3459,n3460,n3461);
and (n3460,n839,n495);
and (n3461,n841,n494);
or (n3462,n950,n3410);
and (n3463,n3448,n3449);
and (n3464,n3438,n3444);
xor (n3465,n3390,n3428);
and (n3466,n3434,n3435);
not (n3467,n3468);
nand (n3468,n3469,n3728);
or (n3469,n3470,n3513);
not (n3470,n3471);
nand (n3471,n3472,n3474);
not (n3472,n3473);
xor (n3473,n3433,n3465);
not (n3474,n3475);
or (n3475,n3476,n3512);
and (n3476,n3477,n3511);
xor (n3477,n3478,n3479);
xor (n3478,n3407,n3421);
or (n3479,n3480,n3510);
and (n3480,n3481,n3497);
xor (n3481,n3482,n3489);
nand (n3482,n3483,n3488);
or (n3483,n3484,n893);
not (n3484,n3485);
nor (n3485,n3486,n3487);
and (n3486,n1002,n859);
and (n3487,n1004,n903);
nand (n3488,n1067,n3401);
nand (n3489,n3490,n3495);
or (n3490,n3491,n853);
not (n3491,n3492);
nand (n3492,n3493,n3494);
or (n3493,n864,n828);
or (n3494,n863,n826);
nand (n3495,n3496,n855);
not (n3496,n3440);
and (n3497,n3498,n3504);
nor (n3498,n3499,n494);
nor (n3499,n3500,n3503);
and (n3500,n3501,n863);
not (n3501,n3502);
and (n3502,n887,n952);
and (n3503,n935,n954);
nand (n3504,n3505,n3509);
or (n3505,n981,n3506);
nor (n3506,n3507,n3508);
and (n3507,n1030,n896);
and (n3508,n1032,n897);
or (n3509,n3453,n982);
and (n3510,n3482,n3489);
xor (n3511,n3437,n3445);
and (n3512,n3478,n3479);
not (n3513,n3514);
nand (n3514,n3515,n3724,n3727);
nand (n3515,n3516,n3704,n3717);
nand (n3516,n3517,n3703);
or (n3517,n3518,n3593);
not (n3518,n3519);
nand (n3519,n3520,n3567);
not (n3520,n3521);
xor (n3521,n3522,n3547);
xor (n3522,n3523,n3524);
xor (n3523,n3498,n3504);
or (n3524,n3525,n3546);
and (n3525,n3526,n3536);
xor (n3526,n3527,n3528);
and (n3527,n963,n887);
nand (n3528,n3529,n3534);
or (n3529,n981,n3530);
not (n3530,n3531);
nor (n3531,n3532,n3533);
and (n3532,n1004,n896);
and (n3533,n1002,n897);
nand (n3534,n3535,n983);
not (n3535,n3506);
nand (n3536,n3537,n3542);
or (n3537,n3538,n893);
not (n3538,n3539);
nor (n3539,n3540,n3541);
and (n3540,n828,n903);
and (n3541,n826,n859);
nand (n3542,n1067,n3543);
nor (n3543,n3544,n3545);
and (n3544,n832,n859);
and (n3545,n834,n903);
and (n3546,n3527,n3528);
xor (n3547,n3548,n3560);
xor (n3548,n3549,n3556);
nand (n3549,n3550,n3555);
or (n3550,n3551,n949);
not (n3551,n3552);
nand (n3552,n3553,n3554);
or (n3553,n494,n887);
or (n3554,n935,n495);
nand (n3555,n963,n3459);
nand (n3556,n3557,n3559);
or (n3557,n3558,n893);
not (n3558,n3543);
nand (n3559,n1067,n3485);
nand (n3560,n3561,n3566);
or (n3561,n3562,n853);
not (n3562,n3563);
nand (n3563,n3564,n3565);
or (n3564,n864,n846);
or (n3565,n863,n847);
nand (n3566,n855,n3492);
not (n3567,n3568);
or (n3568,n3569,n3592);
and (n3569,n3570,n3591);
xor (n3570,n3571,n3578);
nand (n3571,n3572,n3577);
or (n3572,n3573,n853);
not (n3573,n3574);
nor (n3574,n3575,n3576);
and (n3575,n839,n864);
and (n3576,n841,n863);
nand (n3577,n855,n3563);
and (n3578,n3579,n3584);
and (n3579,n3580,n864);
nand (n3580,n3581,n3583);
or (n3581,n3582,n859);
and (n3582,n887,n858);
or (n3583,n887,n858);
nand (n3584,n3585,n3586);
or (n3585,n982,n3530);
nand (n3586,n3587,n1361);
not (n3587,n3588);
nor (n3588,n3589,n3590);
and (n3589,n832,n896);
and (n3590,n834,n897);
xor (n3591,n3526,n3536);
and (n3592,n3571,n3578);
not (n3593,n3594);
nand (n3594,n3595,n3702);
or (n3595,n3596,n3620);
not (n3596,n3597);
nand (n3597,n3598,n3600);
not (n3598,n3599);
xor (n3599,n3570,n3591);
not (n3600,n3601);
or (n3601,n3602,n3619);
and (n3602,n3603,n3618);
xor (n3603,n3604,n3611);
nand (n3604,n3605,n3610);
or (n3605,n3606,n893);
not (n3606,n3607);
nor (n3607,n3608,n3609);
and (n3608,n846,n903);
and (n3609,n847,n859);
nand (n3610,n1067,n3539);
nand (n3611,n3612,n3617);
or (n3612,n3613,n853);
not (n3613,n3614);
nand (n3614,n3615,n3616);
or (n3615,n887,n863);
or (n3616,n864,n935);
nand (n3617,n855,n3574);
xor (n3618,n3579,n3584);
and (n3619,n3604,n3611);
not (n3620,n3621);
nand (n3621,n3622,n3701);
or (n3622,n3623,n3647);
not (n3623,n3624);
nand (n3624,n3625,n3627);
not (n3625,n3626);
xor (n3626,n3603,n3618);
not (n3627,n3628);
or (n3628,n3629,n3646);
and (n3629,n3630,n3639);
xor (n3630,n3631,n3632);
and (n3631,n855,n887);
nand (n3632,n3633,n3638);
or (n3633,n3634,n893);
not (n3634,n3635);
nor (n3635,n3636,n3637);
and (n3636,n839,n859);
and (n3637,n841,n903);
nand (n3638,n1067,n3607);
nand (n3639,n3640,n3645);
or (n3640,n981,n3641);
not (n3641,n3642);
nor (n3642,n3643,n3644);
and (n3643,n828,n896);
and (n3644,n826,n897);
or (n3645,n3588,n982);
and (n3646,n3631,n3632);
not (n3647,n3648);
nand (n3648,n3649,n3700);
or (n3649,n3650,n3665);
nor (n3650,n3651,n3652);
xor (n3651,n3630,n3639);
and (n3652,n3653,n3659);
nor (n3653,n3654,n903);
and (n3654,n3655,n3658);
nand (n3655,n3656,n896);
not (n3656,n3657);
and (n3657,n887,n898);
nand (n3658,n935,n900);
nand (n3659,n3660,n3661);
or (n3660,n982,n3641);
nand (n3661,n3662,n1361);
nand (n3662,n3663,n3664);
or (n3663,n847,n896);
nand (n3664,n896,n847);
not (n3665,n3666);
or (n3666,n3667,n3699);
and (n3667,n3668,n3677);
xor (n3668,n3669,n3676);
nand (n3669,n3670,n3675);
or (n3670,n3671,n893);
not (n3671,n3672);
nand (n3672,n3673,n3674);
or (n3673,n903,n887);
or (n3674,n859,n935);
nand (n3675,n1067,n3635);
xor (n3676,n3653,n3659);
nand (n3677,n3678,n3698);
or (n3678,n3679,n3688);
nor (n3679,n3680,n3687);
nand (n3680,n3681,n3683);
or (n3681,n982,n3682);
not (n3682,n3662);
nand (n3683,n3684,n1361);
nand (n3684,n3685,n3686);
or (n3685,n839,n896);
nand (n3686,n896,n839);
and (n3687,n1067,n887);
nand (n3688,n3689,n3696);
nand (n3689,n3690,n3692);
or (n3690,n982,n3691);
not (n3691,n3684);
nand (n3692,n3693,n1361);
nor (n3693,n3694,n3695);
and (n3694,n935,n896);
and (n3695,n887,n897);
nor (n3696,n3697,n896);
nor (n3697,n935,n982);
nand (n3698,n3680,n3687);
and (n3699,n3669,n3676);
nand (n3700,n3651,n3652);
nand (n3701,n3626,n3628);
nand (n3702,n3599,n3601);
nand (n3703,n3568,n3521);
nand (n3704,n3705,n3707);
not (n3705,n3706);
xor (n3706,n3477,n3511);
not (n3707,n3708);
or (n3708,n3709,n3716);
and (n3709,n3710,n3715);
xor (n3710,n3711,n3714);
or (n3711,n3712,n3713);
and (n3712,n3548,n3560);
and (n3713,n3549,n3556);
xor (n3714,n3447,n3456);
xor (n3715,n3481,n3497);
and (n3716,n3711,n3714);
nand (n3717,n3718,n3720);
not (n3718,n3719);
xor (n3719,n3710,n3715);
not (n3720,n3721);
or (n3721,n3722,n3723);
and (n3722,n3522,n3547);
and (n3723,n3523,n3524);
nand (n3724,n3704,n3725);
not (n3725,n3726);
nand (n3726,n3719,n3721);
nand (n3727,n3706,n3708);
or (n3728,n3472,n3474);
nand (n3729,n3340,n3431);
nor (n3730,n3731,n3742);
nor (n3731,n3732,n3733);
xor (n3732,n3302,n3330);
or (n3733,n3734,n3741);
and (n3734,n3735,n3740);
xor (n3735,n3736,n3737);
xor (n3736,n3188,n3210);
or (n3737,n3738,n3739);
and (n3738,n3344,n3387);
and (n3739,n3345,n3363);
xor (n3740,n3306,n3309);
and (n3741,n3736,n3737);
nor (n3742,n3743,n3744);
xor (n3743,n3735,n3740);
or (n3744,n3745,n3746);
and (n3745,n3341,n3388);
and (n3746,n3342,n3343);
nor (n3747,n3748,n3752);
and (n3748,n3749,n3750);
not (n3749,n3731);
not (n3750,n3751);
nand (n3751,n3743,n3744);
and (n3752,n3732,n3733);
and (n3753,n3300,n3332);
and (n3754,n2992,n3235);
and (n3755,n3756,n3787,n3818);
or (n3756,n3757,n3758);
xor (n3757,n2890,n2969);
or (n3758,n3759,n3786);
and (n3759,n3760,n3785);
xor (n3760,n3761,n3762);
xor (n3761,n2862,n2881);
or (n3762,n3763,n3784);
and (n3763,n3764,n3777);
xor (n3764,n3765,n3776);
or (n3765,n3766,n3775);
and (n3766,n3767,n3772);
xor (n3767,n3768,n3769);
and (n3768,n3282,n3288);
or (n3769,n3770,n3771);
and (n3770,n3254,n3265);
and (n3771,n3255,n3259);
or (n3772,n3773,n3774);
and (n3773,n3243,n3250);
and (n3774,n3244,n3247);
and (n3775,n3768,n3769);
xor (n3776,n2897,n2937);
or (n3777,n3778,n3783);
and (n3778,n3779,n3782);
xor (n3779,n3780,n3781);
xor (n3780,n2917,n2930);
xor (n3781,n2900,n2908);
xor (n3782,n2939,n2952);
and (n3783,n3780,n3781);
and (n3784,n3765,n3776);
xor (n3785,n2894,n2967);
and (n3786,n3761,n3762);
nor (n3787,n3788,n3813);
nor (n3788,n3789,n3804);
xor (n3789,n3790,n3803);
xor (n3790,n3791,n3792);
xor (n3791,n2962,n2965);
or (n3792,n3793,n3802);
and (n3793,n3794,n3799);
xor (n3794,n3795,n3798);
or (n3795,n3796,n3797);
and (n3796,n3277,n3291);
and (n3797,n3278,n3281);
xor (n3798,n3767,n3772);
or (n3799,n3800,n3801);
and (n3800,n3238,n3253);
and (n3801,n3239,n3242);
and (n3802,n3795,n3798);
xor (n3803,n3764,n3777);
or (n3804,n3805,n3812);
and (n3805,n3806,n3811);
xor (n3806,n3807,n3808);
xor (n3807,n3779,n3782);
or (n3808,n3809,n3810);
and (n3809,n3272,n3294);
and (n3810,n3273,n3276);
xor (n3811,n3794,n3799);
and (n3812,n3807,n3808);
nor (n3813,n3814,n3815);
xor (n3814,n3806,n3811);
or (n3815,n3816,n3817);
and (n3816,n3236,n3271);
and (n3817,n3237,n3268);
nand (n3818,n3819,n3821);
not (n3819,n3820);
xor (n3820,n3760,n3785);
not (n3821,n3822);
or (n3822,n3823,n3824);
and (n3823,n3790,n3803);
and (n3824,n3791,n3792);
nand (n3825,n3826,n2984);
nand (n3826,n3827,n3836);
or (n3827,n3828,n3835);
nand (n3828,n3829,n3834);
or (n3829,n3830,n3832);
not (n3830,n3831);
nand (n3831,n2887,n2888);
not (n3832,n3833);
nand (n3833,n2674,n2774);
not (n3834,n2673);
not (n3835,n2971);
nand (n3836,n2973,n2981);
nand (n3837,n2671,n3838);
nand (n3838,n3839,n3849);
nand (n3839,n3840,n3756);
nand (n3840,n3841,n3848);
or (n3841,n3842,n3843);
not (n3842,n3818);
not (n3843,n3844);
nand (n3844,n3845,n3847);
or (n3845,n3788,n3846);
nand (n3846,n3814,n3815);
nand (n3847,n3789,n3804);
nand (n3848,n3820,n3822);
nand (n3849,n3757,n3758);
nand (n3850,n2985,n2988);
nand (n3851,n3852,n3862);
nand (n3852,n3853,n2662);
nand (n3853,n3854,n3861);
or (n3854,n2654,n3855);
not (n3855,n3856);
nand (n3856,n3857,n3860);
or (n3857,n3858,n3859);
not (n3858,n1979);
nand (n3859,n2306,n2308);
nand (n3860,n1981,n2295);
nand (n3861,n2655,n2656);
nand (n3862,n2312,n2645);
nand (n3863,n3864,n5021);
not (n3864,n3865);
nand (n3865,n3866,n4951);
nor (n3866,n3867,n4878);
nand (n3867,n3868,n4702);
not (n3868,n3869);
nor (n3869,n3870,n4619);
xor (n3870,n3871,n4454);
xor (n3871,n3872,n4195);
xor (n3872,n3873,n4134);
xor (n3873,n3874,n3942);
xor (n3874,n3875,n3919);
xor (n3875,n3876,n3896);
xor (n3876,n3877,n3890);
xor (n3877,n3878,n3884);
nand (n3878,n3879,n3881);
or (n3879,n3880,n963);
not (n3880,n949);
nor (n3881,n3882,n3883);
and (n3882,n192,n495);
and (n3883,n194,n494);
nand (n3884,n3885,n3889);
or (n3885,n609,n3886);
nor (n3886,n3887,n3888);
and (n3887,n188,n208);
and (n3888,n185,n210);
or (n3889,n614,n610);
nand (n3890,n3891,n3895);
or (n3891,n197,n3892);
nor (n3892,n3893,n3894);
and (n3893,n149,n230);
and (n3894,n150,n232);
or (n3895,n198,n617);
xor (n3896,n3897,n3913);
xor (n3897,n3898,n3904);
nand (n3898,n3899,n3903);
or (n3899,n18,n3900);
nor (n3900,n3901,n3902);
and (n3901,n28,n111);
and (n3902,n29,n113);
or (n3903,n647,n19);
nand (n3904,n3905,n3909);
or (n3905,n44,n3906);
nor (n3906,n3907,n3908);
and (n3907,n53,n135);
and (n3908,n54,n137);
or (n3909,n45,n3910);
nor (n3910,n3911,n3912);
and (n3911,n53,n141);
and (n3912,n54,n143);
nand (n3913,n3914,n3918);
or (n3914,n389,n3915);
nor (n3915,n3916,n3917);
and (n3916,n179,n161);
and (n3917,n180,n163);
or (n3918,n183,n600);
xor (n3919,n3920,n3936);
xor (n3920,n3921,n3930);
nand (n3921,n3922,n3926);
or (n3922,n296,n3923);
nor (n3923,n3924,n3925);
and (n3924,n305,n33);
and (n3925,n306,n35);
or (n3926,n297,n3927);
nor (n3927,n3928,n3929);
and (n3928,n305,n39);
and (n3929,n306,n41);
nand (n3930,n3931,n3935);
or (n3931,n331,n3932);
nor (n3932,n3933,n3934);
and (n3933,n21,n58);
and (n3934,n22,n60);
or (n3935,n332,n641);
nand (n3936,n3937,n3941);
or (n3937,n146,n3938);
nor (n3938,n3939,n3940);
and (n3939,n156,n84);
and (n3940,n157,n86);
or (n3941,n147,n635);
or (n3942,n3943,n4133);
and (n3943,n3944,n4078);
xor (n3944,n3945,n3979);
or (n3945,n3946,n3978);
and (n3946,n3947,n3966);
xor (n3947,n3948,n3957);
nand (n3948,n3949,n3953);
or (n3949,n219,n3950);
nor (n3950,n3951,n3952);
and (n3951,n74,n356);
and (n3952,n75,n358);
or (n3953,n220,n3954);
nor (n3954,n3955,n3956);
and (n3955,n74,n342);
and (n3956,n75,n344);
nand (n3957,n3958,n3962);
or (n3958,n122,n3959);
nor (n3959,n3960,n3961);
and (n3960,n130,n1002);
and (n3961,n131,n1004);
or (n3962,n123,n3963);
nor (n3963,n3964,n3965);
and (n3964,n1030,n130);
and (n3965,n131,n1032);
not (n3966,n3967);
nor (n3967,n3968,n3973);
and (n3968,n963,n3969);
not (n3969,n3970);
nor (n3970,n3971,n3972);
and (n3971,n494,n208);
and (n3972,n495,n210);
and (n3973,n3880,n3974);
not (n3974,n3975);
nor (n3975,n3976,n3977);
and (n3976,n494,n167);
and (n3977,n495,n169);
and (n3978,n3948,n3957);
or (n3979,n3980,n4077);
and (n3980,n3981,n4045);
xor (n3981,n3982,n4014);
or (n3982,n3983,n4013);
and (n3983,n3984,n4004);
xor (n3984,n3985,n3995);
nand (n3985,n3986,n3990);
or (n3986,n3987,n389);
nor (n3987,n3988,n3989);
and (n3988,n179,n90);
and (n3989,n180,n92);
nand (n3990,n3991,n182);
not (n3991,n3992);
nor (n3992,n3993,n3994);
and (n3993,n179,n230);
and (n3994,n180,n232);
nand (n3995,n3996,n4000);
or (n3996,n69,n3997);
nor (n3997,n3998,n3999);
and (n3998,n64,n79);
and (n3999,n66,n80);
nand (n4000,n71,n4001);
nand (n4001,n4002,n4003);
or (n4002,n80,n35);
or (n4003,n79,n33);
nand (n4004,n4005,n4009);
or (n4005,n296,n4006);
nor (n4006,n4007,n4008);
and (n4007,n305,n117);
and (n4008,n306,n119);
or (n4009,n297,n4010);
nor (n4010,n4011,n4012);
and (n4011,n305,n58);
and (n4012,n306,n60);
and (n4013,n3985,n3995);
or (n4014,n4015,n4044);
and (n4015,n4016,n4035);
xor (n4016,n4017,n4026);
nand (n4017,n4018,n4022);
or (n4018,n197,n4019);
nor (n4019,n4020,n4021);
and (n4020,n312,n150);
and (n4021,n310,n149);
or (n4022,n198,n4023);
nor (n4023,n4024,n4025);
and (n4024,n149,n84);
and (n4025,n150,n86);
nand (n4026,n4027,n4031);
or (n4027,n331,n4028);
nor (n4028,n4029,n4030);
and (n4029,n21,n141);
and (n4030,n143,n22);
or (n4031,n332,n4032);
nor (n4032,n4033,n4034);
and (n4033,n21,n111);
and (n4034,n22,n113);
nand (n4035,n4036,n4040);
or (n4036,n18,n4037);
nor (n4037,n4038,n4039);
and (n4038,n28,n448);
and (n4039,n29,n450);
or (n4040,n19,n4041);
nor (n4041,n4042,n4043);
and (n4042,n28,n135);
and (n4043,n29,n137);
and (n4044,n4017,n4026);
or (n4045,n4046,n4076);
and (n4046,n4047,n4067);
xor (n4047,n4048,n4057);
nand (n4048,n4049,n4053);
or (n4049,n853,n4050);
nor (n4050,n4051,n4052);
and (n4051,n863,n214);
and (n4052,n864,n216);
or (n4053,n870,n4054);
nor (n4054,n4055,n4056);
and (n4055,n863,n192);
and (n4056,n864,n194);
nand (n4057,n4058,n4062);
or (n4058,n146,n4059);
nor (n4059,n4060,n4061);
and (n4060,n156,n342);
and (n4061,n157,n344);
or (n4062,n147,n4063);
not (n4063,n4064);
nand (n4064,n4065,n4066);
or (n4065,n157,n350);
or (n4066,n156,n348);
nand (n4067,n4068,n4072);
or (n4068,n44,n4069);
nor (n4069,n4070,n4071);
and (n4070,n53,n625);
and (n4071,n54,n627);
or (n4072,n45,n4073);
nor (n4073,n4074,n4075);
and (n4074,n53,n474);
and (n4075,n54,n476);
and (n4076,n4048,n4057);
and (n4077,n3982,n4014);
xor (n4078,n4079,n4111);
xor (n4079,n4080,n4087);
not (n4080,n4081);
nand (n4081,n4082,n4086);
or (n4082,n609,n4083);
nor (n4083,n4084,n4085);
and (n4084,n188,n167);
and (n4085,n185,n169);
or (n4086,n614,n3886);
or (n4087,n4088,n4110);
and (n4088,n4089,n4104);
xor (n4089,n4090,n4098);
nand (n4090,n4091,n4093);
or (n4091,n4092,n69);
not (n4092,n4001);
nand (n4093,n4094,n71);
not (n4094,n4095);
nor (n4095,n4096,n4097);
and (n4096,n79,n39);
and (n4097,n80,n41);
nand (n4098,n4099,n4100);
or (n4099,n296,n4010);
or (n4100,n297,n4101);
nor (n4101,n4102,n4103);
and (n4102,n305,n64);
and (n4103,n306,n66);
nand (n4104,n4105,n4106);
or (n4105,n197,n4023);
or (n4106,n198,n4107);
nor (n4107,n4108,n4109);
and (n4108,n149,n90);
and (n4109,n150,n92);
and (n4110,n4090,n4098);
or (n4111,n4112,n4132);
and (n4112,n4113,n4126);
xor (n4113,n4114,n4120);
nand (n4114,n4115,n4116);
or (n4115,n331,n4032);
or (n4116,n332,n4117);
nor (n4117,n4118,n4119);
and (n4118,n21,n117);
and (n4119,n22,n119);
nand (n4120,n4121,n4122);
or (n4121,n18,n4041);
or (n4122,n19,n4123);
nor (n4123,n4124,n4125);
and (n4124,n28,n141);
and (n4125,n29,n143);
nand (n4126,n4127,n4131);
or (n4127,n609,n4128);
nor (n4128,n4129,n4130);
and (n4129,n188,n161);
and (n4130,n185,n163);
or (n4131,n614,n4083);
and (n4132,n4114,n4120);
and (n4133,n3945,n3979);
xor (n4134,n4135,n4192);
xor (n4135,n4136,n4162);
xor (n4136,n4137,n4156);
xor (n4137,n4138,n4147);
nand (n4138,n4139,n4143);
or (n4139,n219,n4140);
nor (n4140,n4141,n4142);
and (n4141,n74,n348);
and (n4142,n75,n350);
or (n4143,n220,n4144);
nor (n4144,n4145,n4146);
and (n4145,n74,n310);
and (n4146,n75,n312);
nand (n4147,n4148,n4152);
or (n4148,n97,n4149);
nor (n4149,n4150,n4151);
and (n4150,n474,n106);
and (n4151,n107,n476);
or (n4152,n99,n4153);
nor (n4153,n4154,n4155);
and (n4154,n448,n106);
and (n4155,n107,n450);
nand (n4156,n4157,n4161);
or (n4157,n122,n4158);
nor (n4158,n4159,n4160);
and (n4159,n1037,n130);
and (n4160,n1036,n131);
or (n4161,n123,n623);
xor (n4162,n4163,n4173);
xor (n4163,n4164,n4081);
nand (n4164,n4165,n4169);
or (n4165,n69,n4166);
nor (n4166,n4167,n4168);
and (n4167,n79,n356);
and (n4168,n80,n358);
or (n4169,n70,n4170);
nor (n4170,n4171,n4172);
and (n4171,n79,n342);
and (n4172,n80,n344);
or (n4173,n4174,n4191);
and (n4174,n4175,n4185);
xor (n4175,n4176,n4182);
nand (n4176,n4177,n4181);
or (n4177,n146,n4178);
nor (n4178,n4179,n4180);
and (n4179,n156,n310);
and (n4180,n157,n312);
or (n4181,n147,n3938);
nand (n4182,n4183,n4184);
or (n4183,n18,n4123);
or (n4184,n19,n3900);
nand (n4185,n4186,n4190);
or (n4186,n44,n4187);
nor (n4187,n4188,n4189);
and (n4188,n53,n448);
and (n4189,n54,n450);
or (n4190,n45,n3906);
and (n4191,n4176,n4182);
or (n4192,n4193,n4194);
and (n4193,n4079,n4111);
and (n4194,n4080,n4087);
xor (n4195,n4196,n4334);
xor (n4196,n4197,n4291);
or (n4197,n4198,n4290);
and (n4198,n4199,n4283);
xor (n4199,n4200,n4255);
xor (n4200,n4201,n4243);
xor (n4201,n4202,n4222);
or (n4202,n4203,n4221);
and (n4203,n4204,n4212);
xor (n4204,n4205,n4209);
nand (n4205,n4206,n4207);
or (n4206,n4063,n146);
nand (n4207,n4208,n790);
not (n4208,n4178);
nand (n4209,n4210,n4211);
or (n4210,n44,n4073);
or (n4211,n45,n4187);
nand (n4212,n4213,n4217);
or (n4213,n97,n4214);
nor (n4214,n4215,n4216);
and (n4215,n1037,n106);
and (n4216,n107,n1036);
or (n4217,n99,n4218);
nor (n4218,n4219,n4220);
and (n4219,n625,n106);
and (n4220,n627,n107);
and (n4221,n4205,n4209);
or (n4222,n4223,n4242);
and (n4223,n4224,n4235);
xor (n4224,n4225,n4228);
nand (n4225,n4226,n4227);
or (n4226,n855,n854);
not (n4227,n4054);
nand (n4228,n4229,n4230);
or (n4229,n949,n3970);
or (n4230,n950,n4231);
not (n4231,n4232);
nor (n4232,n4233,n4234);
and (n4233,n214,n495);
and (n4234,n216,n494);
nand (n4235,n4236,n4237);
or (n4236,n389,n3992);
or (n4237,n183,n4238);
not (n4238,n4239);
nand (n4239,n4240,n4241);
or (n4240,n180,n238);
or (n4241,n179,n236);
and (n4242,n4225,n4228);
xor (n4243,n4244,n4252);
xor (n4244,n4245,n4248);
nand (n4245,n4246,n4247);
or (n4246,n122,n3963);
or (n4247,n4158,n123);
nand (n4248,n4249,n4250);
or (n4249,n4238,n389);
nand (n4250,n4251,n182);
not (n4251,n3915);
nand (n4252,n4253,n4254);
or (n4253,n69,n4095);
or (n4254,n70,n4166);
or (n4255,n4256,n4282);
and (n4256,n4257,n4281);
xor (n4257,n4258,n4280);
or (n4258,n4259,n4279);
and (n4259,n4260,n4273);
xor (n4260,n4261,n4267);
nand (n4261,n4262,n4266);
or (n4262,n97,n4263);
nor (n4263,n4264,n4265);
and (n4264,n1030,n106);
and (n4265,n107,n1032);
or (n4266,n99,n4214);
nand (n4267,n4268,n4272);
or (n4268,n609,n4269);
nor (n4269,n4270,n4271);
and (n4270,n188,n236);
and (n4271,n185,n238);
or (n4272,n614,n4128);
nand (n4273,n4274,n4278);
or (n4274,n122,n4275);
nor (n4275,n4276,n4277);
and (n4276,n832,n130);
and (n4277,n834,n131);
or (n4278,n3959,n123);
and (n4279,n4261,n4267);
xor (n4280,n4089,n4104);
xor (n4281,n4224,n4235);
and (n4282,n4258,n4280);
or (n4283,n4284,n4289);
and (n4284,n4285,n4288);
xor (n4285,n4286,n4287);
xor (n4286,n4204,n4212);
xor (n4287,n4113,n4126);
xor (n4288,n3947,n3966);
and (n4289,n4286,n4287);
and (n4290,n4200,n4255);
xor (n4291,n4292,n4327);
xor (n4292,n4293,n4324);
xor (n4293,n4294,n4311);
xor (n4294,n4295,n4308);
or (n4295,n4296,n4307);
and (n4296,n4297,n4304);
xor (n4297,n4298,n4301);
nand (n4298,n4299,n4300);
or (n4299,n4231,n949);
nand (n4300,n963,n3881);
nand (n4301,n4302,n4303);
or (n4302,n219,n3954);
or (n4303,n220,n4140);
nand (n4304,n4305,n4306);
or (n4305,n97,n4218);
or (n4306,n99,n4149);
and (n4307,n4298,n4301);
or (n4308,n4309,n4310);
and (n4309,n4244,n4252);
and (n4310,n4245,n4248);
or (n4311,n4312,n4323);
and (n4312,n4313,n4320);
xor (n4313,n4314,n4317);
nand (n4314,n4315,n4316);
or (n4315,n197,n4107);
or (n4316,n198,n3892);
nand (n4317,n4318,n4319);
or (n4318,n296,n4101);
or (n4319,n297,n3923);
nand (n4320,n4321,n4322);
or (n4321,n331,n4117);
or (n4322,n332,n3932);
and (n4323,n4314,n4317);
or (n4324,n4325,n4326);
and (n4325,n4201,n4243);
and (n4326,n4202,n4222);
or (n4327,n4328,n4333);
and (n4328,n4329,n4332);
xor (n4329,n4330,n4331);
xor (n4330,n4313,n4320);
xor (n4331,n4297,n4304);
xor (n4332,n4175,n4185);
and (n4333,n4330,n4331);
or (n4334,n4335,n4453);
and (n4335,n4336,n4452);
xor (n4336,n4337,n4338);
xor (n4337,n4329,n4332);
or (n4338,n4339,n4451);
and (n4339,n4340,n4450);
xor (n4340,n4341,n4373);
or (n4341,n4342,n4372);
and (n4342,n4343,n4350);
xor (n4343,n4344,n3967);
nand (n4344,n4345,n4349);
or (n4345,n219,n4346);
nor (n4346,n4347,n4348);
and (n4347,n74,n39);
and (n4348,n75,n41);
or (n4349,n220,n3950);
or (n4350,n4351,n4371);
and (n4351,n4352,n4365);
xor (n4352,n4353,n4359);
nand (n4353,n4354,n4358);
or (n4354,n197,n4355);
nor (n4355,n4356,n4357);
and (n4356,n149,n348);
and (n4357,n150,n350);
or (n4358,n198,n4019);
nand (n4359,n4360,n4364);
or (n4360,n18,n4361);
nor (n4361,n4362,n4363);
and (n4362,n476,n29);
and (n4363,n474,n28);
or (n4364,n4037,n19);
nand (n4365,n4366,n4370);
or (n4366,n44,n4367);
nor (n4367,n4368,n4369);
and (n4368,n1037,n53);
and (n4369,n54,n1036);
or (n4370,n45,n4069);
and (n4371,n4353,n4359);
and (n4372,n4344,n3967);
or (n4373,n4374,n4449);
and (n4374,n4375,n4425);
xor (n4375,n4376,n4400);
or (n4376,n4377,n4399);
and (n4377,n4378,n4393);
xor (n4378,n4379,n4385);
nand (n4379,n4380,n4382);
or (n4380,n1067,n4381);
not (n4381,n893);
nor (n4382,n4383,n4384);
and (n4383,n192,n859);
and (n4384,n194,n903);
nand (n4385,n4386,n4391);
or (n4386,n4387,n853);
not (n4387,n4388);
nand (n4388,n4389,n4390);
or (n4389,n864,n210);
or (n4390,n863,n208);
nand (n4391,n4392,n855);
not (n4392,n4050);
nand (n4393,n4394,n4398);
or (n4394,n609,n4395);
nor (n4395,n4396,n4397);
and (n4396,n188,n230);
and (n4397,n185,n232);
or (n4398,n614,n4269);
and (n4399,n4379,n4385);
or (n4400,n4401,n4424);
and (n4401,n4402,n4418);
xor (n4402,n4403,n4411);
nand (n4403,n4404,n4405);
or (n4404,n4346,n220);
nand (n4405,n4406,n4410);
not (n4406,n4407);
nor (n4407,n4408,n4409);
and (n4408,n74,n33);
and (n4409,n75,n35);
not (n4410,n219);
nand (n4411,n4412,n4416);
or (n4412,n4413,n69);
nor (n4413,n4414,n4415);
and (n4414,n79,n58);
and (n4415,n80,n60);
nand (n4416,n4417,n71);
not (n4417,n3997);
nand (n4418,n4419,n4423);
or (n4419,n389,n4420);
nor (n4420,n4421,n4422);
and (n4421,n179,n84);
and (n4422,n180,n86);
or (n4423,n183,n3987);
and (n4424,n4403,n4411);
or (n4425,n4426,n4448);
and (n4426,n4427,n4442);
xor (n4427,n4428,n4434);
nand (n4428,n4429,n4433);
or (n4429,n296,n4430);
nor (n4430,n4431,n4432);
and (n4431,n305,n111);
and (n4432,n306,n113);
or (n4433,n297,n4006);
nand (n4434,n4435,n4439);
or (n4435,n4436,n331);
nor (n4436,n4437,n4438);
and (n4437,n21,n135);
and (n4438,n22,n137);
nand (n4439,n4440,n4441);
not (n4440,n4028);
not (n4441,n332);
nand (n4442,n4443,n4447);
or (n4443,n949,n4444);
nor (n4444,n4445,n4446);
and (n4445,n494,n161);
and (n4446,n495,n163);
or (n4447,n950,n3975);
and (n4448,n4428,n4434);
and (n4449,n4376,n4400);
xor (n4450,n3981,n4045);
and (n4451,n4341,n4373);
xor (n4452,n3944,n4078);
and (n4453,n4337,n4338);
or (n4454,n4455,n4618);
and (n4455,n4456,n4492);
xor (n4456,n4457,n4458);
xor (n4457,n4199,n4283);
or (n4458,n4459,n4491);
and (n4459,n4460,n4490);
xor (n4460,n4461,n4489);
or (n4461,n4462,n4488);
and (n4462,n4463,n4487);
xor (n4463,n4464,n4486);
or (n4464,n4465,n4485);
and (n4465,n4466,n4479);
xor (n4466,n4467,n4473);
nand (n4467,n4468,n4472);
or (n4468,n146,n4469);
nor (n4469,n4470,n4471);
and (n4470,n156,n356);
and (n4471,n157,n358);
or (n4472,n147,n4059);
nand (n4473,n4474,n4478);
or (n4474,n97,n4475);
nor (n4475,n4476,n4477);
and (n4476,n1002,n106);
and (n4477,n107,n1004);
or (n4478,n99,n4263);
nand (n4479,n4480,n4484);
or (n4480,n122,n4481);
nor (n4481,n4482,n4483);
and (n4482,n826,n130);
and (n4483,n828,n131);
or (n4484,n4275,n123);
and (n4485,n4467,n4473);
xor (n4486,n4260,n4273);
xor (n4487,n3984,n4004);
and (n4488,n4464,n4486);
xor (n4489,n4257,n4281);
xor (n4490,n4285,n4288);
and (n4491,n4461,n4489);
or (n4492,n4493,n4617);
and (n4493,n4494,n4503);
xor (n4494,n4495,n4502);
or (n4495,n4496,n4501);
and (n4496,n4497,n4500);
xor (n4497,n4498,n4499);
xor (n4498,n4047,n4067);
xor (n4499,n4016,n4035);
xor (n4500,n4343,n4350);
and (n4501,n4498,n4499);
xor (n4502,n4340,n4450);
or (n4503,n4504,n4616);
and (n4504,n4505,n4564);
xor (n4505,n4506,n4563);
or (n4506,n4507,n4562);
and (n4507,n4508,n4540);
xor (n4508,n4509,n4517);
not (n4509,n4510);
nor (n4510,n4511,n4516);
and (n4511,n4381,n4512);
not (n4512,n4513);
nor (n4513,n4514,n4515);
and (n4514,n903,n214);
and (n4515,n859,n216);
and (n4516,n1067,n4382);
or (n4517,n4518,n4539);
and (n4518,n4519,n4532);
xor (n4519,n4520,n4526);
nand (n4520,n4521,n4522);
or (n4521,n4387,n870);
nand (n4522,n854,n4523);
nand (n4523,n4524,n4525);
or (n4524,n864,n169);
or (n4525,n863,n167);
nand (n4526,n4527,n4531);
or (n4527,n609,n4528);
nor (n4528,n4529,n4530);
and (n4529,n188,n90);
and (n4530,n185,n92);
or (n4531,n614,n4395);
nand (n4532,n4533,n4538);
or (n4533,n219,n4534);
not (n4534,n4535);
nand (n4535,n4536,n4537);
or (n4536,n75,n66);
or (n4537,n74,n64);
or (n4538,n220,n4407);
and (n4539,n4520,n4526);
or (n4540,n4541,n4561);
and (n4541,n4542,n4555);
xor (n4542,n4543,n4549);
nand (n4543,n4544,n4548);
or (n4544,n69,n4545);
nor (n4545,n4546,n4547);
and (n4546,n79,n117);
and (n4547,n80,n119);
or (n4548,n70,n4413);
nand (n4549,n4550,n4554);
or (n4550,n4551,n389);
nor (n4551,n4552,n4553);
and (n4552,n179,n310);
and (n4553,n180,n312);
or (n4554,n183,n4420);
nand (n4555,n4556,n4560);
or (n4556,n296,n4557);
nor (n4557,n4558,n4559);
and (n4558,n305,n141);
and (n4559,n306,n143);
or (n4560,n297,n4430);
and (n4561,n4543,n4549);
and (n4562,n4509,n4517);
xor (n4563,n4375,n4425);
or (n4564,n4565,n4615);
and (n4565,n4566,n4614);
xor (n4566,n4567,n4591);
or (n4567,n4568,n4590);
and (n4568,n4569,n4584);
xor (n4569,n4570,n4576);
nand (n4570,n4571,n4575);
or (n4571,n331,n4572);
nor (n4572,n4573,n4574);
and (n4573,n21,n448);
and (n4574,n22,n450);
or (n4575,n332,n4436);
nand (n4576,n4577,n4582);
or (n4577,n4578,n949);
not (n4578,n4579);
nand (n4579,n4580,n4581);
or (n4580,n495,n238);
or (n4581,n494,n236);
nand (n4582,n4583,n963);
not (n4583,n4444);
nand (n4584,n4585,n4589);
or (n4585,n197,n4586);
nor (n4586,n4587,n4588);
and (n4587,n149,n342);
and (n4588,n150,n344);
or (n4589,n198,n4355);
and (n4590,n4570,n4576);
or (n4591,n4592,n4613);
and (n4592,n4593,n4607);
xor (n4593,n4594,n4600);
nand (n4594,n4595,n4599);
or (n4595,n18,n4596);
nor (n4596,n4597,n4598);
and (n4597,n28,n625);
and (n4598,n29,n627);
or (n4599,n4361,n19);
nand (n4600,n4601,n4606);
or (n4601,n4602,n44);
not (n4602,n4603);
nand (n4603,n4604,n4605);
or (n4604,n54,n1032);
or (n4605,n53,n1030);
or (n4606,n4367,n45);
nand (n4607,n4608,n4612);
or (n4608,n146,n4609);
nor (n4609,n4610,n4611);
and (n4610,n156,n39);
and (n4611,n157,n41);
or (n4612,n147,n4469);
and (n4613,n4594,n4600);
xor (n4614,n4402,n4418);
and (n4615,n4567,n4591);
and (n4616,n4506,n4563);
and (n4617,n4495,n4502);
and (n4618,n4457,n4458);
or (n4619,n4620,n4701);
and (n4620,n4621,n4624);
xor (n4621,n4622,n4623);
xor (n4622,n4336,n4452);
xor (n4623,n4456,n4492);
or (n4624,n4625,n4700);
and (n4625,n4626,n4699);
xor (n4626,n4627,n4698);
or (n4627,n4628,n4697);
and (n4628,n4629,n4638);
xor (n4629,n4630,n4637);
or (n4630,n4631,n4636);
and (n4631,n4632,n4635);
xor (n4632,n4633,n4634);
xor (n4633,n4466,n4479);
xor (n4634,n4378,n4393);
xor (n4635,n4352,n4365);
and (n4636,n4633,n4634);
xor (n4637,n4463,n4487);
or (n4638,n4639,n4696);
and (n4639,n4640,n4658);
xor (n4640,n4641,n4642);
xor (n4641,n4427,n4442);
or (n4642,n4643,n4657);
and (n4643,n4644,n4510);
xor (n4644,n4645,n4651);
nand (n4645,n4646,n4650);
or (n4646,n97,n4647);
nor (n4647,n4648,n4649);
and (n4648,n832,n106);
and (n4649,n834,n107);
or (n4650,n99,n4475);
nand (n4651,n4652,n4656);
or (n4652,n122,n4653);
nor (n4653,n4654,n4655);
and (n4654,n847,n130);
and (n4655,n846,n131);
or (n4656,n123,n4481);
and (n4657,n4645,n4651);
or (n4658,n4659,n4695);
and (n4659,n4660,n4681);
xor (n4660,n4661,n4668);
or (n4661,n4662,n4665);
nand (n4662,n4663,n4664);
or (n4663,n893,n2584);
or (n4664,n894,n4513);
nand (n4665,n4666,n4667);
or (n4666,n1361,n983);
not (n4667,n2523);
or (n4668,n4669,n4680);
and (n4669,n4670,n4677);
xor (n4670,n4671,n4674);
nand (n4671,n4672,n4673);
or (n4672,n949,n2592);
nand (n4673,n963,n4579);
nand (n4674,n4675,n4676);
or (n4675,n122,n2601);
or (n4676,n4653,n123);
nand (n4677,n4678,n4679);
or (n4678,n146,n2610);
or (n4679,n147,n4609);
and (n4680,n4671,n4674);
or (n4681,n4682,n4694);
and (n4682,n4683,n4691);
xor (n4683,n4684,n4688);
nand (n4684,n4685,n4686);
or (n4685,n4534,n220);
nand (n4686,n4687,n4410);
not (n4687,n2616);
nand (n4688,n4689,n4690);
or (n4689,n609,n2622);
or (n4690,n614,n4528);
nand (n4691,n4692,n4693);
or (n4692,n69,n2326);
or (n4693,n70,n4545);
and (n4694,n4684,n4688);
and (n4695,n4661,n4668);
and (n4696,n4641,n4642);
and (n4697,n4630,n4637);
xor (n4698,n4460,n4490);
xor (n4699,n4494,n4503);
and (n4700,n4627,n4698);
and (n4701,n4622,n4623);
nor (n4702,n4703,n4873);
nor (n4703,n4704,n4864);
or (n4704,n4705,n4863);
and (n4705,n4706,n4820);
xor (n4706,n4707,n4797);
or (n4707,n4708,n4796);
and (n4708,n4709,n4789);
xor (n4709,n4710,n4739);
or (n4710,n4711,n4738);
and (n4711,n4712,n4725);
xor (n4712,n4713,n4714);
xor (n4713,n4644,n4510);
or (n4714,n4715,n4724);
and (n4715,n4716,n4723);
xor (n4716,n4717,n4720);
nand (n4717,n4718,n4719);
or (n4718,n2568,n44);
nand (n4719,n46,n4603);
nand (n4720,n4721,n4722);
or (n4721,n97,n2574);
or (n4722,n99,n4647);
and (n4723,n2510,n2516);
and (n4724,n4717,n4720);
or (n4725,n4726,n4737);
and (n4726,n4727,n4734);
xor (n4727,n4728,n4731);
or (n4728,n4729,n4730);
and (n4729,n2578,n2595);
and (n4730,n2579,n2587);
or (n4731,n4732,n4733);
and (n4732,n2605,n2619);
and (n4733,n2606,n2613);
or (n4734,n4735,n4736);
and (n4735,n2319,n2338);
and (n4736,n2320,n2329);
and (n4737,n4728,n4731);
and (n4738,n4713,n4714);
or (n4739,n4740,n4788);
and (n4740,n4741,n4757);
xor (n4741,n4742,n4756);
or (n4742,n4743,n4755);
and (n4743,n4744,n4751);
xor (n4744,n4745,n4748);
or (n4745,n4746,n4747);
and (n4746,n2348,n2367);
and (n4747,n2349,n2358);
or (n4748,n4749,n4750);
and (n4749,n2558,n2571);
and (n4750,n2559,n2565);
nand (n4751,n4752,n4661);
or (n4752,n4753,n4754);
not (n4753,n4665);
not (n4754,n4662);
and (n4755,n4745,n4748);
xor (n4756,n4660,n4681);
xor (n4757,n4758,n4787);
xor (n4758,n4759,n4773);
or (n4759,n4760,n4772);
and (n4760,n4761,n4769);
xor (n4761,n4762,n4765);
nand (n4762,n4763,n4764);
or (n4763,n296,n2335);
or (n4764,n297,n4557);
nand (n4765,n4766,n4767);
or (n4766,n853,n2344);
or (n4767,n870,n4768);
not (n4768,n4523);
nand (n4769,n4770,n4771);
or (n4770,n389,n2355);
or (n4771,n183,n4551);
and (n4772,n4762,n4765);
or (n4773,n4774,n4786);
and (n4774,n4775,n4782);
xor (n4775,n4776,n4779);
nand (n4776,n4777,n4778);
or (n4777,n331,n2364);
or (n4778,n332,n4572);
nand (n4779,n4780,n4781);
or (n4780,n18,n2373);
or (n4781,n19,n4596);
nand (n4782,n4783,n4785);
or (n4783,n4784,n197);
not (n4784,n2562);
or (n4785,n198,n4586);
and (n4786,n4776,n4779);
xor (n4787,n4519,n4532);
and (n4788,n4742,n4756);
xor (n4789,n4790,n4793);
xor (n4790,n4791,n4792);
xor (n4791,n4508,n4540);
xor (n4792,n4566,n4614);
or (n4793,n4794,n4795);
and (n4794,n4758,n4787);
and (n4795,n4759,n4773);
and (n4796,n4710,n4739);
xor (n4797,n4798,n4813);
xor (n4798,n4799,n4800);
xor (n4799,n4629,n4638);
or (n4800,n4801,n4812);
and (n4801,n4802,n4811);
xor (n4802,n4803,n4810);
or (n4803,n4804,n4809);
and (n4804,n4805,n4808);
xor (n4805,n4806,n4807);
xor (n4806,n4593,n4607);
xor (n4807,n4542,n4555);
xor (n4808,n4569,n4584);
and (n4809,n4806,n4807);
xor (n4810,n4632,n4635);
xor (n4811,n4640,n4658);
and (n4812,n4803,n4810);
xor (n4813,n4814,n4819);
xor (n4814,n4815,n4816);
xor (n4815,n4497,n4500);
or (n4816,n4817,n4818);
and (n4817,n4790,n4793);
and (n4818,n4791,n4792);
xor (n4819,n4505,n4564);
or (n4820,n4821,n4862);
and (n4821,n4822,n4837);
xor (n4822,n4823,n4824);
xor (n4823,n4802,n4811);
or (n4824,n4825,n4836);
and (n4825,n4826,n4835);
xor (n4826,n4827,n4834);
or (n4827,n4828,n4833);
and (n4828,n4829,n4832);
xor (n4829,n4830,n4831);
xor (n4830,n4683,n4691);
xor (n4831,n4761,n4769);
xor (n4832,n4775,n4782);
and (n4833,n4830,n4831);
xor (n4834,n4805,n4808);
xor (n4835,n4712,n4725);
and (n4836,n4827,n4834);
or (n4837,n4838,n4861);
and (n4838,n4839,n4860);
xor (n4839,n4840,n4849);
or (n4840,n4841,n4848);
and (n4841,n4842,n4845);
xor (n4842,n4843,n4844);
xor (n4843,n4670,n4677);
xor (n4844,n4716,n4723);
or (n4845,n4846,n4847);
and (n4846,n2468,n2486);
and (n4847,n2469,n2472);
and (n4848,n4843,n4844);
or (n4849,n4850,n4859);
and (n4850,n4851,n4858);
xor (n4851,n4852,n4855);
or (n4852,n4853,n4854);
and (n4853,n2508,n2540);
and (n4854,n2509,n2526);
or (n4855,n4856,n4857);
and (n4856,n2556,n2604);
and (n4857,n2557,n2577);
xor (n4858,n4744,n4751);
and (n4859,n4852,n4855);
xor (n4860,n4741,n4757);
and (n4861,n4840,n4849);
and (n4862,n4823,n4824);
and (n4863,n4707,n4797);
xor (n4864,n4865,n4870);
xor (n4865,n4866,n4869);
or (n4866,n4867,n4868);
and (n4867,n4814,n4819);
and (n4868,n4815,n4816);
xor (n4869,n4626,n4699);
or (n4870,n4871,n4872);
and (n4871,n4798,n4813);
and (n4872,n4799,n4800);
nor (n4873,n4874,n4875);
xor (n4874,n4621,n4624);
or (n4875,n4876,n4877);
and (n4876,n4865,n4870);
and (n4877,n4866,n4869);
nor (n4878,n4879,n4882);
or (n4879,n4880,n4881);
and (n4880,n3871,n4454);
and (n4881,n3872,n4195);
xor (n4882,n4883,n4948);
xor (n4883,n4884,n4921);
xor (n4884,n4885,n4896);
xor (n4885,n4886,n4893);
xor (n4886,n4887,n4892);
xor (n4887,n4888,n4891);
or (n4888,n4889,n4890);
and (n4889,n3920,n3936);
and (n4890,n3921,n3930);
xor (n4891,n606,n621);
xor (n4892,n632,n645);
or (n4893,n4894,n4895);
and (n4894,n4135,n4192);
and (n4895,n4136,n4162);
xor (n4896,n4897,n4918);
xor (n4897,n4898,n4909);
xor (n4898,n4899,n4906);
xor (n4899,n4900,n4903);
nand (n4900,n4901,n4902);
or (n4901,n219,n4144);
or (n4902,n220,n538);
nand (n4903,n4904,n4905);
or (n4904,n44,n3910);
or (n4905,n45,n556);
nand (n4906,n4907,n4908);
or (n4907,n97,n4153);
or (n4908,n99,n562);
xor (n4909,n4910,n4917);
xor (n4910,n4911,n4914);
nand (n4911,n4912,n4913);
or (n4912,n69,n4170);
or (n4913,n70,n466);
nand (n4914,n4915,n4916);
or (n4915,n296,n3927);
or (n4916,n297,n480);
not (n4917,n598);
or (n4918,n4919,n4920);
and (n4919,n4294,n4311);
and (n4920,n4295,n4308);
xor (n4921,n4922,n4945);
xor (n4922,n4923,n4926);
or (n4923,n4924,n4925);
and (n4924,n4292,n4327);
and (n4925,n4293,n4324);
xor (n4926,n4927,n4942);
xor (n4927,n4928,n4931);
or (n4928,n4929,n4930);
and (n4929,n4163,n4173);
and (n4930,n4164,n4081);
xor (n4931,n4932,n4939);
xor (n4932,n4933,n4936);
or (n4933,n4934,n4935);
and (n4934,n3897,n3913);
and (n4935,n3898,n3904);
or (n4936,n4937,n4938);
and (n4937,n4137,n4156);
and (n4938,n4138,n4147);
or (n4939,n4940,n4941);
and (n4940,n3877,n3890);
and (n4941,n3878,n3884);
or (n4942,n4943,n4944);
and (n4943,n3875,n3919);
and (n4944,n3876,n3896);
or (n4945,n4946,n4947);
and (n4946,n3873,n4134);
and (n4947,n3874,n3942);
or (n4948,n4949,n4950);
and (n4949,n4196,n4334);
and (n4950,n4197,n4291);
nor (n4951,n4952,n5002);
not (n4952,n4953);
nor (n4953,n4954,n4987);
nor (n4954,n4955,n4956);
xor (n4955,n4706,n4820);
or (n4956,n4957,n4986);
and (n4957,n4958,n4961);
xor (n4958,n4959,n4960);
xor (n4959,n4709,n4789);
xor (n4960,n4822,n4837);
or (n4961,n4962,n4985);
and (n4962,n4963,n4974);
xor (n4963,n4964,n4965);
xor (n4964,n4826,n4835);
or (n4965,n4966,n4973);
and (n4966,n4967,n4970);
xor (n4967,n4968,n4969);
xor (n4968,n4727,n4734);
xor (n4969,n4829,n4832);
or (n4970,n4971,n4972);
and (n4971,n2317,n2376);
and (n4972,n2318,n2347);
and (n4973,n4968,n4969);
or (n4974,n4975,n4984);
and (n4975,n4976,n4981);
xor (n4976,n4977,n4978);
xor (n4977,n4842,n4845);
or (n4978,n4979,n4980);
and (n4979,n2463,n2507);
and (n4980,n2464,n2467);
or (n4981,n4982,n4983);
and (n4982,n2544,n2555);
and (n4983,n2545,n2552);
and (n4984,n4977,n4978);
and (n4985,n4964,n4965);
and (n4986,n4959,n4960);
nor (n4987,n4988,n5001);
or (n4988,n4989,n5000);
and (n4989,n4990,n4993);
xor (n4990,n4991,n4992);
xor (n4991,n4839,n4860);
xor (n4992,n4963,n4974);
or (n4993,n4994,n4999);
and (n4994,n4995,n4998);
xor (n4995,n4996,n4997);
xor (n4996,n4851,n4858);
xor (n4997,n4967,n4970);
xor (n4998,n4976,n4981);
and (n4999,n4996,n4997);
and (n5000,n4991,n4992);
xor (n5001,n4958,n4961);
or (n5002,n5003,n5016);
nor (n5003,n5004,n5007);
or (n5004,n5005,n5006);
and (n5005,n2313,n2636);
and (n5006,n2314,n2460);
xor (n5007,n5008,n5015);
xor (n5008,n5009,n5012);
or (n5009,n5010,n5011);
and (n5010,n2315,n2411);
and (n5011,n2316,n2389);
or (n5012,n5013,n5014);
and (n5013,n2461,n2625);
and (n5014,n2462,n2543);
xor (n5015,n4995,n4998);
nor (n5016,n5017,n5018);
xor (n5017,n4990,n4993);
or (n5018,n5019,n5020);
and (n5019,n5008,n5015);
and (n5020,n5009,n5012);
not (n5021,n5022);
nand (n5022,n5023,n5112);
and (n5023,n5024,n5097);
nor (n5024,n5025,n5070);
nor (n5025,n5026,n5029);
or (n5026,n5027,n5028);
and (n5027,n4883,n4948);
and (n5028,n4884,n4921);
xor (n5029,n5030,n5067);
xor (n5030,n5031,n5050);
xor (n5031,n5032,n5047);
xor (n5032,n5033,n5040);
xor (n5033,n5034,n5039);
xor (n5034,n5035,n5038);
or (n5035,n5036,n5037);
and (n5036,n4899,n4906);
and (n5037,n4900,n4903);
xor (n5038,n553,n566);
xor (n5039,n463,n478);
xor (n5040,n5041,n5044);
xor (n5041,n5042,n5043);
xor (n5042,n487,n511);
xor (n5043,n520,n536);
or (n5044,n5045,n5046);
and (n5045,n4910,n4917);
and (n5046,n4911,n4914);
or (n5047,n5048,n5049);
and (n5048,n4897,n4918);
and (n5049,n4898,n4909);
xor (n5050,n5051,n5064);
xor (n5051,n5052,n5055);
or (n5052,n5053,n5054);
and (n5053,n4927,n4942);
and (n5054,n4928,n4931);
xor (n5055,n5056,n5063);
xor (n5056,n5057,n5060);
or (n5057,n5058,n5059);
and (n5058,n4932,n4939);
and (n5059,n4933,n4936);
or (n5060,n5061,n5062);
and (n5061,n4887,n4892);
and (n5062,n4888,n4891);
xor (n5063,n597,n630);
or (n5064,n5065,n5066);
and (n5065,n4885,n4896);
and (n5066,n4886,n4893);
or (n5067,n5068,n5069);
and (n5068,n4922,n4945);
and (n5069,n4923,n4926);
nor (n5070,n5071,n5074);
or (n5071,n5072,n5073);
and (n5072,n5030,n5067);
and (n5073,n5031,n5050);
xor (n5074,n5075,n5094);
xor (n5075,n5076,n5085);
xor (n5076,n5077,n5084);
xor (n5077,n5078,n5081);
or (n5078,n5079,n5080);
and (n5079,n5034,n5039);
and (n5080,n5035,n5038);
or (n5081,n5082,n5083);
and (n5082,n5041,n5044);
and (n5083,n5042,n5043);
xor (n5084,n581,n584);
xor (n5085,n5086,n5091);
xor (n5086,n5087,n5088);
xor (n5087,n594,n654);
or (n5088,n5089,n5090);
and (n5089,n5056,n5063);
and (n5090,n5057,n5060);
or (n5091,n5092,n5093);
and (n5092,n5032,n5047);
and (n5093,n5033,n5040);
or (n5094,n5095,n5096);
and (n5095,n5051,n5064);
and (n5096,n5052,n5055);
nand (n5097,n5098,n5108);
not (n5098,n5099);
xor (n5099,n5100,n5105);
xor (n5100,n5101,n5104);
or (n5101,n5102,n5103);
and (n5102,n5077,n5084);
and (n5103,n5078,n5081);
xor (n5104,n590,n656);
or (n5105,n5106,n5107);
and (n5106,n5086,n5091);
and (n5107,n5087,n5088);
not (n5108,n5109);
or (n5109,n5110,n5111);
and (n5110,n5075,n5094);
and (n5111,n5076,n5085);
nand (n5112,n5113,n5117);
not (n5113,n5114);
or (n5114,n5115,n5116);
and (n5115,n5100,n5105);
and (n5116,n5101,n5104);
not (n5117,n5118);
xor (n5118,n8,n588);
nand (n5119,n5120,n5147);
or (n5120,n5022,n5121);
not (n5121,n5122);
nand (n5122,n5123,n5137,n5146);
nand (n5123,n3866,n5124);
nand (n5124,n5125,n5131);
or (n5125,n4952,n5126);
not (n5126,n5127);
nand (n5127,n5128,n5130);
or (n5128,n5016,n5129);
nand (n5129,n5004,n5007);
nand (n5130,n5017,n5018);
nor (n5131,n5132,n5136);
and (n5132,n5133,n5134);
not (n5133,n4954);
not (n5134,n5135);
nand (n5135,n4988,n5001);
and (n5136,n4955,n4956);
nand (n5137,n5138,n5145);
nand (n5138,n5139,n5144);
or (n5139,n5140,n3869);
nor (n5140,n5141,n5143);
nor (n5141,n4873,n5142);
nand (n5142,n4864,n4704);
and (n5143,n4874,n4875);
nand (n5144,n3870,n4619);
not (n5145,n4878);
nand (n5146,n4879,n4882);
not (n5147,n5148);
nand (n5148,n5149,n5161);
or (n5149,n5150,n5151);
not (n5150,n5112);
not (n5151,n5152);
nand (n5152,n5153,n5160);
or (n5153,n5154,n5155);
not (n5154,n5097);
not (n5155,n5156);
nand (n5156,n5157,n5159);
or (n5157,n5158,n5070);
nand (n5158,n5026,n5029);
nand (n5159,n5071,n5074);
nand (n5160,n5099,n5109);
or (n5161,n5113,n5117);
or (n5162,n762,n3);
xor (n5163,n5164,n10060);
xor (n5164,n5165,n10413);
xor (n5165,n5166,n10055);
xor (n5166,n5167,n10406);
xor (n5167,n5168,n10049);
xor (n5168,n5169,n10394);
xor (n5169,n5170,n10043);
xor (n5170,n5171,n10377);
xor (n5171,n5172,n10037);
xor (n5172,n5173,n10355);
xor (n5173,n5174,n10031);
xor (n5174,n5175,n10328);
xor (n5175,n5176,n10025);
xor (n5176,n5177,n10296);
xor (n5177,n5178,n10019);
xor (n5178,n5179,n10259);
xor (n5179,n5180,n10013);
xor (n5180,n5181,n10217);
xor (n5181,n5182,n10007);
xor (n5182,n5183,n10170);
xor (n5183,n5184,n10001);
xor (n5184,n5185,n10118);
xor (n5185,n5186,n9995);
xor (n5186,n5187,n10061);
xor (n5187,n5188,n9989);
xor (n5188,n5189,n9986);
xor (n5189,n5190,n9985);
xor (n5190,n5191,n9905);
xor (n5191,n5192,n9904);
xor (n5192,n5193,n9817);
xor (n5193,n5194,n9816);
xor (n5194,n5195,n9724);
xor (n5195,n5196,n9723);
xor (n5196,n5197,n9624);
xor (n5197,n5198,n9623);
xor (n5198,n5199,n9519);
xor (n5199,n5200,n9518);
xor (n5200,n5201,n9408);
xor (n5201,n5202,n9407);
xor (n5202,n5203,n9291);
xor (n5203,n5204,n9290);
xor (n5204,n5205,n9167);
xor (n5205,n5206,n9166);
xor (n5206,n5207,n9038);
xor (n5207,n5208,n9037);
xor (n5208,n5209,n8902);
xor (n5209,n5210,n8901);
xor (n5210,n5211,n8761);
xor (n5211,n5212,n8760);
xor (n5212,n5213,n8616);
xor (n5213,n5214,n8615);
xor (n5214,n5215,n8463);
xor (n5215,n5216,n8462);
xor (n5216,n5217,n8303);
xor (n5217,n5218,n8302);
xor (n5218,n5219,n8138);
xor (n5219,n5220,n8137);
xor (n5220,n5221,n7972);
xor (n5221,n5222,n7971);
xor (n5222,n5223,n7795);
xor (n5223,n5224,n7794);
xor (n5224,n5225,n7611);
xor (n5225,n5226,n7610);
xor (n5226,n5227,n7423);
xor (n5227,n5228,n7422);
xor (n5228,n5229,n7230);
xor (n5229,n5230,n7229);
xor (n5230,n5231,n7032);
xor (n5231,n5232,n7031);
xor (n5232,n5233,n6832);
xor (n5233,n5234,n6831);
xor (n5234,n5235,n6265);
xor (n5235,n5236,n6264);
xor (n5236,n5237,n6239);
xor (n5237,n5238,n3882);
xor (n5238,n5239,n6214);
xor (n5239,n5240,n6213);
xor (n5240,n5241,n6007);
xor (n5241,n5242,n6006);
xor (n5242,n5243,n5797);
xor (n5243,n5244,n5796);
xor (n5244,n5245,n5255);
xor (n5245,n5246,n4383);
xor (n5246,n5247,n5254);
xor (n5247,n5248,n5253);
xor (n5248,n5249,n5252);
xor (n5249,n5250,n5251);
and (n5250,n192,n983);
and (n5251,n192,n897);
and (n5252,n5250,n5251);
and (n5253,n192,n898);
and (n5254,n5248,n5253);
or (n5255,n5256,n5257);
and (n5256,n5246,n4383);
and (n5257,n5245,n5258);
or (n5258,n5256,n5259);
and (n5259,n5245,n5260);
or (n5260,n5256,n5261);
and (n5261,n5245,n5262);
or (n5262,n5256,n5263);
and (n5263,n5245,n5264);
or (n5264,n5265,1'b0);
or (n5265,n5256,n5266);
and (n5266,n5245,n5267);
or (n5267,n5268,n5626);
and (n5268,n5269,n5625);
xor (n5269,n5247,n5270);
or (n5270,n5271,n5447);
and (n5271,n5272,n5446);
xor (n5272,n5249,n5273);
or (n5273,n5274,n5275);
and (n5274,n5250,n2521);
and (n5275,n5276,n5277);
xor (n5276,n5250,n2521);
or (n5277,n5278,n5280);
and (n5278,n5279,n2171);
and (n5279,n214,n983);
and (n5280,n5281,n5282);
xor (n5281,n5279,n2171);
or (n5282,n5283,n5286);
and (n5283,n5284,n5285);
and (n5284,n208,n983);
and (n5285,n167,n897);
and (n5286,n5287,n5288);
xor (n5287,n5284,n5285);
or (n5288,n5289,n5292);
and (n5289,n5290,n5291);
and (n5290,n167,n983);
and (n5291,n161,n897);
and (n5292,n5293,n5294);
xor (n5293,n5290,n5291);
or (n5294,n5295,n5298);
and (n5295,n5296,n5297);
and (n5296,n161,n983);
and (n5297,n236,n897);
and (n5298,n5299,n5300);
xor (n5299,n5296,n5297);
or (n5300,n5301,n5304);
and (n5301,n5302,n5303);
and (n5302,n236,n983);
and (n5303,n230,n897);
and (n5304,n5305,n5306);
xor (n5305,n5302,n5303);
or (n5306,n5307,n5310);
and (n5307,n5308,n5309);
and (n5308,n230,n983);
and (n5309,n90,n897);
and (n5310,n5311,n5312);
xor (n5311,n5308,n5309);
or (n5312,n5313,n5315);
and (n5313,n5314,n1248);
and (n5314,n90,n983);
and (n5315,n5316,n5317);
xor (n5316,n5314,n1248);
or (n5317,n5318,n5321);
and (n5318,n5319,n5320);
and (n5319,n84,n983);
and (n5320,n310,n897);
and (n5321,n5322,n5323);
xor (n5322,n5319,n5320);
or (n5323,n5324,n5327);
and (n5324,n5325,n5326);
and (n5325,n310,n983);
and (n5326,n348,n897);
and (n5327,n5328,n5329);
xor (n5328,n5325,n5326);
or (n5329,n5330,n5332);
and (n5330,n5331,n1648);
and (n5331,n348,n983);
and (n5332,n5333,n5334);
xor (n5333,n5331,n1648);
or (n5334,n5335,n5338);
and (n5335,n5336,n5337);
and (n5336,n342,n983);
and (n5337,n356,n897);
and (n5338,n5339,n5340);
xor (n5339,n5336,n5337);
or (n5340,n5341,n5343);
and (n5341,n5342,n1879);
and (n5342,n356,n983);
and (n5343,n5344,n5345);
xor (n5344,n5342,n1879);
or (n5345,n5346,n5348);
and (n5346,n5347,n2692);
and (n5347,n39,n983);
and (n5348,n5349,n5350);
xor (n5349,n5347,n2692);
or (n5350,n5351,n5354);
and (n5351,n5352,n5353);
and (n5352,n33,n983);
and (n5353,n64,n897);
and (n5354,n5355,n5356);
xor (n5355,n5352,n5353);
or (n5356,n5357,n5360);
and (n5357,n5358,n5359);
and (n5358,n64,n983);
and (n5359,n58,n897);
and (n5360,n5361,n5362);
xor (n5361,n5358,n5359);
or (n5362,n5363,n5366);
and (n5363,n5364,n5365);
and (n5364,n58,n983);
and (n5365,n117,n897);
and (n5366,n5367,n5368);
xor (n5367,n5364,n5365);
or (n5368,n5369,n5372);
and (n5369,n5370,n5371);
and (n5370,n117,n983);
and (n5371,n111,n897);
and (n5372,n5373,n5374);
xor (n5373,n5370,n5371);
or (n5374,n5375,n5378);
and (n5375,n5376,n5377);
and (n5376,n111,n983);
and (n5377,n141,n897);
and (n5378,n5379,n5380);
xor (n5379,n5376,n5377);
or (n5380,n5381,n5384);
and (n5381,n5382,n5383);
and (n5382,n141,n983);
and (n5383,n135,n897);
and (n5384,n5385,n5386);
xor (n5385,n5382,n5383);
or (n5386,n5387,n5390);
and (n5387,n5388,n5389);
and (n5388,n135,n983);
and (n5389,n448,n897);
and (n5390,n5391,n5392);
xor (n5391,n5388,n5389);
or (n5392,n5393,n5396);
and (n5393,n5394,n5395);
and (n5394,n448,n983);
and (n5395,n474,n897);
and (n5396,n5397,n5398);
xor (n5397,n5394,n5395);
or (n5398,n5399,n5402);
and (n5399,n5400,n5401);
and (n5400,n474,n983);
and (n5401,n625,n897);
and (n5402,n5403,n5404);
xor (n5403,n5400,n5401);
or (n5404,n5405,n5408);
and (n5405,n5406,n5407);
and (n5406,n625,n983);
and (n5407,n1037,n897);
and (n5408,n5409,n5410);
xor (n5409,n5406,n5407);
or (n5410,n5411,n5414);
and (n5411,n5412,n5413);
and (n5412,n1037,n983);
and (n5413,n1030,n897);
and (n5414,n5415,n5416);
xor (n5415,n5412,n5413);
or (n5416,n5417,n5419);
and (n5417,n5418,n3533);
and (n5418,n1030,n983);
and (n5419,n5420,n5421);
xor (n5420,n5418,n3533);
or (n5421,n5422,n5425);
and (n5422,n5423,n5424);
and (n5423,n1002,n983);
and (n5424,n832,n897);
and (n5425,n5426,n5427);
xor (n5426,n5423,n5424);
or (n5427,n5428,n5430);
and (n5428,n5429,n3644);
and (n5429,n832,n983);
and (n5430,n5431,n5432);
xor (n5431,n5429,n3644);
or (n5432,n5433,n5436);
and (n5433,n5434,n5435);
and (n5434,n826,n983);
and (n5435,n847,n897);
and (n5436,n5437,n5438);
xor (n5437,n5434,n5435);
or (n5438,n5439,n5442);
and (n5439,n5440,n5441);
and (n5440,n847,n983);
and (n5441,n839,n897);
and (n5442,n5443,n5444);
xor (n5443,n5440,n5441);
and (n5444,n5445,n3695);
and (n5445,n839,n983);
and (n5446,n214,n898);
and (n5447,n5448,n5449);
xor (n5448,n5272,n5446);
or (n5449,n5450,n5453);
and (n5450,n5451,n5452);
xor (n5451,n5276,n5277);
and (n5452,n208,n898);
and (n5453,n5454,n5455);
xor (n5454,n5451,n5452);
or (n5455,n5456,n5459);
and (n5456,n5457,n5458);
xor (n5457,n5281,n5282);
and (n5458,n167,n898);
and (n5459,n5460,n5461);
xor (n5460,n5457,n5458);
or (n5461,n5462,n5465);
and (n5462,n5463,n5464);
xor (n5463,n5287,n5288);
and (n5464,n161,n898);
and (n5465,n5466,n5467);
xor (n5466,n5463,n5464);
or (n5467,n5468,n5471);
and (n5468,n5469,n5470);
xor (n5469,n5293,n5294);
and (n5470,n236,n898);
and (n5471,n5472,n5473);
xor (n5472,n5469,n5470);
or (n5473,n5474,n5477);
and (n5474,n5475,n5476);
xor (n5475,n5299,n5300);
and (n5476,n230,n898);
and (n5477,n5478,n5479);
xor (n5478,n5475,n5476);
or (n5479,n5480,n5483);
and (n5480,n5481,n5482);
xor (n5481,n5305,n5306);
and (n5482,n90,n898);
and (n5483,n5484,n5485);
xor (n5484,n5481,n5482);
or (n5485,n5486,n5489);
and (n5486,n5487,n5488);
xor (n5487,n5311,n5312);
and (n5488,n84,n898);
and (n5489,n5490,n5491);
xor (n5490,n5487,n5488);
or (n5491,n5492,n5495);
and (n5492,n5493,n5494);
xor (n5493,n5316,n5317);
and (n5494,n310,n898);
and (n5495,n5496,n5497);
xor (n5496,n5493,n5494);
or (n5497,n5498,n5501);
and (n5498,n5499,n5500);
xor (n5499,n5322,n5323);
and (n5500,n348,n898);
and (n5501,n5502,n5503);
xor (n5502,n5499,n5500);
or (n5503,n5504,n5507);
and (n5504,n5505,n5506);
xor (n5505,n5328,n5329);
and (n5506,n342,n898);
and (n5507,n5508,n5509);
xor (n5508,n5505,n5506);
or (n5509,n5510,n5513);
and (n5510,n5511,n5512);
xor (n5511,n5333,n5334);
and (n5512,n356,n898);
and (n5513,n5514,n5515);
xor (n5514,n5511,n5512);
or (n5515,n5516,n5519);
and (n5516,n5517,n5518);
xor (n5517,n5339,n5340);
and (n5518,n39,n898);
and (n5519,n5520,n5521);
xor (n5520,n5517,n5518);
or (n5521,n5522,n5525);
and (n5522,n5523,n5524);
xor (n5523,n5344,n5345);
and (n5524,n33,n898);
and (n5525,n5526,n5527);
xor (n5526,n5523,n5524);
or (n5527,n5528,n5531);
and (n5528,n5529,n5530);
xor (n5529,n5349,n5350);
and (n5530,n64,n898);
and (n5531,n5532,n5533);
xor (n5532,n5529,n5530);
or (n5533,n5534,n5537);
and (n5534,n5535,n5536);
xor (n5535,n5355,n5356);
and (n5536,n58,n898);
and (n5537,n5538,n5539);
xor (n5538,n5535,n5536);
or (n5539,n5540,n5543);
and (n5540,n5541,n5542);
xor (n5541,n5361,n5362);
and (n5542,n117,n898);
and (n5543,n5544,n5545);
xor (n5544,n5541,n5542);
or (n5545,n5546,n5549);
and (n5546,n5547,n5548);
xor (n5547,n5367,n5368);
and (n5548,n111,n898);
and (n5549,n5550,n5551);
xor (n5550,n5547,n5548);
or (n5551,n5552,n5555);
and (n5552,n5553,n5554);
xor (n5553,n5373,n5374);
and (n5554,n141,n898);
and (n5555,n5556,n5557);
xor (n5556,n5553,n5554);
or (n5557,n5558,n5561);
and (n5558,n5559,n5560);
xor (n5559,n5379,n5380);
and (n5560,n135,n898);
and (n5561,n5562,n5563);
xor (n5562,n5559,n5560);
or (n5563,n5564,n5567);
and (n5564,n5565,n5566);
xor (n5565,n5385,n5386);
and (n5566,n448,n898);
and (n5567,n5568,n5569);
xor (n5568,n5565,n5566);
or (n5569,n5570,n5573);
and (n5570,n5571,n5572);
xor (n5571,n5391,n5392);
and (n5572,n474,n898);
and (n5573,n5574,n5575);
xor (n5574,n5571,n5572);
or (n5575,n5576,n5579);
and (n5576,n5577,n5578);
xor (n5577,n5397,n5398);
and (n5578,n625,n898);
and (n5579,n5580,n5581);
xor (n5580,n5577,n5578);
or (n5581,n5582,n5585);
and (n5582,n5583,n5584);
xor (n5583,n5403,n5404);
and (n5584,n1037,n898);
and (n5585,n5586,n5587);
xor (n5586,n5583,n5584);
or (n5587,n5588,n5591);
and (n5588,n5589,n5590);
xor (n5589,n5409,n5410);
and (n5590,n1030,n898);
and (n5591,n5592,n5593);
xor (n5592,n5589,n5590);
or (n5593,n5594,n5597);
and (n5594,n5595,n5596);
xor (n5595,n5415,n5416);
and (n5596,n1002,n898);
and (n5597,n5598,n5599);
xor (n5598,n5595,n5596);
or (n5599,n5600,n5603);
and (n5600,n5601,n5602);
xor (n5601,n5420,n5421);
and (n5602,n832,n898);
and (n5603,n5604,n5605);
xor (n5604,n5601,n5602);
or (n5605,n5606,n5609);
and (n5606,n5607,n5608);
xor (n5607,n5426,n5427);
and (n5608,n826,n898);
and (n5609,n5610,n5611);
xor (n5610,n5607,n5608);
or (n5611,n5612,n5615);
and (n5612,n5613,n5614);
xor (n5613,n5431,n5432);
and (n5614,n847,n898);
and (n5615,n5616,n5617);
xor (n5616,n5613,n5614);
or (n5617,n5618,n5621);
and (n5618,n5619,n5620);
xor (n5619,n5437,n5438);
and (n5620,n839,n898);
and (n5621,n5622,n5623);
xor (n5622,n5619,n5620);
and (n5623,n5624,n3657);
xor (n5624,n5443,n5444);
and (n5625,n214,n859);
and (n5626,n5627,n5628);
xor (n5627,n5269,n5625);
or (n5628,n5629,n5632);
and (n5629,n5630,n5631);
xor (n5630,n5448,n5449);
and (n5631,n208,n859);
and (n5632,n5633,n5634);
xor (n5633,n5630,n5631);
or (n5634,n5635,n5637);
and (n5635,n5636,n2537);
xor (n5636,n5454,n5455);
and (n5637,n5638,n5639);
xor (n5638,n5636,n2537);
or (n5639,n5640,n5643);
and (n5640,n5641,n5642);
xor (n5641,n5460,n5461);
and (n5642,n161,n859);
and (n5643,n5644,n5645);
xor (n5644,n5641,n5642);
or (n5645,n5646,n5649);
and (n5646,n5647,n5648);
xor (n5647,n5466,n5467);
and (n5648,n236,n859);
and (n5649,n5650,n5651);
xor (n5650,n5647,n5648);
or (n5651,n5652,n5654);
and (n5652,n5653,n1069);
xor (n5653,n5472,n5473);
and (n5654,n5655,n5656);
xor (n5655,n5653,n1069);
or (n5656,n5657,n5660);
and (n5657,n5658,n5659);
xor (n5658,n5478,n5479);
and (n5659,n90,n859);
and (n5660,n5661,n5662);
xor (n5661,n5658,n5659);
or (n5662,n5663,n5666);
and (n5663,n5664,n5665);
xor (n5664,n5484,n5485);
and (n5665,n84,n859);
and (n5666,n5667,n5668);
xor (n5667,n5664,n5665);
or (n5668,n5669,n5672);
and (n5669,n5670,n5671);
xor (n5670,n5490,n5491);
and (n5671,n310,n859);
and (n5672,n5673,n5674);
xor (n5673,n5670,n5671);
or (n5674,n5675,n5678);
and (n5675,n5676,n5677);
xor (n5676,n5496,n5497);
and (n5677,n348,n859);
and (n5678,n5679,n5680);
xor (n5679,n5676,n5677);
or (n5680,n5681,n5683);
and (n5681,n5682,n1115);
xor (n5682,n5502,n5503);
and (n5683,n5684,n5685);
xor (n5684,n5682,n1115);
or (n5685,n5686,n5689);
and (n5686,n5687,n5688);
xor (n5687,n5508,n5509);
and (n5688,n356,n859);
and (n5689,n5690,n5691);
xor (n5690,n5687,n5688);
or (n5691,n5692,n5695);
and (n5692,n5693,n5694);
xor (n5693,n5514,n5515);
and (n5694,n39,n859);
and (n5695,n5696,n5697);
xor (n5696,n5693,n5694);
or (n5697,n5698,n5701);
and (n5698,n5699,n5700);
xor (n5699,n5520,n5521);
and (n5700,n33,n859);
and (n5701,n5702,n5703);
xor (n5702,n5699,n5700);
or (n5703,n5704,n5707);
and (n5704,n5705,n5706);
xor (n5705,n5526,n5527);
and (n5706,n64,n859);
and (n5707,n5708,n5709);
xor (n5708,n5705,n5706);
or (n5709,n5710,n5713);
and (n5710,n5711,n5712);
xor (n5711,n5532,n5533);
and (n5712,n58,n859);
and (n5713,n5714,n5715);
xor (n5714,n5711,n5712);
or (n5715,n5716,n5719);
and (n5716,n5717,n5718);
xor (n5717,n5538,n5539);
and (n5718,n117,n859);
and (n5719,n5720,n5721);
xor (n5720,n5717,n5718);
or (n5721,n5722,n5725);
and (n5722,n5723,n5724);
xor (n5723,n5544,n5545);
and (n5724,n111,n859);
and (n5725,n5726,n5727);
xor (n5726,n5723,n5724);
or (n5727,n5728,n5731);
and (n5728,n5729,n5730);
xor (n5729,n5550,n5551);
and (n5730,n141,n859);
and (n5731,n5732,n5733);
xor (n5732,n5729,n5730);
or (n5733,n5734,n5737);
and (n5734,n5735,n5736);
xor (n5735,n5556,n5557);
and (n5736,n135,n859);
and (n5737,n5738,n5739);
xor (n5738,n5735,n5736);
or (n5739,n5740,n5742);
and (n5740,n5741,n3004);
xor (n5741,n5562,n5563);
and (n5742,n5743,n5744);
xor (n5743,n5741,n3004);
or (n5744,n5745,n5748);
and (n5745,n5746,n5747);
xor (n5746,n5568,n5569);
and (n5747,n474,n859);
and (n5748,n5749,n5750);
xor (n5749,n5746,n5747);
or (n5750,n5751,n5754);
and (n5751,n5752,n5753);
xor (n5752,n5574,n5575);
and (n5753,n625,n859);
and (n5754,n5755,n5756);
xor (n5755,n5752,n5753);
or (n5756,n5757,n5760);
and (n5757,n5758,n5759);
xor (n5758,n5580,n5581);
and (n5759,n1037,n859);
and (n5760,n5761,n5762);
xor (n5761,n5758,n5759);
or (n5762,n5763,n5765);
and (n5763,n5764,n3402);
xor (n5764,n5586,n5587);
and (n5765,n5766,n5767);
xor (n5766,n5764,n3402);
or (n5767,n5768,n5770);
and (n5768,n5769,n3486);
xor (n5769,n5592,n5593);
and (n5770,n5771,n5772);
xor (n5771,n5769,n3486);
or (n5772,n5773,n5775);
and (n5773,n5774,n3544);
xor (n5774,n5598,n5599);
and (n5775,n5776,n5777);
xor (n5776,n5774,n3544);
or (n5777,n5778,n5780);
and (n5778,n5779,n3541);
xor (n5779,n5604,n5605);
and (n5780,n5781,n5782);
xor (n5781,n5779,n3541);
or (n5782,n5783,n5785);
and (n5783,n5784,n3609);
xor (n5784,n5610,n5611);
and (n5785,n5786,n5787);
xor (n5786,n5784,n3609);
or (n5787,n5788,n5790);
and (n5788,n5789,n3636);
xor (n5789,n5616,n5617);
and (n5790,n5791,n5792);
xor (n5791,n5789,n3636);
and (n5792,n5793,n5794);
xor (n5793,n5622,n5623);
and (n5794,n887,n859);
and (n5796,n192,n858);
or (n5797,n5798,n5800);
and (n5798,n5799,n5796);
xor (n5799,n5245,n5258);
and (n5800,n5801,n5802);
xor (n5801,n5799,n5796);
or (n5802,n5803,n5805);
and (n5803,n5804,n5796);
xor (n5804,n5245,n5260);
and (n5805,n5806,n5807);
xor (n5806,n5804,n5796);
or (n5807,n5808,n5810);
and (n5808,n5809,n5796);
xor (n5809,n5245,n5262);
and (n5810,n5811,n5812);
xor (n5811,n5809,n5796);
or (n5812,n5813,n5815);
and (n5813,n5814,n5796);
xor (n5814,n5245,n5264);
and (n5815,n5816,n5817);
xor (n5816,n5814,n5796);
or (n5817,n5818,n6005);
or (n5818,n5819,n5821);
and (n5819,n5820,n5796);
xor (n5820,n5245,n5265);
and (n5821,n5822,n5823);
xor (n5822,n5820,n5796);
or (n5823,n5824,n5827);
and (n5824,n5825,n5826);
xor (n5825,n5245,n5267);
and (n5826,n214,n858);
and (n5827,n5828,n5829);
xor (n5828,n5825,n5826);
or (n5829,n5830,n5833);
and (n5830,n5831,n5832);
xor (n5831,n5627,n5628);
and (n5832,n208,n858);
and (n5833,n5834,n5835);
xor (n5834,n5831,n5832);
or (n5835,n5836,n5839);
and (n5836,n5837,n5838);
xor (n5837,n5633,n5634);
and (n5838,n167,n858);
and (n5839,n5840,n5841);
xor (n5840,n5837,n5838);
or (n5841,n5842,n5845);
and (n5842,n5843,n5844);
xor (n5843,n5638,n5639);
and (n5844,n161,n858);
and (n5845,n5846,n5847);
xor (n5846,n5843,n5844);
or (n5847,n5848,n5851);
and (n5848,n5849,n5850);
xor (n5849,n5644,n5645);
and (n5850,n236,n858);
and (n5851,n5852,n5853);
xor (n5852,n5849,n5850);
or (n5853,n5854,n5857);
and (n5854,n5855,n5856);
xor (n5855,n5650,n5651);
and (n5856,n230,n858);
and (n5857,n5858,n5859);
xor (n5858,n5855,n5856);
or (n5859,n5860,n5863);
and (n5860,n5861,n5862);
xor (n5861,n5655,n5656);
and (n5862,n90,n858);
and (n5863,n5864,n5865);
xor (n5864,n5861,n5862);
or (n5865,n5866,n5869);
and (n5866,n5867,n5868);
xor (n5867,n5661,n5662);
and (n5868,n84,n858);
and (n5869,n5870,n5871);
xor (n5870,n5867,n5868);
or (n5871,n5872,n5875);
and (n5872,n5873,n5874);
xor (n5873,n5667,n5668);
and (n5874,n310,n858);
and (n5875,n5876,n5877);
xor (n5876,n5873,n5874);
or (n5877,n5878,n5881);
and (n5878,n5879,n5880);
xor (n5879,n5673,n5674);
and (n5880,n348,n858);
and (n5881,n5882,n5883);
xor (n5882,n5879,n5880);
or (n5883,n5884,n5887);
and (n5884,n5885,n5886);
xor (n5885,n5679,n5680);
and (n5886,n342,n858);
and (n5887,n5888,n5889);
xor (n5888,n5885,n5886);
or (n5889,n5890,n5893);
and (n5890,n5891,n5892);
xor (n5891,n5684,n5685);
and (n5892,n356,n858);
and (n5893,n5894,n5895);
xor (n5894,n5891,n5892);
or (n5895,n5896,n5899);
and (n5896,n5897,n5898);
xor (n5897,n5690,n5691);
and (n5898,n39,n858);
and (n5899,n5900,n5901);
xor (n5900,n5897,n5898);
or (n5901,n5902,n5905);
and (n5902,n5903,n5904);
xor (n5903,n5696,n5697);
and (n5904,n33,n858);
and (n5905,n5906,n5907);
xor (n5906,n5903,n5904);
or (n5907,n5908,n5911);
and (n5908,n5909,n5910);
xor (n5909,n5702,n5703);
and (n5910,n64,n858);
and (n5911,n5912,n5913);
xor (n5912,n5909,n5910);
or (n5913,n5914,n5917);
and (n5914,n5915,n5916);
xor (n5915,n5708,n5709);
and (n5916,n58,n858);
and (n5917,n5918,n5919);
xor (n5918,n5915,n5916);
or (n5919,n5920,n5923);
and (n5920,n5921,n5922);
xor (n5921,n5714,n5715);
and (n5922,n117,n858);
and (n5923,n5924,n5925);
xor (n5924,n5921,n5922);
or (n5925,n5926,n5929);
and (n5926,n5927,n5928);
xor (n5927,n5720,n5721);
and (n5928,n111,n858);
and (n5929,n5930,n5931);
xor (n5930,n5927,n5928);
or (n5931,n5932,n5935);
and (n5932,n5933,n5934);
xor (n5933,n5726,n5727);
and (n5934,n141,n858);
and (n5935,n5936,n5937);
xor (n5936,n5933,n5934);
or (n5937,n5938,n5941);
and (n5938,n5939,n5940);
xor (n5939,n5732,n5733);
and (n5940,n135,n858);
and (n5941,n5942,n5943);
xor (n5942,n5939,n5940);
or (n5943,n5944,n5947);
and (n5944,n5945,n5946);
xor (n5945,n5738,n5739);
and (n5946,n448,n858);
and (n5947,n5948,n5949);
xor (n5948,n5945,n5946);
or (n5949,n5950,n5953);
and (n5950,n5951,n5952);
xor (n5951,n5743,n5744);
and (n5952,n474,n858);
and (n5953,n5954,n5955);
xor (n5954,n5951,n5952);
or (n5955,n5956,n5959);
and (n5956,n5957,n5958);
xor (n5957,n5749,n5750);
and (n5958,n625,n858);
and (n5959,n5960,n5961);
xor (n5960,n5957,n5958);
or (n5961,n5962,n5965);
and (n5962,n5963,n5964);
xor (n5963,n5755,n5756);
and (n5964,n1037,n858);
and (n5965,n5966,n5967);
xor (n5966,n5963,n5964);
or (n5967,n5968,n5971);
and (n5968,n5969,n5970);
xor (n5969,n5761,n5762);
and (n5970,n1030,n858);
and (n5971,n5972,n5973);
xor (n5972,n5969,n5970);
or (n5973,n5974,n5977);
and (n5974,n5975,n5976);
xor (n5975,n5766,n5767);
and (n5976,n1002,n858);
and (n5977,n5978,n5979);
xor (n5978,n5975,n5976);
or (n5979,n5980,n5983);
and (n5980,n5981,n5982);
xor (n5981,n5771,n5772);
and (n5982,n832,n858);
and (n5983,n5984,n5985);
xor (n5984,n5981,n5982);
or (n5985,n5986,n5989);
and (n5986,n5987,n5988);
xor (n5987,n5776,n5777);
and (n5988,n826,n858);
and (n5989,n5990,n5991);
xor (n5990,n5987,n5988);
or (n5991,n5992,n5995);
and (n5992,n5993,n5994);
xor (n5993,n5781,n5782);
and (n5994,n847,n858);
and (n5995,n5996,n5997);
xor (n5996,n5993,n5994);
or (n5997,n5998,n6001);
and (n5998,n5999,n6000);
xor (n5999,n5786,n5787);
and (n6000,n839,n858);
and (n6001,n6002,n6003);
xor (n6002,n5999,n6000);
and (n6003,n6004,n3582);
xor (n6004,n5791,n5792);
and (n6005,n5822,n5819);
and (n6006,n192,n864);
or (n6007,n6008,n6010);
and (n6008,n6009,n6006);
xor (n6009,n5801,n5802);
and (n6010,n6011,n6012);
xor (n6011,n6009,n6006);
or (n6012,n6013,n6015);
and (n6013,n6014,n6006);
xor (n6014,n5806,n5807);
and (n6015,n6016,n6017);
xor (n6016,n6014,n6006);
or (n6017,n6018,n6020);
and (n6018,n6019,n6006);
xor (n6019,n5811,n5812);
and (n6020,n6021,n6022);
xor (n6021,n6019,n6006);
or (n6022,n6023,n6025);
and (n6023,n6024,n6006);
xor (n6024,n5816,n5817);
and (n6025,n6026,n6027);
xor (n6026,n6024,n6006);
or (n6027,n6028,n6212);
or (n6028,n6029,n6031);
and (n6029,n6030,n6006);
xor (n6030,n5822,n5818);
and (n6031,n6032,n6033);
xor (n6032,n6030,n6006);
or (n6033,n6034,n6037);
and (n6034,n6035,n6036);
xor (n6035,n5822,n5823);
and (n6036,n214,n864);
and (n6037,n6038,n6039);
xor (n6038,n6035,n6036);
or (n6039,n6040,n6043);
and (n6040,n6041,n6042);
xor (n6041,n5828,n5829);
and (n6042,n208,n864);
and (n6043,n6044,n6045);
xor (n6044,n6041,n6042);
or (n6045,n6046,n6049);
and (n6046,n6047,n6048);
xor (n6047,n5834,n5835);
and (n6048,n167,n864);
and (n6049,n6050,n6051);
xor (n6050,n6047,n6048);
or (n6051,n6052,n6055);
and (n6052,n6053,n6054);
xor (n6053,n5840,n5841);
and (n6054,n161,n864);
and (n6055,n6056,n6057);
xor (n6056,n6053,n6054);
or (n6057,n6058,n6061);
and (n6058,n6059,n6060);
xor (n6059,n5846,n5847);
and (n6060,n236,n864);
and (n6061,n6062,n6063);
xor (n6062,n6059,n6060);
or (n6063,n6064,n6067);
and (n6064,n6065,n6066);
xor (n6065,n5852,n5853);
and (n6066,n230,n864);
and (n6067,n6068,n6069);
xor (n6068,n6065,n6066);
or (n6069,n6070,n6073);
and (n6070,n6071,n6072);
xor (n6071,n5858,n5859);
and (n6072,n90,n864);
and (n6073,n6074,n6075);
xor (n6074,n6071,n6072);
or (n6075,n6076,n6079);
and (n6076,n6077,n6078);
xor (n6077,n5864,n5865);
and (n6078,n84,n864);
and (n6079,n6080,n6081);
xor (n6080,n6077,n6078);
or (n6081,n6082,n6085);
and (n6082,n6083,n6084);
xor (n6083,n5870,n5871);
and (n6084,n310,n864);
and (n6085,n6086,n6087);
xor (n6086,n6083,n6084);
or (n6087,n6088,n6091);
and (n6088,n6089,n6090);
xor (n6089,n5876,n5877);
and (n6090,n348,n864);
and (n6091,n6092,n6093);
xor (n6092,n6089,n6090);
or (n6093,n6094,n6097);
and (n6094,n6095,n6096);
xor (n6095,n5882,n5883);
and (n6096,n342,n864);
and (n6097,n6098,n6099);
xor (n6098,n6095,n6096);
or (n6099,n6100,n6102);
and (n6100,n6101,n1165);
xor (n6101,n5888,n5889);
and (n6102,n6103,n6104);
xor (n6103,n6101,n1165);
or (n6104,n6105,n6107);
and (n6105,n6106,n1366);
xor (n6106,n5894,n5895);
and (n6107,n6108,n6109);
xor (n6108,n6106,n1366);
or (n6109,n6110,n6113);
and (n6110,n6111,n6112);
xor (n6111,n5900,n5901);
and (n6112,n33,n864);
and (n6113,n6114,n6115);
xor (n6114,n6111,n6112);
or (n6115,n6116,n6119);
and (n6116,n6117,n6118);
xor (n6117,n5906,n5907);
and (n6118,n64,n864);
and (n6119,n6120,n6121);
xor (n6120,n6117,n6118);
or (n6121,n6122,n6125);
and (n6122,n6123,n6124);
xor (n6123,n5912,n5913);
and (n6124,n58,n864);
and (n6125,n6126,n6127);
xor (n6126,n6123,n6124);
or (n6127,n6128,n6130);
and (n6128,n6129,n1926);
xor (n6129,n5918,n5919);
and (n6130,n6131,n6132);
xor (n6131,n6129,n1926);
or (n6132,n6133,n6136);
and (n6133,n6134,n6135);
xor (n6134,n5924,n5925);
and (n6135,n111,n864);
and (n6136,n6137,n6138);
xor (n6137,n6134,n6135);
or (n6138,n6139,n6142);
and (n6139,n6140,n6141);
xor (n6140,n5930,n5931);
and (n6141,n141,n864);
and (n6142,n6143,n6144);
xor (n6143,n6140,n6141);
or (n6144,n6145,n6148);
and (n6145,n6146,n6147);
xor (n6146,n5936,n5937);
and (n6147,n135,n864);
and (n6148,n6149,n6150);
xor (n6149,n6146,n6147);
or (n6150,n6151,n6154);
and (n6151,n6152,n6153);
xor (n6152,n5942,n5943);
and (n6153,n448,n864);
and (n6154,n6155,n6156);
xor (n6155,n6152,n6153);
or (n6156,n6157,n6160);
and (n6157,n6158,n6159);
xor (n6158,n5948,n5949);
and (n6159,n474,n864);
and (n6160,n6161,n6162);
xor (n6161,n6158,n6159);
or (n6162,n6163,n6166);
and (n6163,n6164,n6165);
xor (n6164,n5954,n5955);
and (n6165,n625,n864);
and (n6166,n6167,n6168);
xor (n6167,n6164,n6165);
or (n6168,n6169,n6172);
and (n6169,n6170,n6171);
xor (n6170,n5960,n5961);
and (n6171,n1037,n864);
and (n6172,n6173,n6174);
xor (n6173,n6170,n6171);
or (n6174,n6175,n6178);
and (n6175,n6176,n6177);
xor (n6176,n5966,n5967);
and (n6177,n1030,n864);
and (n6178,n6179,n6180);
xor (n6179,n6176,n6177);
or (n6180,n6181,n6184);
and (n6181,n6182,n6183);
xor (n6182,n5972,n5973);
and (n6183,n1002,n864);
and (n6184,n6185,n6186);
xor (n6185,n6182,n6183);
or (n6186,n6187,n6190);
and (n6187,n6188,n6189);
xor (n6188,n5978,n5979);
and (n6189,n832,n864);
and (n6190,n6191,n6192);
xor (n6191,n6188,n6189);
or (n6192,n6193,n6196);
and (n6193,n6194,n6195);
xor (n6194,n5984,n5985);
and (n6195,n826,n864);
and (n6196,n6197,n6198);
xor (n6197,n6194,n6195);
or (n6198,n6199,n6202);
and (n6199,n6200,n6201);
xor (n6200,n5990,n5991);
and (n6201,n847,n864);
and (n6202,n6203,n6204);
xor (n6203,n6200,n6201);
or (n6204,n6205,n6207);
and (n6205,n6206,n3575);
xor (n6206,n5996,n5997);
and (n6207,n6208,n6209);
xor (n6208,n6206,n3575);
and (n6209,n6210,n6211);
xor (n6210,n6002,n6003);
and (n6211,n887,n864);
and (n6212,n6032,n6029);
and (n6213,n192,n952);
or (n6214,n6215,n6217);
and (n6215,n6216,n6213);
xor (n6216,n6011,n6012);
and (n6217,n6218,n6219);
xor (n6218,n6216,n6213);
or (n6219,n6220,n6222);
and (n6220,n6221,n6213);
xor (n6221,n6016,n6017);
and (n6222,n6223,n6224);
xor (n6223,n6221,n6213);
or (n6224,n6225,n6227);
and (n6225,n6226,n6213);
xor (n6226,n6021,n6022);
and (n6227,n6228,n6229);
xor (n6228,n6226,n6213);
or (n6229,n6230,n6232);
and (n6230,n6231,n6213);
xor (n6231,n6026,n6027);
and (n6232,n6233,n6234);
xor (n6233,n6231,n6213);
or (n6234,n6235,n6237);
and (n6235,n6236,n6213);
xor (n6236,n6032,n6028);
and (n6237,n6238,n6235);
xor (n6238,n6236,n6213);
or (n6239,n6240,n6242);
and (n6240,n6241,n3882);
xor (n6241,n6218,n6219);
and (n6242,n6243,n6244);
xor (n6243,n6241,n3882);
or (n6244,n6245,n6247);
and (n6245,n6246,n3882);
xor (n6246,n6223,n6224);
and (n6247,n6248,n6249);
xor (n6248,n6246,n3882);
or (n6249,n6250,n6252);
and (n6250,n6251,n3882);
xor (n6251,n6228,n6229);
and (n6252,n6253,n6254);
xor (n6253,n6251,n3882);
or (n6254,n6255,n6257);
and (n6255,n6256,n3882);
xor (n6256,n6233,n6234);
and (n6257,n6258,n6259);
xor (n6258,n6256,n3882);
or (n6259,n6260,n6262);
and (n6260,n6261,n3882);
xor (n6261,n6238,n6235);
and (n6262,n6263,n6260);
xor (n6263,n6261,n3882);
and (n6264,n192,n493);
or (n6265,n6266,n6268);
and (n6266,n6267,n6264);
xor (n6267,n6243,n6244);
and (n6268,n6269,n6270);
xor (n6269,n6267,n6264);
or (n6270,n6271,n6273);
and (n6271,n6272,n6264);
xor (n6272,n6248,n6249);
and (n6273,n6274,n6275);
xor (n6274,n6272,n6264);
or (n6275,n6276,n6278);
and (n6276,n6277,n6264);
xor (n6277,n6253,n6254);
and (n6278,n6279,n6280);
xor (n6279,n6277,n6264);
or (n6280,n6281,n6283);
and (n6281,n6282,n6264);
xor (n6282,n6258,n6259);
and (n6283,n6284,n6285);
xor (n6284,n6282,n6264);
or (n6285,n6286,n6288);
and (n6286,n6287,n6264);
xor (n6287,n6263,n6260);
and (n6288,n6289,n6290);
xor (n6289,n6287,n6264);
or (n6290,n6291,n6653);
and (n6291,n6292,n6652);
xor (n6292,n6263,n6293);
or (n6293,n6294,n6478);
and (n6294,n6295,n4233);
xor (n6295,n6238,n6296);
or (n6296,n6297,n6300);
and (n6297,n6298,n6299);
xor (n6298,n6032,n6033);
and (n6299,n214,n952);
and (n6300,n6301,n6302);
xor (n6301,n6298,n6299);
or (n6302,n6303,n6306);
and (n6303,n6304,n6305);
xor (n6304,n6038,n6039);
and (n6305,n208,n952);
and (n6306,n6307,n6308);
xor (n6307,n6304,n6305);
or (n6308,n6309,n6312);
and (n6309,n6310,n6311);
xor (n6310,n6044,n6045);
and (n6311,n167,n952);
and (n6312,n6313,n6314);
xor (n6313,n6310,n6311);
or (n6314,n6315,n6318);
and (n6315,n6316,n6317);
xor (n6316,n6050,n6051);
and (n6317,n161,n952);
and (n6318,n6319,n6320);
xor (n6319,n6316,n6317);
or (n6320,n6321,n6324);
and (n6321,n6322,n6323);
xor (n6322,n6056,n6057);
and (n6323,n236,n952);
and (n6324,n6325,n6326);
xor (n6325,n6322,n6323);
or (n6326,n6327,n6330);
and (n6327,n6328,n6329);
xor (n6328,n6062,n6063);
and (n6329,n230,n952);
and (n6330,n6331,n6332);
xor (n6331,n6328,n6329);
or (n6332,n6333,n6336);
and (n6333,n6334,n6335);
xor (n6334,n6068,n6069);
and (n6335,n90,n952);
and (n6336,n6337,n6338);
xor (n6337,n6334,n6335);
or (n6338,n6339,n6342);
and (n6339,n6340,n6341);
xor (n6340,n6074,n6075);
and (n6341,n84,n952);
and (n6342,n6343,n6344);
xor (n6343,n6340,n6341);
or (n6344,n6345,n6348);
and (n6345,n6346,n6347);
xor (n6346,n6080,n6081);
and (n6347,n310,n952);
and (n6348,n6349,n6350);
xor (n6349,n6346,n6347);
or (n6350,n6351,n6354);
and (n6351,n6352,n6353);
xor (n6352,n6086,n6087);
and (n6353,n348,n952);
and (n6354,n6355,n6356);
xor (n6355,n6352,n6353);
or (n6356,n6357,n6360);
and (n6357,n6358,n6359);
xor (n6358,n6092,n6093);
and (n6359,n342,n952);
and (n6360,n6361,n6362);
xor (n6361,n6358,n6359);
or (n6362,n6363,n6366);
and (n6363,n6364,n6365);
xor (n6364,n6098,n6099);
and (n6365,n356,n952);
and (n6366,n6367,n6368);
xor (n6367,n6364,n6365);
or (n6368,n6369,n6372);
and (n6369,n6370,n6371);
xor (n6370,n6103,n6104);
and (n6371,n39,n952);
and (n6372,n6373,n6374);
xor (n6373,n6370,n6371);
or (n6374,n6375,n6378);
and (n6375,n6376,n6377);
xor (n6376,n6108,n6109);
and (n6377,n33,n952);
and (n6378,n6379,n6380);
xor (n6379,n6376,n6377);
or (n6380,n6381,n6384);
and (n6381,n6382,n6383);
xor (n6382,n6114,n6115);
and (n6383,n64,n952);
and (n6384,n6385,n6386);
xor (n6385,n6382,n6383);
or (n6386,n6387,n6390);
and (n6387,n6388,n6389);
xor (n6388,n6120,n6121);
and (n6389,n58,n952);
and (n6390,n6391,n6392);
xor (n6391,n6388,n6389);
or (n6392,n6393,n6396);
and (n6393,n6394,n6395);
xor (n6394,n6126,n6127);
and (n6395,n117,n952);
and (n6396,n6397,n6398);
xor (n6397,n6394,n6395);
or (n6398,n6399,n6402);
and (n6399,n6400,n6401);
xor (n6400,n6131,n6132);
and (n6401,n111,n952);
and (n6402,n6403,n6404);
xor (n6403,n6400,n6401);
or (n6404,n6405,n6408);
and (n6405,n6406,n6407);
xor (n6406,n6137,n6138);
and (n6407,n141,n952);
and (n6408,n6409,n6410);
xor (n6409,n6406,n6407);
or (n6410,n6411,n6414);
and (n6411,n6412,n6413);
xor (n6412,n6143,n6144);
and (n6413,n135,n952);
and (n6414,n6415,n6416);
xor (n6415,n6412,n6413);
or (n6416,n6417,n6420);
and (n6417,n6418,n6419);
xor (n6418,n6149,n6150);
and (n6419,n448,n952);
and (n6420,n6421,n6422);
xor (n6421,n6418,n6419);
or (n6422,n6423,n6426);
and (n6423,n6424,n6425);
xor (n6424,n6155,n6156);
and (n6425,n474,n952);
and (n6426,n6427,n6428);
xor (n6427,n6424,n6425);
or (n6428,n6429,n6432);
and (n6429,n6430,n6431);
xor (n6430,n6161,n6162);
and (n6431,n625,n952);
and (n6432,n6433,n6434);
xor (n6433,n6430,n6431);
or (n6434,n6435,n6438);
and (n6435,n6436,n6437);
xor (n6436,n6167,n6168);
and (n6437,n1037,n952);
and (n6438,n6439,n6440);
xor (n6439,n6436,n6437);
or (n6440,n6441,n6444);
and (n6441,n6442,n6443);
xor (n6442,n6173,n6174);
and (n6443,n1030,n952);
and (n6444,n6445,n6446);
xor (n6445,n6442,n6443);
or (n6446,n6447,n6450);
and (n6447,n6448,n6449);
xor (n6448,n6179,n6180);
and (n6449,n1002,n952);
and (n6450,n6451,n6452);
xor (n6451,n6448,n6449);
or (n6452,n6453,n6456);
and (n6453,n6454,n6455);
xor (n6454,n6185,n6186);
and (n6455,n832,n952);
and (n6456,n6457,n6458);
xor (n6457,n6454,n6455);
or (n6458,n6459,n6462);
and (n6459,n6460,n6461);
xor (n6460,n6191,n6192);
and (n6461,n826,n952);
and (n6462,n6463,n6464);
xor (n6463,n6460,n6461);
or (n6464,n6465,n6468);
and (n6465,n6466,n6467);
xor (n6466,n6197,n6198);
and (n6467,n847,n952);
and (n6468,n6469,n6470);
xor (n6469,n6466,n6467);
or (n6470,n6471,n6474);
and (n6471,n6472,n6473);
xor (n6472,n6203,n6204);
and (n6473,n839,n952);
and (n6474,n6475,n6476);
xor (n6475,n6472,n6473);
and (n6476,n6477,n3502);
xor (n6477,n6208,n6209);
and (n6478,n6479,n6480);
xor (n6479,n6295,n4233);
or (n6480,n6481,n6484);
and (n6481,n6482,n6483);
xor (n6482,n6301,n6302);
and (n6483,n208,n495);
and (n6484,n6485,n6486);
xor (n6485,n6482,n6483);
or (n6486,n6487,n6490);
and (n6487,n6488,n6489);
xor (n6488,n6307,n6308);
and (n6489,n167,n495);
and (n6490,n6491,n6492);
xor (n6491,n6488,n6489);
or (n6492,n6493,n6496);
and (n6493,n6494,n6495);
xor (n6494,n6313,n6314);
and (n6495,n161,n495);
and (n6496,n6497,n6498);
xor (n6497,n6494,n6495);
or (n6498,n6499,n6502);
and (n6499,n6500,n6501);
xor (n6500,n6319,n6320);
and (n6501,n236,n495);
and (n6502,n6503,n6504);
xor (n6503,n6500,n6501);
or (n6504,n6505,n6508);
and (n6505,n6506,n6507);
xor (n6506,n6325,n6326);
and (n6507,n230,n495);
and (n6508,n6509,n6510);
xor (n6509,n6506,n6507);
or (n6510,n6511,n6514);
and (n6511,n6512,n6513);
xor (n6512,n6331,n6332);
and (n6513,n90,n495);
and (n6514,n6515,n6516);
xor (n6515,n6512,n6513);
or (n6516,n6517,n6520);
and (n6517,n6518,n6519);
xor (n6518,n6337,n6338);
and (n6519,n84,n495);
and (n6520,n6521,n6522);
xor (n6521,n6518,n6519);
or (n6522,n6523,n6526);
and (n6523,n6524,n6525);
xor (n6524,n6343,n6344);
and (n6525,n310,n495);
and (n6526,n6527,n6528);
xor (n6527,n6524,n6525);
or (n6528,n6529,n6532);
and (n6529,n6530,n6531);
xor (n6530,n6349,n6350);
and (n6531,n348,n495);
and (n6532,n6533,n6534);
xor (n6533,n6530,n6531);
or (n6534,n6535,n6537);
and (n6535,n6536,n947);
xor (n6536,n6355,n6356);
and (n6537,n6538,n6539);
xor (n6538,n6536,n947);
or (n6539,n6540,n6543);
and (n6540,n6541,n6542);
xor (n6541,n6361,n6362);
and (n6542,n356,n495);
and (n6543,n6544,n6545);
xor (n6544,n6541,n6542);
or (n6545,n6546,n6549);
and (n6546,n6547,n6548);
xor (n6547,n6367,n6368);
and (n6548,n39,n495);
and (n6549,n6550,n6551);
xor (n6550,n6547,n6548);
or (n6551,n6552,n6555);
and (n6552,n6553,n6554);
xor (n6553,n6373,n6374);
and (n6554,n33,n495);
and (n6555,n6556,n6557);
xor (n6556,n6553,n6554);
or (n6557,n6558,n6561);
and (n6558,n6559,n6560);
xor (n6559,n6379,n6380);
and (n6560,n64,n495);
and (n6561,n6562,n6563);
xor (n6562,n6559,n6560);
or (n6563,n6564,n6567);
and (n6564,n6565,n6566);
xor (n6565,n6385,n6386);
and (n6566,n58,n495);
and (n6567,n6568,n6569);
xor (n6568,n6565,n6566);
or (n6569,n6570,n6573);
and (n6570,n6571,n6572);
xor (n6571,n6391,n6392);
and (n6572,n117,n495);
and (n6573,n6574,n6575);
xor (n6574,n6571,n6572);
or (n6575,n6576,n6578);
and (n6576,n6577,n1814);
xor (n6577,n6397,n6398);
and (n6578,n6579,n6580);
xor (n6579,n6577,n1814);
or (n6580,n6581,n6583);
and (n6581,n6582,n1902);
xor (n6582,n6403,n6404);
and (n6583,n6584,n6585);
xor (n6584,n6582,n1902);
or (n6585,n6586,n6589);
and (n6586,n6587,n6588);
xor (n6587,n6409,n6410);
and (n6588,n135,n495);
and (n6589,n6590,n6591);
xor (n6590,n6587,n6588);
or (n6591,n6592,n6595);
and (n6592,n6593,n6594);
xor (n6593,n6415,n6416);
and (n6594,n448,n495);
and (n6595,n6596,n6597);
xor (n6596,n6593,n6594);
or (n6597,n6598,n6601);
and (n6598,n6599,n6600);
xor (n6599,n6421,n6422);
and (n6600,n474,n495);
and (n6601,n6602,n6603);
xor (n6602,n6599,n6600);
or (n6603,n6604,n6607);
and (n6604,n6605,n6606);
xor (n6605,n6427,n6428);
and (n6606,n625,n495);
and (n6607,n6608,n6609);
xor (n6608,n6605,n6606);
or (n6609,n6610,n6613);
and (n6610,n6611,n6612);
xor (n6611,n6433,n6434);
and (n6612,n1037,n495);
and (n6613,n6614,n6615);
xor (n6614,n6611,n6612);
or (n6615,n6616,n6619);
and (n6616,n6617,n6618);
xor (n6617,n6439,n6440);
and (n6618,n1030,n495);
and (n6619,n6620,n6621);
xor (n6620,n6617,n6618);
or (n6621,n6622,n6624);
and (n6622,n6623,n3154);
xor (n6623,n6445,n6446);
and (n6624,n6625,n6626);
xor (n6625,n6623,n3154);
or (n6626,n6627,n6630);
and (n6627,n6628,n6629);
xor (n6628,n6451,n6452);
and (n6629,n832,n495);
and (n6630,n6631,n6632);
xor (n6631,n6628,n6629);
or (n6632,n6633,n6636);
and (n6633,n6634,n6635);
xor (n6634,n6457,n6458);
and (n6635,n826,n495);
and (n6636,n6637,n6638);
xor (n6637,n6634,n6635);
or (n6638,n6639,n6642);
and (n6639,n6640,n6641);
xor (n6640,n6463,n6464);
and (n6641,n847,n495);
and (n6642,n6643,n6644);
xor (n6643,n6640,n6641);
or (n6644,n6645,n6647);
and (n6645,n6646,n3460);
xor (n6646,n6469,n6470);
and (n6647,n6648,n6649);
xor (n6648,n6646,n3460);
and (n6649,n6650,n6651);
xor (n6650,n6475,n6476);
and (n6651,n887,n495);
and (n6652,n214,n493);
and (n6653,n6654,n6655);
xor (n6654,n6292,n6652);
or (n6655,n6656,n6659);
and (n6656,n6657,n6658);
xor (n6657,n6479,n6480);
and (n6658,n208,n493);
and (n6659,n6660,n6661);
xor (n6660,n6657,n6658);
or (n6661,n6662,n6665);
and (n6662,n6663,n6664);
xor (n6663,n6485,n6486);
and (n6664,n167,n493);
and (n6665,n6666,n6667);
xor (n6666,n6663,n6664);
or (n6667,n6668,n6671);
and (n6668,n6669,n6670);
xor (n6669,n6491,n6492);
and (n6670,n161,n493);
and (n6671,n6672,n6673);
xor (n6672,n6669,n6670);
or (n6673,n6674,n6677);
and (n6674,n6675,n6676);
xor (n6675,n6497,n6498);
and (n6676,n236,n493);
and (n6677,n6678,n6679);
xor (n6678,n6675,n6676);
or (n6679,n6680,n6683);
and (n6680,n6681,n6682);
xor (n6681,n6503,n6504);
and (n6682,n230,n493);
and (n6683,n6684,n6685);
xor (n6684,n6681,n6682);
or (n6685,n6686,n6689);
and (n6686,n6687,n6688);
xor (n6687,n6509,n6510);
and (n6688,n90,n493);
and (n6689,n6690,n6691);
xor (n6690,n6687,n6688);
or (n6691,n6692,n6695);
and (n6692,n6693,n6694);
xor (n6693,n6515,n6516);
and (n6694,n84,n493);
and (n6695,n6696,n6697);
xor (n6696,n6693,n6694);
or (n6697,n6698,n6701);
and (n6698,n6699,n6700);
xor (n6699,n6521,n6522);
and (n6700,n310,n493);
and (n6701,n6702,n6703);
xor (n6702,n6699,n6700);
or (n6703,n6704,n6707);
and (n6704,n6705,n6706);
xor (n6705,n6527,n6528);
and (n6706,n348,n493);
and (n6707,n6708,n6709);
xor (n6708,n6705,n6706);
or (n6709,n6710,n6713);
and (n6710,n6711,n6712);
xor (n6711,n6533,n6534);
and (n6712,n342,n493);
and (n6713,n6714,n6715);
xor (n6714,n6711,n6712);
or (n6715,n6716,n6719);
and (n6716,n6717,n6718);
xor (n6717,n6538,n6539);
and (n6718,n356,n493);
and (n6719,n6720,n6721);
xor (n6720,n6717,n6718);
or (n6721,n6722,n6725);
and (n6722,n6723,n6724);
xor (n6723,n6544,n6545);
and (n6724,n39,n493);
and (n6725,n6726,n6727);
xor (n6726,n6723,n6724);
or (n6727,n6728,n6731);
and (n6728,n6729,n6730);
xor (n6729,n6550,n6551);
and (n6730,n33,n493);
and (n6731,n6732,n6733);
xor (n6732,n6729,n6730);
or (n6733,n6734,n6737);
and (n6734,n6735,n6736);
xor (n6735,n6556,n6557);
and (n6736,n64,n493);
and (n6737,n6738,n6739);
xor (n6738,n6735,n6736);
or (n6739,n6740,n6743);
and (n6740,n6741,n6742);
xor (n6741,n6562,n6563);
and (n6742,n58,n493);
and (n6743,n6744,n6745);
xor (n6744,n6741,n6742);
or (n6745,n6746,n6749);
and (n6746,n6747,n6748);
xor (n6747,n6568,n6569);
and (n6748,n117,n493);
and (n6749,n6750,n6751);
xor (n6750,n6747,n6748);
or (n6751,n6752,n6755);
and (n6752,n6753,n6754);
xor (n6753,n6574,n6575);
and (n6754,n111,n493);
and (n6755,n6756,n6757);
xor (n6756,n6753,n6754);
or (n6757,n6758,n6761);
and (n6758,n6759,n6760);
xor (n6759,n6579,n6580);
and (n6760,n141,n493);
and (n6761,n6762,n6763);
xor (n6762,n6759,n6760);
or (n6763,n6764,n6767);
and (n6764,n6765,n6766);
xor (n6765,n6584,n6585);
and (n6766,n135,n493);
and (n6767,n6768,n6769);
xor (n6768,n6765,n6766);
or (n6769,n6770,n6773);
and (n6770,n6771,n6772);
xor (n6771,n6590,n6591);
and (n6772,n448,n493);
and (n6773,n6774,n6775);
xor (n6774,n6771,n6772);
or (n6775,n6776,n6779);
and (n6776,n6777,n6778);
xor (n6777,n6596,n6597);
and (n6778,n474,n493);
and (n6779,n6780,n6781);
xor (n6780,n6777,n6778);
or (n6781,n6782,n6785);
and (n6782,n6783,n6784);
xor (n6783,n6602,n6603);
and (n6784,n625,n493);
and (n6785,n6786,n6787);
xor (n6786,n6783,n6784);
or (n6787,n6788,n6791);
and (n6788,n6789,n6790);
xor (n6789,n6608,n6609);
and (n6790,n1037,n493);
and (n6791,n6792,n6793);
xor (n6792,n6789,n6790);
or (n6793,n6794,n6797);
and (n6794,n6795,n6796);
xor (n6795,n6614,n6615);
and (n6796,n1030,n493);
and (n6797,n6798,n6799);
xor (n6798,n6795,n6796);
or (n6799,n6800,n6803);
and (n6800,n6801,n6802);
xor (n6801,n6620,n6621);
and (n6802,n1002,n493);
and (n6803,n6804,n6805);
xor (n6804,n6801,n6802);
or (n6805,n6806,n6809);
and (n6806,n6807,n6808);
xor (n6807,n6625,n6626);
and (n6808,n832,n493);
and (n6809,n6810,n6811);
xor (n6810,n6807,n6808);
or (n6811,n6812,n6815);
and (n6812,n6813,n6814);
xor (n6813,n6631,n6632);
and (n6814,n826,n493);
and (n6815,n6816,n6817);
xor (n6816,n6813,n6814);
or (n6817,n6818,n6821);
and (n6818,n6819,n6820);
xor (n6819,n6637,n6638);
and (n6820,n847,n493);
and (n6821,n6822,n6823);
xor (n6822,n6819,n6820);
or (n6823,n6824,n6827);
and (n6824,n6825,n6826);
xor (n6825,n6643,n6644);
and (n6826,n839,n493);
and (n6827,n6828,n6829);
xor (n6828,n6825,n6826);
and (n6829,n6830,n3397);
xor (n6830,n6648,n6649);
and (n6831,n192,n185);
or (n6832,n6833,n6835);
and (n6833,n6834,n6831);
xor (n6834,n6269,n6270);
and (n6835,n6836,n6837);
xor (n6836,n6834,n6831);
or (n6837,n6838,n6840);
and (n6838,n6839,n6831);
xor (n6839,n6274,n6275);
and (n6840,n6841,n6842);
xor (n6841,n6839,n6831);
or (n6842,n6843,n6845);
and (n6843,n6844,n6831);
xor (n6844,n6279,n6280);
and (n6845,n6846,n6847);
xor (n6846,n6844,n6831);
or (n6847,n6848,n6850);
and (n6848,n6849,n6831);
xor (n6849,n6284,n6285);
and (n6850,n6851,n6852);
xor (n6851,n6849,n6831);
or (n6852,n6853,n6856);
and (n6853,n6854,n6855);
xor (n6854,n6289,n6290);
and (n6855,n214,n185);
and (n6856,n6857,n6858);
xor (n6857,n6854,n6855);
or (n6858,n6859,n6862);
and (n6859,n6860,n6861);
xor (n6860,n6654,n6655);
and (n6861,n208,n185);
and (n6862,n6863,n6864);
xor (n6863,n6860,n6861);
or (n6864,n6865,n6868);
and (n6865,n6866,n6867);
xor (n6866,n6660,n6661);
and (n6867,n167,n185);
and (n6868,n6869,n6870);
xor (n6869,n6866,n6867);
or (n6870,n6871,n6874);
and (n6871,n6872,n6873);
xor (n6872,n6666,n6667);
and (n6873,n161,n185);
and (n6874,n6875,n6876);
xor (n6875,n6872,n6873);
or (n6876,n6877,n6880);
and (n6877,n6878,n6879);
xor (n6878,n6672,n6673);
and (n6879,n236,n185);
and (n6880,n6881,n6882);
xor (n6881,n6878,n6879);
or (n6882,n6883,n6886);
and (n6883,n6884,n6885);
xor (n6884,n6678,n6679);
and (n6885,n230,n185);
and (n6886,n6887,n6888);
xor (n6887,n6884,n6885);
or (n6888,n6889,n6892);
and (n6889,n6890,n6891);
xor (n6890,n6684,n6685);
and (n6891,n90,n185);
and (n6892,n6893,n6894);
xor (n6893,n6890,n6891);
or (n6894,n6895,n6898);
and (n6895,n6896,n6897);
xor (n6896,n6690,n6691);
and (n6897,n84,n185);
and (n6898,n6899,n6900);
xor (n6899,n6896,n6897);
or (n6900,n6901,n6904);
and (n6901,n6902,n6903);
xor (n6902,n6696,n6697);
and (n6903,n310,n185);
and (n6904,n6905,n6906);
xor (n6905,n6902,n6903);
or (n6906,n6907,n6910);
and (n6907,n6908,n6909);
xor (n6908,n6702,n6703);
and (n6909,n348,n185);
and (n6910,n6911,n6912);
xor (n6911,n6908,n6909);
or (n6912,n6913,n6916);
and (n6913,n6914,n6915);
xor (n6914,n6708,n6709);
and (n6915,n342,n185);
and (n6916,n6917,n6918);
xor (n6917,n6914,n6915);
or (n6918,n6919,n6922);
and (n6919,n6920,n6921);
xor (n6920,n6714,n6715);
and (n6921,n356,n185);
and (n6922,n6923,n6924);
xor (n6923,n6920,n6921);
or (n6924,n6925,n6927);
and (n6925,n6926,n804);
xor (n6926,n6720,n6721);
and (n6927,n6928,n6929);
xor (n6928,n6926,n804);
or (n6929,n6930,n6933);
and (n6930,n6931,n6932);
xor (n6931,n6726,n6727);
and (n6932,n33,n185);
and (n6933,n6934,n6935);
xor (n6934,n6931,n6932);
or (n6935,n6936,n6939);
and (n6936,n6937,n6938);
xor (n6937,n6732,n6733);
and (n6938,n64,n185);
and (n6939,n6940,n6941);
xor (n6940,n6937,n6938);
or (n6941,n6942,n6945);
and (n6942,n6943,n6944);
xor (n6943,n6738,n6739);
and (n6944,n58,n185);
and (n6945,n6946,n6947);
xor (n6946,n6943,n6944);
or (n6947,n6948,n6951);
and (n6948,n6949,n6950);
xor (n6949,n6744,n6745);
and (n6950,n117,n185);
and (n6951,n6952,n6953);
xor (n6952,n6949,n6950);
or (n6953,n6954,n6957);
and (n6954,n6955,n6956);
xor (n6955,n6750,n6751);
and (n6956,n111,n185);
and (n6957,n6958,n6959);
xor (n6958,n6955,n6956);
or (n6959,n6960,n6963);
and (n6960,n6961,n6962);
xor (n6961,n6756,n6757);
and (n6962,n141,n185);
and (n6963,n6964,n6965);
xor (n6964,n6961,n6962);
or (n6965,n6966,n6969);
and (n6966,n6967,n6968);
xor (n6967,n6762,n6763);
and (n6968,n135,n185);
and (n6969,n6970,n6971);
xor (n6970,n6967,n6968);
or (n6971,n6972,n6975);
and (n6972,n6973,n6974);
xor (n6973,n6768,n6769);
and (n6974,n448,n185);
and (n6975,n6976,n6977);
xor (n6976,n6973,n6974);
or (n6977,n6978,n6981);
and (n6978,n6979,n6980);
xor (n6979,n6774,n6775);
and (n6980,n474,n185);
and (n6981,n6982,n6983);
xor (n6982,n6979,n6980);
or (n6983,n6984,n6987);
and (n6984,n6985,n6986);
xor (n6985,n6780,n6781);
and (n6986,n625,n185);
and (n6987,n6988,n6989);
xor (n6988,n6985,n6986);
or (n6989,n6990,n6993);
and (n6990,n6991,n6992);
xor (n6991,n6786,n6787);
and (n6992,n1037,n185);
and (n6993,n6994,n6995);
xor (n6994,n6991,n6992);
or (n6995,n6996,n6999);
and (n6996,n6997,n6998);
xor (n6997,n6792,n6793);
and (n6998,n1030,n185);
and (n6999,n7000,n7001);
xor (n7000,n6997,n6998);
or (n7001,n7002,n7005);
and (n7002,n7003,n7004);
xor (n7003,n6798,n6799);
and (n7004,n1002,n185);
and (n7005,n7006,n7007);
xor (n7006,n7003,n7004);
or (n7007,n7008,n7010);
and (n7008,n7009,n3026);
xor (n7009,n6804,n6805);
and (n7010,n7011,n7012);
xor (n7011,n7009,n3026);
or (n7012,n7013,n7015);
and (n7013,n7014,n3165);
xor (n7014,n6810,n6811);
and (n7015,n7016,n7017);
xor (n7016,n7014,n3165);
or (n7017,n7018,n7020);
and (n7018,n7019,n3222);
xor (n7019,n6816,n6817);
and (n7020,n7021,n7022);
xor (n7021,n7019,n3222);
or (n7022,n7023,n7026);
and (n7023,n7024,n7025);
xor (n7024,n6822,n6823);
and (n7025,n839,n185);
and (n7026,n7027,n7028);
xor (n7027,n7024,n7025);
and (n7028,n7029,n7030);
xor (n7029,n6828,n6829);
and (n7030,n887,n185);
and (n7031,n192,n178);
or (n7032,n7033,n7035);
and (n7033,n7034,n7031);
xor (n7034,n6836,n6837);
and (n7035,n7036,n7037);
xor (n7036,n7034,n7031);
or (n7037,n7038,n7040);
and (n7038,n7039,n7031);
xor (n7039,n6841,n6842);
and (n7040,n7041,n7042);
xor (n7041,n7039,n7031);
or (n7042,n7043,n7045);
and (n7043,n7044,n7031);
xor (n7044,n6846,n6847);
and (n7045,n7046,n7047);
xor (n7046,n7044,n7031);
or (n7047,n7048,n7051);
and (n7048,n7049,n7050);
xor (n7049,n6851,n6852);
and (n7050,n214,n178);
and (n7051,n7052,n7053);
xor (n7052,n7049,n7050);
or (n7053,n7054,n7057);
and (n7054,n7055,n7056);
xor (n7055,n6857,n6858);
and (n7056,n208,n178);
and (n7057,n7058,n7059);
xor (n7058,n7055,n7056);
or (n7059,n7060,n7063);
and (n7060,n7061,n7062);
xor (n7061,n6863,n6864);
and (n7062,n167,n178);
and (n7063,n7064,n7065);
xor (n7064,n7061,n7062);
or (n7065,n7066,n7069);
and (n7066,n7067,n7068);
xor (n7067,n6869,n6870);
and (n7068,n161,n178);
and (n7069,n7070,n7071);
xor (n7070,n7067,n7068);
or (n7071,n7072,n7075);
and (n7072,n7073,n7074);
xor (n7073,n6875,n6876);
and (n7074,n236,n178);
and (n7075,n7076,n7077);
xor (n7076,n7073,n7074);
or (n7077,n7078,n7081);
and (n7078,n7079,n7080);
xor (n7079,n6881,n6882);
and (n7080,n230,n178);
and (n7081,n7082,n7083);
xor (n7082,n7079,n7080);
or (n7083,n7084,n7087);
and (n7084,n7085,n7086);
xor (n7085,n6887,n6888);
and (n7086,n90,n178);
and (n7087,n7088,n7089);
xor (n7088,n7085,n7086);
or (n7089,n7090,n7093);
and (n7090,n7091,n7092);
xor (n7091,n6893,n6894);
and (n7092,n84,n178);
and (n7093,n7094,n7095);
xor (n7094,n7091,n7092);
or (n7095,n7096,n7099);
and (n7096,n7097,n7098);
xor (n7097,n6899,n6900);
and (n7098,n310,n178);
and (n7099,n7100,n7101);
xor (n7100,n7097,n7098);
or (n7101,n7102,n7105);
and (n7102,n7103,n7104);
xor (n7103,n6905,n6906);
and (n7104,n348,n178);
and (n7105,n7106,n7107);
xor (n7106,n7103,n7104);
or (n7107,n7108,n7111);
and (n7108,n7109,n7110);
xor (n7109,n6911,n6912);
and (n7110,n342,n178);
and (n7111,n7112,n7113);
xor (n7112,n7109,n7110);
or (n7113,n7114,n7117);
and (n7114,n7115,n7116);
xor (n7115,n6917,n6918);
and (n7116,n356,n178);
and (n7117,n7118,n7119);
xor (n7118,n7115,n7116);
or (n7119,n7120,n7123);
and (n7120,n7121,n7122);
xor (n7121,n6923,n6924);
and (n7122,n39,n178);
and (n7123,n7124,n7125);
xor (n7124,n7121,n7122);
or (n7125,n7126,n7129);
and (n7126,n7127,n7128);
xor (n7127,n6928,n6929);
and (n7128,n33,n178);
and (n7129,n7130,n7131);
xor (n7130,n7127,n7128);
or (n7131,n7132,n7135);
and (n7132,n7133,n7134);
xor (n7133,n6934,n6935);
and (n7134,n64,n178);
and (n7135,n7136,n7137);
xor (n7136,n7133,n7134);
or (n7137,n7138,n7141);
and (n7138,n7139,n7140);
xor (n7139,n6940,n6941);
and (n7140,n58,n178);
and (n7141,n7142,n7143);
xor (n7142,n7139,n7140);
or (n7143,n7144,n7147);
and (n7144,n7145,n7146);
xor (n7145,n6946,n6947);
and (n7146,n117,n178);
and (n7147,n7148,n7149);
xor (n7148,n7145,n7146);
or (n7149,n7150,n7153);
and (n7150,n7151,n7152);
xor (n7151,n6952,n6953);
and (n7152,n111,n178);
and (n7153,n7154,n7155);
xor (n7154,n7151,n7152);
or (n7155,n7156,n7159);
and (n7156,n7157,n7158);
xor (n7157,n6958,n6959);
and (n7158,n141,n178);
and (n7159,n7160,n7161);
xor (n7160,n7157,n7158);
or (n7161,n7162,n7165);
and (n7162,n7163,n7164);
xor (n7163,n6964,n6965);
and (n7164,n135,n178);
and (n7165,n7166,n7167);
xor (n7166,n7163,n7164);
or (n7167,n7168,n7171);
and (n7168,n7169,n7170);
xor (n7169,n6970,n6971);
and (n7170,n448,n178);
and (n7171,n7172,n7173);
xor (n7172,n7169,n7170);
or (n7173,n7174,n7177);
and (n7174,n7175,n7176);
xor (n7175,n6976,n6977);
and (n7176,n474,n178);
and (n7177,n7178,n7179);
xor (n7178,n7175,n7176);
or (n7179,n7180,n7183);
and (n7180,n7181,n7182);
xor (n7181,n6982,n6983);
and (n7182,n625,n178);
and (n7183,n7184,n7185);
xor (n7184,n7181,n7182);
or (n7185,n7186,n7189);
and (n7186,n7187,n7188);
xor (n7187,n6988,n6989);
and (n7188,n1037,n178);
and (n7189,n7190,n7191);
xor (n7190,n7187,n7188);
or (n7191,n7192,n7195);
and (n7192,n7193,n7194);
xor (n7193,n6994,n6995);
and (n7194,n1030,n178);
and (n7195,n7196,n7197);
xor (n7196,n7193,n7194);
or (n7197,n7198,n7201);
and (n7198,n7199,n7200);
xor (n7199,n7000,n7001);
and (n7200,n1002,n178);
and (n7201,n7202,n7203);
xor (n7202,n7199,n7200);
or (n7203,n7204,n7207);
and (n7204,n7205,n7206);
xor (n7205,n7006,n7007);
and (n7206,n832,n178);
and (n7207,n7208,n7209);
xor (n7208,n7205,n7206);
or (n7209,n7210,n7213);
and (n7210,n7211,n7212);
xor (n7211,n7011,n7012);
and (n7212,n826,n178);
and (n7213,n7214,n7215);
xor (n7214,n7211,n7212);
or (n7215,n7216,n7219);
and (n7216,n7217,n7218);
xor (n7217,n7016,n7017);
and (n7218,n847,n178);
and (n7219,n7220,n7221);
xor (n7220,n7217,n7218);
or (n7221,n7222,n7225);
and (n7222,n7223,n7224);
xor (n7223,n7021,n7022);
and (n7224,n839,n178);
and (n7225,n7226,n7227);
xor (n7226,n7223,n7224);
and (n7227,n7228,n3209);
xor (n7228,n7027,n7028);
and (n7229,n192,n180);
or (n7230,n7231,n7233);
and (n7231,n7232,n7229);
xor (n7232,n7036,n7037);
and (n7233,n7234,n7235);
xor (n7234,n7232,n7229);
or (n7235,n7236,n7238);
and (n7236,n7237,n7229);
xor (n7237,n7041,n7042);
and (n7238,n7239,n7240);
xor (n7239,n7237,n7229);
or (n7240,n7241,n7244);
and (n7241,n7242,n7243);
xor (n7242,n7046,n7047);
and (n7243,n214,n180);
and (n7244,n7245,n7246);
xor (n7245,n7242,n7243);
or (n7246,n7247,n7250);
and (n7247,n7248,n7249);
xor (n7248,n7052,n7053);
and (n7249,n208,n180);
and (n7250,n7251,n7252);
xor (n7251,n7248,n7249);
or (n7252,n7253,n7256);
and (n7253,n7254,n7255);
xor (n7254,n7058,n7059);
and (n7255,n167,n180);
and (n7256,n7257,n7258);
xor (n7257,n7254,n7255);
or (n7258,n7259,n7262);
and (n7259,n7260,n7261);
xor (n7260,n7064,n7065);
and (n7261,n161,n180);
and (n7262,n7263,n7264);
xor (n7263,n7260,n7261);
or (n7264,n7265,n7268);
and (n7265,n7266,n7267);
xor (n7266,n7070,n7071);
and (n7267,n236,n180);
and (n7268,n7269,n7270);
xor (n7269,n7266,n7267);
or (n7270,n7271,n7274);
and (n7271,n7272,n7273);
xor (n7272,n7076,n7077);
and (n7273,n230,n180);
and (n7274,n7275,n7276);
xor (n7275,n7272,n7273);
or (n7276,n7277,n7280);
and (n7277,n7278,n7279);
xor (n7278,n7082,n7083);
and (n7279,n90,n180);
and (n7280,n7281,n7282);
xor (n7281,n7278,n7279);
or (n7282,n7283,n7286);
and (n7283,n7284,n7285);
xor (n7284,n7088,n7089);
and (n7285,n84,n180);
and (n7286,n7287,n7288);
xor (n7287,n7284,n7285);
or (n7288,n7289,n7292);
and (n7289,n7290,n7291);
xor (n7290,n7094,n7095);
and (n7291,n310,n180);
and (n7292,n7293,n7294);
xor (n7293,n7290,n7291);
or (n7294,n7295,n7298);
and (n7295,n7296,n7297);
xor (n7296,n7100,n7101);
and (n7297,n348,n180);
and (n7298,n7299,n7300);
xor (n7299,n7296,n7297);
or (n7300,n7301,n7304);
and (n7301,n7302,n7303);
xor (n7302,n7106,n7107);
and (n7303,n342,n180);
and (n7304,n7305,n7306);
xor (n7305,n7302,n7303);
or (n7306,n7307,n7310);
and (n7307,n7308,n7309);
xor (n7308,n7112,n7113);
and (n7309,n356,n180);
and (n7310,n7311,n7312);
xor (n7311,n7308,n7309);
or (n7312,n7313,n7316);
and (n7313,n7314,n7315);
xor (n7314,n7118,n7119);
and (n7315,n39,n180);
and (n7316,n7317,n7318);
xor (n7317,n7314,n7315);
or (n7318,n7319,n7322);
and (n7319,n7320,n7321);
xor (n7320,n7124,n7125);
and (n7321,n33,n180);
and (n7322,n7323,n7324);
xor (n7323,n7320,n7321);
or (n7324,n7325,n7327);
and (n7325,n7326,n820);
xor (n7326,n7130,n7131);
and (n7327,n7328,n7329);
xor (n7328,n7326,n820);
or (n7329,n7330,n7333);
and (n7330,n7331,n7332);
xor (n7331,n7136,n7137);
and (n7332,n58,n180);
and (n7333,n7334,n7335);
xor (n7334,n7331,n7332);
or (n7335,n7336,n7339);
and (n7336,n7337,n7338);
xor (n7337,n7142,n7143);
and (n7338,n117,n180);
and (n7339,n7340,n7341);
xor (n7340,n7337,n7338);
or (n7341,n7342,n7345);
and (n7342,n7343,n7344);
xor (n7343,n7148,n7149);
and (n7344,n111,n180);
and (n7345,n7346,n7347);
xor (n7346,n7343,n7344);
or (n7347,n7348,n7351);
and (n7348,n7349,n7350);
xor (n7349,n7154,n7155);
and (n7350,n141,n180);
and (n7351,n7352,n7353);
xor (n7352,n7349,n7350);
or (n7353,n7354,n7357);
and (n7354,n7355,n7356);
xor (n7355,n7160,n7161);
and (n7356,n135,n180);
and (n7357,n7358,n7359);
xor (n7358,n7355,n7356);
or (n7359,n7360,n7363);
and (n7360,n7361,n7362);
xor (n7361,n7166,n7167);
and (n7362,n448,n180);
and (n7363,n7364,n7365);
xor (n7364,n7361,n7362);
or (n7365,n7366,n7369);
and (n7366,n7367,n7368);
xor (n7367,n7172,n7173);
and (n7368,n474,n180);
and (n7369,n7370,n7371);
xor (n7370,n7367,n7368);
or (n7371,n7372,n7375);
and (n7372,n7373,n7374);
xor (n7373,n7178,n7179);
and (n7374,n625,n180);
and (n7375,n7376,n7377);
xor (n7376,n7373,n7374);
or (n7377,n7378,n7381);
and (n7378,n7379,n7380);
xor (n7379,n7184,n7185);
and (n7380,n1037,n180);
and (n7381,n7382,n7383);
xor (n7382,n7379,n7380);
or (n7383,n7384,n7387);
and (n7384,n7385,n7386);
xor (n7385,n7190,n7191);
and (n7386,n1030,n180);
and (n7387,n7388,n7389);
xor (n7388,n7385,n7386);
or (n7389,n7390,n7393);
and (n7390,n7391,n7392);
xor (n7391,n7196,n7197);
and (n7392,n1002,n180);
and (n7393,n7394,n7395);
xor (n7394,n7391,n7392);
or (n7395,n7396,n7399);
and (n7396,n7397,n7398);
xor (n7397,n7202,n7203);
and (n7398,n832,n180);
and (n7399,n7400,n7401);
xor (n7400,n7397,n7398);
or (n7401,n7402,n7405);
and (n7402,n7403,n7404);
xor (n7403,n7208,n7209);
and (n7404,n826,n180);
and (n7405,n7406,n7407);
xor (n7406,n7403,n7404);
or (n7407,n7408,n7411);
and (n7408,n7409,n7410);
xor (n7409,n7214,n7215);
and (n7410,n847,n180);
and (n7411,n7412,n7413);
xor (n7412,n7409,n7410);
or (n7413,n7414,n7417);
and (n7414,n7415,n7416);
xor (n7415,n7220,n7221);
and (n7416,n839,n180);
and (n7417,n7418,n7419);
xor (n7418,n7415,n7416);
and (n7419,n7420,n7421);
xor (n7420,n7226,n7227);
and (n7421,n887,n180);
and (n7422,n192,n200);
or (n7423,n7424,n7426);
and (n7424,n7425,n7422);
xor (n7425,n7234,n7235);
and (n7426,n7427,n7428);
xor (n7427,n7425,n7422);
or (n7428,n7429,n7432);
and (n7429,n7430,n7431);
xor (n7430,n7239,n7240);
and (n7431,n214,n200);
and (n7432,n7433,n7434);
xor (n7433,n7430,n7431);
or (n7434,n7435,n7438);
and (n7435,n7436,n7437);
xor (n7436,n7245,n7246);
and (n7437,n208,n200);
and (n7438,n7439,n7440);
xor (n7439,n7436,n7437);
or (n7440,n7441,n7444);
and (n7441,n7442,n7443);
xor (n7442,n7251,n7252);
and (n7443,n167,n200);
and (n7444,n7445,n7446);
xor (n7445,n7442,n7443);
or (n7446,n7447,n7450);
and (n7447,n7448,n7449);
xor (n7448,n7257,n7258);
and (n7449,n161,n200);
and (n7450,n7451,n7452);
xor (n7451,n7448,n7449);
or (n7452,n7453,n7456);
and (n7453,n7454,n7455);
xor (n7454,n7263,n7264);
and (n7455,n236,n200);
and (n7456,n7457,n7458);
xor (n7457,n7454,n7455);
or (n7458,n7459,n7462);
and (n7459,n7460,n7461);
xor (n7460,n7269,n7270);
and (n7461,n230,n200);
and (n7462,n7463,n7464);
xor (n7463,n7460,n7461);
or (n7464,n7465,n7468);
and (n7465,n7466,n7467);
xor (n7466,n7275,n7276);
and (n7467,n90,n200);
and (n7468,n7469,n7470);
xor (n7469,n7466,n7467);
or (n7470,n7471,n7474);
and (n7471,n7472,n7473);
xor (n7472,n7281,n7282);
and (n7473,n84,n200);
and (n7474,n7475,n7476);
xor (n7475,n7472,n7473);
or (n7476,n7477,n7480);
and (n7477,n7478,n7479);
xor (n7478,n7287,n7288);
and (n7479,n310,n200);
and (n7480,n7481,n7482);
xor (n7481,n7478,n7479);
or (n7482,n7483,n7486);
and (n7483,n7484,n7485);
xor (n7484,n7293,n7294);
and (n7485,n348,n200);
and (n7486,n7487,n7488);
xor (n7487,n7484,n7485);
or (n7488,n7489,n7492);
and (n7489,n7490,n7491);
xor (n7490,n7299,n7300);
and (n7491,n342,n200);
and (n7492,n7493,n7494);
xor (n7493,n7490,n7491);
or (n7494,n7495,n7498);
and (n7495,n7496,n7497);
xor (n7496,n7305,n7306);
and (n7497,n356,n200);
and (n7498,n7499,n7500);
xor (n7499,n7496,n7497);
or (n7500,n7501,n7504);
and (n7501,n7502,n7503);
xor (n7502,n7311,n7312);
and (n7503,n39,n200);
and (n7504,n7505,n7506);
xor (n7505,n7502,n7503);
or (n7506,n7507,n7510);
and (n7507,n7508,n7509);
xor (n7508,n7317,n7318);
and (n7509,n33,n200);
and (n7510,n7511,n7512);
xor (n7511,n7508,n7509);
or (n7512,n7513,n7516);
and (n7513,n7514,n7515);
xor (n7514,n7323,n7324);
and (n7515,n64,n200);
and (n7516,n7517,n7518);
xor (n7517,n7514,n7515);
or (n7518,n7519,n7522);
and (n7519,n7520,n7521);
xor (n7520,n7328,n7329);
and (n7521,n58,n200);
and (n7522,n7523,n7524);
xor (n7523,n7520,n7521);
or (n7524,n7525,n7528);
and (n7525,n7526,n7527);
xor (n7526,n7334,n7335);
and (n7527,n117,n200);
and (n7528,n7529,n7530);
xor (n7529,n7526,n7527);
or (n7530,n7531,n7534);
and (n7531,n7532,n7533);
xor (n7532,n7340,n7341);
and (n7533,n111,n200);
and (n7534,n7535,n7536);
xor (n7535,n7532,n7533);
or (n7536,n7537,n7540);
and (n7537,n7538,n7539);
xor (n7538,n7346,n7347);
and (n7539,n141,n200);
and (n7540,n7541,n7542);
xor (n7541,n7538,n7539);
or (n7542,n7543,n7546);
and (n7543,n7544,n7545);
xor (n7544,n7352,n7353);
and (n7545,n135,n200);
and (n7546,n7547,n7548);
xor (n7547,n7544,n7545);
or (n7548,n7549,n7552);
and (n7549,n7550,n7551);
xor (n7550,n7358,n7359);
and (n7551,n448,n200);
and (n7552,n7553,n7554);
xor (n7553,n7550,n7551);
or (n7554,n7555,n7558);
and (n7555,n7556,n7557);
xor (n7556,n7364,n7365);
and (n7557,n474,n200);
and (n7558,n7559,n7560);
xor (n7559,n7556,n7557);
or (n7560,n7561,n7564);
and (n7561,n7562,n7563);
xor (n7562,n7370,n7371);
and (n7563,n625,n200);
and (n7564,n7565,n7566);
xor (n7565,n7562,n7563);
or (n7566,n7567,n7570);
and (n7567,n7568,n7569);
xor (n7568,n7376,n7377);
and (n7569,n1037,n200);
and (n7570,n7571,n7572);
xor (n7571,n7568,n7569);
or (n7572,n7573,n7576);
and (n7573,n7574,n7575);
xor (n7574,n7382,n7383);
and (n7575,n1030,n200);
and (n7576,n7577,n7578);
xor (n7577,n7574,n7575);
or (n7578,n7579,n7582);
and (n7579,n7580,n7581);
xor (n7580,n7388,n7389);
and (n7581,n1002,n200);
and (n7582,n7583,n7584);
xor (n7583,n7580,n7581);
or (n7584,n7585,n7588);
and (n7585,n7586,n7587);
xor (n7586,n7394,n7395);
and (n7587,n832,n200);
and (n7588,n7589,n7590);
xor (n7589,n7586,n7587);
or (n7590,n7591,n7594);
and (n7591,n7592,n7593);
xor (n7592,n7400,n7401);
and (n7593,n826,n200);
and (n7594,n7595,n7596);
xor (n7595,n7592,n7593);
or (n7596,n7597,n7600);
and (n7597,n7598,n7599);
xor (n7598,n7406,n7407);
and (n7599,n847,n200);
and (n7600,n7601,n7602);
xor (n7601,n7598,n7599);
or (n7602,n7603,n7606);
and (n7603,n7604,n7605);
xor (n7604,n7412,n7413);
and (n7605,n839,n200);
and (n7606,n7607,n7608);
xor (n7607,n7604,n7605);
and (n7608,n7609,n3126);
xor (n7609,n7418,n7419);
and (n7610,n192,n150);
or (n7611,n7612,n7615);
and (n7612,n7613,n7614);
xor (n7613,n7427,n7428);
and (n7614,n214,n150);
and (n7615,n7616,n7617);
xor (n7616,n7613,n7614);
or (n7617,n7618,n7621);
and (n7618,n7619,n7620);
xor (n7619,n7433,n7434);
and (n7620,n208,n150);
and (n7621,n7622,n7623);
xor (n7622,n7619,n7620);
or (n7623,n7624,n7627);
and (n7624,n7625,n7626);
xor (n7625,n7439,n7440);
and (n7626,n167,n150);
and (n7627,n7628,n7629);
xor (n7628,n7625,n7626);
or (n7629,n7630,n7633);
and (n7630,n7631,n7632);
xor (n7631,n7445,n7446);
and (n7632,n161,n150);
and (n7633,n7634,n7635);
xor (n7634,n7631,n7632);
or (n7635,n7636,n7639);
and (n7636,n7637,n7638);
xor (n7637,n7451,n7452);
and (n7638,n236,n150);
and (n7639,n7640,n7641);
xor (n7640,n7637,n7638);
or (n7641,n7642,n7645);
and (n7642,n7643,n7644);
xor (n7643,n7457,n7458);
and (n7644,n230,n150);
and (n7645,n7646,n7647);
xor (n7646,n7643,n7644);
or (n7647,n7648,n7651);
and (n7648,n7649,n7650);
xor (n7649,n7463,n7464);
and (n7650,n90,n150);
and (n7651,n7652,n7653);
xor (n7652,n7649,n7650);
or (n7653,n7654,n7657);
and (n7654,n7655,n7656);
xor (n7655,n7469,n7470);
and (n7656,n84,n150);
and (n7657,n7658,n7659);
xor (n7658,n7655,n7656);
or (n7659,n7660,n7663);
and (n7660,n7661,n7662);
xor (n7661,n7475,n7476);
and (n7662,n310,n150);
and (n7663,n7664,n7665);
xor (n7664,n7661,n7662);
or (n7665,n7666,n7669);
and (n7666,n7667,n7668);
xor (n7667,n7481,n7482);
and (n7668,n348,n150);
and (n7669,n7670,n7671);
xor (n7670,n7667,n7668);
or (n7671,n7672,n7675);
and (n7672,n7673,n7674);
xor (n7673,n7487,n7488);
and (n7674,n342,n150);
and (n7675,n7676,n7677);
xor (n7676,n7673,n7674);
or (n7677,n7678,n7681);
and (n7678,n7679,n7680);
xor (n7679,n7493,n7494);
and (n7680,n356,n150);
and (n7681,n7682,n7683);
xor (n7682,n7679,n7680);
or (n7683,n7684,n7687);
and (n7684,n7685,n7686);
xor (n7685,n7499,n7500);
and (n7686,n39,n150);
and (n7687,n7688,n7689);
xor (n7688,n7685,n7686);
or (n7689,n7690,n7693);
and (n7690,n7691,n7692);
xor (n7691,n7505,n7506);
and (n7692,n33,n150);
and (n7693,n7694,n7695);
xor (n7694,n7691,n7692);
or (n7695,n7696,n7699);
and (n7696,n7697,n7698);
xor (n7697,n7511,n7512);
and (n7698,n64,n150);
and (n7699,n7700,n7701);
xor (n7700,n7697,n7698);
or (n7701,n7702,n7705);
and (n7702,n7703,n7704);
xor (n7703,n7517,n7518);
and (n7704,n58,n150);
and (n7705,n7706,n7707);
xor (n7706,n7703,n7704);
or (n7707,n7708,n7711);
and (n7708,n7709,n7710);
xor (n7709,n7523,n7524);
and (n7710,n117,n150);
and (n7711,n7712,n7713);
xor (n7712,n7709,n7710);
or (n7713,n7714,n7717);
and (n7714,n7715,n7716);
xor (n7715,n7529,n7530);
and (n7716,n111,n150);
and (n7717,n7718,n7719);
xor (n7718,n7715,n7716);
or (n7719,n7720,n7723);
and (n7720,n7721,n7722);
xor (n7721,n7535,n7536);
and (n7722,n141,n150);
and (n7723,n7724,n7725);
xor (n7724,n7721,n7722);
or (n7725,n7726,n7729);
and (n7726,n7727,n7728);
xor (n7727,n7541,n7542);
and (n7728,n135,n150);
and (n7729,n7730,n7731);
xor (n7730,n7727,n7728);
or (n7731,n7732,n7735);
and (n7732,n7733,n7734);
xor (n7733,n7547,n7548);
and (n7734,n448,n150);
and (n7735,n7736,n7737);
xor (n7736,n7733,n7734);
or (n7737,n7738,n7741);
and (n7738,n7739,n7740);
xor (n7739,n7553,n7554);
and (n7740,n474,n150);
and (n7741,n7742,n7743);
xor (n7742,n7739,n7740);
or (n7743,n7744,n7747);
and (n7744,n7745,n7746);
xor (n7745,n7559,n7560);
and (n7746,n625,n150);
and (n7747,n7748,n7749);
xor (n7748,n7745,n7746);
or (n7749,n7750,n7753);
and (n7750,n7751,n7752);
xor (n7751,n7565,n7566);
and (n7752,n1037,n150);
and (n7753,n7754,n7755);
xor (n7754,n7751,n7752);
or (n7755,n7756,n7759);
and (n7756,n7757,n7758);
xor (n7757,n7571,n7572);
and (n7758,n1030,n150);
and (n7759,n7760,n7761);
xor (n7760,n7757,n7758);
or (n7761,n7762,n7765);
and (n7762,n7763,n7764);
xor (n7763,n7577,n7578);
and (n7764,n1002,n150);
and (n7765,n7766,n7767);
xor (n7766,n7763,n7764);
or (n7767,n7768,n7771);
and (n7768,n7769,n7770);
xor (n7769,n7583,n7584);
and (n7770,n832,n150);
and (n7771,n7772,n7773);
xor (n7772,n7769,n7770);
or (n7773,n7774,n7777);
and (n7774,n7775,n7776);
xor (n7775,n7589,n7590);
and (n7776,n826,n150);
and (n7777,n7778,n7779);
xor (n7778,n7775,n7776);
or (n7779,n7780,n7783);
and (n7780,n7781,n7782);
xor (n7781,n7595,n7596);
and (n7782,n847,n150);
and (n7783,n7784,n7785);
xor (n7784,n7781,n7782);
or (n7785,n7786,n7789);
and (n7786,n7787,n7788);
xor (n7787,n7601,n7602);
and (n7788,n839,n150);
and (n7789,n7790,n7791);
xor (n7790,n7787,n7788);
and (n7791,n7792,n7793);
xor (n7792,n7607,n7608);
and (n7793,n887,n150);
and (n7794,n214,n151);
or (n7795,n7796,n7799);
and (n7796,n7797,n7798);
xor (n7797,n7616,n7617);
and (n7798,n208,n151);
and (n7799,n7800,n7801);
xor (n7800,n7797,n7798);
or (n7801,n7802,n7805);
and (n7802,n7803,n7804);
xor (n7803,n7622,n7623);
and (n7804,n167,n151);
and (n7805,n7806,n7807);
xor (n7806,n7803,n7804);
or (n7807,n7808,n7811);
and (n7808,n7809,n7810);
xor (n7809,n7628,n7629);
and (n7810,n161,n151);
and (n7811,n7812,n7813);
xor (n7812,n7809,n7810);
or (n7813,n7814,n7817);
and (n7814,n7815,n7816);
xor (n7815,n7634,n7635);
and (n7816,n236,n151);
and (n7817,n7818,n7819);
xor (n7818,n7815,n7816);
or (n7819,n7820,n7823);
and (n7820,n7821,n7822);
xor (n7821,n7640,n7641);
and (n7822,n230,n151);
and (n7823,n7824,n7825);
xor (n7824,n7821,n7822);
or (n7825,n7826,n7829);
and (n7826,n7827,n7828);
xor (n7827,n7646,n7647);
and (n7828,n90,n151);
and (n7829,n7830,n7831);
xor (n7830,n7827,n7828);
or (n7831,n7832,n7835);
and (n7832,n7833,n7834);
xor (n7833,n7652,n7653);
and (n7834,n84,n151);
and (n7835,n7836,n7837);
xor (n7836,n7833,n7834);
or (n7837,n7838,n7841);
and (n7838,n7839,n7840);
xor (n7839,n7658,n7659);
and (n7840,n310,n151);
and (n7841,n7842,n7843);
xor (n7842,n7839,n7840);
or (n7843,n7844,n7847);
and (n7844,n7845,n7846);
xor (n7845,n7664,n7665);
and (n7846,n348,n151);
and (n7847,n7848,n7849);
xor (n7848,n7845,n7846);
or (n7849,n7850,n7853);
and (n7850,n7851,n7852);
xor (n7851,n7670,n7671);
and (n7852,n342,n151);
and (n7853,n7854,n7855);
xor (n7854,n7851,n7852);
or (n7855,n7856,n7859);
and (n7856,n7857,n7858);
xor (n7857,n7676,n7677);
and (n7858,n356,n151);
and (n7859,n7860,n7861);
xor (n7860,n7857,n7858);
or (n7861,n7862,n7865);
and (n7862,n7863,n7864);
xor (n7863,n7682,n7683);
and (n7864,n39,n151);
and (n7865,n7866,n7867);
xor (n7866,n7863,n7864);
or (n7867,n7868,n7871);
and (n7868,n7869,n7870);
xor (n7869,n7688,n7689);
and (n7870,n33,n151);
and (n7871,n7872,n7873);
xor (n7872,n7869,n7870);
or (n7873,n7874,n7877);
and (n7874,n7875,n7876);
xor (n7875,n7694,n7695);
and (n7876,n64,n151);
and (n7877,n7878,n7879);
xor (n7878,n7875,n7876);
or (n7879,n7880,n7883);
and (n7880,n7881,n7882);
xor (n7881,n7700,n7701);
and (n7882,n58,n151);
and (n7883,n7884,n7885);
xor (n7884,n7881,n7882);
or (n7885,n7886,n7889);
and (n7886,n7887,n7888);
xor (n7887,n7706,n7707);
and (n7888,n117,n151);
and (n7889,n7890,n7891);
xor (n7890,n7887,n7888);
or (n7891,n7892,n7895);
and (n7892,n7893,n7894);
xor (n7893,n7712,n7713);
and (n7894,n111,n151);
and (n7895,n7896,n7897);
xor (n7896,n7893,n7894);
or (n7897,n7898,n7901);
and (n7898,n7899,n7900);
xor (n7899,n7718,n7719);
and (n7900,n141,n151);
and (n7901,n7902,n7903);
xor (n7902,n7899,n7900);
or (n7903,n7904,n7907);
and (n7904,n7905,n7906);
xor (n7905,n7724,n7725);
and (n7906,n135,n151);
and (n7907,n7908,n7909);
xor (n7908,n7905,n7906);
or (n7909,n7910,n7913);
and (n7910,n7911,n7912);
xor (n7911,n7730,n7731);
and (n7912,n448,n151);
and (n7913,n7914,n7915);
xor (n7914,n7911,n7912);
or (n7915,n7916,n7919);
and (n7916,n7917,n7918);
xor (n7917,n7736,n7737);
and (n7918,n474,n151);
and (n7919,n7920,n7921);
xor (n7920,n7917,n7918);
or (n7921,n7922,n7925);
and (n7922,n7923,n7924);
xor (n7923,n7742,n7743);
and (n7924,n625,n151);
and (n7925,n7926,n7927);
xor (n7926,n7923,n7924);
or (n7927,n7928,n7931);
and (n7928,n7929,n7930);
xor (n7929,n7748,n7749);
and (n7930,n1037,n151);
and (n7931,n7932,n7933);
xor (n7932,n7929,n7930);
or (n7933,n7934,n7937);
and (n7934,n7935,n7936);
xor (n7935,n7754,n7755);
and (n7936,n1030,n151);
and (n7937,n7938,n7939);
xor (n7938,n7935,n7936);
or (n7939,n7940,n7943);
and (n7940,n7941,n7942);
xor (n7941,n7760,n7761);
and (n7942,n1002,n151);
and (n7943,n7944,n7945);
xor (n7944,n7941,n7942);
or (n7945,n7946,n7949);
and (n7946,n7947,n7948);
xor (n7947,n7766,n7767);
and (n7948,n832,n151);
and (n7949,n7950,n7951);
xor (n7950,n7947,n7948);
or (n7951,n7952,n7955);
and (n7952,n7953,n7954);
xor (n7953,n7772,n7773);
and (n7954,n826,n151);
and (n7955,n7956,n7957);
xor (n7956,n7953,n7954);
or (n7957,n7958,n7961);
and (n7958,n7959,n7960);
xor (n7959,n7778,n7779);
and (n7960,n847,n151);
and (n7961,n7962,n7963);
xor (n7962,n7959,n7960);
or (n7963,n7964,n7967);
and (n7964,n7965,n7966);
xor (n7965,n7784,n7785);
and (n7966,n839,n151);
and (n7967,n7968,n7969);
xor (n7968,n7965,n7966);
and (n7969,n7970,n3286);
xor (n7970,n7790,n7791);
and (n7971,n208,n157);
or (n7972,n7973,n7976);
and (n7973,n7974,n7975);
xor (n7974,n7800,n7801);
and (n7975,n167,n157);
and (n7976,n7977,n7978);
xor (n7977,n7974,n7975);
or (n7978,n7979,n7982);
and (n7979,n7980,n7981);
xor (n7980,n7806,n7807);
and (n7981,n161,n157);
and (n7982,n7983,n7984);
xor (n7983,n7980,n7981);
or (n7984,n7985,n7988);
and (n7985,n7986,n7987);
xor (n7986,n7812,n7813);
and (n7987,n236,n157);
and (n7988,n7989,n7990);
xor (n7989,n7986,n7987);
or (n7990,n7991,n7994);
and (n7991,n7992,n7993);
xor (n7992,n7818,n7819);
and (n7993,n230,n157);
and (n7994,n7995,n7996);
xor (n7995,n7992,n7993);
or (n7996,n7997,n8000);
and (n7997,n7998,n7999);
xor (n7998,n7824,n7825);
and (n7999,n90,n157);
and (n8000,n8001,n8002);
xor (n8001,n7998,n7999);
or (n8002,n8003,n8006);
and (n8003,n8004,n8005);
xor (n8004,n7830,n7831);
and (n8005,n84,n157);
and (n8006,n8007,n8008);
xor (n8007,n8004,n8005);
or (n8008,n8009,n8012);
and (n8009,n8010,n8011);
xor (n8010,n7836,n7837);
and (n8011,n310,n157);
and (n8012,n8013,n8014);
xor (n8013,n8010,n8011);
or (n8014,n8015,n8018);
and (n8015,n8016,n8017);
xor (n8016,n7842,n7843);
and (n8017,n348,n157);
and (n8018,n8019,n8020);
xor (n8019,n8016,n8017);
or (n8020,n8021,n8024);
and (n8021,n8022,n8023);
xor (n8022,n7848,n7849);
and (n8023,n342,n157);
and (n8024,n8025,n8026);
xor (n8025,n8022,n8023);
or (n8026,n8027,n8030);
and (n8027,n8028,n8029);
xor (n8028,n7854,n7855);
and (n8029,n356,n157);
and (n8030,n8031,n8032);
xor (n8031,n8028,n8029);
or (n8032,n8033,n8036);
and (n8033,n8034,n8035);
xor (n8034,n7860,n7861);
and (n8035,n39,n157);
and (n8036,n8037,n8038);
xor (n8037,n8034,n8035);
or (n8038,n8039,n8042);
and (n8039,n8040,n8041);
xor (n8040,n7866,n7867);
and (n8041,n33,n157);
and (n8042,n8043,n8044);
xor (n8043,n8040,n8041);
or (n8044,n8045,n8048);
and (n8045,n8046,n8047);
xor (n8046,n7872,n7873);
and (n8047,n64,n157);
and (n8048,n8049,n8050);
xor (n8049,n8046,n8047);
or (n8050,n8051,n8054);
and (n8051,n8052,n8053);
xor (n8052,n7878,n7879);
and (n8053,n58,n157);
and (n8054,n8055,n8056);
xor (n8055,n8052,n8053);
or (n8056,n8057,n8060);
and (n8057,n8058,n8059);
xor (n8058,n7884,n7885);
and (n8059,n117,n157);
and (n8060,n8061,n8062);
xor (n8061,n8058,n8059);
or (n8062,n8063,n8066);
and (n8063,n8064,n8065);
xor (n8064,n7890,n7891);
and (n8065,n111,n157);
and (n8066,n8067,n8068);
xor (n8067,n8064,n8065);
or (n8068,n8069,n8071);
and (n8069,n8070,n789);
xor (n8070,n7896,n7897);
and (n8071,n8072,n8073);
xor (n8072,n8070,n789);
or (n8073,n8074,n8076);
and (n8074,n8075,n785);
xor (n8075,n7902,n7903);
and (n8076,n8077,n8078);
xor (n8077,n8075,n785);
or (n8078,n8079,n8082);
and (n8079,n8080,n8081);
xor (n8080,n7908,n7909);
and (n8081,n448,n157);
and (n8082,n8083,n8084);
xor (n8083,n8080,n8081);
or (n8084,n8085,n8088);
and (n8085,n8086,n8087);
xor (n8086,n7914,n7915);
and (n8087,n474,n157);
and (n8088,n8089,n8090);
xor (n8089,n8086,n8087);
or (n8090,n8091,n8093);
and (n8091,n8092,n1391);
xor (n8092,n7920,n7921);
and (n8093,n8094,n8095);
xor (n8094,n8092,n1391);
or (n8095,n8096,n8099);
and (n8096,n8097,n8098);
xor (n8097,n7926,n7927);
and (n8098,n1037,n157);
and (n8099,n8100,n8101);
xor (n8100,n8097,n8098);
or (n8101,n8102,n8104);
and (n8102,n8103,n1711);
xor (n8103,n7932,n7933);
and (n8104,n8105,n8106);
xor (n8105,n8103,n1711);
or (n8106,n8107,n8109);
and (n8107,n8108,n1764);
xor (n8108,n7938,n7939);
and (n8109,n8110,n8111);
xor (n8110,n8108,n1764);
or (n8111,n8112,n8114);
and (n8112,n8113,n1910);
xor (n8113,n7944,n7945);
and (n8114,n8115,n8116);
xor (n8115,n8113,n1910);
or (n8116,n8117,n8120);
and (n8117,n8118,n8119);
xor (n8118,n7950,n7951);
and (n8119,n826,n157);
and (n8120,n8121,n8122);
xor (n8121,n8118,n8119);
or (n8122,n8123,n8126);
and (n8123,n8124,n8125);
xor (n8124,n7956,n7957);
and (n8125,n847,n157);
and (n8126,n8127,n8128);
xor (n8127,n8124,n8125);
or (n8128,n8129,n8132);
and (n8129,n8130,n8131);
xor (n8130,n7962,n7963);
and (n8131,n839,n157);
and (n8132,n8133,n8134);
xor (n8133,n8130,n8131);
and (n8134,n8135,n8136);
xor (n8135,n7968,n7969);
and (n8136,n887,n157);
and (n8137,n167,n222);
or (n8138,n8139,n8142);
and (n8139,n8140,n8141);
xor (n8140,n7977,n7978);
and (n8141,n161,n222);
and (n8142,n8143,n8144);
xor (n8143,n8140,n8141);
or (n8144,n8145,n8148);
and (n8145,n8146,n8147);
xor (n8146,n7983,n7984);
and (n8147,n236,n222);
and (n8148,n8149,n8150);
xor (n8149,n8146,n8147);
or (n8150,n8151,n8154);
and (n8151,n8152,n8153);
xor (n8152,n7989,n7990);
and (n8153,n230,n222);
and (n8154,n8155,n8156);
xor (n8155,n8152,n8153);
or (n8156,n8157,n8160);
and (n8157,n8158,n8159);
xor (n8158,n7995,n7996);
and (n8159,n90,n222);
and (n8160,n8161,n8162);
xor (n8161,n8158,n8159);
or (n8162,n8163,n8166);
and (n8163,n8164,n8165);
xor (n8164,n8001,n8002);
and (n8165,n84,n222);
and (n8166,n8167,n8168);
xor (n8167,n8164,n8165);
or (n8168,n8169,n8172);
and (n8169,n8170,n8171);
xor (n8170,n8007,n8008);
and (n8171,n310,n222);
and (n8172,n8173,n8174);
xor (n8173,n8170,n8171);
or (n8174,n8175,n8178);
and (n8175,n8176,n8177);
xor (n8176,n8013,n8014);
and (n8177,n348,n222);
and (n8178,n8179,n8180);
xor (n8179,n8176,n8177);
or (n8180,n8181,n8184);
and (n8181,n8182,n8183);
xor (n8182,n8019,n8020);
and (n8183,n342,n222);
and (n8184,n8185,n8186);
xor (n8185,n8182,n8183);
or (n8186,n8187,n8190);
and (n8187,n8188,n8189);
xor (n8188,n8025,n8026);
and (n8189,n356,n222);
and (n8190,n8191,n8192);
xor (n8191,n8188,n8189);
or (n8192,n8193,n8196);
and (n8193,n8194,n8195);
xor (n8194,n8031,n8032);
and (n8195,n39,n222);
and (n8196,n8197,n8198);
xor (n8197,n8194,n8195);
or (n8198,n8199,n8202);
and (n8199,n8200,n8201);
xor (n8200,n8037,n8038);
and (n8201,n33,n222);
and (n8202,n8203,n8204);
xor (n8203,n8200,n8201);
or (n8204,n8205,n8208);
and (n8205,n8206,n8207);
xor (n8206,n8043,n8044);
and (n8207,n64,n222);
and (n8208,n8209,n8210);
xor (n8209,n8206,n8207);
or (n8210,n8211,n8214);
and (n8211,n8212,n8213);
xor (n8212,n8049,n8050);
and (n8213,n58,n222);
and (n8214,n8215,n8216);
xor (n8215,n8212,n8213);
or (n8216,n8217,n8220);
and (n8217,n8218,n8219);
xor (n8218,n8055,n8056);
and (n8219,n117,n222);
and (n8220,n8221,n8222);
xor (n8221,n8218,n8219);
or (n8222,n8223,n8226);
and (n8223,n8224,n8225);
xor (n8224,n8061,n8062);
and (n8225,n111,n222);
and (n8226,n8227,n8228);
xor (n8227,n8224,n8225);
or (n8228,n8229,n8232);
and (n8229,n8230,n8231);
xor (n8230,n8067,n8068);
and (n8231,n141,n222);
and (n8232,n8233,n8234);
xor (n8233,n8230,n8231);
or (n8234,n8235,n8238);
and (n8235,n8236,n8237);
xor (n8236,n8072,n8073);
and (n8237,n135,n222);
and (n8238,n8239,n8240);
xor (n8239,n8236,n8237);
or (n8240,n8241,n8244);
and (n8241,n8242,n8243);
xor (n8242,n8077,n8078);
and (n8243,n448,n222);
and (n8244,n8245,n8246);
xor (n8245,n8242,n8243);
or (n8246,n8247,n8250);
and (n8247,n8248,n8249);
xor (n8248,n8083,n8084);
and (n8249,n474,n222);
and (n8250,n8251,n8252);
xor (n8251,n8248,n8249);
or (n8252,n8253,n8256);
and (n8253,n8254,n8255);
xor (n8254,n8089,n8090);
and (n8255,n625,n222);
and (n8256,n8257,n8258);
xor (n8257,n8254,n8255);
or (n8258,n8259,n8262);
and (n8259,n8260,n8261);
xor (n8260,n8094,n8095);
and (n8261,n1037,n222);
and (n8262,n8263,n8264);
xor (n8263,n8260,n8261);
or (n8264,n8265,n8268);
and (n8265,n8266,n8267);
xor (n8266,n8100,n8101);
and (n8267,n1030,n222);
and (n8268,n8269,n8270);
xor (n8269,n8266,n8267);
or (n8270,n8271,n8274);
and (n8271,n8272,n8273);
xor (n8272,n8105,n8106);
and (n8273,n1002,n222);
and (n8274,n8275,n8276);
xor (n8275,n8272,n8273);
or (n8276,n8277,n8280);
and (n8277,n8278,n8279);
xor (n8278,n8110,n8111);
and (n8279,n832,n222);
and (n8280,n8281,n8282);
xor (n8281,n8278,n8279);
or (n8282,n8283,n8286);
and (n8283,n8284,n8285);
xor (n8284,n8115,n8116);
and (n8285,n826,n222);
and (n8286,n8287,n8288);
xor (n8287,n8284,n8285);
or (n8288,n8289,n8292);
and (n8289,n8290,n8291);
xor (n8290,n8121,n8122);
and (n8291,n847,n222);
and (n8292,n8293,n8294);
xor (n8293,n8290,n8291);
or (n8294,n8295,n8298);
and (n8295,n8296,n8297);
xor (n8296,n8127,n8128);
and (n8297,n839,n222);
and (n8298,n8299,n8300);
xor (n8299,n8296,n8297);
and (n8300,n8301,n2795);
xor (n8301,n8133,n8134);
and (n8302,n161,n75);
or (n8303,n8304,n8307);
and (n8304,n8305,n8306);
xor (n8305,n8143,n8144);
and (n8306,n236,n75);
and (n8307,n8308,n8309);
xor (n8308,n8305,n8306);
or (n8309,n8310,n8313);
and (n8310,n8311,n8312);
xor (n8311,n8149,n8150);
and (n8312,n230,n75);
and (n8313,n8314,n8315);
xor (n8314,n8311,n8312);
or (n8315,n8316,n8319);
and (n8316,n8317,n8318);
xor (n8317,n8155,n8156);
and (n8318,n90,n75);
and (n8319,n8320,n8321);
xor (n8320,n8317,n8318);
or (n8321,n8322,n8325);
and (n8322,n8323,n8324);
xor (n8323,n8161,n8162);
and (n8324,n84,n75);
and (n8325,n8326,n8327);
xor (n8326,n8323,n8324);
or (n8327,n8328,n8331);
and (n8328,n8329,n8330);
xor (n8329,n8167,n8168);
and (n8330,n310,n75);
and (n8331,n8332,n8333);
xor (n8332,n8329,n8330);
or (n8333,n8334,n8337);
and (n8334,n8335,n8336);
xor (n8335,n8173,n8174);
and (n8336,n348,n75);
and (n8337,n8338,n8339);
xor (n8338,n8335,n8336);
or (n8339,n8340,n8343);
and (n8340,n8341,n8342);
xor (n8341,n8179,n8180);
and (n8342,n342,n75);
and (n8343,n8344,n8345);
xor (n8344,n8341,n8342);
or (n8345,n8346,n8349);
and (n8346,n8347,n8348);
xor (n8347,n8185,n8186);
and (n8348,n356,n75);
and (n8349,n8350,n8351);
xor (n8350,n8347,n8348);
or (n8351,n8352,n8355);
and (n8352,n8353,n8354);
xor (n8353,n8191,n8192);
and (n8354,n39,n75);
and (n8355,n8356,n8357);
xor (n8356,n8353,n8354);
or (n8357,n8358,n8361);
and (n8358,n8359,n8360);
xor (n8359,n8197,n8198);
and (n8360,n33,n75);
and (n8361,n8362,n8363);
xor (n8362,n8359,n8360);
or (n8363,n8364,n8367);
and (n8364,n8365,n8366);
xor (n8365,n8203,n8204);
and (n8366,n64,n75);
and (n8367,n8368,n8369);
xor (n8368,n8365,n8366);
or (n8369,n8370,n8373);
and (n8370,n8371,n8372);
xor (n8371,n8209,n8210);
and (n8372,n58,n75);
and (n8373,n8374,n8375);
xor (n8374,n8371,n8372);
or (n8375,n8376,n8379);
and (n8376,n8377,n8378);
xor (n8377,n8215,n8216);
and (n8378,n117,n75);
and (n8379,n8380,n8381);
xor (n8380,n8377,n8378);
or (n8381,n8382,n8385);
and (n8382,n8383,n8384);
xor (n8383,n8221,n8222);
and (n8384,n111,n75);
and (n8385,n8386,n8387);
xor (n8386,n8383,n8384);
or (n8387,n8388,n8391);
and (n8388,n8389,n8390);
xor (n8389,n8227,n8228);
and (n8390,n141,n75);
and (n8391,n8392,n8393);
xor (n8392,n8389,n8390);
or (n8393,n8394,n8397);
and (n8394,n8395,n8396);
xor (n8395,n8233,n8234);
and (n8396,n135,n75);
and (n8397,n8398,n8399);
xor (n8398,n8395,n8396);
or (n8399,n8400,n8403);
and (n8400,n8401,n8402);
xor (n8401,n8239,n8240);
and (n8402,n448,n75);
and (n8403,n8404,n8405);
xor (n8404,n8401,n8402);
or (n8405,n8406,n8409);
and (n8406,n8407,n8408);
xor (n8407,n8245,n8246);
and (n8408,n474,n75);
and (n8409,n8410,n8411);
xor (n8410,n8407,n8408);
or (n8411,n8412,n8415);
and (n8412,n8413,n8414);
xor (n8413,n8251,n8252);
and (n8414,n625,n75);
and (n8415,n8416,n8417);
xor (n8416,n8413,n8414);
or (n8417,n8418,n8421);
and (n8418,n8419,n8420);
xor (n8419,n8257,n8258);
and (n8420,n1037,n75);
and (n8421,n8422,n8423);
xor (n8422,n8419,n8420);
or (n8423,n8424,n8427);
and (n8424,n8425,n8426);
xor (n8425,n8263,n8264);
and (n8426,n1030,n75);
and (n8427,n8428,n8429);
xor (n8428,n8425,n8426);
or (n8429,n8430,n8433);
and (n8430,n8431,n8432);
xor (n8431,n8269,n8270);
and (n8432,n1002,n75);
and (n8433,n8434,n8435);
xor (n8434,n8431,n8432);
or (n8435,n8436,n8439);
and (n8436,n8437,n8438);
xor (n8437,n8275,n8276);
and (n8438,n832,n75);
and (n8439,n8440,n8441);
xor (n8440,n8437,n8438);
or (n8441,n8442,n8445);
and (n8442,n8443,n8444);
xor (n8443,n8281,n8282);
and (n8444,n826,n75);
and (n8445,n8446,n8447);
xor (n8446,n8443,n8444);
or (n8447,n8448,n8451);
and (n8448,n8449,n8450);
xor (n8449,n8287,n8288);
and (n8450,n847,n75);
and (n8451,n8452,n8453);
xor (n8452,n8449,n8450);
or (n8453,n8454,n8457);
and (n8454,n8455,n8456);
xor (n8455,n8293,n8294);
and (n8456,n839,n75);
and (n8457,n8458,n8459);
xor (n8458,n8455,n8456);
and (n8459,n8460,n8461);
xor (n8460,n8299,n8300);
and (n8461,n887,n75);
and (n8462,n236,n73);
or (n8463,n8464,n8467);
and (n8464,n8465,n8466);
xor (n8465,n8308,n8309);
and (n8466,n230,n73);
and (n8467,n8468,n8469);
xor (n8468,n8465,n8466);
or (n8469,n8470,n8473);
and (n8470,n8471,n8472);
xor (n8471,n8314,n8315);
and (n8472,n90,n73);
and (n8473,n8474,n8475);
xor (n8474,n8471,n8472);
or (n8475,n8476,n8479);
and (n8476,n8477,n8478);
xor (n8477,n8320,n8321);
and (n8478,n84,n73);
and (n8479,n8480,n8481);
xor (n8480,n8477,n8478);
or (n8481,n8482,n8485);
and (n8482,n8483,n8484);
xor (n8483,n8326,n8327);
and (n8484,n310,n73);
and (n8485,n8486,n8487);
xor (n8486,n8483,n8484);
or (n8487,n8488,n8491);
and (n8488,n8489,n8490);
xor (n8489,n8332,n8333);
and (n8490,n348,n73);
and (n8491,n8492,n8493);
xor (n8492,n8489,n8490);
or (n8493,n8494,n8497);
and (n8494,n8495,n8496);
xor (n8495,n8338,n8339);
and (n8496,n342,n73);
and (n8497,n8498,n8499);
xor (n8498,n8495,n8496);
or (n8499,n8500,n8503);
and (n8500,n8501,n8502);
xor (n8501,n8344,n8345);
and (n8502,n356,n73);
and (n8503,n8504,n8505);
xor (n8504,n8501,n8502);
or (n8505,n8506,n8509);
and (n8506,n8507,n8508);
xor (n8507,n8350,n8351);
and (n8508,n39,n73);
and (n8509,n8510,n8511);
xor (n8510,n8507,n8508);
or (n8511,n8512,n8515);
and (n8512,n8513,n8514);
xor (n8513,n8356,n8357);
and (n8514,n33,n73);
and (n8515,n8516,n8517);
xor (n8516,n8513,n8514);
or (n8517,n8518,n8521);
and (n8518,n8519,n8520);
xor (n8519,n8362,n8363);
and (n8520,n64,n73);
and (n8521,n8522,n8523);
xor (n8522,n8519,n8520);
or (n8523,n8524,n8527);
and (n8524,n8525,n8526);
xor (n8525,n8368,n8369);
and (n8526,n58,n73);
and (n8527,n8528,n8529);
xor (n8528,n8525,n8526);
or (n8529,n8530,n8533);
and (n8530,n8531,n8532);
xor (n8531,n8374,n8375);
and (n8532,n117,n73);
and (n8533,n8534,n8535);
xor (n8534,n8531,n8532);
or (n8535,n8536,n8539);
and (n8536,n8537,n8538);
xor (n8537,n8380,n8381);
and (n8538,n111,n73);
and (n8539,n8540,n8541);
xor (n8540,n8537,n8538);
or (n8541,n8542,n8545);
and (n8542,n8543,n8544);
xor (n8543,n8386,n8387);
and (n8544,n141,n73);
and (n8545,n8546,n8547);
xor (n8546,n8543,n8544);
or (n8547,n8548,n8551);
and (n8548,n8549,n8550);
xor (n8549,n8392,n8393);
and (n8550,n135,n73);
and (n8551,n8552,n8553);
xor (n8552,n8549,n8550);
or (n8553,n8554,n8557);
and (n8554,n8555,n8556);
xor (n8555,n8398,n8399);
and (n8556,n448,n73);
and (n8557,n8558,n8559);
xor (n8558,n8555,n8556);
or (n8559,n8560,n8563);
and (n8560,n8561,n8562);
xor (n8561,n8404,n8405);
and (n8562,n474,n73);
and (n8563,n8564,n8565);
xor (n8564,n8561,n8562);
or (n8565,n8566,n8569);
and (n8566,n8567,n8568);
xor (n8567,n8410,n8411);
and (n8568,n625,n73);
and (n8569,n8570,n8571);
xor (n8570,n8567,n8568);
or (n8571,n8572,n8575);
and (n8572,n8573,n8574);
xor (n8573,n8416,n8417);
and (n8574,n1037,n73);
and (n8575,n8576,n8577);
xor (n8576,n8573,n8574);
or (n8577,n8578,n8581);
and (n8578,n8579,n8580);
xor (n8579,n8422,n8423);
and (n8580,n1030,n73);
and (n8581,n8582,n8583);
xor (n8582,n8579,n8580);
or (n8583,n8584,n8587);
and (n8584,n8585,n8586);
xor (n8585,n8428,n8429);
and (n8586,n1002,n73);
and (n8587,n8588,n8589);
xor (n8588,n8585,n8586);
or (n8589,n8590,n8593);
and (n8590,n8591,n8592);
xor (n8591,n8434,n8435);
and (n8592,n832,n73);
and (n8593,n8594,n8595);
xor (n8594,n8591,n8592);
or (n8595,n8596,n8599);
and (n8596,n8597,n8598);
xor (n8597,n8440,n8441);
and (n8598,n826,n73);
and (n8599,n8600,n8601);
xor (n8600,n8597,n8598);
or (n8601,n8602,n8605);
and (n8602,n8603,n8604);
xor (n8603,n8446,n8447);
and (n8604,n847,n73);
and (n8605,n8606,n8607);
xor (n8606,n8603,n8604);
or (n8607,n8608,n8611);
and (n8608,n8609,n8610);
xor (n8609,n8452,n8453);
and (n8610,n839,n73);
and (n8611,n8612,n8613);
xor (n8612,n8609,n8610);
and (n8613,n8614,n1871);
xor (n8614,n8458,n8459);
and (n8615,n230,n80);
or (n8616,n8617,n8620);
and (n8617,n8618,n8619);
xor (n8618,n8468,n8469);
and (n8619,n90,n80);
and (n8620,n8621,n8622);
xor (n8621,n8618,n8619);
or (n8622,n8623,n8626);
and (n8623,n8624,n8625);
xor (n8624,n8474,n8475);
and (n8625,n84,n80);
and (n8626,n8627,n8628);
xor (n8627,n8624,n8625);
or (n8628,n8629,n8632);
and (n8629,n8630,n8631);
xor (n8630,n8480,n8481);
and (n8631,n310,n80);
and (n8632,n8633,n8634);
xor (n8633,n8630,n8631);
or (n8634,n8635,n8638);
and (n8635,n8636,n8637);
xor (n8636,n8486,n8487);
and (n8637,n348,n80);
and (n8638,n8639,n8640);
xor (n8639,n8636,n8637);
or (n8640,n8641,n8644);
and (n8641,n8642,n8643);
xor (n8642,n8492,n8493);
and (n8643,n342,n80);
and (n8644,n8645,n8646);
xor (n8645,n8642,n8643);
or (n8646,n8647,n8650);
and (n8647,n8648,n8649);
xor (n8648,n8498,n8499);
and (n8649,n356,n80);
and (n8650,n8651,n8652);
xor (n8651,n8648,n8649);
or (n8652,n8653,n8656);
and (n8653,n8654,n8655);
xor (n8654,n8504,n8505);
and (n8655,n39,n80);
and (n8656,n8657,n8658);
xor (n8657,n8654,n8655);
or (n8658,n8659,n8662);
and (n8659,n8660,n8661);
xor (n8660,n8510,n8511);
and (n8661,n33,n80);
and (n8662,n8663,n8664);
xor (n8663,n8660,n8661);
or (n8664,n8665,n8668);
and (n8665,n8666,n8667);
xor (n8666,n8516,n8517);
and (n8667,n64,n80);
and (n8668,n8669,n8670);
xor (n8669,n8666,n8667);
or (n8670,n8671,n8674);
and (n8671,n8672,n8673);
xor (n8672,n8522,n8523);
and (n8673,n58,n80);
and (n8674,n8675,n8676);
xor (n8675,n8672,n8673);
or (n8676,n8677,n8680);
and (n8677,n8678,n8679);
xor (n8678,n8528,n8529);
and (n8679,n117,n80);
and (n8680,n8681,n8682);
xor (n8681,n8678,n8679);
or (n8682,n8683,n8686);
and (n8683,n8684,n8685);
xor (n8684,n8534,n8535);
and (n8685,n111,n80);
and (n8686,n8687,n8688);
xor (n8687,n8684,n8685);
or (n8688,n8689,n8692);
and (n8689,n8690,n8691);
xor (n8690,n8540,n8541);
and (n8691,n141,n80);
and (n8692,n8693,n8694);
xor (n8693,n8690,n8691);
or (n8694,n8695,n8698);
and (n8695,n8696,n8697);
xor (n8696,n8546,n8547);
and (n8697,n135,n80);
and (n8698,n8699,n8700);
xor (n8699,n8696,n8697);
or (n8700,n8701,n8704);
and (n8701,n8702,n8703);
xor (n8702,n8552,n8553);
and (n8703,n448,n80);
and (n8704,n8705,n8706);
xor (n8705,n8702,n8703);
or (n8706,n8707,n8710);
and (n8707,n8708,n8709);
xor (n8708,n8558,n8559);
and (n8709,n474,n80);
and (n8710,n8711,n8712);
xor (n8711,n8708,n8709);
or (n8712,n8713,n8715);
and (n8713,n8714,n1021);
xor (n8714,n8564,n8565);
and (n8715,n8716,n8717);
xor (n8716,n8714,n1021);
or (n8717,n8718,n8721);
and (n8718,n8719,n8720);
xor (n8719,n8570,n8571);
and (n8720,n1037,n80);
and (n8721,n8722,n8723);
xor (n8722,n8719,n8720);
or (n8723,n8724,n8727);
and (n8724,n8725,n8726);
xor (n8725,n8576,n8577);
and (n8726,n1030,n80);
and (n8727,n8728,n8729);
xor (n8728,n8725,n8726);
or (n8729,n8730,n8733);
and (n8730,n8731,n8732);
xor (n8731,n8582,n8583);
and (n8732,n1002,n80);
and (n8733,n8734,n8735);
xor (n8734,n8731,n8732);
or (n8735,n8736,n8738);
and (n8736,n8737,n1139);
xor (n8737,n8588,n8589);
and (n8738,n8739,n8740);
xor (n8739,n8737,n1139);
or (n8740,n8741,n8743);
and (n8741,n8742,n1505);
xor (n8742,n8594,n8595);
and (n8743,n8744,n8745);
xor (n8744,n8742,n1505);
or (n8745,n8746,n8749);
and (n8746,n8747,n8748);
xor (n8747,n8600,n8601);
and (n8748,n847,n80);
and (n8749,n8750,n8751);
xor (n8750,n8747,n8748);
or (n8751,n8752,n8755);
and (n8752,n8753,n8754);
xor (n8753,n8606,n8607);
and (n8754,n839,n80);
and (n8755,n8756,n8757);
xor (n8756,n8753,n8754);
and (n8757,n8758,n8759);
xor (n8758,n8612,n8613);
and (n8759,n887,n80);
and (n8760,n90,n301);
or (n8761,n8762,n8765);
and (n8762,n8763,n8764);
xor (n8763,n8621,n8622);
and (n8764,n84,n301);
and (n8765,n8766,n8767);
xor (n8766,n8763,n8764);
or (n8767,n8768,n8771);
and (n8768,n8769,n8770);
xor (n8769,n8627,n8628);
and (n8770,n310,n301);
and (n8771,n8772,n8773);
xor (n8772,n8769,n8770);
or (n8773,n8774,n8777);
and (n8774,n8775,n8776);
xor (n8775,n8633,n8634);
and (n8776,n348,n301);
and (n8777,n8778,n8779);
xor (n8778,n8775,n8776);
or (n8779,n8780,n8783);
and (n8780,n8781,n8782);
xor (n8781,n8639,n8640);
and (n8782,n342,n301);
and (n8783,n8784,n8785);
xor (n8784,n8781,n8782);
or (n8785,n8786,n8789);
and (n8786,n8787,n8788);
xor (n8787,n8645,n8646);
and (n8788,n356,n301);
and (n8789,n8790,n8791);
xor (n8790,n8787,n8788);
or (n8791,n8792,n8795);
and (n8792,n8793,n8794);
xor (n8793,n8651,n8652);
and (n8794,n39,n301);
and (n8795,n8796,n8797);
xor (n8796,n8793,n8794);
or (n8797,n8798,n8801);
and (n8798,n8799,n8800);
xor (n8799,n8657,n8658);
and (n8800,n33,n301);
and (n8801,n8802,n8803);
xor (n8802,n8799,n8800);
or (n8803,n8804,n8807);
and (n8804,n8805,n8806);
xor (n8805,n8663,n8664);
and (n8806,n64,n301);
and (n8807,n8808,n8809);
xor (n8808,n8805,n8806);
or (n8809,n8810,n8813);
and (n8810,n8811,n8812);
xor (n8811,n8669,n8670);
and (n8812,n58,n301);
and (n8813,n8814,n8815);
xor (n8814,n8811,n8812);
or (n8815,n8816,n8819);
and (n8816,n8817,n8818);
xor (n8817,n8675,n8676);
and (n8818,n117,n301);
and (n8819,n8820,n8821);
xor (n8820,n8817,n8818);
or (n8821,n8822,n8825);
and (n8822,n8823,n8824);
xor (n8823,n8681,n8682);
and (n8824,n111,n301);
and (n8825,n8826,n8827);
xor (n8826,n8823,n8824);
or (n8827,n8828,n8831);
and (n8828,n8829,n8830);
xor (n8829,n8687,n8688);
and (n8830,n141,n301);
and (n8831,n8832,n8833);
xor (n8832,n8829,n8830);
or (n8833,n8834,n8837);
and (n8834,n8835,n8836);
xor (n8835,n8693,n8694);
and (n8836,n135,n301);
and (n8837,n8838,n8839);
xor (n8838,n8835,n8836);
or (n8839,n8840,n8843);
and (n8840,n8841,n8842);
xor (n8841,n8699,n8700);
and (n8842,n448,n301);
and (n8843,n8844,n8845);
xor (n8844,n8841,n8842);
or (n8845,n8846,n8849);
and (n8846,n8847,n8848);
xor (n8847,n8705,n8706);
and (n8848,n474,n301);
and (n8849,n8850,n8851);
xor (n8850,n8847,n8848);
or (n8851,n8852,n8855);
and (n8852,n8853,n8854);
xor (n8853,n8711,n8712);
and (n8854,n625,n301);
and (n8855,n8856,n8857);
xor (n8856,n8853,n8854);
or (n8857,n8858,n8861);
and (n8858,n8859,n8860);
xor (n8859,n8716,n8717);
and (n8860,n1037,n301);
and (n8861,n8862,n8863);
xor (n8862,n8859,n8860);
or (n8863,n8864,n8867);
and (n8864,n8865,n8866);
xor (n8865,n8722,n8723);
and (n8866,n1030,n301);
and (n8867,n8868,n8869);
xor (n8868,n8865,n8866);
or (n8869,n8870,n8873);
and (n8870,n8871,n8872);
xor (n8871,n8728,n8729);
and (n8872,n1002,n301);
and (n8873,n8874,n8875);
xor (n8874,n8871,n8872);
or (n8875,n8876,n8879);
and (n8876,n8877,n8878);
xor (n8877,n8734,n8735);
and (n8878,n832,n301);
and (n8879,n8880,n8881);
xor (n8880,n8877,n8878);
or (n8881,n8882,n8885);
and (n8882,n8883,n8884);
xor (n8883,n8739,n8740);
and (n8884,n826,n301);
and (n8885,n8886,n8887);
xor (n8886,n8883,n8884);
or (n8887,n8888,n8891);
and (n8888,n8889,n8890);
xor (n8889,n8744,n8745);
and (n8890,n847,n301);
and (n8891,n8892,n8893);
xor (n8892,n8889,n8890);
or (n8893,n8894,n8897);
and (n8894,n8895,n8896);
xor (n8895,n8750,n8751);
and (n8896,n839,n301);
and (n8897,n8898,n8899);
xor (n8898,n8895,n8896);
and (n8899,n8900,n1633);
xor (n8900,n8756,n8757);
and (n8901,n84,n306);
or (n8902,n8903,n8906);
and (n8903,n8904,n8905);
xor (n8904,n8766,n8767);
and (n8905,n310,n306);
and (n8906,n8907,n8908);
xor (n8907,n8904,n8905);
or (n8908,n8909,n8912);
and (n8909,n8910,n8911);
xor (n8910,n8772,n8773);
and (n8911,n348,n306);
and (n8912,n8913,n8914);
xor (n8913,n8910,n8911);
or (n8914,n8915,n8918);
and (n8915,n8916,n8917);
xor (n8916,n8778,n8779);
and (n8917,n342,n306);
and (n8918,n8919,n8920);
xor (n8919,n8916,n8917);
or (n8920,n8921,n8924);
and (n8921,n8922,n8923);
xor (n8922,n8784,n8785);
and (n8923,n356,n306);
and (n8924,n8925,n8926);
xor (n8925,n8922,n8923);
or (n8926,n8927,n8930);
and (n8927,n8928,n8929);
xor (n8928,n8790,n8791);
and (n8929,n39,n306);
and (n8930,n8931,n8932);
xor (n8931,n8928,n8929);
or (n8932,n8933,n8936);
and (n8933,n8934,n8935);
xor (n8934,n8796,n8797);
and (n8935,n33,n306);
and (n8936,n8937,n8938);
xor (n8937,n8934,n8935);
or (n8938,n8939,n8942);
and (n8939,n8940,n8941);
xor (n8940,n8802,n8803);
and (n8941,n64,n306);
and (n8942,n8943,n8944);
xor (n8943,n8940,n8941);
or (n8944,n8945,n8948);
and (n8945,n8946,n8947);
xor (n8946,n8808,n8809);
and (n8947,n58,n306);
and (n8948,n8949,n8950);
xor (n8949,n8946,n8947);
or (n8950,n8951,n8954);
and (n8951,n8952,n8953);
xor (n8952,n8814,n8815);
and (n8953,n117,n306);
and (n8954,n8955,n8956);
xor (n8955,n8952,n8953);
or (n8956,n8957,n8960);
and (n8957,n8958,n8959);
xor (n8958,n8820,n8821);
and (n8959,n111,n306);
and (n8960,n8961,n8962);
xor (n8961,n8958,n8959);
or (n8962,n8963,n8966);
and (n8963,n8964,n8965);
xor (n8964,n8826,n8827);
and (n8965,n141,n306);
and (n8966,n8967,n8968);
xor (n8967,n8964,n8965);
or (n8968,n8969,n8972);
and (n8969,n8970,n8971);
xor (n8970,n8832,n8833);
and (n8971,n135,n306);
and (n8972,n8973,n8974);
xor (n8973,n8970,n8971);
or (n8974,n8975,n8978);
and (n8975,n8976,n8977);
xor (n8976,n8838,n8839);
and (n8977,n448,n306);
and (n8978,n8979,n8980);
xor (n8979,n8976,n8977);
or (n8980,n8981,n8984);
and (n8981,n8982,n8983);
xor (n8982,n8844,n8845);
and (n8983,n474,n306);
and (n8984,n8985,n8986);
xor (n8985,n8982,n8983);
or (n8986,n8987,n8990);
and (n8987,n8988,n8989);
xor (n8988,n8850,n8851);
and (n8989,n625,n306);
and (n8990,n8991,n8992);
xor (n8991,n8988,n8989);
or (n8992,n8993,n8996);
and (n8993,n8994,n8995);
xor (n8994,n8856,n8857);
and (n8995,n1037,n306);
and (n8996,n8997,n8998);
xor (n8997,n8994,n8995);
or (n8998,n8999,n9002);
and (n8999,n9000,n9001);
xor (n9000,n8862,n8863);
and (n9001,n1030,n306);
and (n9002,n9003,n9004);
xor (n9003,n9000,n9001);
or (n9004,n9005,n9008);
and (n9005,n9006,n9007);
xor (n9006,n8868,n8869);
and (n9007,n1002,n306);
and (n9008,n9009,n9010);
xor (n9009,n9006,n9007);
or (n9010,n9011,n9014);
and (n9011,n9012,n9013);
xor (n9012,n8874,n8875);
and (n9013,n832,n306);
and (n9014,n9015,n9016);
xor (n9015,n9012,n9013);
or (n9016,n9017,n9020);
and (n9017,n9018,n9019);
xor (n9018,n8880,n8881);
and (n9019,n826,n306);
and (n9020,n9021,n9022);
xor (n9021,n9018,n9019);
or (n9022,n9023,n9026);
and (n9023,n9024,n9025);
xor (n9024,n8886,n8887);
and (n9025,n847,n306);
and (n9026,n9027,n9028);
xor (n9027,n9024,n9025);
or (n9028,n9029,n9032);
and (n9029,n9030,n9031);
xor (n9030,n8892,n8893);
and (n9031,n839,n306);
and (n9032,n9033,n9034);
xor (n9033,n9030,n9031);
and (n9034,n9035,n9036);
xor (n9035,n8898,n8899);
and (n9036,n887,n306);
and (n9037,n310,n335);
or (n9038,n9039,n9042);
and (n9039,n9040,n9041);
xor (n9040,n8907,n8908);
and (n9041,n348,n335);
and (n9042,n9043,n9044);
xor (n9043,n9040,n9041);
or (n9044,n9045,n9048);
and (n9045,n9046,n9047);
xor (n9046,n8913,n8914);
and (n9047,n342,n335);
and (n9048,n9049,n9050);
xor (n9049,n9046,n9047);
or (n9050,n9051,n9054);
and (n9051,n9052,n9053);
xor (n9052,n8919,n8920);
and (n9053,n356,n335);
and (n9054,n9055,n9056);
xor (n9055,n9052,n9053);
or (n9056,n9057,n9060);
and (n9057,n9058,n9059);
xor (n9058,n8925,n8926);
and (n9059,n39,n335);
and (n9060,n9061,n9062);
xor (n9061,n9058,n9059);
or (n9062,n9063,n9066);
and (n9063,n9064,n9065);
xor (n9064,n8931,n8932);
and (n9065,n33,n335);
and (n9066,n9067,n9068);
xor (n9067,n9064,n9065);
or (n9068,n9069,n9072);
and (n9069,n9070,n9071);
xor (n9070,n8937,n8938);
and (n9071,n64,n335);
and (n9072,n9073,n9074);
xor (n9073,n9070,n9071);
or (n9074,n9075,n9078);
and (n9075,n9076,n9077);
xor (n9076,n8943,n8944);
and (n9077,n58,n335);
and (n9078,n9079,n9080);
xor (n9079,n9076,n9077);
or (n9080,n9081,n9084);
and (n9081,n9082,n9083);
xor (n9082,n8949,n8950);
and (n9083,n117,n335);
and (n9084,n9085,n9086);
xor (n9085,n9082,n9083);
or (n9086,n9087,n9090);
and (n9087,n9088,n9089);
xor (n9088,n8955,n8956);
and (n9089,n111,n335);
and (n9090,n9091,n9092);
xor (n9091,n9088,n9089);
or (n9092,n9093,n9096);
and (n9093,n9094,n9095);
xor (n9094,n8961,n8962);
and (n9095,n141,n335);
and (n9096,n9097,n9098);
xor (n9097,n9094,n9095);
or (n9098,n9099,n9102);
and (n9099,n9100,n9101);
xor (n9100,n8967,n8968);
and (n9101,n135,n335);
and (n9102,n9103,n9104);
xor (n9103,n9100,n9101);
or (n9104,n9105,n9108);
and (n9105,n9106,n9107);
xor (n9106,n8973,n8974);
and (n9107,n448,n335);
and (n9108,n9109,n9110);
xor (n9109,n9106,n9107);
or (n9110,n9111,n9114);
and (n9111,n9112,n9113);
xor (n9112,n8979,n8980);
and (n9113,n474,n335);
and (n9114,n9115,n9116);
xor (n9115,n9112,n9113);
or (n9116,n9117,n9120);
and (n9117,n9118,n9119);
xor (n9118,n8985,n8986);
and (n9119,n625,n335);
and (n9120,n9121,n9122);
xor (n9121,n9118,n9119);
or (n9122,n9123,n9126);
and (n9123,n9124,n9125);
xor (n9124,n8991,n8992);
and (n9125,n1037,n335);
and (n9126,n9127,n9128);
xor (n9127,n9124,n9125);
or (n9128,n9129,n9132);
and (n9129,n9130,n9131);
xor (n9130,n8997,n8998);
and (n9131,n1030,n335);
and (n9132,n9133,n9134);
xor (n9133,n9130,n9131);
or (n9134,n9135,n9138);
and (n9135,n9136,n9137);
xor (n9136,n9003,n9004);
and (n9137,n1002,n335);
and (n9138,n9139,n9140);
xor (n9139,n9136,n9137);
or (n9140,n9141,n9144);
and (n9141,n9142,n9143);
xor (n9142,n9009,n9010);
and (n9143,n832,n335);
and (n9144,n9145,n9146);
xor (n9145,n9142,n9143);
or (n9146,n9147,n9150);
and (n9147,n9148,n9149);
xor (n9148,n9015,n9016);
and (n9149,n826,n335);
and (n9150,n9151,n9152);
xor (n9151,n9148,n9149);
or (n9152,n9153,n9156);
and (n9153,n9154,n9155);
xor (n9154,n9021,n9022);
and (n9155,n847,n335);
and (n9156,n9157,n9158);
xor (n9157,n9154,n9155);
or (n9158,n9159,n9162);
and (n9159,n9160,n9161);
xor (n9160,n9027,n9028);
and (n9161,n839,n335);
and (n9162,n9163,n9164);
xor (n9163,n9160,n9161);
and (n9164,n9165,n1110);
xor (n9165,n9033,n9034);
and (n9166,n348,n22);
or (n9167,n9168,n9171);
and (n9168,n9169,n9170);
xor (n9169,n9043,n9044);
and (n9170,n342,n22);
and (n9171,n9172,n9173);
xor (n9172,n9169,n9170);
or (n9173,n9174,n9177);
and (n9174,n9175,n9176);
xor (n9175,n9049,n9050);
and (n9176,n356,n22);
and (n9177,n9178,n9179);
xor (n9178,n9175,n9176);
or (n9179,n9180,n9183);
and (n9180,n9181,n9182);
xor (n9181,n9055,n9056);
and (n9182,n39,n22);
and (n9183,n9184,n9185);
xor (n9184,n9181,n9182);
or (n9185,n9186,n9189);
and (n9186,n9187,n9188);
xor (n9187,n9061,n9062);
and (n9188,n33,n22);
and (n9189,n9190,n9191);
xor (n9190,n9187,n9188);
or (n9191,n9192,n9195);
and (n9192,n9193,n9194);
xor (n9193,n9067,n9068);
and (n9194,n64,n22);
and (n9195,n9196,n9197);
xor (n9196,n9193,n9194);
or (n9197,n9198,n9201);
and (n9198,n9199,n9200);
xor (n9199,n9073,n9074);
and (n9200,n58,n22);
and (n9201,n9202,n9203);
xor (n9202,n9199,n9200);
or (n9203,n9204,n9207);
and (n9204,n9205,n9206);
xor (n9205,n9079,n9080);
and (n9206,n117,n22);
and (n9207,n9208,n9209);
xor (n9208,n9205,n9206);
or (n9209,n9210,n9213);
and (n9210,n9211,n9212);
xor (n9211,n9085,n9086);
and (n9212,n111,n22);
and (n9213,n9214,n9215);
xor (n9214,n9211,n9212);
or (n9215,n9216,n9219);
and (n9216,n9217,n9218);
xor (n9217,n9091,n9092);
and (n9218,n141,n22);
and (n9219,n9220,n9221);
xor (n9220,n9217,n9218);
or (n9221,n9222,n9225);
and (n9222,n9223,n9224);
xor (n9223,n9097,n9098);
and (n9224,n135,n22);
and (n9225,n9226,n9227);
xor (n9226,n9223,n9224);
or (n9227,n9228,n9231);
and (n9228,n9229,n9230);
xor (n9229,n9103,n9104);
and (n9230,n448,n22);
and (n9231,n9232,n9233);
xor (n9232,n9229,n9230);
or (n9233,n9234,n9237);
and (n9234,n9235,n9236);
xor (n9235,n9109,n9110);
and (n9236,n474,n22);
and (n9237,n9238,n9239);
xor (n9238,n9235,n9236);
or (n9239,n9240,n9243);
and (n9240,n9241,n9242);
xor (n9241,n9115,n9116);
and (n9242,n625,n22);
and (n9243,n9244,n9245);
xor (n9244,n9241,n9242);
or (n9245,n9246,n9249);
and (n9246,n9247,n9248);
xor (n9247,n9121,n9122);
and (n9248,n1037,n22);
and (n9249,n9250,n9251);
xor (n9250,n9247,n9248);
or (n9251,n9252,n9255);
and (n9252,n9253,n9254);
xor (n9253,n9127,n9128);
and (n9254,n1030,n22);
and (n9255,n9256,n9257);
xor (n9256,n9253,n9254);
or (n9257,n9258,n9261);
and (n9258,n9259,n9260);
xor (n9259,n9133,n9134);
and (n9260,n1002,n22);
and (n9261,n9262,n9263);
xor (n9262,n9259,n9260);
or (n9263,n9264,n9267);
and (n9264,n9265,n9266);
xor (n9265,n9139,n9140);
and (n9266,n832,n22);
and (n9267,n9268,n9269);
xor (n9268,n9265,n9266);
or (n9269,n9270,n9273);
and (n9270,n9271,n9272);
xor (n9271,n9145,n9146);
and (n9272,n826,n22);
and (n9273,n9274,n9275);
xor (n9274,n9271,n9272);
or (n9275,n9276,n9279);
and (n9276,n9277,n9278);
xor (n9277,n9151,n9152);
and (n9278,n847,n22);
and (n9279,n9280,n9281);
xor (n9280,n9277,n9278);
or (n9281,n9282,n9285);
and (n9282,n9283,n9284);
xor (n9283,n9157,n9158);
and (n9284,n839,n22);
and (n9285,n9286,n9287);
xor (n9286,n9283,n9284);
and (n9287,n9288,n9289);
xor (n9288,n9163,n9164);
and (n9289,n887,n22);
and (n9290,n342,n23);
or (n9291,n9292,n9295);
and (n9292,n9293,n9294);
xor (n9293,n9172,n9173);
and (n9294,n356,n23);
and (n9295,n9296,n9297);
xor (n9296,n9293,n9294);
or (n9297,n9298,n9301);
and (n9298,n9299,n9300);
xor (n9299,n9178,n9179);
and (n9300,n39,n23);
and (n9301,n9302,n9303);
xor (n9302,n9299,n9300);
or (n9303,n9304,n9307);
and (n9304,n9305,n9306);
xor (n9305,n9184,n9185);
and (n9306,n33,n23);
and (n9307,n9308,n9309);
xor (n9308,n9305,n9306);
or (n9309,n9310,n9313);
and (n9310,n9311,n9312);
xor (n9311,n9190,n9191);
and (n9312,n64,n23);
and (n9313,n9314,n9315);
xor (n9314,n9311,n9312);
or (n9315,n9316,n9319);
and (n9316,n9317,n9318);
xor (n9317,n9196,n9197);
and (n9318,n58,n23);
and (n9319,n9320,n9321);
xor (n9320,n9317,n9318);
or (n9321,n9322,n9325);
and (n9322,n9323,n9324);
xor (n9323,n9202,n9203);
and (n9324,n117,n23);
and (n9325,n9326,n9327);
xor (n9326,n9323,n9324);
or (n9327,n9328,n9331);
and (n9328,n9329,n9330);
xor (n9329,n9208,n9209);
and (n9330,n111,n23);
and (n9331,n9332,n9333);
xor (n9332,n9329,n9330);
or (n9333,n9334,n9337);
and (n9334,n9335,n9336);
xor (n9335,n9214,n9215);
and (n9336,n141,n23);
and (n9337,n9338,n9339);
xor (n9338,n9335,n9336);
or (n9339,n9340,n9343);
and (n9340,n9341,n9342);
xor (n9341,n9220,n9221);
and (n9342,n135,n23);
and (n9343,n9344,n9345);
xor (n9344,n9341,n9342);
or (n9345,n9346,n9349);
and (n9346,n9347,n9348);
xor (n9347,n9226,n9227);
and (n9348,n448,n23);
and (n9349,n9350,n9351);
xor (n9350,n9347,n9348);
or (n9351,n9352,n9355);
and (n9352,n9353,n9354);
xor (n9353,n9232,n9233);
and (n9354,n474,n23);
and (n9355,n9356,n9357);
xor (n9356,n9353,n9354);
or (n9357,n9358,n9361);
and (n9358,n9359,n9360);
xor (n9359,n9238,n9239);
and (n9360,n625,n23);
and (n9361,n9362,n9363);
xor (n9362,n9359,n9360);
or (n9363,n9364,n9367);
and (n9364,n9365,n9366);
xor (n9365,n9244,n9245);
and (n9366,n1037,n23);
and (n9367,n9368,n9369);
xor (n9368,n9365,n9366);
or (n9369,n9370,n9373);
and (n9370,n9371,n9372);
xor (n9371,n9250,n9251);
and (n9372,n1030,n23);
and (n9373,n9374,n9375);
xor (n9374,n9371,n9372);
or (n9375,n9376,n9379);
and (n9376,n9377,n9378);
xor (n9377,n9256,n9257);
and (n9378,n1002,n23);
and (n9379,n9380,n9381);
xor (n9380,n9377,n9378);
or (n9381,n9382,n9385);
and (n9382,n9383,n9384);
xor (n9383,n9262,n9263);
and (n9384,n832,n23);
and (n9385,n9386,n9387);
xor (n9386,n9383,n9384);
or (n9387,n9388,n9391);
and (n9388,n9389,n9390);
xor (n9389,n9268,n9269);
and (n9390,n826,n23);
and (n9391,n9392,n9393);
xor (n9392,n9389,n9390);
or (n9393,n9394,n9397);
and (n9394,n9395,n9396);
xor (n9395,n9274,n9275);
and (n9396,n847,n23);
and (n9397,n9398,n9399);
xor (n9398,n9395,n9396);
or (n9399,n9400,n9403);
and (n9400,n9401,n9402);
xor (n9401,n9280,n9281);
and (n9402,n839,n23);
and (n9403,n9404,n9405);
xor (n9404,n9401,n9402);
and (n9405,n9406,n890);
xor (n9406,n9286,n9287);
and (n9407,n356,n29);
or (n9408,n9409,n9412);
and (n9409,n9410,n9411);
xor (n9410,n9296,n9297);
and (n9411,n39,n29);
and (n9412,n9413,n9414);
xor (n9413,n9410,n9411);
or (n9414,n9415,n9418);
and (n9415,n9416,n9417);
xor (n9416,n9302,n9303);
and (n9417,n33,n29);
and (n9418,n9419,n9420);
xor (n9419,n9416,n9417);
or (n9420,n9421,n9424);
and (n9421,n9422,n9423);
xor (n9422,n9308,n9309);
and (n9423,n64,n29);
and (n9424,n9425,n9426);
xor (n9425,n9422,n9423);
or (n9426,n9427,n9430);
and (n9427,n9428,n9429);
xor (n9428,n9314,n9315);
and (n9429,n58,n29);
and (n9430,n9431,n9432);
xor (n9431,n9428,n9429);
or (n9432,n9433,n9436);
and (n9433,n9434,n9435);
xor (n9434,n9320,n9321);
and (n9435,n117,n29);
and (n9436,n9437,n9438);
xor (n9437,n9434,n9435);
or (n9438,n9439,n9442);
and (n9439,n9440,n9441);
xor (n9440,n9326,n9327);
and (n9441,n111,n29);
and (n9442,n9443,n9444);
xor (n9443,n9440,n9441);
or (n9444,n9445,n9448);
and (n9445,n9446,n9447);
xor (n9446,n9332,n9333);
and (n9447,n141,n29);
and (n9448,n9449,n9450);
xor (n9449,n9446,n9447);
or (n9450,n9451,n9454);
and (n9451,n9452,n9453);
xor (n9452,n9338,n9339);
and (n9453,n135,n29);
and (n9454,n9455,n9456);
xor (n9455,n9452,n9453);
or (n9456,n9457,n9460);
and (n9457,n9458,n9459);
xor (n9458,n9344,n9345);
and (n9459,n448,n29);
and (n9460,n9461,n9462);
xor (n9461,n9458,n9459);
or (n9462,n9463,n9466);
and (n9463,n9464,n9465);
xor (n9464,n9350,n9351);
and (n9465,n474,n29);
and (n9466,n9467,n9468);
xor (n9467,n9464,n9465);
or (n9468,n9469,n9472);
and (n9469,n9470,n9471);
xor (n9470,n9356,n9357);
and (n9471,n625,n29);
and (n9472,n9473,n9474);
xor (n9473,n9470,n9471);
or (n9474,n9475,n9478);
and (n9475,n9476,n9477);
xor (n9476,n9362,n9363);
and (n9477,n1037,n29);
and (n9478,n9479,n9480);
xor (n9479,n9476,n9477);
or (n9480,n9481,n9484);
and (n9481,n9482,n9483);
xor (n9482,n9368,n9369);
and (n9483,n1030,n29);
and (n9484,n9485,n9486);
xor (n9485,n9482,n9483);
or (n9486,n9487,n9490);
and (n9487,n9488,n9489);
xor (n9488,n9374,n9375);
and (n9489,n1002,n29);
and (n9490,n9491,n9492);
xor (n9491,n9488,n9489);
or (n9492,n9493,n9496);
and (n9493,n9494,n9495);
xor (n9494,n9380,n9381);
and (n9495,n832,n29);
and (n9496,n9497,n9498);
xor (n9497,n9494,n9495);
or (n9498,n9499,n9501);
and (n9499,n9500,n922);
xor (n9500,n9386,n9387);
and (n9501,n9502,n9503);
xor (n9502,n9500,n922);
or (n9503,n9504,n9507);
and (n9504,n9505,n9506);
xor (n9505,n9392,n9393);
and (n9506,n847,n29);
and (n9507,n9508,n9509);
xor (n9508,n9505,n9506);
or (n9509,n9510,n9513);
and (n9510,n9511,n9512);
xor (n9511,n9398,n9399);
and (n9512,n839,n29);
and (n9513,n9514,n9515);
xor (n9514,n9511,n9512);
and (n9515,n9516,n9517);
xor (n9516,n9404,n9405);
and (n9517,n887,n29);
and (n9518,n39,n49);
or (n9519,n9520,n9523);
and (n9520,n9521,n9522);
xor (n9521,n9413,n9414);
and (n9522,n33,n49);
and (n9523,n9524,n9525);
xor (n9524,n9521,n9522);
or (n9525,n9526,n9529);
and (n9526,n9527,n9528);
xor (n9527,n9419,n9420);
and (n9528,n64,n49);
and (n9529,n9530,n9531);
xor (n9530,n9527,n9528);
or (n9531,n9532,n9535);
and (n9532,n9533,n9534);
xor (n9533,n9425,n9426);
and (n9534,n58,n49);
and (n9535,n9536,n9537);
xor (n9536,n9533,n9534);
or (n9537,n9538,n9541);
and (n9538,n9539,n9540);
xor (n9539,n9431,n9432);
and (n9540,n117,n49);
and (n9541,n9542,n9543);
xor (n9542,n9539,n9540);
or (n9543,n9544,n9547);
and (n9544,n9545,n9546);
xor (n9545,n9437,n9438);
and (n9546,n111,n49);
and (n9547,n9548,n9549);
xor (n9548,n9545,n9546);
or (n9549,n9550,n9553);
and (n9550,n9551,n9552);
xor (n9551,n9443,n9444);
and (n9552,n141,n49);
and (n9553,n9554,n9555);
xor (n9554,n9551,n9552);
or (n9555,n9556,n9559);
and (n9556,n9557,n9558);
xor (n9557,n9449,n9450);
and (n9558,n135,n49);
and (n9559,n9560,n9561);
xor (n9560,n9557,n9558);
or (n9561,n9562,n9565);
and (n9562,n9563,n9564);
xor (n9563,n9455,n9456);
and (n9564,n448,n49);
and (n9565,n9566,n9567);
xor (n9566,n9563,n9564);
or (n9567,n9568,n9571);
and (n9568,n9569,n9570);
xor (n9569,n9461,n9462);
and (n9570,n474,n49);
and (n9571,n9572,n9573);
xor (n9572,n9569,n9570);
or (n9573,n9574,n9577);
and (n9574,n9575,n9576);
xor (n9575,n9467,n9468);
and (n9576,n625,n49);
and (n9577,n9578,n9579);
xor (n9578,n9575,n9576);
or (n9579,n9580,n9583);
and (n9580,n9581,n9582);
xor (n9581,n9473,n9474);
and (n9582,n1037,n49);
and (n9583,n9584,n9585);
xor (n9584,n9581,n9582);
or (n9585,n9586,n9589);
and (n9586,n9587,n9588);
xor (n9587,n9479,n9480);
and (n9588,n1030,n49);
and (n9589,n9590,n9591);
xor (n9590,n9587,n9588);
or (n9591,n9592,n9595);
and (n9592,n9593,n9594);
xor (n9593,n9485,n9486);
and (n9594,n1002,n49);
and (n9595,n9596,n9597);
xor (n9596,n9593,n9594);
or (n9597,n9598,n9601);
and (n9598,n9599,n9600);
xor (n9599,n9491,n9492);
and (n9600,n832,n49);
and (n9601,n9602,n9603);
xor (n9602,n9599,n9600);
or (n9603,n9604,n9607);
and (n9604,n9605,n9606);
xor (n9605,n9497,n9498);
and (n9606,n826,n49);
and (n9607,n9608,n9609);
xor (n9608,n9605,n9606);
or (n9609,n9610,n9613);
and (n9610,n9611,n9612);
xor (n9611,n9502,n9503);
and (n9612,n847,n49);
and (n9613,n9614,n9615);
xor (n9614,n9611,n9612);
or (n9615,n9616,n9619);
and (n9616,n9617,n9618);
xor (n9617,n9508,n9509);
and (n9618,n839,n49);
and (n9619,n9620,n9621);
xor (n9620,n9617,n9618);
and (n9621,n9622,n1058);
xor (n9622,n9514,n9515);
and (n9623,n33,n54);
or (n9624,n9625,n9628);
and (n9625,n9626,n9627);
xor (n9626,n9524,n9525);
and (n9627,n64,n54);
and (n9628,n9629,n9630);
xor (n9629,n9626,n9627);
or (n9630,n9631,n9634);
and (n9631,n9632,n9633);
xor (n9632,n9530,n9531);
and (n9633,n58,n54);
and (n9634,n9635,n9636);
xor (n9635,n9632,n9633);
or (n9636,n9637,n9640);
and (n9637,n9638,n9639);
xor (n9638,n9536,n9537);
and (n9639,n117,n54);
and (n9640,n9641,n9642);
xor (n9641,n9638,n9639);
or (n9642,n9643,n9646);
and (n9643,n9644,n9645);
xor (n9644,n9542,n9543);
and (n9645,n111,n54);
and (n9646,n9647,n9648);
xor (n9647,n9644,n9645);
or (n9648,n9649,n9652);
and (n9649,n9650,n9651);
xor (n9650,n9548,n9549);
and (n9651,n141,n54);
and (n9652,n9653,n9654);
xor (n9653,n9650,n9651);
or (n9654,n9655,n9658);
and (n9655,n9656,n9657);
xor (n9656,n9554,n9555);
and (n9657,n135,n54);
and (n9658,n9659,n9660);
xor (n9659,n9656,n9657);
or (n9660,n9661,n9664);
and (n9661,n9662,n9663);
xor (n9662,n9560,n9561);
and (n9663,n448,n54);
and (n9664,n9665,n9666);
xor (n9665,n9662,n9663);
or (n9666,n9667,n9670);
and (n9667,n9668,n9669);
xor (n9668,n9566,n9567);
and (n9669,n474,n54);
and (n9670,n9671,n9672);
xor (n9671,n9668,n9669);
or (n9672,n9673,n9676);
and (n9673,n9674,n9675);
xor (n9674,n9572,n9573);
and (n9675,n625,n54);
and (n9676,n9677,n9678);
xor (n9677,n9674,n9675);
or (n9678,n9679,n9682);
and (n9679,n9680,n9681);
xor (n9680,n9578,n9579);
and (n9681,n1037,n54);
and (n9682,n9683,n9684);
xor (n9683,n9680,n9681);
or (n9684,n9685,n9688);
and (n9685,n9686,n9687);
xor (n9686,n9584,n9585);
and (n9687,n1030,n54);
and (n9688,n9689,n9690);
xor (n9689,n9686,n9687);
or (n9690,n9691,n9694);
and (n9691,n9692,n9693);
xor (n9692,n9590,n9591);
and (n9693,n1002,n54);
and (n9694,n9695,n9696);
xor (n9695,n9692,n9693);
or (n9696,n9697,n9700);
and (n9697,n9698,n9699);
xor (n9698,n9596,n9597);
and (n9699,n832,n54);
and (n9700,n9701,n9702);
xor (n9701,n9698,n9699);
or (n9702,n9703,n9706);
and (n9703,n9704,n9705);
xor (n9704,n9602,n9603);
and (n9705,n826,n54);
and (n9706,n9707,n9708);
xor (n9707,n9704,n9705);
or (n9708,n9709,n9712);
and (n9709,n9710,n9711);
xor (n9710,n9608,n9609);
and (n9711,n847,n54);
and (n9712,n9713,n9714);
xor (n9713,n9710,n9711);
or (n9714,n9715,n9718);
and (n9715,n9716,n9717);
xor (n9716,n9614,n9615);
and (n9717,n839,n54);
and (n9718,n9719,n9720);
xor (n9719,n9716,n9717);
and (n9720,n9721,n9722);
xor (n9721,n9620,n9621);
and (n9722,n887,n54);
and (n9723,n64,n102);
or (n9724,n9725,n9728);
and (n9725,n9726,n9727);
xor (n9726,n9629,n9630);
and (n9727,n58,n102);
and (n9728,n9729,n9730);
xor (n9729,n9726,n9727);
or (n9730,n9731,n9734);
and (n9731,n9732,n9733);
xor (n9732,n9635,n9636);
and (n9733,n117,n102);
and (n9734,n9735,n9736);
xor (n9735,n9732,n9733);
or (n9736,n9737,n9740);
and (n9737,n9738,n9739);
xor (n9738,n9641,n9642);
and (n9739,n111,n102);
and (n9740,n9741,n9742);
xor (n9741,n9738,n9739);
or (n9742,n9743,n9746);
and (n9743,n9744,n9745);
xor (n9744,n9647,n9648);
and (n9745,n141,n102);
and (n9746,n9747,n9748);
xor (n9747,n9744,n9745);
or (n9748,n9749,n9752);
and (n9749,n9750,n9751);
xor (n9750,n9653,n9654);
and (n9751,n135,n102);
and (n9752,n9753,n9754);
xor (n9753,n9750,n9751);
or (n9754,n9755,n9758);
and (n9755,n9756,n9757);
xor (n9756,n9659,n9660);
and (n9757,n448,n102);
and (n9758,n9759,n9760);
xor (n9759,n9756,n9757);
or (n9760,n9761,n9764);
and (n9761,n9762,n9763);
xor (n9762,n9665,n9666);
and (n9763,n474,n102);
and (n9764,n9765,n9766);
xor (n9765,n9762,n9763);
or (n9766,n9767,n9770);
and (n9767,n9768,n9769);
xor (n9768,n9671,n9672);
and (n9769,n625,n102);
and (n9770,n9771,n9772);
xor (n9771,n9768,n9769);
or (n9772,n9773,n9776);
and (n9773,n9774,n9775);
xor (n9774,n9677,n9678);
and (n9775,n1037,n102);
and (n9776,n9777,n9778);
xor (n9777,n9774,n9775);
or (n9778,n9779,n9782);
and (n9779,n9780,n9781);
xor (n9780,n9683,n9684);
and (n9781,n1030,n102);
and (n9782,n9783,n9784);
xor (n9783,n9780,n9781);
or (n9784,n9785,n9788);
and (n9785,n9786,n9787);
xor (n9786,n9689,n9690);
and (n9787,n1002,n102);
and (n9788,n9789,n9790);
xor (n9789,n9786,n9787);
or (n9790,n9791,n9794);
and (n9791,n9792,n9793);
xor (n9792,n9695,n9696);
and (n9793,n832,n102);
and (n9794,n9795,n9796);
xor (n9795,n9792,n9793);
or (n9796,n9797,n9800);
and (n9797,n9798,n9799);
xor (n9798,n9701,n9702);
and (n9799,n826,n102);
and (n9800,n9801,n9802);
xor (n9801,n9798,n9799);
or (n9802,n9803,n9806);
and (n9803,n9804,n9805);
xor (n9804,n9707,n9708);
and (n9805,n847,n102);
and (n9806,n9807,n9808);
xor (n9807,n9804,n9805);
or (n9808,n9809,n9812);
and (n9809,n9810,n9811);
xor (n9810,n9713,n9714);
and (n9811,n839,n102);
and (n9812,n9813,n9814);
xor (n9813,n9810,n9811);
and (n9814,n9815,n2164);
xor (n9815,n9719,n9720);
and (n9816,n58,n107);
or (n9817,n9818,n9821);
and (n9818,n9819,n9820);
xor (n9819,n9729,n9730);
and (n9820,n117,n107);
and (n9821,n9822,n9823);
xor (n9822,n9819,n9820);
or (n9823,n9824,n9827);
and (n9824,n9825,n9826);
xor (n9825,n9735,n9736);
and (n9826,n111,n107);
and (n9827,n9828,n9829);
xor (n9828,n9825,n9826);
or (n9829,n9830,n9833);
and (n9830,n9831,n9832);
xor (n9831,n9741,n9742);
and (n9832,n141,n107);
and (n9833,n9834,n9835);
xor (n9834,n9831,n9832);
or (n9835,n9836,n9839);
and (n9836,n9837,n9838);
xor (n9837,n9747,n9748);
and (n9838,n135,n107);
and (n9839,n9840,n9841);
xor (n9840,n9837,n9838);
or (n9841,n9842,n9845);
and (n9842,n9843,n9844);
xor (n9843,n9753,n9754);
and (n9844,n448,n107);
and (n9845,n9846,n9847);
xor (n9846,n9843,n9844);
or (n9847,n9848,n9851);
and (n9848,n9849,n9850);
xor (n9849,n9759,n9760);
and (n9850,n474,n107);
and (n9851,n9852,n9853);
xor (n9852,n9849,n9850);
or (n9853,n9854,n9857);
and (n9854,n9855,n9856);
xor (n9855,n9765,n9766);
and (n9856,n625,n107);
and (n9857,n9858,n9859);
xor (n9858,n9855,n9856);
or (n9859,n9860,n9863);
and (n9860,n9861,n9862);
xor (n9861,n9771,n9772);
and (n9862,n1037,n107);
and (n9863,n9864,n9865);
xor (n9864,n9861,n9862);
or (n9865,n9866,n9869);
and (n9866,n9867,n9868);
xor (n9867,n9777,n9778);
and (n9868,n1030,n107);
and (n9869,n9870,n9871);
xor (n9870,n9867,n9868);
or (n9871,n9872,n9875);
and (n9872,n9873,n9874);
xor (n9873,n9783,n9784);
and (n9874,n1002,n107);
and (n9875,n9876,n9877);
xor (n9876,n9873,n9874);
or (n9877,n9878,n9881);
and (n9878,n9879,n9880);
xor (n9879,n9789,n9790);
and (n9880,n832,n107);
and (n9881,n9882,n9883);
xor (n9882,n9879,n9880);
or (n9883,n9884,n9887);
and (n9884,n9885,n9886);
xor (n9885,n9795,n9796);
and (n9886,n826,n107);
and (n9887,n9888,n9889);
xor (n9888,n9885,n9886);
or (n9889,n9890,n9893);
and (n9890,n9891,n9892);
xor (n9891,n9801,n9802);
and (n9892,n847,n107);
and (n9893,n9894,n9895);
xor (n9894,n9891,n9892);
or (n9895,n9896,n9899);
and (n9896,n9897,n9898);
xor (n9897,n9807,n9808);
and (n9898,n839,n107);
and (n9899,n9900,n9901);
xor (n9900,n9897,n9898);
and (n9901,n9902,n9903);
xor (n9902,n9813,n9814);
and (n9903,n887,n107);
and (n9904,n117,n125);
or (n9905,n9906,n9909);
and (n9906,n9907,n9908);
xor (n9907,n9822,n9823);
and (n9908,n111,n125);
and (n9909,n9910,n9911);
xor (n9910,n9907,n9908);
or (n9911,n9912,n9915);
and (n9912,n9913,n9914);
xor (n9913,n9828,n9829);
and (n9914,n141,n125);
and (n9915,n9916,n9917);
xor (n9916,n9913,n9914);
or (n9917,n9918,n9921);
and (n9918,n9919,n9920);
xor (n9919,n9834,n9835);
and (n9920,n135,n125);
and (n9921,n9922,n9923);
xor (n9922,n9919,n9920);
or (n9923,n9924,n9927);
and (n9924,n9925,n9926);
xor (n9925,n9840,n9841);
and (n9926,n448,n125);
and (n9927,n9928,n9929);
xor (n9928,n9925,n9926);
or (n9929,n9930,n9933);
and (n9930,n9931,n9932);
xor (n9931,n9846,n9847);
and (n9932,n474,n125);
and (n9933,n9934,n9935);
xor (n9934,n9931,n9932);
or (n9935,n9936,n9939);
and (n9936,n9937,n9938);
xor (n9937,n9852,n9853);
and (n9938,n625,n125);
and (n9939,n9940,n9941);
xor (n9940,n9937,n9938);
or (n9941,n9942,n9945);
and (n9942,n9943,n9944);
xor (n9943,n9858,n9859);
and (n9944,n1037,n125);
and (n9945,n9946,n9947);
xor (n9946,n9943,n9944);
or (n9947,n9948,n9951);
and (n9948,n9949,n9950);
xor (n9949,n9864,n9865);
and (n9950,n1030,n125);
and (n9951,n9952,n9953);
xor (n9952,n9949,n9950);
or (n9953,n9954,n9957);
and (n9954,n9955,n9956);
xor (n9955,n9870,n9871);
and (n9956,n1002,n125);
and (n9957,n9958,n9959);
xor (n9958,n9955,n9956);
or (n9959,n9960,n9963);
and (n9960,n9961,n9962);
xor (n9961,n9876,n9877);
and (n9962,n832,n125);
and (n9963,n9964,n9965);
xor (n9964,n9961,n9962);
or (n9965,n9966,n9969);
and (n9966,n9967,n9968);
xor (n9967,n9882,n9883);
and (n9968,n826,n125);
and (n9969,n9970,n9971);
xor (n9970,n9967,n9968);
or (n9971,n9972,n9975);
and (n9972,n9973,n9974);
xor (n9973,n9888,n9889);
and (n9974,n847,n125);
and (n9975,n9976,n9977);
xor (n9976,n9973,n9974);
or (n9977,n9978,n9981);
and (n9978,n9979,n9980);
xor (n9979,n9894,n9895);
and (n9980,n839,n125);
and (n9981,n9982,n9983);
xor (n9982,n9979,n9980);
and (n9983,n9984,n2514);
xor (n9984,n9900,n9901);
and (n9985,n111,n131);
or (n9986,n9987,n9990);
and (n9987,n9988,n9989);
xor (n9988,n9910,n9911);
and (n9989,n141,n131);
and (n9990,n9991,n9992);
xor (n9991,n9988,n9989);
or (n9992,n9993,n9996);
and (n9993,n9994,n9995);
xor (n9994,n9916,n9917);
and (n9995,n135,n131);
and (n9996,n9997,n9998);
xor (n9997,n9994,n9995);
or (n9998,n9999,n10002);
and (n9999,n10000,n10001);
xor (n10000,n9922,n9923);
and (n10001,n448,n131);
and (n10002,n10003,n10004);
xor (n10003,n10000,n10001);
or (n10004,n10005,n10008);
and (n10005,n10006,n10007);
xor (n10006,n9928,n9929);
and (n10007,n474,n131);
and (n10008,n10009,n10010);
xor (n10009,n10006,n10007);
or (n10010,n10011,n10014);
and (n10011,n10012,n10013);
xor (n10012,n9934,n9935);
and (n10013,n625,n131);
and (n10014,n10015,n10016);
xor (n10015,n10012,n10013);
or (n10016,n10017,n10020);
and (n10017,n10018,n10019);
xor (n10018,n9940,n9941);
and (n10019,n1037,n131);
and (n10020,n10021,n10022);
xor (n10021,n10018,n10019);
or (n10022,n10023,n10026);
and (n10023,n10024,n10025);
xor (n10024,n9946,n9947);
and (n10025,n1030,n131);
and (n10026,n10027,n10028);
xor (n10027,n10024,n10025);
or (n10028,n10029,n10032);
and (n10029,n10030,n10031);
xor (n10030,n9952,n9953);
and (n10031,n1002,n131);
and (n10032,n10033,n10034);
xor (n10033,n10030,n10031);
or (n10034,n10035,n10038);
and (n10035,n10036,n10037);
xor (n10036,n9958,n9959);
and (n10037,n832,n131);
and (n10038,n10039,n10040);
xor (n10039,n10036,n10037);
or (n10040,n10041,n10044);
and (n10041,n10042,n10043);
xor (n10042,n9964,n9965);
and (n10043,n826,n131);
and (n10044,n10045,n10046);
xor (n10045,n10042,n10043);
or (n10046,n10047,n10050);
and (n10047,n10048,n10049);
xor (n10048,n9970,n9971);
and (n10049,n847,n131);
and (n10050,n10051,n10052);
xor (n10051,n10048,n10049);
or (n10052,n10053,n10056);
and (n10053,n10054,n10055);
xor (n10054,n9976,n9977);
and (n10055,n839,n131);
and (n10056,n10057,n10058);
xor (n10057,n10054,n10055);
and (n10058,n10059,n10060);
xor (n10059,n9982,n9983);
and (n10060,n887,n131);
or (n10061,n10062,n10064);
and (n10062,n10063,n9995);
xor (n10063,n9991,n9992);
and (n10064,n10065,n10066);
xor (n10065,n10063,n9995);
or (n10066,n10067,n10069);
and (n10067,n10068,n10001);
xor (n10068,n9997,n9998);
and (n10069,n10070,n10071);
xor (n10070,n10068,n10001);
or (n10071,n10072,n10074);
and (n10072,n10073,n10007);
xor (n10073,n10003,n10004);
and (n10074,n10075,n10076);
xor (n10075,n10073,n10007);
or (n10076,n10077,n10079);
and (n10077,n10078,n10013);
xor (n10078,n10009,n10010);
and (n10079,n10080,n10081);
xor (n10080,n10078,n10013);
or (n10081,n10082,n10084);
and (n10082,n10083,n10019);
xor (n10083,n10015,n10016);
and (n10084,n10085,n10086);
xor (n10085,n10083,n10019);
or (n10086,n10087,n10089);
and (n10087,n10088,n10025);
xor (n10088,n10021,n10022);
and (n10089,n10090,n10091);
xor (n10090,n10088,n10025);
or (n10091,n10092,n10094);
and (n10092,n10093,n10031);
xor (n10093,n10027,n10028);
and (n10094,n10095,n10096);
xor (n10095,n10093,n10031);
or (n10096,n10097,n10099);
and (n10097,n10098,n10037);
xor (n10098,n10033,n10034);
and (n10099,n10100,n10101);
xor (n10100,n10098,n10037);
or (n10101,n10102,n10104);
and (n10102,n10103,n10043);
xor (n10103,n10039,n10040);
and (n10104,n10105,n10106);
xor (n10105,n10103,n10043);
or (n10106,n10107,n10109);
and (n10107,n10108,n10049);
xor (n10108,n10045,n10046);
and (n10109,n10110,n10111);
xor (n10110,n10108,n10049);
or (n10111,n10112,n10114);
and (n10112,n10113,n10055);
xor (n10113,n10051,n10052);
and (n10114,n10115,n10116);
xor (n10115,n10113,n10055);
and (n10116,n10117,n10060);
xor (n10117,n10057,n10058);
or (n10118,n10119,n10121);
and (n10119,n10120,n10001);
xor (n10120,n10065,n10066);
and (n10121,n10122,n10123);
xor (n10122,n10120,n10001);
or (n10123,n10124,n10126);
and (n10124,n10125,n10007);
xor (n10125,n10070,n10071);
and (n10126,n10127,n10128);
xor (n10127,n10125,n10007);
or (n10128,n10129,n10131);
and (n10129,n10130,n10013);
xor (n10130,n10075,n10076);
and (n10131,n10132,n10133);
xor (n10132,n10130,n10013);
or (n10133,n10134,n10136);
and (n10134,n10135,n10019);
xor (n10135,n10080,n10081);
and (n10136,n10137,n10138);
xor (n10137,n10135,n10019);
or (n10138,n10139,n10141);
and (n10139,n10140,n10025);
xor (n10140,n10085,n10086);
and (n10141,n10142,n10143);
xor (n10142,n10140,n10025);
or (n10143,n10144,n10146);
and (n10144,n10145,n10031);
xor (n10145,n10090,n10091);
and (n10146,n10147,n10148);
xor (n10147,n10145,n10031);
or (n10148,n10149,n10151);
and (n10149,n10150,n10037);
xor (n10150,n10095,n10096);
and (n10151,n10152,n10153);
xor (n10152,n10150,n10037);
or (n10153,n10154,n10156);
and (n10154,n10155,n10043);
xor (n10155,n10100,n10101);
and (n10156,n10157,n10158);
xor (n10157,n10155,n10043);
or (n10158,n10159,n10161);
and (n10159,n10160,n10049);
xor (n10160,n10105,n10106);
and (n10161,n10162,n10163);
xor (n10162,n10160,n10049);
or (n10163,n10164,n10166);
and (n10164,n10165,n10055);
xor (n10165,n10110,n10111);
and (n10166,n10167,n10168);
xor (n10167,n10165,n10055);
and (n10168,n10169,n10060);
xor (n10169,n10115,n10116);
or (n10170,n10171,n10173);
and (n10171,n10172,n10007);
xor (n10172,n10122,n10123);
and (n10173,n10174,n10175);
xor (n10174,n10172,n10007);
or (n10175,n10176,n10178);
and (n10176,n10177,n10013);
xor (n10177,n10127,n10128);
and (n10178,n10179,n10180);
xor (n10179,n10177,n10013);
or (n10180,n10181,n10183);
and (n10181,n10182,n10019);
xor (n10182,n10132,n10133);
and (n10183,n10184,n10185);
xor (n10184,n10182,n10019);
or (n10185,n10186,n10188);
and (n10186,n10187,n10025);
xor (n10187,n10137,n10138);
and (n10188,n10189,n10190);
xor (n10189,n10187,n10025);
or (n10190,n10191,n10193);
and (n10191,n10192,n10031);
xor (n10192,n10142,n10143);
and (n10193,n10194,n10195);
xor (n10194,n10192,n10031);
or (n10195,n10196,n10198);
and (n10196,n10197,n10037);
xor (n10197,n10147,n10148);
and (n10198,n10199,n10200);
xor (n10199,n10197,n10037);
or (n10200,n10201,n10203);
and (n10201,n10202,n10043);
xor (n10202,n10152,n10153);
and (n10203,n10204,n10205);
xor (n10204,n10202,n10043);
or (n10205,n10206,n10208);
and (n10206,n10207,n10049);
xor (n10207,n10157,n10158);
and (n10208,n10209,n10210);
xor (n10209,n10207,n10049);
or (n10210,n10211,n10213);
and (n10211,n10212,n10055);
xor (n10212,n10162,n10163);
and (n10213,n10214,n10215);
xor (n10214,n10212,n10055);
and (n10215,n10216,n10060);
xor (n10216,n10167,n10168);
or (n10217,n10218,n10220);
and (n10218,n10219,n10013);
xor (n10219,n10174,n10175);
and (n10220,n10221,n10222);
xor (n10221,n10219,n10013);
or (n10222,n10223,n10225);
and (n10223,n10224,n10019);
xor (n10224,n10179,n10180);
and (n10225,n10226,n10227);
xor (n10226,n10224,n10019);
or (n10227,n10228,n10230);
and (n10228,n10229,n10025);
xor (n10229,n10184,n10185);
and (n10230,n10231,n10232);
xor (n10231,n10229,n10025);
or (n10232,n10233,n10235);
and (n10233,n10234,n10031);
xor (n10234,n10189,n10190);
and (n10235,n10236,n10237);
xor (n10236,n10234,n10031);
or (n10237,n10238,n10240);
and (n10238,n10239,n10037);
xor (n10239,n10194,n10195);
and (n10240,n10241,n10242);
xor (n10241,n10239,n10037);
or (n10242,n10243,n10245);
and (n10243,n10244,n10043);
xor (n10244,n10199,n10200);
and (n10245,n10246,n10247);
xor (n10246,n10244,n10043);
or (n10247,n10248,n10250);
and (n10248,n10249,n10049);
xor (n10249,n10204,n10205);
and (n10250,n10251,n10252);
xor (n10251,n10249,n10049);
or (n10252,n10253,n10255);
and (n10253,n10254,n10055);
xor (n10254,n10209,n10210);
and (n10255,n10256,n10257);
xor (n10256,n10254,n10055);
and (n10257,n10258,n10060);
xor (n10258,n10214,n10215);
or (n10259,n10260,n10262);
and (n10260,n10261,n10019);
xor (n10261,n10221,n10222);
and (n10262,n10263,n10264);
xor (n10263,n10261,n10019);
or (n10264,n10265,n10267);
and (n10265,n10266,n10025);
xor (n10266,n10226,n10227);
and (n10267,n10268,n10269);
xor (n10268,n10266,n10025);
or (n10269,n10270,n10272);
and (n10270,n10271,n10031);
xor (n10271,n10231,n10232);
and (n10272,n10273,n10274);
xor (n10273,n10271,n10031);
or (n10274,n10275,n10277);
and (n10275,n10276,n10037);
xor (n10276,n10236,n10237);
and (n10277,n10278,n10279);
xor (n10278,n10276,n10037);
or (n10279,n10280,n10282);
and (n10280,n10281,n10043);
xor (n10281,n10241,n10242);
and (n10282,n10283,n10284);
xor (n10283,n10281,n10043);
or (n10284,n10285,n10287);
and (n10285,n10286,n10049);
xor (n10286,n10246,n10247);
and (n10287,n10288,n10289);
xor (n10288,n10286,n10049);
or (n10289,n10290,n10292);
and (n10290,n10291,n10055);
xor (n10291,n10251,n10252);
and (n10292,n10293,n10294);
xor (n10293,n10291,n10055);
and (n10294,n10295,n10060);
xor (n10295,n10256,n10257);
or (n10296,n10297,n10299);
and (n10297,n10298,n10025);
xor (n10298,n10263,n10264);
and (n10299,n10300,n10301);
xor (n10300,n10298,n10025);
or (n10301,n10302,n10304);
and (n10302,n10303,n10031);
xor (n10303,n10268,n10269);
and (n10304,n10305,n10306);
xor (n10305,n10303,n10031);
or (n10306,n10307,n10309);
and (n10307,n10308,n10037);
xor (n10308,n10273,n10274);
and (n10309,n10310,n10311);
xor (n10310,n10308,n10037);
or (n10311,n10312,n10314);
and (n10312,n10313,n10043);
xor (n10313,n10278,n10279);
and (n10314,n10315,n10316);
xor (n10315,n10313,n10043);
or (n10316,n10317,n10319);
and (n10317,n10318,n10049);
xor (n10318,n10283,n10284);
and (n10319,n10320,n10321);
xor (n10320,n10318,n10049);
or (n10321,n10322,n10324);
and (n10322,n10323,n10055);
xor (n10323,n10288,n10289);
and (n10324,n10325,n10326);
xor (n10325,n10323,n10055);
and (n10326,n10327,n10060);
xor (n10327,n10293,n10294);
or (n10328,n10329,n10331);
and (n10329,n10330,n10031);
xor (n10330,n10300,n10301);
and (n10331,n10332,n10333);
xor (n10332,n10330,n10031);
or (n10333,n10334,n10336);
and (n10334,n10335,n10037);
xor (n10335,n10305,n10306);
and (n10336,n10337,n10338);
xor (n10337,n10335,n10037);
or (n10338,n10339,n10341);
and (n10339,n10340,n10043);
xor (n10340,n10310,n10311);
and (n10341,n10342,n10343);
xor (n10342,n10340,n10043);
or (n10343,n10344,n10346);
and (n10344,n10345,n10049);
xor (n10345,n10315,n10316);
and (n10346,n10347,n10348);
xor (n10347,n10345,n10049);
or (n10348,n10349,n10351);
and (n10349,n10350,n10055);
xor (n10350,n10320,n10321);
and (n10351,n10352,n10353);
xor (n10352,n10350,n10055);
and (n10353,n10354,n10060);
xor (n10354,n10325,n10326);
or (n10355,n10356,n10358);
and (n10356,n10357,n10037);
xor (n10357,n10332,n10333);
and (n10358,n10359,n10360);
xor (n10359,n10357,n10037);
or (n10360,n10361,n10363);
and (n10361,n10362,n10043);
xor (n10362,n10337,n10338);
and (n10363,n10364,n10365);
xor (n10364,n10362,n10043);
or (n10365,n10366,n10368);
and (n10366,n10367,n10049);
xor (n10367,n10342,n10343);
and (n10368,n10369,n10370);
xor (n10369,n10367,n10049);
or (n10370,n10371,n10373);
and (n10371,n10372,n10055);
xor (n10372,n10347,n10348);
and (n10373,n10374,n10375);
xor (n10374,n10372,n10055);
and (n10375,n10376,n10060);
xor (n10376,n10352,n10353);
or (n10377,n10378,n10380);
and (n10378,n10379,n10043);
xor (n10379,n10359,n10360);
and (n10380,n10381,n10382);
xor (n10381,n10379,n10043);
or (n10382,n10383,n10385);
and (n10383,n10384,n10049);
xor (n10384,n10364,n10365);
and (n10385,n10386,n10387);
xor (n10386,n10384,n10049);
or (n10387,n10388,n10390);
and (n10388,n10389,n10055);
xor (n10389,n10369,n10370);
and (n10390,n10391,n10392);
xor (n10391,n10389,n10055);
and (n10392,n10393,n10060);
xor (n10393,n10374,n10375);
or (n10394,n10395,n10397);
and (n10395,n10396,n10049);
xor (n10396,n10381,n10382);
and (n10397,n10398,n10399);
xor (n10398,n10396,n10049);
or (n10399,n10400,n10402);
and (n10400,n10401,n10055);
xor (n10401,n10386,n10387);
and (n10402,n10403,n10404);
xor (n10403,n10401,n10055);
and (n10404,n10405,n10060);
xor (n10405,n10391,n10392);
or (n10406,n10407,n10409);
and (n10407,n10408,n10055);
xor (n10408,n10398,n10399);
and (n10409,n10410,n10411);
xor (n10410,n10408,n10055);
and (n10411,n10412,n10060);
xor (n10412,n10403,n10404);
and (n10413,n10414,n10060);
xor (n10414,n10410,n10411);
endmodule
