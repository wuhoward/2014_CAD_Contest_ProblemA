module top (out,n3,n4,n5,n23,n24,n29,n33,n40,n49
        ,n50,n56,n60,n66,n84,n91,n92,n102,n122,n124
        ,n130,n140,n158,n167,n177,n181,n188,n213);
output out;
input n3;
input n4;
input n5;
input n23;
input n24;
input n29;
input n33;
input n40;
input n49;
input n50;
input n56;
input n60;
input n66;
input n84;
input n91;
input n92;
input n102;
input n122;
input n124;
input n130;
input n140;
input n158;
input n167;
input n177;
input n181;
input n188;
input n213;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
xnor (out,n0,n550);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n547);
nand (n7,n8,n546);
or (n8,n9,n296);
not (n9,n10);
nand (n10,n11,n295);
nand (n11,n12,n260);
not (n12,n13);
xor (n13,n14,n216);
xor (n14,n15,n105);
xor (n15,n16,n69);
xor (n16,n17,n43);
nand (n17,n18,n37);
or (n18,n19,n31);
nand (n19,n20,n27);
nor (n20,n21,n25);
and (n21,n22,n24);
not (n22,n23);
and (n25,n23,n26);
not (n26,n24);
nand (n27,n28,n30);
or (n28,n26,n29);
nand (n30,n26,n29);
nor (n31,n32,n35);
and (n32,n33,n34);
not (n34,n29);
and (n35,n36,n29);
not (n36,n33);
or (n37,n20,n38);
nor (n38,n39,n41);
and (n39,n34,n40);
and (n41,n29,n42);
not (n42,n40);
nand (n43,n44,n63);
or (n44,n45,n58);
nand (n45,n46,n53);
nor (n46,n47,n51);
and (n47,n48,n50);
not (n48,n49);
and (n51,n49,n52);
not (n52,n50);
nand (n53,n54,n57);
or (n54,n50,n55);
not (n55,n56);
nand (n57,n55,n50);
nor (n58,n59,n61);
and (n59,n55,n60);
and (n61,n56,n62);
not (n62,n60);
or (n63,n46,n64);
nor (n64,n65,n67);
and (n65,n55,n66);
and (n67,n56,n68);
not (n68,n66);
nand (n69,n70,n104);
or (n70,n71,n77);
not (n71,n72);
nand (n72,n73,n29);
nand (n73,n74,n75);
or (n74,n23,n24);
nand (n75,n76,n36);
or (n76,n26,n22);
not (n77,n78);
nand (n78,n79,n98);
or (n79,n80,n86);
not (n80,n81);
nand (n81,n82,n85);
or (n82,n49,n83);
not (n83,n84);
or (n85,n48,n84);
not (n86,n87);
nor (n87,n88,n94);
nand (n88,n89,n93);
or (n89,n90,n92);
not (n90,n91);
nand (n93,n90,n92);
nor (n94,n95,n96);
and (n95,n48,n92);
and (n96,n49,n97);
not (n97,n92);
nand (n98,n88,n99);
nand (n99,n100,n103);
or (n100,n49,n101);
not (n101,n102);
or (n103,n48,n102);
or (n104,n78,n72);
xor (n105,n106,n193);
xor (n106,n107,n144);
or (n107,n108,n143);
and (n108,n109,n117);
xor (n109,n110,n111);
nor (n110,n20,n36);
nand (n111,n112,n116);
or (n112,n113,n86);
nor (n113,n114,n115);
and (n114,n68,n49);
and (n115,n66,n48);
nand (n116,n81,n88);
nand (n117,n118,n136);
or (n118,n119,n127);
not (n119,n120);
nand (n120,n121,n125);
or (n121,n122,n123);
not (n123,n124);
or (n125,n126,n124);
not (n126,n122);
nand (n127,n128,n132);
nand (n128,n129,n131);
or (n129,n130,n126);
nand (n131,n126,n130);
not (n132,n133);
nand (n133,n134,n135);
or (n134,n55,n130);
nand (n135,n55,n130);
nand (n136,n137,n133);
not (n137,n138);
nor (n138,n139,n141);
and (n139,n126,n140);
and (n141,n122,n142);
not (n142,n140);
and (n143,n110,n111);
or (n144,n145,n192);
and (n145,n146,n184);
xor (n146,n147,n170);
nand (n147,n148,n163);
or (n148,n149,n153);
not (n149,n150);
nand (n150,n151,n152);
or (n151,n23,n42);
or (n152,n22,n40);
not (n153,n154);
and (n154,n155,n160);
not (n155,n156);
nand (n156,n157,n159);
or (n157,n158,n126);
nand (n159,n158,n126);
nand (n160,n161,n162);
or (n161,n158,n22);
nand (n162,n22,n158);
nand (n163,n164,n156);
not (n164,n165);
nor (n165,n166,n168);
and (n166,n22,n167);
and (n168,n23,n169);
not (n169,n167);
nand (n170,n171,n178);
or (n171,n172,n175);
nor (n172,n173,n174);
and (n173,n90,n102);
and (n174,n91,n101);
nand (n175,n91,n176);
not (n176,n177);
or (n178,n179,n176);
nor (n179,n180,n182);
and (n180,n90,n181);
and (n182,n91,n183);
not (n183,n181);
nand (n184,n185,n191);
or (n185,n45,n186);
nor (n186,n187,n189);
and (n187,n55,n188);
and (n189,n56,n190);
not (n190,n188);
or (n191,n46,n58);
and (n192,n147,n170);
xor (n193,n194,n208);
xor (n194,n195,n201);
nand (n195,n196,n197);
or (n196,n127,n138);
or (n197,n132,n198);
nor (n198,n199,n200);
and (n199,n126,n188);
and (n200,n122,n190);
nand (n201,n202,n203);
or (n202,n153,n165);
or (n203,n155,n204);
not (n204,n205);
nor (n205,n206,n207);
and (n206,n123,n22);
and (n207,n23,n124);
nand (n208,n209,n210);
or (n209,n179,n175);
or (n210,n211,n176);
nor (n211,n212,n214);
and (n212,n90,n213);
and (n214,n91,n215);
not (n215,n213);
or (n216,n217,n259);
and (n217,n218,n258);
xor (n218,n219,n234);
and (n219,n220,n226);
and (n220,n221,n23);
nand (n221,n222,n223);
or (n222,n122,n158);
nand (n223,n224,n36);
or (n224,n225,n126);
not (n225,n158);
nand (n226,n227,n232);
or (n227,n228,n86);
not (n228,n229);
nand (n229,n230,n231);
or (n230,n49,n62);
or (n231,n48,n60);
or (n232,n233,n113);
not (n233,n88);
or (n234,n235,n257);
and (n235,n236,n250);
xor (n236,n237,n243);
nand (n237,n238,n239);
or (n238,n132,n119);
or (n239,n240,n127);
nor (n240,n241,n242);
and (n241,n169,n122);
and (n242,n167,n126);
nand (n243,n244,n249);
or (n244,n245,n153);
not (n245,n246);
nand (n246,n247,n248);
or (n247,n23,n36);
or (n248,n22,n33);
nand (n249,n150,n156);
nand (n250,n251,n256);
or (n251,n252,n175);
not (n252,n253);
nor (n253,n254,n255);
and (n254,n83,n90);
and (n255,n91,n84);
or (n256,n172,n176);
and (n257,n237,n243);
xor (n258,n109,n117);
and (n259,n219,n234);
not (n260,n261);
or (n261,n262,n294);
and (n262,n263,n293);
xor (n263,n264,n265);
xor (n264,n146,n184);
or (n265,n266,n292);
and (n266,n267,n275);
xor (n267,n268,n274);
nand (n268,n269,n273);
or (n269,n45,n270);
nor (n270,n271,n272);
and (n271,n55,n140);
and (n272,n56,n142);
or (n273,n186,n46);
xor (n274,n220,n226);
or (n275,n276,n291);
and (n276,n277,n285);
xor (n277,n278,n279);
and (n278,n156,n33);
nand (n279,n280,n281);
or (n280,n176,n252);
or (n281,n282,n175);
nor (n282,n283,n284);
and (n283,n90,n66);
and (n284,n91,n68);
nand (n285,n286,n290);
or (n286,n127,n287);
nor (n287,n288,n289);
and (n288,n126,n40);
and (n289,n122,n42);
or (n290,n132,n240);
and (n291,n278,n279);
and (n292,n268,n274);
xor (n293,n218,n258);
and (n294,n264,n265);
nand (n295,n13,n261);
not (n296,n297);
nand (n297,n298,n545);
or (n298,n299,n540);
nor (n299,n300,n532);
and (n300,n301,n501);
or (n301,n302,n500);
and (n302,n303,n391);
xor (n303,n304,n355);
or (n304,n305,n354);
and (n305,n306,n333);
xor (n306,n307,n316);
nand (n307,n308,n312);
or (n308,n45,n309);
nor (n309,n310,n311);
and (n310,n55,n40);
and (n311,n56,n42);
or (n312,n46,n313);
nor (n313,n314,n315);
and (n314,n55,n167);
and (n315,n56,n169);
and (n316,n317,n327);
nand (n317,n318,n323);
or (n318,n175,n319);
not (n319,n320);
nor (n320,n321,n322);
and (n321,n91,n140);
and (n322,n142,n90);
nand (n323,n324,n177);
nand (n324,n325,n326);
or (n325,n188,n90);
nand (n326,n90,n188);
not (n327,n328);
nand (n328,n329,n56);
nand (n329,n330,n331);
or (n330,n49,n50);
nand (n331,n332,n36);
or (n332,n52,n48);
xor (n333,n334,n344);
xor (n334,n335,n336);
and (n335,n133,n33);
nand (n336,n337,n342);
or (n337,n176,n338);
not (n338,n339);
nor (n339,n340,n341);
and (n340,n91,n60);
and (n341,n62,n90);
or (n342,n343,n175);
not (n343,n324);
nand (n344,n345,n350);
or (n345,n346,n86);
not (n346,n347);
nor (n347,n348,n349);
and (n348,n49,n124);
and (n349,n123,n48);
nand (n350,n88,n351);
nand (n351,n352,n353);
or (n352,n49,n142);
or (n353,n48,n140);
and (n354,n307,n316);
xor (n355,n356,n370);
xor (n356,n357,n367);
xor (n357,n358,n364);
nor (n358,n359,n126);
nor (n359,n360,n362);
and (n360,n361,n36);
nand (n361,n56,n130);
and (n362,n55,n363);
not (n363,n130);
nand (n364,n365,n366);
or (n365,n175,n338);
or (n366,n282,n176);
or (n367,n368,n369);
and (n368,n334,n344);
and (n369,n335,n336);
xor (n370,n371,n385);
xor (n371,n372,n378);
nand (n372,n373,n377);
or (n373,n127,n374);
nor (n374,n375,n376);
and (n375,n126,n33);
and (n376,n122,n36);
or (n377,n287,n132);
nand (n378,n379,n384);
or (n379,n380,n233);
not (n380,n381);
nand (n381,n382,n383);
or (n382,n49,n190);
or (n383,n48,n188);
nand (n384,n87,n351);
nand (n385,n386,n387);
or (n386,n45,n313);
or (n387,n46,n388);
nor (n388,n389,n390);
and (n389,n124,n55);
and (n390,n56,n123);
or (n391,n392,n499);
and (n392,n393,n417);
xor (n393,n394,n416);
or (n394,n395,n415);
and (n395,n396,n411);
xor (n396,n397,n404);
nand (n397,n398,n403);
or (n398,n399,n86);
not (n399,n400);
nand (n400,n401,n402);
or (n401,n49,n169);
or (n402,n48,n167);
nand (n403,n88,n347);
nand (n404,n405,n410);
or (n405,n406,n45);
not (n406,n407);
nand (n407,n408,n409);
or (n408,n36,n56);
or (n409,n55,n33);
or (n410,n46,n309);
nand (n411,n412,n414);
or (n412,n327,n413);
not (n413,n317);
or (n414,n317,n328);
and (n415,n397,n404);
xor (n416,n306,n333);
or (n417,n418,n498);
and (n418,n419,n440);
xor (n419,n420,n439);
or (n420,n421,n438);
and (n421,n422,n431);
xor (n422,n423,n424);
nor (n423,n46,n36);
nand (n424,n425,n430);
or (n425,n426,n86);
not (n426,n427);
nor (n427,n428,n429);
and (n428,n42,n48);
and (n429,n49,n40);
nand (n430,n88,n400);
nand (n431,n432,n437);
or (n432,n175,n433);
not (n433,n434);
nor (n434,n435,n436);
and (n435,n123,n90);
and (n436,n91,n124);
or (n437,n319,n176);
and (n438,n423,n424);
xor (n439,n396,n411);
or (n440,n441,n497);
and (n441,n442,n496);
xor (n442,n443,n457);
nor (n443,n444,n452);
not (n444,n445);
nand (n445,n446,n447);
or (n446,n176,n433);
nand (n447,n448,n451);
nor (n448,n449,n450);
and (n449,n169,n90);
and (n450,n91,n167);
not (n451,n175);
nand (n452,n453,n49);
nand (n453,n454,n455);
or (n454,n92,n91);
or (n455,n456,n33);
and (n456,n91,n92);
nand (n457,n458,n495);
or (n458,n459,n483);
not (n459,n460);
nand (n460,n461,n482);
or (n461,n462,n471);
nor (n462,n463,n464);
and (n463,n88,n33);
nand (n464,n465,n467);
or (n465,n176,n466);
not (n466,n448);
nand (n467,n468,n451);
nand (n468,n469,n470);
or (n469,n42,n91);
or (n470,n90,n40);
nand (n471,n472,n475);
not (n472,n473);
nand (n473,n474,n91);
nand (n474,n33,n177);
nand (n475,n476,n478);
or (n476,n176,n477);
not (n477,n468);
nand (n478,n479,n451);
nor (n479,n480,n481);
and (n480,n36,n90);
and (n481,n91,n33);
nand (n482,n463,n464);
not (n483,n484);
nand (n484,n485,n489);
nor (n485,n486,n487);
and (n486,n452,n445);
and (n487,n488,n444);
not (n488,n452);
nor (n489,n490,n494);
and (n490,n87,n491);
nand (n491,n492,n493);
or (n492,n49,n36);
or (n493,n48,n33);
and (n494,n88,n427);
or (n495,n485,n489);
xor (n496,n422,n431);
and (n497,n443,n457);
and (n498,n420,n439);
and (n499,n394,n416);
and (n500,n304,n355);
nor (n501,n502,n527);
nor (n502,n503,n518);
xor (n503,n504,n517);
xor (n504,n505,n506);
xor (n505,n236,n250);
or (n506,n507,n516);
and (n507,n508,n515);
xor (n508,n509,n512);
nand (n509,n510,n511);
or (n510,n380,n86);
nand (n511,n88,n229);
nand (n512,n513,n514);
or (n513,n45,n388);
or (n514,n46,n270);
and (n515,n358,n364);
and (n516,n509,n512);
xor (n517,n267,n275);
or (n518,n519,n526);
and (n519,n520,n525);
xor (n520,n521,n524);
or (n521,n522,n523);
and (n522,n371,n385);
and (n523,n372,n378);
xor (n524,n277,n285);
xor (n525,n508,n515);
and (n526,n521,n524);
nor (n527,n528,n529);
xor (n528,n520,n525);
or (n529,n530,n531);
and (n530,n356,n370);
and (n531,n357,n367);
not (n532,n533);
nand (n533,n534,n539);
or (n534,n535,n537);
not (n535,n536);
nand (n536,n528,n529);
not (n537,n538);
nand (n538,n503,n518);
not (n539,n502);
nor (n540,n541,n542);
xor (n541,n263,n293);
or (n542,n543,n544);
and (n543,n504,n517);
and (n544,n505,n506);
nand (n545,n541,n542);
or (n546,n297,n10);
not (n547,n548);
nand (n548,n549,n3);
not (n549,n4);
wire s0n550,s1n550,notn550;
or (n550,s0n550,s1n550);
not(notn550,n4);
and (s0n550,notn550,n551);
and (s1n550,n4,1'b0);
wire s0n551,s1n551,notn551;
or (n551,s0n551,s1n551);
not(notn551,n3);
and (s0n551,notn551,n5);
and (s1n551,n3,n552);
xor (n552,n553,n876);
xor (n553,n554,n873);
xor (n554,n555,n872);
xor (n555,n556,n863);
xor (n556,n557,n862);
xor (n557,n558,n848);
xor (n558,n559,n847);
xor (n559,n560,n826);
xor (n560,n561,n825);
xor (n561,n562,n799);
xor (n562,n563,n798);
xor (n563,n564,n765);
xor (n564,n565,n764);
xor (n565,n566,n726);
xor (n566,n567,n725);
xor (n567,n568,n682);
xor (n568,n569,n681);
xor (n569,n570,n631);
xor (n570,n571,n630);
xor (n571,n572,n575);
xor (n572,n573,n574);
and (n573,n29,n33);
and (n574,n24,n40);
or (n575,n576,n579);
and (n576,n577,n578);
and (n577,n24,n33);
and (n578,n23,n40);
and (n579,n580,n581);
xor (n580,n577,n578);
or (n581,n582,n585);
and (n582,n583,n584);
and (n583,n23,n33);
and (n584,n158,n40);
and (n585,n586,n587);
xor (n586,n583,n584);
or (n587,n588,n591);
and (n588,n589,n590);
and (n589,n158,n33);
and (n590,n122,n40);
and (n591,n592,n593);
xor (n592,n589,n590);
or (n593,n594,n597);
and (n594,n595,n596);
and (n595,n122,n33);
and (n596,n130,n40);
and (n597,n598,n599);
xor (n598,n595,n596);
or (n599,n600,n603);
and (n600,n601,n602);
and (n601,n130,n33);
and (n602,n56,n40);
and (n603,n604,n605);
xor (n604,n601,n602);
or (n605,n606,n609);
and (n606,n607,n608);
and (n607,n56,n33);
and (n608,n50,n40);
and (n609,n610,n611);
xor (n610,n607,n608);
or (n611,n612,n614);
and (n612,n613,n429);
and (n613,n50,n33);
and (n614,n615,n616);
xor (n615,n613,n429);
or (n616,n617,n620);
and (n617,n618,n619);
and (n618,n49,n33);
and (n619,n92,n40);
and (n620,n621,n622);
xor (n621,n618,n619);
or (n622,n623,n626);
and (n623,n624,n625);
and (n624,n92,n33);
and (n625,n91,n40);
and (n626,n627,n628);
xor (n627,n624,n625);
and (n628,n481,n629);
and (n629,n177,n40);
and (n630,n23,n167);
or (n631,n632,n635);
and (n632,n633,n634);
xor (n633,n580,n581);
and (n634,n158,n167);
and (n635,n636,n637);
xor (n636,n633,n634);
or (n637,n638,n641);
and (n638,n639,n640);
xor (n639,n586,n587);
and (n640,n122,n167);
and (n641,n642,n643);
xor (n642,n639,n640);
or (n643,n644,n647);
and (n644,n645,n646);
xor (n645,n592,n593);
and (n646,n130,n167);
and (n647,n648,n649);
xor (n648,n645,n646);
or (n649,n650,n653);
and (n650,n651,n652);
xor (n651,n598,n599);
and (n652,n56,n167);
and (n653,n654,n655);
xor (n654,n651,n652);
or (n655,n656,n659);
and (n656,n657,n658);
xor (n657,n604,n605);
and (n658,n50,n167);
and (n659,n660,n661);
xor (n660,n657,n658);
or (n661,n662,n665);
and (n662,n663,n664);
xor (n663,n610,n611);
and (n664,n49,n167);
and (n665,n666,n667);
xor (n666,n663,n664);
or (n667,n668,n671);
and (n668,n669,n670);
xor (n669,n615,n616);
and (n670,n92,n167);
and (n671,n672,n673);
xor (n672,n669,n670);
or (n673,n674,n676);
and (n674,n675,n450);
xor (n675,n621,n622);
and (n676,n677,n678);
xor (n677,n675,n450);
and (n678,n679,n680);
xor (n679,n627,n628);
and (n680,n177,n167);
and (n681,n158,n124);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n636,n637);
and (n685,n122,n124);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n642,n643);
and (n691,n130,n124);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n698);
and (n695,n696,n697);
xor (n696,n648,n649);
and (n697,n56,n124);
and (n698,n699,n700);
xor (n699,n696,n697);
or (n700,n701,n704);
and (n701,n702,n703);
xor (n702,n654,n655);
and (n703,n50,n124);
and (n704,n705,n706);
xor (n705,n702,n703);
or (n706,n707,n709);
and (n707,n708,n348);
xor (n708,n660,n661);
and (n709,n710,n711);
xor (n710,n708,n348);
or (n711,n712,n715);
and (n712,n713,n714);
xor (n713,n666,n667);
and (n714,n92,n124);
and (n715,n716,n717);
xor (n716,n713,n714);
or (n717,n718,n720);
and (n718,n719,n436);
xor (n719,n672,n673);
and (n720,n721,n722);
xor (n721,n719,n436);
and (n722,n723,n724);
xor (n723,n677,n678);
and (n724,n177,n124);
and (n725,n122,n140);
or (n726,n727,n730);
and (n727,n728,n729);
xor (n728,n687,n688);
and (n729,n130,n140);
and (n730,n731,n732);
xor (n731,n728,n729);
or (n732,n733,n736);
and (n733,n734,n735);
xor (n734,n693,n694);
and (n735,n56,n140);
and (n736,n737,n738);
xor (n737,n734,n735);
or (n738,n739,n742);
and (n739,n740,n741);
xor (n740,n699,n700);
and (n741,n50,n140);
and (n742,n743,n744);
xor (n743,n740,n741);
or (n744,n745,n748);
and (n745,n746,n747);
xor (n746,n705,n706);
and (n747,n49,n140);
and (n748,n749,n750);
xor (n749,n746,n747);
or (n750,n751,n754);
and (n751,n752,n753);
xor (n752,n710,n711);
and (n753,n92,n140);
and (n754,n755,n756);
xor (n755,n752,n753);
or (n756,n757,n759);
and (n757,n758,n321);
xor (n758,n716,n717);
and (n759,n760,n761);
xor (n760,n758,n321);
and (n761,n762,n763);
xor (n762,n721,n722);
and (n763,n177,n140);
and (n764,n130,n188);
or (n765,n766,n769);
and (n766,n767,n768);
xor (n767,n731,n732);
and (n768,n56,n188);
and (n769,n770,n771);
xor (n770,n767,n768);
or (n771,n772,n775);
and (n772,n773,n774);
xor (n773,n737,n738);
and (n774,n50,n188);
and (n775,n776,n777);
xor (n776,n773,n774);
or (n777,n778,n781);
and (n778,n779,n780);
xor (n779,n743,n744);
and (n780,n49,n188);
and (n781,n782,n783);
xor (n782,n779,n780);
or (n783,n784,n787);
and (n784,n785,n786);
xor (n785,n749,n750);
and (n786,n92,n188);
and (n787,n788,n789);
xor (n788,n785,n786);
or (n789,n790,n793);
and (n790,n791,n792);
xor (n791,n755,n756);
and (n792,n91,n188);
and (n793,n794,n795);
xor (n794,n791,n792);
and (n795,n796,n797);
xor (n796,n760,n761);
and (n797,n177,n188);
and (n798,n56,n60);
or (n799,n800,n803);
and (n800,n801,n802);
xor (n801,n770,n771);
and (n802,n50,n60);
and (n803,n804,n805);
xor (n804,n801,n802);
or (n805,n806,n809);
and (n806,n807,n808);
xor (n807,n776,n777);
and (n808,n49,n60);
and (n809,n810,n811);
xor (n810,n807,n808);
or (n811,n812,n815);
and (n812,n813,n814);
xor (n813,n782,n783);
and (n814,n92,n60);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n820);
and (n818,n819,n340);
xor (n819,n788,n789);
and (n820,n821,n822);
xor (n821,n819,n340);
and (n822,n823,n824);
xor (n823,n794,n795);
and (n824,n177,n60);
and (n825,n50,n66);
or (n826,n827,n830);
and (n827,n828,n829);
xor (n828,n804,n805);
and (n829,n49,n66);
and (n830,n831,n832);
xor (n831,n828,n829);
or (n832,n833,n836);
and (n833,n834,n835);
xor (n834,n810,n811);
and (n835,n92,n66);
and (n836,n837,n838);
xor (n837,n834,n835);
or (n838,n839,n842);
and (n839,n840,n841);
xor (n840,n816,n817);
and (n841,n91,n66);
and (n842,n843,n844);
xor (n843,n840,n841);
and (n844,n845,n846);
xor (n845,n821,n822);
and (n846,n177,n66);
and (n847,n49,n84);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n831,n832);
and (n851,n92,n84);
and (n852,n853,n854);
xor (n853,n850,n851);
or (n854,n855,n857);
and (n855,n856,n255);
xor (n856,n837,n838);
and (n857,n858,n859);
xor (n858,n856,n255);
and (n859,n860,n861);
xor (n860,n843,n844);
and (n861,n177,n84);
and (n862,n92,n102);
or (n863,n864,n867);
and (n864,n865,n866);
xor (n865,n853,n854);
and (n866,n91,n102);
and (n867,n868,n869);
xor (n868,n865,n866);
and (n869,n870,n871);
xor (n870,n858,n859);
and (n871,n177,n102);
and (n872,n91,n181);
and (n873,n874,n875);
xor (n874,n868,n869);
and (n875,n177,n181);
and (n876,n177,n213);
endmodule
