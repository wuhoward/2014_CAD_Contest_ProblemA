module top (out,n14,n16,n17,n19,n22,n26,n28,n30,n33
        ,n37,n39,n41,n44,n50,n52,n54,n57,n61,n63
        ,n65,n68,n73,n75,n76,n90,n104,n105,n177,n186
        ,n187,n223,n295,n325,n326,n530,n534,n536,n562,n563
        ,n670,n687,n688,n855,n859,n861,n872,n884,n898);
output out;
input n14;
input n16;
input n17;
input n19;
input n22;
input n26;
input n28;
input n30;
input n33;
input n37;
input n39;
input n41;
input n44;
input n50;
input n52;
input n54;
input n57;
input n61;
input n63;
input n65;
input n68;
input n73;
input n75;
input n76;
input n90;
input n104;
input n105;
input n177;
input n186;
input n187;
input n223;
input n295;
input n325;
input n326;
input n530;
input n534;
input n536;
input n562;
input n563;
input n670;
input n687;
input n688;
input n855;
input n859;
input n861;
input n872;
input n884;
input n898;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n18;
wire n20;
wire n21;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n38;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n53;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n62;
wire n64;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n531;
wire n532;
wire n533;
wire n535;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n856;
wire n857;
wire n858;
wire n860;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
xor (out,n0,n2857);
xnor (n0,n1,n2798);
nand (n1,n2,n425);
nor (n2,n3,n423);
nor (n3,n4,n368);
nand (n4,n5,n245);
xor (n5,n6,n202);
xor (n6,n7,n93);
xor (n7,n8,n80);
xor (n8,n9,n45);
xor (n9,n10,n34);
xor (n10,n11,n23);
xor (n11,n12,n22);
or (n12,n13,n18);
and (n13,n14,n15);
xor (n15,n16,n17);
and (n18,n19,n20);
nor (n20,n15,n21);
xnor (n21,n22,n16);
xor (n23,n24,n33);
or (n24,n25,n29);
and (n25,n26,n27);
xor (n27,n28,n22);
and (n29,n30,n31);
nor (n31,n27,n32);
xnor (n32,n33,n28);
xor (n34,n35,n44);
or (n35,n36,n40);
and (n36,n37,n38);
xor (n38,n39,n33);
and (n40,n41,n42);
nor (n42,n38,n43);
xnor (n43,n44,n39);
xor (n45,n46,n69);
xor (n46,n47,n58);
xor (n47,n48,n57);
or (n48,n49,n53);
and (n49,n50,n51);
xor (n51,n52,n44);
and (n53,n54,n55);
nor (n55,n51,n56);
xnor (n56,n57,n52);
xor (n58,n59,n68);
or (n59,n60,n64);
and (n60,n61,n62);
xor (n62,n63,n57);
and (n64,n65,n66);
nor (n66,n62,n67);
xnor (n67,n68,n63);
not (n69,n70);
xor (n70,n71,n17);
or (n71,n72,n77);
and (n72,n73,n74);
xor (n74,n75,n76);
and (n77,n73,n78);
nor (n78,n74,n79);
xnor (n79,n17,n75);
nand (n80,n81,n91,n92);
nand (n81,n82,n86);
xor (n82,n83,n57);
or (n83,n84,n85);
and (n84,n54,n51);
and (n85,n61,n55);
xor (n86,n87,n68);
or (n87,n88,n89);
and (n88,n65,n62);
and (n89,n90,n66);
nand (n91,n68,n86);
nand (n92,n82,n68);
xor (n93,n94,n164);
xor (n94,n95,n130);
xor (n95,n96,n118);
xor (n96,n68,n97);
nand (n97,n98,n112,n117);
nand (n98,n99,n109);
not (n99,n100);
xor (n100,n101,n76);
or (n101,n102,n106);
and (n102,n73,n103);
xor (n103,n104,n105);
and (n106,n73,n107);
nor (n107,n103,n108);
xnor (n108,n76,n104);
xor (n109,n110,n17);
or (n110,n72,n111);
and (n111,n14,n78);
nand (n112,n113,n109);
xor (n113,n114,n33);
or (n114,n115,n116);
and (n115,n30,n27);
and (n116,n37,n31);
nand (n117,n99,n113);
nand (n118,n119,n124,n129);
nand (n119,n120,n100);
xor (n120,n121,n22);
or (n121,n122,n123);
and (n122,n19,n15);
and (n123,n26,n20);
nand (n124,n125,n100);
xor (n125,n126,n44);
or (n126,n127,n128);
and (n127,n41,n38);
and (n128,n50,n42);
nand (n129,n120,n125);
nand (n130,n131,n150,n163);
nand (n131,n132,n134);
xor (n132,n133,n113);
xor (n133,n99,n109);
nand (n134,n135,n144,n149);
nand (n135,n136,n140);
xor (n136,n137,n17);
or (n137,n138,n139);
and (n138,n14,n74);
and (n139,n19,n78);
xor (n140,n141,n33);
or (n141,n142,n143);
and (n142,n37,n27);
and (n143,n41,n31);
nand (n144,n145,n140);
xor (n145,n146,n22);
or (n146,n147,n148);
and (n147,n26,n15);
and (n148,n30,n20);
nand (n149,n136,n145);
nand (n150,n151,n134);
nand (n151,n152,n157,n162);
nand (n152,n99,n153);
xor (n153,n154,n44);
or (n154,n155,n156);
and (n155,n50,n38);
and (n156,n54,n42);
nand (n157,n158,n153);
xor (n158,n159,n57);
or (n159,n160,n161);
and (n160,n61,n51);
and (n161,n65,n55);
nand (n162,n99,n158);
nand (n163,n132,n151);
nand (n164,n165,n170,n201);
nand (n165,n166,n168);
xor (n166,n167,n68);
xor (n167,n82,n86);
xor (n168,n169,n125);
xor (n169,n120,n100);
nand (n170,n171,n168);
nand (n171,n172,n178,n200);
nand (n172,n173,n68);
xor (n173,n174,n68);
or (n174,n175,n176);
and (n175,n90,n62);
and (n176,n177,n66);
nand (n178,n179,n68);
nand (n179,n180,n194,n199);
nand (n180,n181,n191);
not (n181,n182);
xor (n182,n183,n105);
or (n183,n184,n188);
and (n184,n73,n185);
xor (n185,n186,n187);
and (n188,n73,n189);
nor (n189,n185,n190);
xnor (n190,n105,n186);
xor (n191,n192,n76);
or (n192,n102,n193);
and (n193,n14,n107);
nand (n194,n195,n191);
xor (n195,n196,n17);
or (n196,n197,n198);
and (n197,n19,n74);
and (n198,n26,n78);
nand (n199,n181,n195);
nand (n200,n173,n179);
nand (n201,n166,n171);
nand (n202,n203,n241,n244);
nand (n203,n204,n239);
nand (n204,n205,n225,n238);
nand (n205,n206,n208);
xor (n206,n207,n145);
xor (n207,n136,n140);
nand (n208,n209,n218,n224);
nand (n209,n210,n214);
xor (n210,n211,n22);
or (n211,n212,n213);
and (n212,n30,n15);
and (n213,n37,n20);
xor (n214,n215,n33);
or (n215,n216,n217);
and (n216,n41,n27);
and (n217,n50,n31);
nand (n218,n219,n214);
xor (n219,n220,n68);
or (n220,n221,n222);
and (n221,n177,n62);
and (n222,n223,n66);
nand (n224,n210,n219);
nand (n225,n226,n208);
nand (n226,n227,n232,n237);
nand (n227,n182,n228);
xor (n228,n229,n44);
or (n229,n230,n231);
and (n230,n54,n38);
and (n231,n61,n42);
nand (n232,n233,n228);
xor (n233,n234,n57);
or (n234,n235,n236);
and (n235,n65,n51);
and (n236,n90,n55);
nand (n237,n182,n233);
nand (n238,n206,n226);
xor (n239,n240,n151);
xor (n240,n132,n134);
nand (n241,n242,n239);
xor (n242,n243,n171);
xor (n243,n166,n168);
nand (n244,n204,n242);
nand (n245,n246,n278,n367);
nand (n246,n247,n276);
nand (n247,n248,n252,n275);
nand (n248,n249,n251);
xor (n249,n250,n158);
xor (n250,n99,n153);
xor (n251,n174,n179);
nand (n252,n253,n251);
nand (n253,n254,n257,n274);
nand (n254,n68,n255);
xor (n255,n256,n195);
xor (n256,n181,n191);
nand (n257,n258,n255);
nand (n258,n259,n268,n273);
nand (n259,n260,n264);
xor (n260,n261,n76);
or (n261,n262,n263);
and (n262,n14,n103);
and (n263,n19,n107);
xor (n264,n265,n17);
or (n265,n266,n267);
and (n266,n26,n74);
and (n267,n30,n78);
nand (n268,n269,n264);
xor (n269,n270,n22);
or (n270,n271,n272);
and (n271,n37,n15);
and (n272,n41,n20);
nand (n273,n260,n269);
nand (n274,n68,n258);
nand (n275,n249,n253);
xor (n276,n277,n242);
xor (n277,n204,n239);
nand (n278,n279,n276);
nand (n279,n280,n304,n366);
nand (n280,n281,n283);
xor (n281,n282,n226);
xor (n282,n206,n208);
nand (n283,n284,n300,n303);
nand (n284,n285,n298);
nand (n285,n286,n296,n297);
nand (n286,n287,n291);
xor (n287,n288,n33);
or (n288,n289,n290);
and (n289,n50,n27);
and (n290,n54,n31);
xor (n291,n292,n68);
or (n292,n293,n294);
and (n293,n223,n62);
and (n294,n295,n66);
nand (n296,n181,n291);
nand (n297,n287,n181);
xor (n298,n299,n219);
xor (n299,n210,n214);
nand (n300,n301,n298);
xor (n301,n302,n233);
xor (n302,n182,n228);
nand (n303,n285,n301);
nand (n304,n305,n283);
nand (n305,n306,n362,n365);
nand (n306,n307,n340);
nand (n307,n308,n317,n339);
nand (n308,n309,n313);
xor (n309,n310,n44);
or (n310,n311,n312);
and (n311,n61,n38);
and (n312,n65,n42);
xor (n313,n314,n57);
or (n314,n315,n316);
and (n315,n90,n51);
and (n316,n177,n55);
nand (n317,n318,n313);
nand (n318,n319,n333,n338);
nand (n319,n320,n330);
not (n320,n321);
xor (n321,n322,n187);
or (n322,n323,n327);
and (n323,n73,n324);
xor (n324,n325,n326);
and (n327,n73,n328);
nor (n328,n324,n329);
xnor (n329,n187,n325);
xor (n330,n331,n105);
or (n331,n184,n332);
and (n332,n14,n189);
nand (n333,n334,n330);
xor (n334,n335,n17);
or (n335,n336,n337);
and (n336,n30,n74);
and (n337,n37,n78);
nand (n338,n320,n334);
nand (n339,n309,n318);
nand (n340,n341,n344,n361);
nand (n341,n68,n342);
xor (n342,n343,n269);
xor (n343,n260,n264);
nand (n344,n345,n342);
nand (n345,n346,n355,n360);
nand (n346,n347,n351);
xor (n347,n348,n76);
or (n348,n349,n350);
and (n349,n19,n103);
and (n350,n26,n107);
xor (n351,n352,n22);
or (n352,n353,n354);
and (n353,n41,n15);
and (n354,n50,n20);
nand (n355,n356,n351);
xor (n356,n357,n33);
or (n357,n358,n359);
and (n358,n54,n27);
and (n359,n61,n31);
nand (n360,n347,n356);
nand (n361,n68,n345);
nand (n362,n363,n340);
xor (n363,n364,n258);
xor (n364,n68,n255);
nand (n365,n307,n363);
nand (n366,n281,n305);
nand (n367,n247,n279);
nor (n368,n369,n373);
nand (n369,n370,n371,n372);
nand (n370,n7,n93);
nand (n371,n202,n93);
nand (n372,n7,n202);
xor (n373,n374,n419);
xor (n374,n375,n379);
nand (n375,n376,n377,n378);
nand (n376,n9,n45);
nand (n377,n80,n45);
nand (n378,n9,n80);
xor (n379,n380,n393);
xor (n380,n381,n385);
nand (n381,n382,n383,n384);
nand (n382,n68,n97);
nand (n383,n118,n97);
nand (n384,n68,n118);
xor (n385,n386,n389);
or (n386,n387,n388);
and (n387,n54,n62);
and (n388,n61,n66);
nand (n389,n390,n391,n392);
nand (n390,n11,n23);
nand (n391,n34,n23);
nand (n392,n11,n34);
xor (n393,n394,n409);
xor (n394,n395,n399);
nand (n395,n396,n397,n398);
nand (n396,n47,n58);
nand (n397,n69,n58);
nand (n398,n47,n69);
xor (n399,n400,n405);
xor (n400,n69,n401);
xor (n401,n402,n22);
or (n402,n403,n404);
and (n403,n73,n15);
and (n404,n14,n20);
xor (n405,n406,n33);
or (n406,n407,n408);
and (n407,n19,n27);
and (n408,n26,n31);
xor (n409,n410,n415);
xor (n410,n411,n70);
xor (n411,n412,n44);
or (n412,n413,n414);
and (n413,n30,n38);
and (n414,n37,n42);
xor (n415,n416,n57);
or (n416,n417,n418);
and (n417,n41,n51);
and (n418,n50,n55);
nand (n419,n420,n421,n422);
nand (n420,n95,n130);
nand (n421,n164,n130);
nand (n422,n95,n164);
not (n423,n424);
nand (n424,n369,n373);
nand (n425,n426,n428);
nor (n426,n427,n368);
nor (n427,n5,n245);
nand (n428,n429,n836);
nor (n429,n430,n830);
nor (n430,n431,n806);
nor (n431,n432,n804);
nor (n432,n433,n779);
nand (n433,n434,n741);
nand (n434,n435,n657,n740);
nand (n435,n436,n520);
xor (n436,n437,n510);
xor (n437,n438,n460);
xor (n438,n439,n444);
xor (n439,n440,n68);
xor (n440,n441,n44);
or (n441,n442,n443);
and (n442,n65,n38);
and (n443,n90,n42);
nand (n444,n445,n454,n459);
nand (n445,n446,n450);
xor (n446,n447,n17);
or (n447,n448,n449);
and (n448,n37,n74);
and (n449,n41,n78);
xor (n450,n451,n105);
or (n451,n452,n453);
and (n452,n14,n185);
and (n453,n19,n189);
nand (n454,n455,n450);
xor (n455,n456,n76);
or (n456,n457,n458);
and (n457,n26,n103);
and (n458,n30,n107);
nand (n459,n446,n455);
nand (n460,n461,n492,n509);
nand (n461,n462,n478);
nand (n462,n463,n472,n477);
nand (n463,n464,n468);
xor (n464,n465,n17);
or (n465,n466,n467);
and (n466,n41,n74);
and (n467,n50,n78);
xor (n468,n469,n105);
or (n469,n470,n471);
and (n470,n19,n185);
and (n471,n26,n189);
nand (n472,n473,n468);
xor (n473,n474,n22);
or (n474,n475,n476);
and (n475,n54,n15);
and (n476,n61,n20);
nand (n477,n464,n473);
xor (n478,n479,n488);
xor (n479,n480,n484);
xor (n480,n481,n22);
or (n481,n482,n483);
and (n482,n50,n15);
and (n483,n54,n20);
xor (n484,n485,n33);
or (n485,n486,n487);
and (n486,n61,n27);
and (n487,n65,n31);
xor (n488,n489,n57);
or (n489,n490,n491);
and (n490,n223,n51);
and (n491,n295,n55);
nand (n492,n493,n478);
nand (n493,n494,n503,n508);
nand (n494,n495,n499);
xor (n495,n496,n187);
or (n496,n497,n498);
and (n497,n14,n324);
and (n498,n19,n328);
xor (n499,n500,n33);
or (n500,n501,n502);
and (n501,n65,n27);
and (n502,n90,n31);
nand (n503,n504,n499);
xor (n504,n505,n44);
or (n505,n506,n507);
and (n506,n177,n38);
and (n507,n223,n42);
nand (n508,n495,n504);
nand (n509,n462,n493);
xor (n510,n511,n516);
xor (n511,n512,n514);
xor (n512,n513,n334);
xor (n513,n320,n330);
xor (n514,n515,n356);
xor (n515,n347,n351);
nand (n516,n517,n518,n519);
nand (n517,n480,n484);
nand (n518,n488,n484);
nand (n519,n480,n488);
xor (n520,n521,n596);
xor (n521,n522,n576);
nand (n522,n523,n549,n575);
nand (n523,n524,n539);
nand (n524,n525,n537,n538);
nand (n525,n526,n531);
xor (n526,n527,n57);
or (n527,n528,n529);
and (n528,n295,n51);
and (n529,n530,n55);
xor (n531,n532,n68);
or (n532,n533,n535);
and (n533,n534,n62);
and (n535,n536,n66);
nand (n537,n68,n531);
nand (n538,n526,n68);
xor (n539,n540,n545);
xor (n540,n541,n320);
xor (n541,n542,n68);
or (n542,n543,n544);
and (n543,n530,n62);
and (n544,n534,n66);
xor (n545,n546,n44);
or (n546,n547,n548);
and (n547,n90,n38);
and (n548,n177,n42);
nand (n549,n550,n539);
xor (n550,n551,n573);
xor (n551,n68,n552);
nand (n552,n553,n567,n572);
nand (n553,n554,n557);
xor (n554,n555,n187);
or (n555,n323,n556);
and (n556,n14,n328);
not (n557,n558);
xor (n558,n559,n326);
or (n559,n560,n564);
and (n560,n73,n561);
xor (n561,n562,n563);
and (n564,n73,n565);
nor (n565,n561,n566);
xnor (n566,n326,n562);
nand (n567,n568,n557);
xor (n568,n569,n76);
or (n569,n570,n571);
and (n570,n30,n103);
and (n571,n37,n107);
nand (n572,n554,n568);
xor (n573,n574,n455);
xor (n574,n446,n450);
nand (n575,n524,n550);
xor (n576,n577,n592);
xor (n577,n578,n582);
nand (n578,n579,n580,n581);
nand (n579,n541,n320);
nand (n580,n545,n320);
nand (n581,n541,n545);
xor (n582,n583,n321);
xor (n583,n584,n588);
xor (n584,n585,n57);
or (n585,n586,n587);
and (n586,n177,n51);
and (n587,n223,n55);
xor (n588,n589,n68);
or (n589,n590,n591);
and (n590,n295,n62);
and (n591,n530,n66);
nand (n592,n593,n594,n595);
nand (n593,n68,n552);
nand (n594,n573,n552);
nand (n595,n68,n573);
nand (n596,n597,n653,n656);
nand (n597,n598,n618);
nand (n598,n599,n614,n617);
nand (n599,n600,n612);
nand (n600,n601,n606,n611);
nand (n601,n558,n602);
xor (n602,n603,n76);
or (n603,n604,n605);
and (n604,n37,n103);
and (n605,n41,n107);
nand (n606,n607,n602);
xor (n607,n608,n17);
or (n608,n609,n610);
and (n609,n50,n74);
and (n610,n54,n78);
nand (n611,n558,n607);
xor (n612,n613,n473);
xor (n613,n464,n468);
nand (n614,n615,n612);
xor (n615,n616,n568);
xor (n616,n554,n557);
nand (n617,n600,n615);
nand (n618,n619,n649,n652);
nand (n619,n620,n633);
nand (n620,n621,n627,n632);
nand (n621,n622,n626);
xor (n622,n623,n105);
or (n623,n624,n625);
and (n624,n26,n185);
and (n625,n30,n189);
not (n626,n495);
nand (n627,n628,n626);
xor (n628,n629,n22);
or (n629,n630,n631);
and (n630,n61,n15);
and (n631,n65,n20);
nand (n632,n622,n628);
nand (n633,n634,n643,n648);
nand (n634,n635,n639);
xor (n635,n636,n33);
or (n636,n637,n638);
and (n637,n90,n27);
and (n638,n177,n31);
xor (n639,n640,n44);
or (n640,n641,n642);
and (n641,n223,n38);
and (n642,n295,n42);
nand (n643,n644,n639);
xor (n644,n645,n57);
or (n645,n646,n647);
and (n646,n530,n51);
and (n647,n534,n55);
nand (n648,n635,n644);
nand (n649,n650,n633);
xor (n650,n651,n504);
xor (n651,n495,n499);
nand (n652,n620,n650);
nand (n653,n654,n618);
xor (n654,n655,n493);
xor (n655,n462,n478);
nand (n656,n598,n654);
nand (n657,n658,n520);
nand (n658,n659,n736,n739);
nand (n659,n660,n662);
xor (n660,n661,n550);
xor (n661,n524,n539);
nand (n662,n663,n696,n735);
nand (n663,n664,n694);
nand (n664,n665,n671,n693);
nand (n665,n666,n68);
xor (n666,n667,n68);
or (n667,n668,n669);
and (n668,n536,n62);
and (n669,n670,n66);
nand (n671,n672,n68);
nand (n672,n673,n681,n692);
nand (n673,n674,n677);
xor (n674,n675,n326);
or (n675,n560,n676);
and (n676,n14,n565);
xor (n677,n678,n187);
or (n678,n679,n680);
and (n679,n19,n324);
and (n680,n26,n328);
nand (n681,n682,n677);
not (n682,n683);
xor (n683,n684,n563);
or (n684,n685,n689);
and (n685,n73,n686);
xor (n686,n687,n688);
and (n689,n73,n690);
nor (n690,n686,n691);
xnor (n691,n563,n687);
nand (n692,n674,n682);
nand (n693,n666,n672);
xor (n694,n695,n68);
xor (n695,n526,n531);
nand (n696,n697,n694);
nand (n697,n698,n717,n734);
nand (n698,n699,n715);
nand (n699,n700,n709,n714);
nand (n700,n701,n705);
xor (n701,n702,n105);
or (n702,n703,n704);
and (n703,n30,n185);
and (n704,n37,n189);
xor (n705,n706,n76);
or (n706,n707,n708);
and (n707,n41,n103);
and (n708,n50,n107);
nand (n709,n710,n705);
xor (n710,n711,n17);
or (n711,n712,n713);
and (n712,n54,n74);
and (n713,n61,n78);
nand (n714,n701,n710);
xor (n715,n716,n607);
xor (n716,n558,n602);
nand (n717,n718,n715);
nand (n718,n719,n728,n733);
nand (n719,n720,n724);
xor (n720,n721,n33);
or (n721,n722,n723);
and (n722,n177,n27);
and (n723,n223,n31);
xor (n724,n725,n326);
or (n725,n726,n727);
and (n726,n14,n561);
and (n727,n19,n565);
nand (n728,n729,n724);
xor (n729,n730,n22);
or (n730,n731,n732);
and (n731,n65,n15);
and (n732,n90,n20);
nand (n733,n720,n729);
nand (n734,n699,n718);
nand (n735,n664,n697);
nand (n736,n737,n662);
xor (n737,n738,n654);
xor (n738,n598,n618);
nand (n739,n660,n737);
nand (n740,n436,n658);
xor (n741,n742,n775);
xor (n742,n743,n747);
nand (n743,n744,n745,n746);
nand (n744,n438,n460);
nand (n745,n510,n460);
nand (n746,n438,n510);
xor (n747,n748,n763);
xor (n748,n749,n753);
nand (n749,n750,n751,n752);
nand (n750,n578,n582);
nand (n751,n592,n582);
nand (n752,n578,n592);
xor (n753,n754,n761);
xor (n754,n755,n759);
nand (n755,n756,n757,n758);
nand (n756,n584,n588);
nand (n757,n321,n588);
nand (n758,n584,n321);
xor (n759,n760,n318);
xor (n760,n309,n313);
xor (n761,n762,n181);
xor (n762,n287,n291);
xor (n763,n764,n771);
xor (n764,n765,n769);
nand (n765,n766,n767,n768);
nand (n766,n440,n68);
nand (n767,n444,n68);
nand (n768,n440,n444);
xor (n769,n770,n345);
xor (n770,n68,n342);
nand (n771,n772,n773,n774);
nand (n772,n512,n514);
nand (n773,n516,n514);
nand (n774,n512,n516);
nand (n775,n776,n777,n778);
nand (n776,n522,n576);
nand (n777,n596,n576);
nand (n778,n522,n596);
nor (n779,n780,n784);
nand (n780,n781,n782,n783);
nand (n781,n743,n747);
nand (n782,n775,n747);
nand (n783,n743,n775);
xor (n784,n785,n800);
xor (n785,n786,n788);
xor (n786,n787,n363);
xor (n787,n307,n340);
xor (n788,n789,n796);
xor (n789,n790,n792);
xor (n790,n791,n301);
xor (n791,n285,n298);
nand (n792,n793,n794,n795);
nand (n793,n755,n759);
nand (n794,n761,n759);
nand (n795,n755,n761);
nand (n796,n797,n798,n799);
nand (n797,n765,n769);
nand (n798,n771,n769);
nand (n799,n765,n771);
nand (n800,n801,n802,n803);
nand (n801,n749,n753);
nand (n802,n763,n753);
nand (n803,n749,n763);
not (n804,n805);
nand (n805,n780,n784);
not (n806,n807);
nor (n807,n808,n823);
nor (n808,n809,n813);
nand (n809,n810,n811,n812);
nand (n810,n786,n788);
nand (n811,n800,n788);
nand (n812,n786,n800);
xor (n813,n814,n819);
xor (n814,n815,n817);
xor (n815,n816,n253);
xor (n816,n249,n251);
xor (n817,n818,n305);
xor (n818,n281,n283);
nand (n819,n820,n821,n822);
nand (n820,n790,n792);
nand (n821,n796,n792);
nand (n822,n790,n796);
nor (n823,n824,n828);
nand (n824,n825,n826,n827);
nand (n825,n815,n817);
nand (n826,n819,n817);
nand (n827,n815,n819);
xor (n828,n829,n279);
xor (n829,n247,n276);
not (n830,n831);
nor (n831,n832,n834);
nor (n832,n833,n823);
nand (n833,n809,n813);
not (n834,n835);
nand (n835,n824,n828);
nand (n836,n837,n2794);
nand (n837,n838,n2368);
nor (n838,n839,n2336);
nor (n839,n840,n1809);
nor (n840,n841,n1794);
nor (n841,n842,n1515);
nand (n842,n843,n1298);
nor (n843,n844,n1197);
nor (n844,n845,n1107);
nand (n845,n846,n1022,n1106);
nand (n846,n847,n924);
xor (n847,n848,n900);
xor (n848,n849,n874);
xor (n849,n850,n862);
xor (n850,n851,n856);
xor (n851,n852,n22);
or (n852,n853,n854);
and (n853,n670,n15);
and (n854,n855,n20);
xor (n856,n857,n33);
or (n857,n858,n860);
and (n858,n859,n27);
and (n860,n861,n31);
xor (n862,n863,n867);
xor (n863,n864,n563);
or (n864,n865,n866);
and (n865,n41,n686);
and (n866,n50,n690);
xnor (n867,n868,n688);
nor (n868,n869,n873);
and (n869,n37,n870);
and (n870,n871,n688);
not (n871,n872);
and (n873,n30,n872);
nand (n874,n875,n885,n899);
nand (n875,n876,n880);
xor (n876,n877,n22);
or (n877,n878,n879);
and (n878,n855,n15);
and (n879,n859,n20);
xor (n880,n881,n33);
or (n881,n882,n883);
and (n882,n861,n27);
and (n883,n884,n31);
nand (n885,n886,n880);
xor (n886,n887,n896);
xor (n887,n888,n892);
xor (n888,n889,n563);
or (n889,n890,n891);
and (n890,n50,n686);
and (n891,n54,n690);
xor (n892,n893,n187);
or (n893,n894,n895);
and (n894,n90,n324);
and (n895,n177,n328);
xnor (n896,n897,n44);
nand (n897,n898,n38);
nand (n899,n876,n886);
xor (n900,n901,n910);
xor (n901,n902,n906);
xor (n902,n903,n44);
or (n903,n904,n905);
and (n904,n884,n38);
and (n905,n898,n42);
nand (n906,n907,n908,n909);
nand (n907,n888,n892);
nand (n908,n896,n892);
nand (n909,n888,n896);
xor (n910,n911,n920);
xor (n911,n912,n916);
xor (n912,n913,n187);
or (n913,n914,n915);
and (n914,n65,n324);
and (n915,n90,n328);
xor (n916,n917,n326);
or (n917,n918,n919);
and (n918,n54,n561);
and (n919,n61,n565);
xor (n920,n921,n105);
or (n921,n922,n923);
and (n922,n177,n185);
and (n923,n223,n189);
nand (n924,n925,n979,n1021);
nand (n925,n926,n928);
xor (n926,n927,n886);
xor (n927,n876,n880);
xor (n928,n929,n968);
xor (n929,n930,n946);
nand (n930,n931,n940,n945);
nand (n931,n932,n936);
xor (n932,n933,n187);
or (n933,n934,n935);
and (n934,n177,n324);
and (n935,n223,n328);
xor (n936,n937,n326);
or (n937,n938,n939);
and (n938,n65,n561);
and (n939,n90,n565);
nand (n940,n941,n936);
xor (n941,n942,n105);
or (n942,n943,n944);
and (n943,n295,n185);
and (n944,n530,n189);
nand (n945,n932,n941);
nand (n946,n947,n962,n967);
nand (n947,n948,n957);
xor (n948,n949,n953);
xnor (n949,n950,n688);
nor (n950,n951,n952);
and (n951,n50,n870);
and (n952,n41,n872);
xor (n953,n954,n563);
or (n954,n955,n956);
and (n955,n54,n686);
and (n956,n61,n690);
and (n957,n958,n33);
xnor (n958,n959,n688);
nor (n959,n960,n961);
and (n960,n54,n870);
and (n961,n50,n872);
nand (n962,n963,n957);
xor (n963,n964,n76);
or (n964,n965,n966);
and (n965,n534,n103);
and (n966,n536,n107);
nand (n967,n948,n963);
xor (n968,n969,n975);
xor (n969,n970,n974);
xor (n970,n971,n76);
or (n971,n972,n973);
and (n972,n530,n103);
and (n973,n534,n107);
and (n974,n949,n953);
xor (n975,n976,n17);
or (n976,n977,n978);
and (n977,n536,n74);
and (n978,n670,n78);
nand (n979,n980,n928);
nand (n980,n981,n1005,n1020);
nand (n981,n982,n1003);
nand (n982,n983,n997,n1002);
nand (n983,n984,n993);
and (n984,n985,n989);
xnor (n985,n986,n688);
nor (n986,n987,n988);
and (n987,n61,n870);
and (n988,n54,n872);
xor (n989,n990,n563);
or (n990,n991,n992);
and (n991,n65,n686);
and (n992,n90,n690);
xor (n993,n994,n76);
or (n994,n995,n996);
and (n995,n536,n103);
and (n996,n670,n107);
nand (n997,n998,n993);
xor (n998,n999,n17);
or (n999,n1000,n1001);
and (n1000,n855,n74);
and (n1001,n859,n78);
nand (n1002,n984,n998);
xor (n1003,n1004,n963);
xor (n1004,n948,n957);
nand (n1005,n1006,n1003);
xor (n1006,n1007,n1016);
xor (n1007,n1008,n1012);
xor (n1008,n1009,n17);
or (n1009,n1010,n1011);
and (n1010,n670,n74);
and (n1011,n855,n78);
xor (n1012,n1013,n22);
or (n1013,n1014,n1015);
and (n1014,n859,n15);
and (n1015,n861,n20);
xor (n1016,n1017,n33);
or (n1017,n1018,n1019);
and (n1018,n884,n27);
and (n1019,n898,n31);
nand (n1020,n982,n1006);
nand (n1021,n926,n980);
nand (n1022,n1023,n924);
xor (n1023,n1024,n1063);
xor (n1024,n1025,n1029);
nand (n1025,n1026,n1027,n1028);
nand (n1026,n930,n946);
nand (n1027,n968,n946);
nand (n1028,n930,n968);
xor (n1029,n1030,n1052);
xor (n1030,n1031,n1048);
nand (n1031,n1032,n1042,n1047);
nand (n1032,n1033,n1037);
xor (n1033,n1034,n326);
or (n1034,n1035,n1036);
and (n1035,n61,n561);
and (n1036,n65,n565);
xor (n1037,n1038,n44);
xnor (n1038,n1039,n688);
nor (n1039,n1040,n1041);
and (n1040,n41,n870);
and (n1041,n37,n872);
nand (n1042,n1043,n1037);
xor (n1043,n1044,n105);
or (n1044,n1045,n1046);
and (n1045,n223,n185);
and (n1046,n295,n189);
nand (n1047,n1033,n1043);
nand (n1048,n1049,n1050,n1051);
nand (n1049,n970,n974);
nand (n1050,n975,n974);
nand (n1051,n970,n975);
xor (n1052,n1053,n1059);
xor (n1053,n1054,n1055);
and (n1054,n1038,n44);
xor (n1055,n1056,n76);
or (n1056,n1057,n1058);
and (n1057,n295,n103);
and (n1058,n530,n107);
xor (n1059,n1060,n17);
or (n1060,n1061,n1062);
and (n1061,n534,n74);
and (n1062,n536,n78);
nand (n1063,n1064,n1071,n1105);
nand (n1064,n1065,n1069);
nand (n1065,n1066,n1067,n1068);
nand (n1066,n1008,n1012);
nand (n1067,n1016,n1012);
nand (n1068,n1008,n1016);
xor (n1069,n1070,n1043);
xor (n1070,n1033,n1037);
nand (n1071,n1072,n1069);
nand (n1072,n1073,n1090,n1104);
nand (n1073,n1074,n1088);
nand (n1074,n1075,n1084,n1087);
nand (n1075,n1076,n1080);
xor (n1076,n1077,n563);
or (n1077,n1078,n1079);
and (n1078,n61,n686);
and (n1079,n65,n690);
xor (n1080,n1081,n187);
or (n1081,n1082,n1083);
and (n1082,n223,n324);
and (n1083,n295,n328);
nand (n1084,n1085,n1080);
xnor (n1085,n1086,n33);
nand (n1086,n898,n27);
nand (n1087,n1076,n1085);
xor (n1088,n1089,n941);
xor (n1089,n932,n936);
nand (n1090,n1091,n1088);
nand (n1091,n1092,n1098,n1103);
nand (n1092,n1093,n1097);
xor (n1093,n1094,n326);
or (n1094,n1095,n1096);
and (n1095,n90,n561);
and (n1096,n177,n565);
xor (n1097,n958,n33);
nand (n1098,n1099,n1097);
xor (n1099,n1100,n105);
or (n1100,n1101,n1102);
and (n1101,n530,n185);
and (n1102,n534,n189);
nand (n1103,n1093,n1099);
nand (n1104,n1074,n1091);
nand (n1105,n1065,n1072);
nand (n1106,n847,n1023);
xor (n1107,n1108,n1193);
xor (n1108,n1109,n1130);
xor (n1109,n1110,n1126);
xor (n1110,n1111,n1122);
xor (n1111,n1112,n1118);
xor (n1112,n1113,n1117);
xor (n1113,n1114,n33);
or (n1114,n1115,n1116);
and (n1115,n855,n27);
and (n1116,n859,n31);
and (n1117,n863,n867);
xor (n1118,n1119,n44);
or (n1119,n1120,n1121);
and (n1120,n861,n38);
and (n1121,n884,n42);
nand (n1122,n1123,n1124,n1125);
nand (n1123,n902,n906);
nand (n1124,n910,n906);
nand (n1125,n902,n910);
nand (n1126,n1127,n1128,n1129);
nand (n1127,n1031,n1048);
nand (n1128,n1052,n1048);
nand (n1129,n1031,n1052);
xor (n1130,n1131,n1189);
xor (n1131,n1132,n1156);
xor (n1132,n1133,n1152);
xor (n1133,n1134,n1138);
nand (n1134,n1135,n1136,n1137);
nand (n1135,n1054,n1055);
nand (n1136,n1059,n1055);
nand (n1137,n1054,n1059);
xor (n1138,n1139,n1148);
xor (n1139,n1140,n1144);
xnor (n1140,n1141,n688);
nor (n1141,n1142,n1143);
and (n1142,n30,n870);
and (n1143,n26,n872);
xor (n1144,n1145,n187);
or (n1145,n1146,n1147);
and (n1146,n61,n324);
and (n1147,n65,n328);
xor (n1148,n1149,n326);
or (n1149,n1150,n1151);
and (n1150,n50,n561);
and (n1151,n54,n565);
nand (n1152,n1153,n1154,n1155);
nand (n1153,n912,n916);
nand (n1154,n920,n916);
nand (n1155,n912,n920);
xor (n1156,n1157,n1175);
xor (n1157,n1158,n1162);
nand (n1158,n1159,n1160,n1161);
nand (n1159,n851,n856);
nand (n1160,n862,n856);
nand (n1161,n851,n862);
xor (n1162,n1163,n1173);
xor (n1163,n1164,n1168);
xor (n1164,n1165,n105);
or (n1165,n1166,n1167);
and (n1166,n90,n185);
and (n1167,n177,n189);
xor (n1168,n57,n1169);
xor (n1169,n1170,n563);
or (n1170,n1171,n1172);
and (n1171,n37,n686);
and (n1172,n41,n690);
xnor (n1173,n1174,n57);
nand (n1174,n898,n51);
xor (n1175,n1176,n1185);
xor (n1176,n1177,n1181);
xor (n1177,n1178,n76);
or (n1178,n1179,n1180);
and (n1179,n223,n103);
and (n1180,n295,n107);
xor (n1181,n1182,n17);
or (n1182,n1183,n1184);
and (n1183,n530,n74);
and (n1184,n534,n78);
xor (n1185,n1186,n22);
or (n1186,n1187,n1188);
and (n1187,n536,n15);
and (n1188,n670,n20);
nand (n1189,n1190,n1191,n1192);
nand (n1190,n849,n874);
nand (n1191,n900,n874);
nand (n1192,n849,n900);
nand (n1193,n1194,n1195,n1196);
nand (n1194,n1025,n1029);
nand (n1195,n1063,n1029);
nand (n1196,n1025,n1063);
nor (n1197,n1198,n1202);
nand (n1198,n1199,n1200,n1201);
nand (n1199,n1109,n1130);
nand (n1200,n1193,n1130);
nand (n1201,n1109,n1193);
xor (n1202,n1203,n1212);
xor (n1203,n1204,n1208);
nand (n1204,n1205,n1206,n1207);
nand (n1205,n1111,n1122);
nand (n1206,n1126,n1122);
nand (n1207,n1111,n1126);
nand (n1208,n1209,n1210,n1211);
nand (n1209,n1132,n1156);
nand (n1210,n1189,n1156);
nand (n1211,n1132,n1189);
xor (n1212,n1213,n1274);
xor (n1213,n1214,n1245);
xor (n1214,n1215,n1234);
xor (n1215,n1216,n1230);
xor (n1216,n1217,n1226);
xor (n1217,n1218,n1222);
xor (n1218,n1219,n187);
or (n1219,n1220,n1221);
and (n1220,n54,n324);
and (n1221,n61,n328);
xor (n1222,n1223,n326);
or (n1223,n1224,n1225);
and (n1224,n41,n561);
and (n1225,n50,n565);
xor (n1226,n1227,n105);
or (n1227,n1228,n1229);
and (n1228,n65,n185);
and (n1229,n90,n189);
nand (n1230,n1231,n1232,n1233);
nand (n1231,n1164,n1168);
nand (n1232,n1173,n1168);
nand (n1233,n1164,n1173);
xor (n1234,n1235,n1241);
xor (n1235,n1236,n1240);
xor (n1236,n1237,n76);
or (n1237,n1238,n1239);
and (n1238,n177,n103);
and (n1239,n223,n107);
and (n1240,n57,n1169);
xor (n1241,n1242,n17);
or (n1242,n1243,n1244);
and (n1243,n295,n74);
and (n1244,n530,n78);
xor (n1245,n1246,n1270);
xor (n1246,n1247,n1251);
nand (n1247,n1248,n1249,n1250);
nand (n1248,n1177,n1181);
nand (n1249,n1185,n1181);
nand (n1250,n1177,n1185);
xor (n1251,n1252,n1261);
xor (n1252,n1253,n1257);
xor (n1253,n1254,n22);
or (n1254,n1255,n1256);
and (n1255,n534,n15);
and (n1256,n536,n20);
xor (n1257,n1258,n33);
or (n1258,n1259,n1260);
and (n1259,n670,n27);
and (n1260,n855,n31);
xor (n1261,n1262,n1266);
xnor (n1262,n1263,n688);
nor (n1263,n1264,n1265);
and (n1264,n26,n870);
and (n1265,n19,n872);
xor (n1266,n1267,n563);
or (n1267,n1268,n1269);
and (n1268,n30,n686);
and (n1269,n37,n690);
nand (n1270,n1271,n1272,n1273);
nand (n1271,n1113,n1117);
nand (n1272,n1118,n1117);
nand (n1273,n1113,n1118);
xor (n1274,n1275,n1294);
xor (n1275,n1276,n1290);
xor (n1276,n1277,n1286);
xor (n1277,n1278,n1282);
xor (n1278,n1279,n44);
or (n1279,n1280,n1281);
and (n1280,n859,n38);
and (n1281,n861,n42);
xor (n1282,n1283,n57);
or (n1283,n1284,n1285);
and (n1284,n884,n51);
and (n1285,n898,n55);
nand (n1286,n1287,n1288,n1289);
nand (n1287,n1140,n1144);
nand (n1288,n1148,n1144);
nand (n1289,n1140,n1148);
nand (n1290,n1291,n1292,n1293);
nand (n1291,n1134,n1138);
nand (n1292,n1152,n1138);
nand (n1293,n1134,n1152);
nand (n1294,n1295,n1296,n1297);
nand (n1295,n1158,n1162);
nand (n1296,n1175,n1162);
nand (n1297,n1158,n1175);
nor (n1298,n1299,n1404);
nor (n1299,n1300,n1304);
nand (n1300,n1301,n1302,n1303);
nand (n1301,n1204,n1208);
nand (n1302,n1212,n1208);
nand (n1303,n1204,n1212);
xor (n1304,n1305,n1400);
xor (n1305,n1306,n1340);
xor (n1306,n1307,n1336);
xor (n1307,n1308,n1312);
nand (n1308,n1309,n1310,n1311);
nand (n1309,n1216,n1230);
nand (n1310,n1234,n1230);
nand (n1311,n1216,n1234);
xor (n1312,n1313,n1322);
xor (n1313,n1314,n1318);
xor (n1314,n1315,n57);
or (n1315,n1316,n1317);
and (n1316,n861,n51);
and (n1317,n884,n55);
nand (n1318,n1319,n1320,n1321);
nand (n1319,n1236,n1240);
nand (n1320,n1241,n1240);
nand (n1321,n1236,n1241);
xor (n1322,n1323,n1332);
xor (n1323,n1324,n1328);
xor (n1324,n1325,n187);
or (n1325,n1326,n1327);
and (n1326,n50,n324);
and (n1327,n54,n328);
xnor (n1328,n1329,n688);
nor (n1329,n1330,n1331);
and (n1330,n19,n870);
and (n1331,n14,n872);
xor (n1332,n1333,n326);
or (n1333,n1334,n1335);
and (n1334,n37,n561);
and (n1335,n41,n565);
nand (n1336,n1337,n1338,n1339);
nand (n1337,n1247,n1251);
nand (n1338,n1270,n1251);
nand (n1339,n1247,n1270);
xor (n1340,n1341,n1396);
xor (n1341,n1342,n1364);
xor (n1342,n1343,n1352);
xor (n1343,n1344,n1348);
nand (n1344,n1345,n1346,n1347);
nand (n1345,n1218,n1222);
nand (n1346,n1226,n1222);
nand (n1347,n1218,n1226);
nand (n1348,n1349,n1350,n1351);
nand (n1349,n1253,n1257);
nand (n1350,n1261,n1257);
nand (n1351,n1253,n1261);
xor (n1352,n1353,n1360);
xor (n1353,n1354,n1358);
xor (n1354,n1355,n105);
or (n1355,n1356,n1357);
and (n1356,n61,n185);
and (n1357,n65,n189);
xnor (n1358,n1359,n68);
nand (n1359,n898,n62);
xor (n1360,n1361,n76);
or (n1361,n1362,n1363);
and (n1362,n90,n103);
and (n1363,n177,n107);
xor (n1364,n1365,n1384);
xor (n1365,n1366,n1370);
nand (n1366,n1367,n1368,n1369);
nand (n1367,n1278,n1282);
nand (n1368,n1286,n1282);
nand (n1369,n1278,n1286);
xor (n1370,n1371,n1380);
xor (n1371,n1372,n1376);
xor (n1372,n1373,n17);
or (n1373,n1374,n1375);
and (n1374,n223,n74);
and (n1375,n295,n78);
xor (n1376,n1377,n22);
or (n1377,n1378,n1379);
and (n1378,n530,n15);
and (n1379,n534,n20);
xor (n1380,n1381,n33);
or (n1381,n1382,n1383);
and (n1382,n536,n27);
and (n1383,n670,n31);
xor (n1384,n1385,n1392);
xor (n1385,n1386,n1391);
xor (n1386,n68,n1387);
xor (n1387,n1388,n563);
or (n1388,n1389,n1390);
and (n1389,n26,n686);
and (n1390,n30,n690);
and (n1391,n1262,n1266);
xor (n1392,n1393,n44);
or (n1393,n1394,n1395);
and (n1394,n855,n38);
and (n1395,n859,n42);
nand (n1396,n1397,n1398,n1399);
nand (n1397,n1276,n1290);
nand (n1398,n1294,n1290);
nand (n1399,n1276,n1294);
nand (n1400,n1401,n1402,n1403);
nand (n1401,n1214,n1245);
nand (n1402,n1274,n1245);
nand (n1403,n1214,n1274);
nor (n1404,n1405,n1409);
nand (n1405,n1406,n1407,n1408);
nand (n1406,n1306,n1340);
nand (n1407,n1400,n1340);
nand (n1408,n1306,n1400);
xor (n1409,n1410,n1419);
xor (n1410,n1411,n1415);
nand (n1411,n1412,n1413,n1414);
nand (n1412,n1308,n1312);
nand (n1413,n1336,n1312);
nand (n1414,n1308,n1336);
nand (n1415,n1416,n1417,n1418);
nand (n1416,n1342,n1364);
nand (n1417,n1396,n1364);
nand (n1418,n1342,n1396);
xor (n1419,n1420,n1481);
xor (n1420,n1421,n1445);
xor (n1421,n1422,n1441);
xor (n1422,n1423,n1427);
nand (n1423,n1424,n1425,n1426);
nand (n1424,n1372,n1376);
nand (n1425,n1380,n1376);
nand (n1426,n1372,n1380);
xor (n1427,n1428,n1437);
xor (n1428,n1429,n1433);
xor (n1429,n1430,n76);
or (n1430,n1431,n1432);
and (n1431,n65,n103);
and (n1432,n90,n107);
xor (n1433,n1434,n17);
or (n1434,n1435,n1436);
and (n1435,n177,n74);
and (n1436,n223,n78);
xor (n1437,n1438,n22);
or (n1438,n1439,n1440);
and (n1439,n295,n15);
and (n1440,n530,n20);
nand (n1441,n1442,n1443,n1444);
nand (n1442,n1386,n1391);
nand (n1443,n1392,n1391);
nand (n1444,n1386,n1392);
xor (n1445,n1446,n1467);
xor (n1446,n1447,n1463);
xor (n1447,n1448,n1462);
xor (n1448,n1449,n1453);
xor (n1449,n1450,n33);
or (n1450,n1451,n1452);
and (n1451,n534,n27);
and (n1452,n536,n31);
xor (n1453,n1454,n1458);
xnor (n1454,n1455,n688);
nor (n1455,n1456,n1457);
and (n1456,n14,n870);
and (n1457,n73,n872);
xor (n1458,n1459,n563);
or (n1459,n1460,n1461);
and (n1460,n19,n686);
and (n1461,n26,n690);
and (n1462,n68,n1387);
nand (n1463,n1464,n1465,n1466);
nand (n1464,n1314,n1318);
nand (n1465,n1322,n1318);
nand (n1466,n1314,n1322);
xor (n1467,n1468,n1477);
xor (n1468,n1469,n1473);
xor (n1469,n1470,n44);
or (n1470,n1471,n1472);
and (n1471,n670,n38);
and (n1472,n855,n42);
xor (n1473,n1474,n68);
or (n1474,n1475,n1476);
and (n1475,n884,n62);
and (n1476,n898,n66);
xor (n1477,n1478,n57);
or (n1478,n1479,n1480);
and (n1479,n859,n51);
and (n1480,n861,n55);
xor (n1481,n1482,n1511);
xor (n1482,n1483,n1507);
xor (n1483,n1484,n1503);
xor (n1484,n1485,n1489);
nand (n1485,n1486,n1487,n1488);
nand (n1486,n1324,n1328);
nand (n1487,n1332,n1328);
nand (n1488,n1324,n1332);
xor (n1489,n1490,n1499);
xor (n1490,n1491,n1495);
xor (n1491,n1492,n187);
or (n1492,n1493,n1494);
and (n1493,n41,n324);
and (n1494,n50,n328);
xor (n1495,n1496,n326);
or (n1496,n1497,n1498);
and (n1497,n30,n561);
and (n1498,n37,n565);
xor (n1499,n1500,n105);
or (n1500,n1501,n1502);
and (n1501,n54,n185);
and (n1502,n61,n189);
nand (n1503,n1504,n1505,n1506);
nand (n1504,n1354,n1358);
nand (n1505,n1360,n1358);
nand (n1506,n1354,n1360);
nand (n1507,n1508,n1509,n1510);
nand (n1508,n1344,n1348);
nand (n1509,n1352,n1348);
nand (n1510,n1344,n1352);
nand (n1511,n1512,n1513,n1514);
nand (n1512,n1366,n1370);
nand (n1513,n1384,n1370);
nand (n1514,n1366,n1384);
nor (n1515,n1516,n1788);
nor (n1516,n1517,n1764);
nor (n1517,n1518,n1762);
nor (n1518,n1519,n1737);
nand (n1519,n1520,n1699);
nand (n1520,n1521,n1646,n1698);
nand (n1521,n1522,n1573);
xor (n1522,n1523,n1560);
xor (n1523,n1524,n1545);
nand (n1524,n1525,n1539,n1544);
nand (n1525,n1526,n1535);
and (n1526,n1527,n1531);
xnor (n1527,n1528,n688);
nor (n1528,n1529,n1530);
and (n1529,n90,n870);
and (n1530,n65,n872);
xor (n1531,n1532,n563);
or (n1532,n1533,n1534);
and (n1533,n177,n686);
and (n1534,n223,n690);
xor (n1535,n1536,n76);
or (n1536,n1537,n1538);
and (n1537,n855,n103);
and (n1538,n859,n107);
nand (n1539,n1540,n1535);
xor (n1540,n1541,n17);
or (n1541,n1542,n1543);
and (n1542,n861,n74);
and (n1543,n884,n78);
nand (n1544,n1526,n1540);
xor (n1545,n1546,n1555);
xor (n1546,n1547,n1551);
xor (n1547,n1548,n187);
or (n1548,n1549,n1550);
and (n1549,n295,n324);
and (n1550,n530,n328);
xor (n1551,n1552,n326);
or (n1552,n1553,n1554);
and (n1553,n177,n561);
and (n1554,n223,n565);
and (n1555,n1556,n22);
xnor (n1556,n1557,n688);
nor (n1557,n1558,n1559);
and (n1558,n65,n870);
and (n1559,n61,n872);
nand (n1560,n1561,n1567,n1572);
nand (n1561,n1562,n1566);
xor (n1562,n1563,n326);
or (n1563,n1564,n1565);
and (n1564,n223,n561);
and (n1565,n295,n565);
xor (n1566,n1556,n22);
nand (n1567,n1568,n1566);
xor (n1568,n1569,n105);
or (n1569,n1570,n1571);
and (n1570,n536,n185);
and (n1571,n670,n189);
nand (n1572,n1562,n1568);
xor (n1573,n1574,n1610);
xor (n1574,n1575,n1586);
xor (n1575,n1576,n1582);
xor (n1576,n1577,n1581);
xor (n1577,n1578,n105);
or (n1578,n1579,n1580);
and (n1579,n534,n185);
and (n1580,n536,n189);
xor (n1581,n985,n989);
xor (n1582,n1583,n76);
or (n1583,n1584,n1585);
and (n1584,n670,n103);
and (n1585,n855,n107);
xor (n1586,n1587,n1596);
xor (n1587,n1588,n1592);
xor (n1588,n1589,n17);
or (n1589,n1590,n1591);
and (n1590,n859,n74);
and (n1591,n861,n78);
xor (n1592,n1593,n22);
or (n1593,n1594,n1595);
and (n1594,n884,n15);
and (n1595,n898,n20);
nand (n1596,n1597,n1604,n1609);
nand (n1597,n1598,n1602);
xor (n1598,n1599,n563);
or (n1599,n1600,n1601);
and (n1600,n90,n686);
and (n1601,n177,n690);
xnor (n1602,n1603,n22);
nand (n1603,n898,n15);
nand (n1604,n1605,n1602);
xor (n1605,n1606,n187);
or (n1606,n1607,n1608);
and (n1607,n530,n324);
and (n1608,n534,n328);
nand (n1609,n1598,n1605);
nand (n1610,n1611,n1631,n1645);
nand (n1611,n1612,n1614);
xor (n1612,n1613,n1605);
xor (n1613,n1598,n1602);
nand (n1614,n1615,n1624,n1630);
nand (n1615,n1616,n1620);
xor (n1616,n1617,n187);
or (n1617,n1618,n1619);
and (n1618,n534,n324);
and (n1619,n536,n328);
xor (n1620,n1621,n326);
or (n1621,n1622,n1623);
and (n1622,n295,n561);
and (n1623,n530,n565);
nand (n1624,n1625,n1620);
and (n1625,n1626,n17);
xnor (n1626,n1627,n688);
nor (n1627,n1628,n1629);
and (n1628,n177,n870);
and (n1629,n90,n872);
nand (n1630,n1616,n1625);
nand (n1631,n1632,n1614);
nand (n1632,n1633,n1639,n1644);
nand (n1633,n1634,n1638);
xor (n1634,n1635,n105);
or (n1635,n1636,n1637);
and (n1636,n670,n185);
and (n1637,n855,n189);
xor (n1638,n1527,n1531);
nand (n1639,n1640,n1638);
xor (n1640,n1641,n76);
or (n1641,n1642,n1643);
and (n1642,n859,n103);
and (n1643,n861,n107);
nand (n1644,n1634,n1640);
nand (n1645,n1612,n1632);
nand (n1646,n1647,n1573);
nand (n1647,n1648,n1653,n1697);
nand (n1648,n1649,n1651);
xor (n1649,n1650,n1540);
xor (n1650,n1526,n1535);
xor (n1651,n1652,n1568);
xor (n1652,n1562,n1566);
nand (n1653,n1654,n1651);
nand (n1654,n1655,n1674,n1696);
nand (n1655,n1656,n1660);
xor (n1656,n1657,n17);
or (n1657,n1658,n1659);
and (n1658,n884,n74);
and (n1659,n898,n78);
nand (n1660,n1661,n1668,n1673);
nand (n1661,n1662,n1666);
xor (n1662,n1663,n563);
or (n1663,n1664,n1665);
and (n1664,n223,n686);
and (n1665,n295,n690);
xnor (n1666,n1667,n17);
nand (n1667,n898,n74);
nand (n1668,n1669,n1666);
xor (n1669,n1670,n187);
or (n1670,n1671,n1672);
and (n1671,n536,n324);
and (n1672,n670,n328);
nand (n1673,n1662,n1669);
nand (n1674,n1675,n1660);
nand (n1675,n1676,n1690,n1695);
nand (n1676,n1677,n1681);
xor (n1677,n1678,n326);
or (n1678,n1679,n1680);
and (n1679,n530,n561);
and (n1680,n534,n565);
and (n1681,n1682,n1686);
xnor (n1682,n1683,n688);
nor (n1683,n1684,n1685);
and (n1684,n223,n870);
and (n1685,n177,n872);
xor (n1686,n1687,n563);
or (n1687,n1688,n1689);
and (n1688,n295,n686);
and (n1689,n530,n690);
nand (n1690,n1691,n1681);
xor (n1691,n1692,n105);
or (n1692,n1693,n1694);
and (n1693,n855,n185);
and (n1694,n859,n189);
nand (n1695,n1677,n1691);
nand (n1696,n1656,n1675);
nand (n1697,n1649,n1654);
nand (n1698,n1522,n1647);
xor (n1699,n1700,n1715);
xor (n1700,n1701,n1711);
xor (n1701,n1702,n1709);
xor (n1702,n1703,n1707);
nand (n1703,n1704,n1705,n1706);
nand (n1704,n1547,n1551);
nand (n1705,n1555,n1551);
nand (n1706,n1547,n1555);
xor (n1707,n1708,n998);
xor (n1708,n984,n993);
xor (n1709,n1710,n1099);
xor (n1710,n1093,n1097);
nand (n1711,n1712,n1713,n1714);
nand (n1712,n1575,n1586);
nand (n1713,n1610,n1586);
nand (n1714,n1575,n1610);
xor (n1715,n1716,n1725);
xor (n1716,n1717,n1721);
nand (n1717,n1718,n1719,n1720);
nand (n1718,n1588,n1592);
nand (n1719,n1596,n1592);
nand (n1720,n1588,n1596);
nand (n1721,n1722,n1723,n1724);
nand (n1722,n1524,n1545);
nand (n1723,n1560,n1545);
nand (n1724,n1524,n1560);
xor (n1725,n1726,n1735);
xor (n1726,n1727,n1731);
xor (n1727,n1728,n22);
or (n1728,n1729,n1730);
and (n1729,n861,n15);
and (n1730,n884,n20);
nand (n1731,n1732,n1733,n1734);
nand (n1732,n1577,n1581);
nand (n1733,n1582,n1581);
nand (n1734,n1577,n1582);
xor (n1735,n1736,n1085);
xor (n1736,n1076,n1080);
nor (n1737,n1738,n1742);
nand (n1738,n1739,n1740,n1741);
nand (n1739,n1701,n1711);
nand (n1740,n1715,n1711);
nand (n1741,n1701,n1715);
xor (n1742,n1743,n1750);
xor (n1743,n1744,n1746);
xor (n1744,n1745,n1006);
xor (n1745,n982,n1003);
nand (n1746,n1747,n1748,n1749);
nand (n1747,n1717,n1721);
nand (n1748,n1725,n1721);
nand (n1749,n1717,n1725);
xor (n1750,n1751,n1760);
xor (n1751,n1752,n1756);
nand (n1752,n1753,n1754,n1755);
nand (n1753,n1727,n1731);
nand (n1754,n1735,n1731);
nand (n1755,n1727,n1735);
nand (n1756,n1757,n1758,n1759);
nand (n1757,n1703,n1707);
nand (n1758,n1709,n1707);
nand (n1759,n1703,n1709);
xor (n1760,n1761,n1091);
xor (n1761,n1074,n1088);
not (n1762,n1763);
nand (n1763,n1738,n1742);
not (n1764,n1765);
nor (n1765,n1766,n1781);
nor (n1766,n1767,n1771);
nand (n1767,n1768,n1769,n1770);
nand (n1768,n1744,n1746);
nand (n1769,n1750,n1746);
nand (n1770,n1744,n1750);
xor (n1771,n1772,n1779);
xor (n1772,n1773,n1775);
xor (n1773,n1774,n1072);
xor (n1774,n1065,n1069);
nand (n1775,n1776,n1777,n1778);
nand (n1776,n1752,n1756);
nand (n1777,n1760,n1756);
nand (n1778,n1752,n1760);
xor (n1779,n1780,n980);
xor (n1780,n926,n928);
nor (n1781,n1782,n1786);
nand (n1782,n1783,n1784,n1785);
nand (n1783,n1773,n1775);
nand (n1784,n1779,n1775);
nand (n1785,n1773,n1779);
xor (n1786,n1787,n1023);
xor (n1787,n847,n924);
not (n1788,n1789);
nor (n1789,n1790,n1792);
nor (n1790,n1791,n1781);
nand (n1791,n1767,n1771);
not (n1792,n1793);
nand (n1793,n1782,n1786);
not (n1794,n1795);
nor (n1795,n1796,n1803);
nor (n1796,n1797,n1802);
nor (n1797,n1798,n1800);
nor (n1798,n1799,n1197);
nand (n1799,n845,n1107);
not (n1800,n1801);
nand (n1801,n1198,n1202);
not (n1802,n1298);
not (n1803,n1804);
nor (n1804,n1805,n1807);
nor (n1805,n1806,n1404);
nand (n1806,n1300,n1304);
not (n1807,n1808);
nand (n1808,n1405,n1409);
not (n1809,n1810);
nor (n1810,n1811,n2226);
nand (n1811,n1812,n2039);
nor (n1812,n1813,n1925);
nor (n1813,n1814,n1818);
nand (n1814,n1815,n1816,n1817);
nand (n1815,n1411,n1415);
nand (n1816,n1419,n1415);
nand (n1817,n1411,n1419);
xor (n1818,n1819,n1921);
xor (n1819,n1820,n1853);
xor (n1820,n1821,n1849);
xor (n1821,n1822,n1845);
xor (n1822,n1823,n1841);
xor (n1823,n1824,n1837);
xor (n1824,n1825,n1834);
xor (n1825,n1826,n1830);
xor (n1826,n1827,n563);
or (n1827,n1828,n1829);
and (n1828,n14,n686);
and (n1829,n19,n690);
xor (n1830,n1831,n326);
or (n1831,n1832,n1833);
and (n1832,n26,n561);
and (n1833,n30,n565);
xnor (n1834,n1835,n688);
nor (n1835,n1836,n1457);
and (n1836,n73,n870);
nand (n1837,n1838,n1839,n1840);
nand (n1838,n1429,n1433);
nand (n1839,n1437,n1433);
nand (n1840,n1429,n1437);
nand (n1841,n1842,n1843,n1844);
nand (n1842,n1449,n1453);
nand (n1843,n1462,n1453);
nand (n1844,n1449,n1462);
nand (n1845,n1846,n1847,n1848);
nand (n1846,n1423,n1427);
nand (n1847,n1441,n1427);
nand (n1848,n1423,n1441);
nand (n1849,n1850,n1851,n1852);
nand (n1850,n1447,n1463);
nand (n1851,n1467,n1463);
nand (n1852,n1447,n1467);
xor (n1853,n1854,n1917);
xor (n1854,n1855,n1893);
xor (n1855,n1856,n1878);
xor (n1856,n1857,n1871);
xor (n1857,n1858,n1867);
xor (n1858,n1859,n1863);
xor (n1859,n1860,n105);
or (n1860,n1861,n1862);
and (n1861,n50,n185);
and (n1862,n54,n189);
xor (n1863,n1864,n76);
or (n1864,n1865,n1866);
and (n1865,n61,n103);
and (n1866,n65,n107);
xor (n1867,n1868,n17);
or (n1868,n1869,n1870);
and (n1869,n90,n74);
and (n1870,n177,n78);
xor (n1871,n1872,n1874);
xor (n1872,n68,n1873);
and (n1873,n1454,n1458);
xor (n1874,n1875,n44);
or (n1875,n1876,n1877);
and (n1876,n536,n38);
and (n1877,n670,n42);
xor (n1878,n1879,n1888);
xor (n1879,n1880,n1884);
xor (n1880,n1881,n22);
or (n1881,n1882,n1883);
and (n1882,n223,n15);
and (n1883,n295,n20);
xor (n1884,n1885,n33);
or (n1885,n1886,n1887);
and (n1886,n530,n27);
and (n1887,n534,n31);
xor (n1888,n68,n1889);
xor (n1889,n1890,n187);
or (n1890,n1891,n1892);
and (n1891,n37,n324);
and (n1892,n41,n328);
xor (n1893,n1894,n1903);
xor (n1894,n1895,n1899);
nand (n1895,n1896,n1897,n1898);
nand (n1896,n1469,n1473);
nand (n1897,n1477,n1473);
nand (n1898,n1469,n1477);
nand (n1899,n1900,n1901,n1902);
nand (n1900,n1485,n1489);
nand (n1901,n1503,n1489);
nand (n1902,n1485,n1503);
xor (n1903,n1904,n1913);
xor (n1904,n1905,n1909);
xor (n1905,n1906,n57);
or (n1906,n1907,n1908);
and (n1907,n855,n51);
and (n1908,n859,n55);
xor (n1909,n1910,n68);
or (n1910,n1911,n1912);
and (n1911,n861,n62);
and (n1912,n884,n66);
nand (n1913,n1914,n1915,n1916);
nand (n1914,n1491,n1495);
nand (n1915,n1499,n1495);
nand (n1916,n1491,n1499);
nand (n1917,n1918,n1919,n1920);
nand (n1918,n1483,n1507);
nand (n1919,n1511,n1507);
nand (n1920,n1483,n1511);
nand (n1921,n1922,n1923,n1924);
nand (n1922,n1421,n1445);
nand (n1923,n1481,n1445);
nand (n1924,n1421,n1481);
nor (n1925,n1926,n1930);
nand (n1926,n1927,n1928,n1929);
nand (n1927,n1820,n1853);
nand (n1928,n1921,n1853);
nand (n1929,n1820,n1921);
xor (n1930,n1931,n1940);
xor (n1931,n1932,n1936);
nand (n1932,n1933,n1934,n1935);
nand (n1933,n1822,n1845);
nand (n1934,n1849,n1845);
nand (n1935,n1822,n1849);
nand (n1936,n1937,n1938,n1939);
nand (n1937,n1855,n1893);
nand (n1938,n1917,n1893);
nand (n1939,n1855,n1917);
xor (n1940,n1941,n1998);
xor (n1941,n1942,n1973);
xor (n1942,n1943,n1959);
xor (n1943,n1944,n1948);
nand (n1944,n1945,n1946,n1947);
nand (n1945,n68,n1873);
nand (n1946,n1874,n1873);
nand (n1947,n68,n1874);
xor (n1948,n1949,n1955);
xor (n1949,n1950,n1954);
xor (n1950,n1951,n33);
or (n1951,n1952,n1953);
and (n1952,n295,n27);
and (n1953,n530,n31);
and (n1954,n68,n1889);
xor (n1955,n1956,n44);
or (n1956,n1957,n1958);
and (n1957,n534,n38);
and (n1958,n536,n42);
xor (n1959,n1960,n1969);
xor (n1960,n1961,n1965);
xor (n1961,n1962,n57);
or (n1962,n1963,n1964);
and (n1963,n670,n51);
and (n1964,n855,n55);
xor (n1965,n1966,n68);
or (n1966,n1967,n1968);
and (n1967,n859,n62);
and (n1968,n861,n66);
nand (n1969,n1970,n1971,n1972);
nand (n1970,n1826,n1830);
nand (n1971,n1834,n1830);
nand (n1972,n1826,n1834);
xor (n1973,n1974,n1983);
xor (n1974,n1975,n1979);
nand (n1975,n1976,n1977,n1978);
nand (n1976,n1905,n1909);
nand (n1977,n1913,n1909);
nand (n1978,n1905,n1913);
nand (n1979,n1980,n1981,n1982);
nand (n1980,n1824,n1837);
nand (n1981,n1841,n1837);
nand (n1982,n1824,n1841);
xor (n1983,n1984,n68);
xor (n1984,n1985,n1989);
nand (n1985,n1986,n1987,n1988);
nand (n1986,n1859,n1863);
nand (n1987,n1867,n1863);
nand (n1988,n1859,n1867);
xor (n1989,n1990,n1995);
not (n1990,n1991);
xor (n1991,n1992,n187);
or (n1992,n1993,n1994);
and (n1993,n30,n324);
and (n1994,n37,n328);
xor (n1995,n1996,n563);
or (n1996,n685,n1997);
and (n1997,n14,n690);
xor (n1998,n1999,n2035);
xor (n1999,n2000,n2004);
nand (n2000,n2001,n2002,n2003);
nand (n2001,n1857,n1871);
nand (n2002,n1878,n1871);
nand (n2003,n1857,n1878);
xor (n2004,n2005,n2024);
xor (n2005,n2006,n2010);
nand (n2006,n2007,n2008,n2009);
nand (n2007,n1880,n1884);
nand (n2008,n1888,n1884);
nand (n2009,n1880,n1888);
xor (n2010,n2011,n2020);
xor (n2011,n2012,n2016);
xor (n2012,n2013,n76);
or (n2013,n2014,n2015);
and (n2014,n54,n103);
and (n2015,n61,n107);
xor (n2016,n2017,n17);
or (n2017,n2018,n2019);
and (n2018,n65,n74);
and (n2019,n90,n78);
xor (n2020,n2021,n22);
or (n2021,n2022,n2023);
and (n2022,n177,n15);
and (n2023,n223,n20);
xor (n2024,n2025,n2031);
xor (n2025,n2026,n2030);
xor (n2026,n2027,n326);
or (n2027,n2028,n2029);
and (n2028,n19,n561);
and (n2029,n26,n565);
not (n2030,n1834);
xor (n2031,n2032,n105);
or (n2032,n2033,n2034);
and (n2033,n41,n185);
and (n2034,n50,n189);
nand (n2035,n2036,n2037,n2038);
nand (n2036,n1895,n1899);
nand (n2037,n1903,n1899);
nand (n2038,n1895,n1903);
nor (n2039,n2040,n2147);
nor (n2040,n2041,n2045);
nand (n2041,n2042,n2043,n2044);
nand (n2042,n1932,n1936);
nand (n2043,n1940,n1936);
nand (n2044,n1932,n1940);
xor (n2045,n2046,n2143);
xor (n2046,n2047,n2087);
xor (n2047,n2048,n2083);
xor (n2048,n2049,n2079);
xor (n2049,n2050,n2075);
xor (n2050,n2051,n2065);
xor (n2051,n2052,n2061);
xor (n2052,n2053,n2057);
xor (n2053,n2054,n76);
or (n2054,n2055,n2056);
and (n2055,n50,n103);
and (n2056,n54,n107);
xor (n2057,n2058,n17);
or (n2058,n2059,n2060);
and (n2059,n61,n74);
and (n2060,n65,n78);
xor (n2061,n2062,n33);
or (n2062,n2063,n2064);
and (n2063,n223,n27);
and (n2064,n295,n31);
xor (n2065,n2066,n2071);
xor (n2066,n2067,n683);
xor (n2067,n2068,n187);
or (n2068,n2069,n2070);
and (n2069,n26,n324);
and (n2070,n30,n328);
xor (n2071,n2072,n105);
or (n2072,n2073,n2074);
and (n2073,n37,n185);
and (n2074,n41,n189);
nand (n2075,n2076,n2077,n2078);
nand (n2076,n1950,n1954);
nand (n2077,n1955,n1954);
nand (n2078,n1950,n1955);
nand (n2079,n2080,n2081,n2082);
nand (n2080,n1944,n1948);
nand (n2081,n1959,n1948);
nand (n2082,n1944,n1959);
nand (n2083,n2084,n2085,n2086);
nand (n2084,n1975,n1979);
nand (n2085,n1983,n1979);
nand (n2086,n1975,n1983);
xor (n2087,n2088,n2139);
xor (n2088,n2089,n2110);
xor (n2089,n2090,n2106);
xor (n2090,n2091,n2102);
xor (n2091,n2092,n2098);
xor (n2092,n2093,n2094);
not (n2093,n724);
xor (n2094,n2095,n22);
or (n2095,n2096,n2097);
and (n2096,n90,n15);
and (n2097,n177,n20);
xor (n2098,n2099,n44);
or (n2099,n2100,n2101);
and (n2100,n530,n38);
and (n2101,n534,n42);
nand (n2102,n2103,n2104,n2105);
nand (n2103,n1961,n1965);
nand (n2104,n1969,n1965);
nand (n2105,n1961,n1969);
nand (n2106,n2107,n2108,n2109);
nand (n2107,n1985,n1989);
nand (n2108,n68,n1989);
nand (n2109,n1985,n68);
xor (n2110,n2111,n2135);
xor (n2111,n2112,n2125);
xor (n2112,n2113,n2122);
xor (n2113,n2114,n2118);
xor (n2114,n2115,n57);
or (n2115,n2116,n2117);
and (n2116,n536,n51);
and (n2117,n670,n55);
xor (n2118,n2119,n68);
or (n2119,n2120,n2121);
and (n2120,n855,n62);
and (n2121,n859,n66);
nand (n2122,n1990,n2123,n2124);
nand (n2123,n1995,n1991);
not (n2124,n1995);
xor (n2125,n2126,n2131);
xor (n2126,n68,n2127);
nand (n2127,n2128,n2129,n2130);
nand (n2128,n2026,n2030);
nand (n2129,n2031,n2030);
nand (n2130,n2026,n2031);
nand (n2131,n2132,n2133,n2134);
nand (n2132,n2012,n2016);
nand (n2133,n2020,n2016);
nand (n2134,n2012,n2020);
nand (n2135,n2136,n2137,n2138);
nand (n2136,n2006,n2010);
nand (n2137,n2024,n2010);
nand (n2138,n2006,n2024);
nand (n2139,n2140,n2141,n2142);
nand (n2140,n2000,n2004);
nand (n2141,n2035,n2004);
nand (n2142,n2000,n2035);
nand (n2143,n2144,n2145,n2146);
nand (n2144,n1942,n1973);
nand (n2145,n1998,n1973);
nand (n2146,n1942,n1998);
nor (n2147,n2148,n2152);
nand (n2148,n2149,n2150,n2151);
nand (n2149,n2047,n2087);
nand (n2150,n2143,n2087);
nand (n2151,n2047,n2143);
xor (n2152,n2153,n2162);
xor (n2153,n2154,n2158);
nand (n2154,n2155,n2156,n2157);
nand (n2155,n2049,n2079);
nand (n2156,n2083,n2079);
nand (n2157,n2049,n2083);
nand (n2158,n2159,n2160,n2161);
nand (n2159,n2089,n2110);
nand (n2160,n2139,n2110);
nand (n2161,n2089,n2139);
xor (n2162,n2163,n2194);
xor (n2163,n2164,n2168);
nand (n2164,n2165,n2166,n2167);
nand (n2165,n2112,n2125);
nand (n2166,n2135,n2125);
nand (n2167,n2112,n2135);
xor (n2168,n2169,n2182);
xor (n2169,n2170,n2174);
nand (n2170,n2171,n2172,n2173);
nand (n2171,n68,n2127);
nand (n2172,n2131,n2127);
nand (n2173,n68,n2131);
xor (n2174,n2175,n2178);
xor (n2175,n2176,n68);
xor (n2176,n2177,n682);
xor (n2177,n674,n677);
nand (n2178,n2179,n2180,n2181);
nand (n2179,n2067,n683);
nand (n2180,n2071,n683);
nand (n2181,n2067,n2071);
xor (n2182,n2183,n2190);
xor (n2183,n2184,n2186);
xor (n2184,n2185,n710);
xor (n2185,n701,n705);
nand (n2186,n2187,n2188,n2189);
nand (n2187,n2053,n2057);
nand (n2188,n2061,n2057);
nand (n2189,n2053,n2061);
nand (n2190,n2191,n2192,n2193);
nand (n2191,n2114,n2118);
nand (n2192,n2122,n2118);
nand (n2193,n2114,n2122);
xor (n2194,n2195,n2204);
xor (n2195,n2196,n2200);
nand (n2196,n2197,n2198,n2199);
nand (n2197,n2051,n2065);
nand (n2198,n2075,n2065);
nand (n2199,n2051,n2075);
nand (n2200,n2201,n2202,n2203);
nand (n2201,n2091,n2102);
nand (n2202,n2106,n2102);
nand (n2203,n2091,n2106);
xor (n2204,n2205,n2212);
xor (n2205,n2206,n2210);
nand (n2206,n2207,n2208,n2209);
nand (n2207,n2093,n2094);
nand (n2208,n2098,n2094);
nand (n2209,n2093,n2098);
xor (n2210,n2211,n729);
xor (n2211,n720,n724);
xor (n2212,n2213,n2222);
xor (n2213,n2214,n2218);
xor (n2214,n2215,n44);
or (n2215,n2216,n2217);
and (n2216,n295,n38);
and (n2217,n530,n42);
xor (n2218,n2219,n57);
or (n2219,n2220,n2221);
and (n2220,n534,n51);
and (n2221,n536,n55);
xor (n2222,n2223,n68);
or (n2223,n2224,n2225);
and (n2224,n670,n62);
and (n2225,n855,n66);
nand (n2226,n2227,n2311);
nor (n2227,n2228,n2278);
nor (n2228,n2229,n2233);
nand (n2229,n2230,n2231,n2232);
nand (n2230,n2154,n2158);
nand (n2231,n2162,n2158);
nand (n2232,n2154,n2162);
xor (n2233,n2234,n2274);
xor (n2234,n2235,n2255);
xor (n2235,n2236,n2243);
xor (n2236,n2237,n2239);
xor (n2237,n2238,n718);
xor (n2238,n699,n715);
nand (n2239,n2240,n2241,n2242);
nand (n2240,n2206,n2210);
nand (n2241,n2212,n2210);
nand (n2242,n2206,n2212);
xor (n2243,n2244,n2251);
xor (n2244,n2245,n2249);
nand (n2245,n2246,n2247,n2248);
nand (n2246,n2214,n2218);
nand (n2247,n2222,n2218);
nand (n2248,n2214,n2222);
xor (n2249,n2250,n628);
xor (n2250,n622,n626);
nand (n2251,n2252,n2253,n2254);
nand (n2252,n2176,n68);
nand (n2253,n2178,n68);
nand (n2254,n2176,n2178);
xor (n2255,n2256,n2270);
xor (n2256,n2257,n2261);
nand (n2257,n2258,n2259,n2260);
nand (n2258,n2170,n2174);
nand (n2259,n2182,n2174);
nand (n2260,n2170,n2182);
xor (n2261,n2262,n2266);
xor (n2262,n2263,n2265);
xor (n2263,n2264,n644);
xor (n2264,n635,n639);
xor (n2265,n667,n672);
nand (n2266,n2267,n2268,n2269);
nand (n2267,n2184,n2186);
nand (n2268,n2190,n2186);
nand (n2269,n2184,n2190);
nand (n2270,n2271,n2272,n2273);
nand (n2271,n2196,n2200);
nand (n2272,n2204,n2200);
nand (n2273,n2196,n2204);
nand (n2274,n2275,n2276,n2277);
nand (n2275,n2164,n2168);
nand (n2276,n2194,n2168);
nand (n2277,n2164,n2194);
nor (n2278,n2279,n2283);
nand (n2279,n2280,n2281,n2282);
nand (n2280,n2235,n2255);
nand (n2281,n2274,n2255);
nand (n2282,n2235,n2274);
xor (n2283,n2284,n2307);
xor (n2284,n2285,n2295);
xor (n2285,n2286,n2293);
xor (n2286,n2287,n2289);
xor (n2287,n2288,n615);
xor (n2288,n600,n612);
nand (n2289,n2290,n2291,n2292);
nand (n2290,n2245,n2249);
nand (n2291,n2251,n2249);
nand (n2292,n2245,n2251);
xor (n2293,n2294,n650);
xor (n2294,n620,n633);
xor (n2295,n2296,n2303);
xor (n2296,n2297,n2299);
xor (n2297,n2298,n697);
xor (n2298,n664,n694);
nand (n2299,n2300,n2301,n2302);
nand (n2300,n2263,n2265);
nand (n2301,n2266,n2265);
nand (n2302,n2263,n2266);
nand (n2303,n2304,n2305,n2306);
nand (n2304,n2237,n2239);
nand (n2305,n2243,n2239);
nand (n2306,n2237,n2243);
nand (n2307,n2308,n2309,n2310);
nand (n2308,n2257,n2261);
nand (n2309,n2270,n2261);
nand (n2310,n2257,n2270);
nor (n2311,n2312,n2329);
nor (n2312,n2313,n2317);
nand (n2313,n2314,n2315,n2316);
nand (n2314,n2285,n2295);
nand (n2315,n2307,n2295);
nand (n2316,n2285,n2307);
xor (n2317,n2318,n2325);
xor (n2318,n2319,n2323);
nand (n2319,n2320,n2321,n2322);
nand (n2320,n2287,n2289);
nand (n2321,n2293,n2289);
nand (n2322,n2287,n2293);
xor (n2323,n2324,n737);
xor (n2324,n660,n662);
nand (n2325,n2326,n2327,n2328);
nand (n2326,n2297,n2299);
nand (n2327,n2303,n2299);
nand (n2328,n2297,n2303);
nor (n2329,n2330,n2334);
nand (n2330,n2331,n2332,n2333);
nand (n2331,n2319,n2323);
nand (n2332,n2325,n2323);
nand (n2333,n2319,n2325);
xor (n2334,n2335,n658);
xor (n2335,n436,n520);
not (n2336,n2337);
nor (n2337,n2338,n2353);
nor (n2338,n2226,n2339);
nor (n2339,n2340,n2347);
nor (n2340,n2341,n2346);
nor (n2341,n2342,n2344);
nor (n2342,n2343,n1925);
nand (n2343,n1814,n1818);
not (n2344,n2345);
nand (n2345,n1926,n1930);
not (n2346,n2039);
not (n2347,n2348);
nor (n2348,n2349,n2351);
nor (n2349,n2350,n2147);
nand (n2350,n2041,n2045);
not (n2351,n2352);
nand (n2352,n2148,n2152);
not (n2353,n2354);
nor (n2354,n2355,n2362);
nor (n2355,n2356,n2361);
nor (n2356,n2357,n2359);
nor (n2357,n2358,n2278);
nand (n2358,n2229,n2233);
not (n2359,n2360);
nand (n2360,n2279,n2283);
not (n2361,n2311);
not (n2362,n2363);
nor (n2363,n2364,n2366);
nor (n2364,n2365,n2329);
nand (n2365,n2313,n2317);
not (n2366,n2367);
nand (n2367,n2330,n2334);
nand (n2368,n2369,n2788);
nand (n2369,n2370,n2681);
nor (n2370,n2371,n2666);
nor (n2371,n2372,n2537);
nand (n2372,n2373,n2514);
nor (n2373,n2374,n2491);
nor (n2374,n2375,n2464);
nand (n2375,n2376,n2421,n2463);
nand (n2376,n2377,n2389);
xor (n2377,n2378,n2384);
xor (n2378,n2379,n2380);
xor (n2379,n1682,n1686);
xor (n2380,n2381,n76);
or (n2381,n2382,n2383);
and (n2382,n884,n103);
and (n2383,n898,n107);
and (n2384,n76,n2385);
xor (n2385,n2386,n563);
or (n2386,n2387,n2388);
and (n2387,n530,n686);
and (n2388,n534,n690);
nand (n2389,n2390,n2407,n2420);
nand (n2390,n2391,n2392);
xor (n2391,n76,n2385);
nand (n2392,n2393,n2402,n2406);
nand (n2393,n2394,n2398);
xor (n2394,n2395,n187);
or (n2395,n2396,n2397);
and (n2396,n859,n324);
and (n2397,n861,n328);
xor (n2398,n2399,n326);
or (n2399,n2400,n2401);
and (n2400,n670,n561);
and (n2401,n855,n565);
nand (n2402,n2403,n2398);
and (n2403,n105,n2404);
xnor (n2404,n2405,n105);
nand (n2405,n898,n185);
nand (n2406,n2394,n2403);
nand (n2407,n2408,n2392);
xor (n2408,n2409,n2416);
xor (n2409,n2410,n2414);
xnor (n2410,n2411,n688);
nor (n2411,n2412,n2413);
and (n2412,n295,n870);
and (n2413,n223,n872);
xnor (n2414,n2415,n76);
nand (n2415,n898,n103);
xor (n2416,n2417,n187);
or (n2417,n2418,n2419);
and (n2418,n855,n324);
and (n2419,n859,n328);
nand (n2420,n2391,n2408);
nand (n2421,n2422,n2389);
xor (n2422,n2423,n2442);
xor (n2423,n2424,n2428);
nand (n2424,n2425,n2426,n2427);
nand (n2425,n2410,n2414);
nand (n2426,n2416,n2414);
nand (n2427,n2410,n2416);
xor (n2428,n2429,n2438);
xor (n2429,n2430,n2434);
xor (n2430,n2431,n187);
or (n2431,n2432,n2433);
and (n2432,n670,n324);
and (n2433,n855,n328);
xor (n2434,n2435,n326);
or (n2435,n2436,n2437);
and (n2436,n534,n561);
and (n2437,n536,n565);
xor (n2438,n2439,n105);
or (n2439,n2440,n2441);
and (n2440,n859,n185);
and (n2441,n861,n189);
nand (n2442,n2443,n2457,n2462);
nand (n2443,n2444,n2448);
xor (n2444,n2445,n326);
or (n2445,n2446,n2447);
and (n2446,n536,n561);
and (n2447,n670,n565);
and (n2448,n2449,n2453);
xnor (n2449,n2450,n688);
nor (n2450,n2451,n2452);
and (n2451,n530,n870);
and (n2452,n295,n872);
xor (n2453,n2454,n563);
or (n2454,n2455,n2456);
and (n2455,n534,n686);
and (n2456,n536,n690);
nand (n2457,n2458,n2448);
xor (n2458,n2459,n105);
or (n2459,n2460,n2461);
and (n2460,n861,n185);
and (n2461,n884,n189);
nand (n2462,n2444,n2458);
nand (n2463,n2377,n2422);
xor (n2464,n2465,n2479);
xor (n2465,n2466,n2475);
xor (n2466,n2467,n2473);
xor (n2467,n2468,n2472);
xor (n2468,n2469,n76);
or (n2469,n2470,n2471);
and (n2470,n861,n103);
and (n2471,n884,n107);
xor (n2472,n1626,n17);
xor (n2473,n2474,n1669);
xor (n2474,n1662,n1666);
nand (n2475,n2476,n2477,n2478);
nand (n2476,n2424,n2428);
nand (n2477,n2442,n2428);
nand (n2478,n2424,n2442);
xor (n2479,n2480,n2489);
xor (n2480,n2481,n2485);
nand (n2481,n2482,n2483,n2484);
nand (n2482,n2379,n2380);
nand (n2483,n2384,n2380);
nand (n2484,n2379,n2384);
nand (n2485,n2486,n2487,n2488);
nand (n2486,n2430,n2434);
nand (n2487,n2438,n2434);
nand (n2488,n2430,n2438);
xor (n2489,n2490,n1691);
xor (n2490,n1677,n1681);
nor (n2491,n2492,n2496);
nand (n2492,n2493,n2494,n2495);
nand (n2493,n2466,n2475);
nand (n2494,n2479,n2475);
nand (n2495,n2466,n2479);
xor (n2496,n2497,n2504);
xor (n2497,n2498,n2500);
xor (n2498,n2499,n1675);
xor (n2499,n1656,n1660);
nand (n2500,n2501,n2502,n2503);
nand (n2501,n2481,n2485);
nand (n2502,n2489,n2485);
nand (n2503,n2481,n2489);
xor (n2504,n2505,n2510);
xor (n2505,n2506,n2508);
xor (n2506,n2507,n1625);
xor (n2507,n1616,n1620);
xor (n2508,n2509,n1640);
xor (n2509,n1634,n1638);
nand (n2510,n2511,n2512,n2513);
nand (n2511,n2468,n2472);
nand (n2512,n2473,n2472);
nand (n2513,n2468,n2473);
nor (n2514,n2515,n2530);
nor (n2515,n2516,n2520);
nand (n2516,n2517,n2518,n2519);
nand (n2517,n2498,n2500);
nand (n2518,n2504,n2500);
nand (n2519,n2498,n2504);
xor (n2520,n2521,n2528);
xor (n2521,n2522,n2524);
xor (n2522,n2523,n1632);
xor (n2523,n1612,n1614);
nand (n2524,n2525,n2526,n2527);
nand (n2525,n2506,n2508);
nand (n2526,n2510,n2508);
nand (n2527,n2506,n2510);
xor (n2528,n2529,n1654);
xor (n2529,n1649,n1651);
nor (n2530,n2531,n2535);
nand (n2531,n2532,n2533,n2534);
nand (n2532,n2522,n2524);
nand (n2533,n2528,n2524);
nand (n2534,n2522,n2528);
xor (n2535,n2536,n1647);
xor (n2536,n1522,n1573);
nor (n2537,n2538,n2660);
nor (n2538,n2539,n2636);
nor (n2539,n2540,n2633);
nor (n2540,n2541,n2609);
nand (n2541,n2542,n2581);
or (n2542,n2543,n2567,n2580);
and (n2543,n2544,n2553);
xor (n2544,n2545,n2549);
xnor (n2545,n2546,n688);
nor (n2546,n2547,n2548);
and (n2547,n536,n870);
and (n2548,n534,n872);
xnor (n2549,n2550,n563);
nor (n2550,n2551,n2552);
and (n2551,n855,n690);
and (n2552,n670,n686);
or (n2553,n2554,n2561,n2566);
and (n2554,n2555,n2557);
not (n2555,n2556);
nand (n2556,n898,n324);
xnor (n2557,n2558,n688);
nor (n2558,n2559,n2560);
and (n2559,n670,n870);
and (n2560,n536,n872);
and (n2561,n2557,n2562);
xnor (n2562,n2563,n563);
nor (n2563,n2564,n2565);
and (n2564,n859,n690);
and (n2565,n855,n686);
and (n2566,n2555,n2562);
and (n2567,n2553,n2568);
xor (n2568,n2569,n2576);
xor (n2569,n2570,n2572);
and (n2570,n187,n2571);
xnor (n2571,n2556,n187);
xnor (n2572,n2573,n326);
nor (n2573,n2574,n2575);
and (n2574,n861,n565);
and (n2575,n859,n561);
xnor (n2576,n2577,n187);
nor (n2577,n2578,n2579);
and (n2578,n898,n328);
and (n2579,n884,n324);
and (n2580,n2544,n2568);
xor (n2581,n2582,n2598);
xor (n2582,n2583,n2587);
or (n2583,n2584,n2585,n2586);
and (n2584,n2570,n2572);
and (n2585,n2572,n2576);
and (n2586,n2570,n2576);
xor (n2587,n2588,n2594);
xor (n2588,n2589,n2590);
and (n2589,n2545,n2549);
xnor (n2590,n2591,n326);
nor (n2591,n2592,n2593);
and (n2592,n859,n565);
and (n2593,n855,n561);
xnor (n2594,n2595,n187);
nor (n2595,n2596,n2597);
and (n2596,n884,n328);
and (n2597,n861,n324);
xor (n2598,n2599,n2605);
xor (n2599,n2600,n2601);
not (n2600,n2405);
xnor (n2601,n2602,n688);
nor (n2602,n2603,n2604);
and (n2603,n534,n870);
and (n2604,n530,n872);
xnor (n2605,n2606,n563);
nor (n2606,n2607,n2608);
and (n2607,n670,n690);
and (n2608,n536,n686);
nor (n2609,n2610,n2614);
or (n2610,n2611,n2612,n2613);
and (n2611,n2583,n2587);
and (n2612,n2587,n2598);
and (n2613,n2583,n2598);
xor (n2614,n2615,n2622);
xor (n2615,n2616,n2620);
or (n2616,n2617,n2618,n2619);
and (n2617,n2589,n2590);
and (n2618,n2590,n2594);
and (n2619,n2589,n2594);
xor (n2620,n2621,n2403);
xor (n2621,n2394,n2398);
xor (n2622,n2623,n2629);
xor (n2623,n2624,n2628);
xor (n2624,n2625,n105);
or (n2625,n2626,n2627);
and (n2626,n884,n185);
and (n2627,n898,n189);
xor (n2628,n2449,n2453);
or (n2629,n2630,n2631,n2632);
and (n2630,n2600,n2601);
and (n2631,n2601,n2605);
and (n2632,n2600,n2605);
not (n2633,n2634);
not (n2634,n2635);
and (n2635,n2610,n2614);
not (n2636,n2637);
nor (n2637,n2638,n2653);
nor (n2638,n2639,n2643);
nand (n2639,n2640,n2641,n2642);
nand (n2640,n2616,n2620);
nand (n2641,n2622,n2620);
nand (n2642,n2616,n2622);
xor (n2643,n2644,n2651);
xor (n2644,n2645,n2647);
xor (n2645,n2646,n2458);
xor (n2646,n2444,n2448);
nand (n2647,n2648,n2649,n2650);
nand (n2648,n2624,n2628);
nand (n2649,n2629,n2628);
nand (n2650,n2624,n2629);
xor (n2651,n2652,n2408);
xor (n2652,n2391,n2392);
nor (n2653,n2654,n2658);
nand (n2654,n2655,n2656,n2657);
nand (n2655,n2645,n2647);
nand (n2656,n2651,n2647);
nand (n2657,n2645,n2651);
xor (n2658,n2659,n2422);
xor (n2659,n2377,n2389);
not (n2660,n2661);
nor (n2661,n2662,n2664);
nor (n2662,n2663,n2653);
nand (n2663,n2639,n2643);
not (n2664,n2665);
nand (n2665,n2654,n2658);
not (n2666,n2667);
nor (n2667,n2668,n2675);
nor (n2668,n2669,n2674);
nor (n2669,n2670,n2672);
nor (n2670,n2671,n2491);
nand (n2671,n2375,n2464);
not (n2672,n2673);
nand (n2673,n2492,n2496);
not (n2674,n2514);
not (n2675,n2676);
nor (n2676,n2677,n2679);
nor (n2677,n2678,n2530);
nand (n2678,n2516,n2520);
not (n2679,n2680);
nand (n2680,n2531,n2535);
nand (n2681,n2682,n2686);
nor (n2682,n2683,n2372);
nand (n2683,n2684,n2637);
nor (n2684,n2685,n2609);
nor (n2685,n2542,n2581);
or (n2686,n2687,n2709);
and (n2687,n2688,n2690);
xor (n2688,n2689,n2568);
xor (n2689,n2544,n2553);
or (n2690,n2691,n2705,n2708);
and (n2691,n2692,n2701);
and (n2692,n2693,n2697);
xnor (n2693,n2694,n688);
nor (n2694,n2695,n2696);
and (n2695,n855,n870);
and (n2696,n670,n872);
xnor (n2697,n2698,n563);
nor (n2698,n2699,n2700);
and (n2699,n861,n690);
and (n2700,n859,n686);
xnor (n2701,n2702,n326);
nor (n2702,n2703,n2704);
and (n2703,n884,n565);
and (n2704,n861,n561);
and (n2705,n2701,n2706);
xor (n2706,n2707,n2562);
xor (n2707,n2555,n2557);
and (n2708,n2692,n2706);
and (n2709,n2710,n2711);
xor (n2710,n2688,n2690);
or (n2711,n2712,n2727);
and (n2712,n2713,n2725);
or (n2713,n2714,n2719,n2724);
and (n2714,n2715,n2716);
xor (n2715,n2693,n2697);
and (n2716,n326,n2717);
xnor (n2717,n2718,n326);
nand (n2718,n898,n561);
and (n2719,n2716,n2720);
xnor (n2720,n2721,n326);
nor (n2721,n2722,n2723);
and (n2722,n898,n565);
and (n2723,n884,n561);
and (n2724,n2715,n2720);
xor (n2725,n2726,n2706);
xor (n2726,n2692,n2701);
and (n2727,n2728,n2729);
xor (n2728,n2713,n2725);
or (n2729,n2730,n2746);
and (n2730,n2731,n2733);
xor (n2731,n2732,n2720);
xor (n2732,n2715,n2716);
or (n2733,n2734,n2740,n2745);
and (n2734,n2735,n2736);
not (n2735,n2718);
xnor (n2736,n2737,n688);
nor (n2737,n2738,n2739);
and (n2738,n859,n870);
and (n2739,n855,n872);
and (n2740,n2736,n2741);
xnor (n2741,n2742,n563);
nor (n2742,n2743,n2744);
and (n2743,n884,n690);
and (n2744,n861,n686);
and (n2745,n2735,n2741);
and (n2746,n2747,n2748);
xor (n2747,n2731,n2733);
or (n2748,n2749,n2760);
and (n2749,n2750,n2752);
xor (n2750,n2751,n2741);
xor (n2751,n2735,n2736);
and (n2752,n2753,n2756);
and (n2753,n563,n2754);
xnor (n2754,n2755,n563);
nand (n2755,n898,n686);
xnor (n2756,n2757,n688);
nor (n2757,n2758,n2759);
and (n2758,n861,n870);
and (n2759,n859,n872);
and (n2760,n2761,n2762);
xor (n2761,n2750,n2752);
or (n2762,n2763,n2769);
and (n2763,n2764,n2768);
xnor (n2764,n2765,n563);
nor (n2765,n2766,n2767);
and (n2766,n898,n690);
and (n2767,n884,n686);
xor (n2768,n2753,n2756);
and (n2769,n2770,n2771);
xor (n2770,n2764,n2768);
or (n2771,n2772,n2778);
and (n2772,n2773,n2777);
xnor (n2773,n2774,n688);
nor (n2774,n2775,n2776);
and (n2775,n884,n870);
and (n2776,n861,n872);
not (n2777,n2755);
and (n2778,n2779,n2780);
xor (n2779,n2773,n2777);
and (n2780,n2781,n2785);
xnor (n2781,n2782,n688);
nor (n2782,n2783,n2784);
and (n2783,n898,n870);
and (n2784,n884,n872);
and (n2785,n2786,n688);
xnor (n2786,n2787,n688);
nand (n2787,n898,n872);
not (n2788,n2789);
nand (n2789,n2790,n1810);
nor (n2790,n2791,n842);
nand (n2791,n2792,n1765);
nor (n2792,n2793,n1737);
nor (n2793,n1520,n1699);
not (n2794,n2795);
nand (n2795,n2796,n807);
nor (n2796,n2797,n779);
nor (n2797,n434,n741);
nand (n2798,n2799,n2856);
not (n2799,n2800);
nor (n2800,n2801,n2805);
nand (n2801,n2802,n2803,n2804);
nand (n2802,n375,n379);
nand (n2803,n419,n379);
nand (n2804,n375,n419);
xor (n2805,n2806,n2852);
xor (n2806,n2807,n2830);
xor (n2807,n2808,n2817);
xor (n2808,n2809,n2813);
nand (n2809,n2810,n2811,n2812);
nand (n2810,n69,n401);
nand (n2811,n405,n401);
nand (n2812,n69,n405);
nand (n2813,n2814,n2815,n2816);
nand (n2814,n411,n70);
nand (n2815,n415,n70);
nand (n2816,n411,n415);
xor (n2817,n2818,n2826);
xor (n2818,n2819,n2822);
xor (n2819,n2820,n22);
or (n2820,n403,n2821);
and (n2821,n73,n20);
xor (n2822,n2823,n57);
or (n2823,n2824,n2825);
and (n2824,n37,n51);
and (n2825,n41,n55);
xor (n2826,n2827,n68);
or (n2827,n2828,n2829);
and (n2828,n50,n62);
and (n2829,n54,n66);
xor (n2830,n2831,n2848);
xor (n2831,n2832,n2843);
xor (n2832,n2833,n68);
xor (n2833,n2834,n2838);
xor (n2834,n2835,n44);
or (n2835,n2836,n2837);
and (n2836,n26,n38);
and (n2837,n30,n42);
not (n2838,n2839);
xor (n2839,n2840,n33);
or (n2840,n2841,n2842);
and (n2841,n14,n27);
and (n2842,n19,n31);
nand (n2843,n2844,n2846,n2847);
nand (n2844,n2845,n68);
xor (n2845,n386,n68);
nand (n2846,n389,n68);
nand (n2847,n2845,n389);
nand (n2848,n2849,n2850,n2851);
nand (n2849,n395,n399);
nand (n2850,n409,n399);
nand (n2851,n395,n409);
nand (n2852,n2853,n2854,n2855);
nand (n2853,n381,n385);
nand (n2854,n393,n385);
nand (n2855,n381,n393);
nand (n2856,n2801,n2805);
xor (n2857,n2858,n3039);
xnor (n2858,n2859,n2933);
xor (n2859,n2860,n2888);
xor (n2860,n2861,n2875);
or (n2861,n2862,n2867,n2874);
and (n2862,n2863,n2865);
xor (n2863,n2864,n2845);
xor (n2864,n411,n415);
and (n2865,n9,n2866);
not (n2866,n45);
and (n2867,n2865,n2868);
xor (n2868,n2869,n399);
xor (n2869,n389,n2870);
or (n2870,n2871,n2872,n2873);
and (n2871,n70,n47);
not (n2872,n396);
and (n2873,n70,n58);
and (n2874,n2863,n2868);
xor (n2875,n2876,n2885);
xor (n2876,n2877,n2881);
or (n2877,n2878,n2879,n2880);
not (n2878,n2816);
and (n2879,n415,n2845);
and (n2880,n411,n2845);
or (n2881,n2882,n2883,n2884);
and (n2882,n389,n2870);
and (n2883,n2870,n399);
and (n2884,n389,n399);
xor (n2885,n2886,n2809);
xor (n2886,n2887,n2833);
not (n2887,n2817);
or (n2888,n2889,n2902,n2932);
and (n2889,n2890,n2900);
or (n2890,n2891,n2897,n2899);
and (n2891,n2892,n2893);
not (n2892,n81);
or (n2893,n2894,n2895,n2896);
not (n2894,n98);
and (n2895,n109,n120);
and (n2896,n99,n120);
and (n2897,n2893,n2898);
not (n2898,n8);
and (n2899,n2892,n2898);
xor (n2900,n2901,n2868);
xor (n2901,n2863,n2865);
and (n2902,n2900,n2903);
or (n2903,n2904,n2918,n2931);
and (n2904,n2905,n2909);
or (n2905,n2906,n2907,n2908);
and (n2906,n113,n125);
and (n2907,n125,n167);
and (n2908,n113,n167);
or (n2909,n2910,n2915,n2917);
and (n2910,n134,n2911);
or (n2911,n2912,n2913,n2914);
and (n2912,n100,n153);
not (n2913,n157);
and (n2914,n100,n158);
and (n2915,n2911,n2916);
xor (n2916,n133,n120);
and (n2917,n134,n2916);
and (n2918,n2909,n2919);
or (n2919,n2920,n2927,n2930);
and (n2920,n2921,n2922);
not (n2921,n205);
or (n2922,n2923,n2925,n2926);
and (n2923,n173,n2924);
not (n2924,n249);
and (n2925,n2924,n179);
not (n2926,n200);
and (n2927,n2922,n2928);
xor (n2928,n2929,n167);
xor (n2929,n113,n125);
and (n2930,n2921,n2928);
and (n2931,n2905,n2919);
and (n2932,n2890,n2903);
or (n2933,n2934,n2966,n3038);
and (n2934,n2935,n2964);
or (n2935,n2936,n2960,n2963);
and (n2936,n2937,n2939);
xor (n2937,n2938,n2898);
xor (n2938,n2892,n2893);
or (n2939,n2940,n2956,n2959);
and (n2940,n2941,n2943);
xor (n2941,n2942,n2916);
xor (n2942,n134,n2911);
or (n2943,n2944,n2950,n2955);
and (n2944,n282,n2945);
and (n2945,n2946,n298);
or (n2946,n2947,n2948,n2949);
and (n2947,n182,n287);
not (n2948,n286);
and (n2949,n182,n291);
and (n2950,n2945,n2951);
or (n2951,n2952,n2953,n2954);
not (n2952,n232);
and (n2953,n233,n258);
and (n2954,n228,n258);
and (n2955,n282,n2951);
and (n2956,n2943,n2957);
xor (n2957,n2958,n2928);
xor (n2958,n2921,n2922);
and (n2959,n2941,n2957);
and (n2960,n2939,n2961);
xor (n2961,n2962,n2919);
xor (n2962,n2905,n2909);
and (n2963,n2937,n2961);
xor (n2964,n2965,n2903);
xor (n2965,n2890,n2900);
and (n2966,n2964,n2967);
or (n2967,n2968,n2970);
xor (n2968,n2969,n2961);
xor (n2969,n2937,n2939);
or (n2970,n2971,n3002,n3037);
and (n2971,n2972,n3000);
or (n2972,n2973,n2982,n2999);
and (n2973,n2974,n2976);
xor (n2974,n2975,n179);
xor (n2975,n173,n2924);
or (n2976,n2977,n2979,n2981);
and (n2977,n2978,n255);
not (n2978,n308);
and (n2979,n255,n2980);
xor (n2980,n2946,n298);
and (n2981,n2978,n2980);
and (n2982,n2976,n2983);
or (n2983,n2984,n2995,n2998);
and (n2984,n2985,n2990);
or (n2985,n2986,n2988,n2989);
and (n2986,n342,n2987);
not (n2987,n761);
and (n2988,n2987,n760);
and (n2989,n342,n760);
or (n2990,n2991,n2993,n2994);
and (n2991,n345,n2992);
not (n2992,n756);
and (n2993,n2992,n318);
and (n2994,n345,n318);
and (n2995,n2990,n2996);
xor (n2996,n2997,n258);
xor (n2997,n228,n233);
and (n2998,n2985,n2996);
and (n2999,n2974,n2983);
xor (n3000,n3001,n2957);
xor (n3001,n2941,n2943);
and (n3002,n3000,n3003);
or (n3003,n3004,n3033,n3036);
and (n3004,n3005,n3007);
xor (n3005,n3006,n2951);
xor (n3006,n282,n2945);
or (n3007,n3008,n3029,n3032);
and (n3008,n3009,n3027);
or (n3009,n3010,n3023,n3026);
and (n3010,n3011,n3015);
or (n3011,n3012,n3013,n3014);
and (n3012,n440,n514);
and (n3013,n514,n583);
and (n3014,n440,n583);
or (n3015,n3016,n3017,n3022);
and (n3016,n444,n516);
and (n3017,n516,n3018);
or (n3018,n3019,n3020,n3021);
and (n3019,n321,n545);
not (n3020,n581);
and (n3021,n321,n541);
and (n3022,n444,n3018);
and (n3023,n3015,n3024);
xor (n3024,n3025,n760);
xor (n3025,n342,n2987);
and (n3026,n3011,n3024);
xor (n3027,n3028,n2980);
xor (n3028,n2978,n255);
and (n3029,n3027,n3030);
xor (n3030,n3031,n2996);
xor (n3031,n2985,n2990);
and (n3032,n3009,n3030);
and (n3033,n3007,n3034);
xor (n3034,n3035,n2983);
xor (n3035,n2974,n2976);
and (n3036,n3005,n3034);
and (n3037,n2972,n3003);
and (n3038,n2935,n2967);
and (n3039,n3040,n3042);
xor (n3040,n3041,n2967);
xor (n3041,n2935,n2964);
and (n3042,n3043,n3044);
xnor (n3043,n2968,n2970);
or (n3044,n3045,n3125);
and (n3045,n3046,n3048);
xor (n3046,n3047,n3003);
xor (n3047,n2972,n3000);
or (n3048,n3049,n3051);
xor (n3049,n3050,n3034);
xor (n3050,n3005,n3007);
or (n3051,n3052,n3075,n3124);
and (n3052,n3053,n3073);
or (n3053,n3054,n3069,n3072);
and (n3054,n3055,n3057);
xor (n3055,n3056,n318);
xor (n3056,n345,n2992);
or (n3057,n3058,n3065,n3068);
and (n3058,n512,n3059);
or (n3059,n3060,n3062,n3064);
and (n3060,n573,n3061);
not (n3061,n539);
and (n3062,n3061,n3063);
not (n3063,n525);
and (n3064,n573,n3063);
and (n3065,n3059,n3066);
xor (n3066,n3067,n583);
xor (n3067,n440,n514);
and (n3068,n512,n3066);
and (n3069,n3057,n3070);
xor (n3070,n3071,n3024);
xor (n3071,n3011,n3015);
and (n3072,n3055,n3070);
xor (n3073,n3074,n3030);
xor (n3074,n3009,n3027);
and (n3075,n3073,n3076);
or (n3076,n3077,n3088,n3123);
and (n3077,n3078,n3086);
or (n3078,n3079,n3082,n3085);
and (n3079,n3080,n460);
xor (n3080,n3081,n3018);
xor (n3081,n444,n516);
and (n3082,n460,n3083);
xor (n3083,n3084,n3066);
xor (n3084,n512,n3059);
and (n3085,n3080,n3083);
xor (n3086,n3087,n3070);
xor (n3087,n3055,n3057);
and (n3088,n3086,n3089);
or (n3089,n3090,n3119,n3122);
and (n3090,n3091,n3104);
or (n3091,n3092,n3102,n3103);
and (n3092,n3093,n618);
or (n3093,n3094,n3099,n3101);
and (n3094,n3095,n612);
or (n3095,n3096,n3097,n3098);
and (n3096,n557,n602);
not (n3097,n606);
and (n3098,n557,n607);
and (n3099,n612,n3100);
not (n3100,n615);
and (n3101,n3095,n3100);
not (n3102,n653);
and (n3103,n3093,n654);
or (n3104,n3105,n3112,n3118);
and (n3105,n3106,n3110);
or (n3106,n3107,n3108,n3109);
and (n3107,n558,n554);
not (n3108,n572);
and (n3109,n558,n568);
xor (n3110,n3111,n3063);
xor (n3111,n573,n3061);
and (n3112,n3110,n3113);
or (n3113,n3114,n3115,n3117);
and (n3114,n557,n695);
and (n3115,n695,n3116);
not (n3116,n2290);
and (n3117,n557,n3116);
and (n3118,n3106,n3113);
and (n3119,n3104,n3120);
xor (n3120,n3121,n3083);
xor (n3121,n3080,n460);
and (n3122,n3091,n3120);
and (n3123,n3078,n3089);
and (n3124,n3053,n3076);
and (n3125,n3126,n3127);
xor (n3126,n3046,n3048);
and (n3127,n3128,n3129);
xnor (n3128,n3049,n3051);
or (n3129,n3130,n3215);
and (n3130,n3131,n3133);
xor (n3131,n3132,n3076);
xor (n3132,n3053,n3073);
or (n3133,n3134,n3136);
xor (n3134,n3135,n3089);
xor (n3135,n3078,n3086);
or (n3136,n3137,n3159,n3214);
and (n3137,n3138,n3157);
or (n3138,n3139,n3153,n3156);
and (n3139,n3140,n3142);
xor (n3140,n3141,n654);
xor (n3141,n3093,n618);
or (n3142,n3143,n3146,n3152);
and (n3143,n3144,n2293);
xor (n3144,n3145,n3100);
xor (n3145,n3095,n612);
and (n3146,n2293,n3147);
or (n3147,n3148,n3149,n3151);
not (n3148,n734);
and (n3149,n718,n3150);
not (n3150,n715);
and (n3151,n699,n3150);
and (n3152,n3144,n3147);
and (n3153,n3142,n3154);
xor (n3154,n3155,n3113);
xor (n3155,n3106,n3110);
and (n3156,n3140,n3154);
xor (n3157,n3158,n3120);
xor (n3158,n3091,n3104);
and (n3159,n3157,n3160);
or (n3160,n3161,n3176,n3213);
and (n3161,n3162,n3174);
or (n3162,n3163,n3170,n3173);
and (n3163,n3164,n3168);
or (n3164,n3165,n3166,n3167);
and (n3165,n666,n2263);
and (n3166,n2263,n2244);
and (n3167,n666,n2244);
xor (n3168,n3169,n3116);
xor (n3169,n557,n695);
and (n3170,n3168,n3171);
and (n3171,n2239,n3172);
not (n3172,n2237);
and (n3173,n3164,n3171);
xor (n3174,n3175,n3154);
xor (n3175,n3140,n3142);
and (n3176,n3174,n3177);
or (n3177,n3178,n3198,n3212);
and (n3178,n3179,n3196);
or (n3179,n3180,n3185,n3195);
and (n3180,n3181,n2266);
or (n3181,n3182,n3183,n3184);
and (n3182,n683,n674);
not (n3183,n673);
and (n3184,n683,n677);
and (n3185,n2266,n3186);
or (n3186,n3187,n3192,n3194);
and (n3187,n682,n3188);
or (n3188,n3189,n3190,n3191);
and (n3189,n682,n2067);
not (n3190,n2181);
and (n3191,n682,n2071);
and (n3192,n3188,n3193);
not (n3193,n2176);
and (n3194,n682,n3193);
and (n3195,n3181,n3186);
xor (n3196,n3197,n3147);
xor (n3197,n3144,n2293);
and (n3198,n3196,n3199);
or (n3199,n3200,n3204,n3211);
and (n3200,n3201,n3203);
xor (n3201,n3202,n2244);
xor (n3202,n666,n2263);
not (n3203,n2236);
and (n3204,n3203,n3205);
or (n3205,n3206,n3209,n3210);
and (n3206,n3207,n2182);
and (n3207,n2051,n3208);
not (n3208,n2065);
and (n3209,n2182,n2204);
and (n3210,n3207,n2204);
and (n3211,n3201,n3205);
and (n3212,n3179,n3199);
and (n3213,n3162,n3177);
and (n3214,n3138,n3160);
and (n3215,n3216,n3217);
xor (n3216,n3131,n3133);
and (n3217,n3218,n3219);
xnor (n3218,n3134,n3136);
or (n3219,n3220,n3424);
and (n3220,n3221,n3223);
xor (n3221,n3222,n3160);
xor (n3222,n3138,n3157);
or (n3223,n3224,n3299,n3423);
and (n3224,n3225,n3297);
or (n3225,n3226,n3293,n3296);
and (n3226,n3227,n3229);
xor (n3227,n3228,n3171);
xor (n3228,n3164,n3168);
or (n3229,n3230,n3264,n3292);
and (n3230,n3231,n3262);
or (n3231,n3232,n3250,n3261);
and (n3232,n3233,n3242);
and (n3233,n3234,n2091);
or (n3234,n3235,n3240,n3241);
and (n3235,n3236,n1961);
or (n3236,n3237,n3238,n3239);
and (n3237,n2030,n1826);
not (n3238,n1970);
and (n3239,n2030,n1830);
not (n3240,n2103);
and (n3241,n3236,n1965);
or (n3242,n3243,n3248,n3249);
and (n3243,n2131,n3244);
or (n3244,n3245,n3246,n3247);
and (n3245,n2030,n1950);
not (n3246,n2078);
and (n3247,n2030,n1955);
and (n3248,n3244,n2112);
and (n3249,n2131,n2112);
and (n3250,n3242,n3251);
or (n3251,n3252,n3258,n3260);
and (n3252,n3253,n3254);
not (n3253,n2050);
or (n3254,n3255,n3256,n3257);
and (n3255,n1834,n2026);
not (n3256,n2130);
and (n3257,n1834,n2031);
and (n3258,n3254,n3259);
not (n3259,n2107);
and (n3260,n3253,n3259);
and (n3261,n3233,n3251);
xor (n3262,n3263,n3186);
xor (n3263,n3181,n2266);
and (n3264,n3262,n3265);
or (n3265,n3266,n3288,n3291);
and (n3266,n3267,n3269);
xor (n3267,n3268,n3193);
xor (n3268,n682,n3188);
or (n3269,n3270,n3279,n3287);
and (n3270,n3271,n3278);
or (n3271,n3272,n3274,n3277);
and (n3272,n2010,n3273);
not (n3273,n2007);
and (n3274,n3273,n3275);
xor (n3275,n3276,n1955);
xor (n3276,n2030,n1950);
and (n3277,n2010,n3275);
xor (n3278,n3234,n2091);
and (n3279,n3278,n3280);
or (n3280,n3281,n3285,n3286);
and (n3281,n3282,n3283);
not (n3282,n2024);
xor (n3283,n3284,n1965);
xor (n3284,n3236,n1961);
and (n3285,n3283,n1984);
and (n3286,n3282,n1984);
and (n3287,n3271,n3280);
and (n3288,n3269,n3289);
xor (n3289,n3290,n2204);
xor (n3290,n3207,n2182);
and (n3291,n3267,n3289);
and (n3292,n3231,n3265);
and (n3293,n3229,n3294);
xor (n3294,n3295,n3199);
xor (n3295,n3179,n3196);
and (n3296,n3227,n3294);
xor (n3297,n3298,n3177);
xor (n3298,n3162,n3174);
and (n3299,n3297,n3300);
or (n3300,n3301,n3334,n3422);
and (n3301,n3302,n3332);
or (n3302,n3303,n3328,n3331);
and (n3303,n3304,n3306);
xor (n3304,n3305,n3205);
xor (n3305,n3201,n3203);
or (n3306,n3307,n3324,n3327);
and (n3307,n3308,n3310);
xor (n3308,n3309,n3251);
xor (n3309,n3233,n3242);
or (n3310,n3311,n3316,n3323);
and (n3311,n3312,n3314);
xor (n3312,n3313,n2112);
xor (n3313,n2131,n3244);
xor (n3314,n3315,n3259);
xor (n3315,n3253,n3254);
and (n3316,n3314,n3317);
and (n3317,n1975,n3318);
or (n3318,n3319,n3320,n3322);
not (n3319,n1981);
and (n3320,n1841,n3321);
not (n3321,n1824);
and (n3322,n1837,n3321);
and (n3323,n3312,n3317);
and (n3324,n3310,n3325);
xor (n3325,n3326,n3289);
xor (n3326,n3267,n3269);
and (n3327,n3308,n3325);
and (n3328,n3306,n3329);
xor (n3329,n3330,n3265);
xor (n3330,n3231,n3262);
and (n3331,n3304,n3329);
xor (n3332,n3333,n3294);
xor (n3333,n3227,n3229);
and (n3334,n3332,n3335);
or (n3335,n3336,n3393,n3421);
and (n3336,n3337,n3339);
xor (n3337,n3338,n3329);
xor (n3338,n3304,n3306);
or (n3339,n3340,n3372,n3392);
and (n3340,n3341,n3370);
or (n3341,n3342,n3355,n3369);
and (n3342,n3343,n3353);
or (n3343,n3344,n3351,n3352);
and (n3344,n3345,n3349);
or (n3345,n3346,n3347,n3348);
and (n3346,n1889,n1874);
and (n3347,n1874,n1857);
and (n3348,n1889,n1857);
xor (n3349,n3350,n3275);
xor (n3350,n2010,n3273);
and (n3351,n3349,n2035);
and (n3352,n3345,n2035);
xor (n3353,n3354,n3280);
xor (n3354,n3271,n3278);
and (n3355,n3353,n3356);
or (n3356,n3357,n3366,n3368);
and (n3357,n3358,n3364);
or (n3358,n3359,n3360,n3363);
and (n3359,n1879,n1873);
and (n3360,n1873,n3361);
xor (n3361,n3362,n1857);
xor (n3362,n1889,n1874);
and (n3363,n1879,n3361);
xor (n3364,n3365,n1984);
xor (n3365,n3282,n3283);
and (n3366,n3364,n3367);
xor (n3367,n1975,n3318);
and (n3368,n3358,n3367);
and (n3369,n3343,n3356);
xor (n3370,n3371,n3325);
xor (n3371,n3308,n3310);
and (n3372,n3370,n3373);
or (n3373,n3374,n3388,n3391);
and (n3374,n3375,n3377);
xor (n3375,n3376,n3317);
xor (n3376,n3312,n3314);
or (n3377,n3378,n3386,n3387);
and (n3378,n3379,n3381);
xor (n3379,n3380,n2035);
xor (n3380,n3345,n3349);
or (n3381,n3382,n3383,n3385);
not (n3382,n1934);
and (n3383,n1849,n3384);
not (n3384,n1822);
and (n3385,n1845,n3384);
and (n3386,n3381,n1936);
and (n3387,n3379,n1936);
and (n3388,n3377,n3389);
xor (n3389,n3390,n3356);
xor (n3390,n3343,n3353);
and (n3391,n3375,n3389);
and (n3392,n3341,n3373);
and (n3393,n3339,n3394);
or (n3394,n3395,n3397);
xor (n3395,n3396,n3373);
xor (n3396,n3341,n3370);
or (n3397,n3398,n3414,n3420);
and (n3398,n3399,n3412);
or (n3399,n3400,n3408,n3411);
and (n3400,n3401,n3403);
xor (n3401,n3402,n3367);
xor (n3402,n3358,n3364);
or (n3403,n3404,n3406,n3407);
and (n3404,n3405,n1921);
not (n3405,n1820);
not (n3406,n1928);
and (n3407,n3405,n1853);
and (n3408,n3403,n3409);
xor (n3409,n3410,n1936);
xor (n3410,n3379,n3381);
and (n3411,n3401,n3409);
xor (n3412,n3413,n3389);
xor (n3413,n3375,n3377);
and (n3414,n3412,n3415);
or (n3415,n3416,n3418);
or (n3416,n1814,n3417);
not (n3417,n1818);
xor (n3418,n3419,n3409);
xor (n3419,n3401,n3403);
and (n3420,n3399,n3415);
and (n3421,n3337,n3394);
and (n3422,n3302,n3335);
and (n3423,n3225,n3300);
and (n3424,n3425,n3426);
xor (n3425,n3221,n3223);
and (n3426,n3427,n3429);
xor (n3427,n3428,n3300);
xor (n3428,n3225,n3297);
or (n3429,n3430,n3432);
xor (n3430,n3431,n3335);
xor (n3431,n3302,n3332);
and (n3432,n3433,n3434);
not (n3433,n3430);
and (n3434,n3435,n3437);
xor (n3435,n3436,n3394);
xor (n3436,n3337,n3339);
and (n3437,n3438,n3439);
xnor (n3438,n3395,n3397);
and (n3439,n3440,n3442);
xor (n3440,n3441,n3415);
xor (n3441,n3399,n3412);
and (n3442,n3443,n3444);
xnor (n3443,n3416,n3418);
and (n3444,n3445,n3448);
not (n3445,n3446);
nand (n3446,n3447,n2343);
not (n3447,n1813);
nand (n3448,n840,n3449);
nand (n3449,n2790,n2369);
endmodule
