module top (out,n4,n8,n10,n11,n13,n15,n16,n36,n37
        ,n45,n46,n48,n49,n66,n67,n69,n78,n79,n88
        ,n99,n100,n107,n113,n126,n135,n140,n158,n202,n396);
output out;
input n4;
input n8;
input n10;
input n11;
input n13;
input n15;
input n16;
input n36;
input n37;
input n45;
input n46;
input n48;
input n49;
input n66;
input n67;
input n69;
input n78;
input n79;
input n88;
input n99;
input n100;
input n107;
input n113;
input n126;
input n135;
input n140;
input n158;
input n202;
input n396;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n9;
wire n12;
wire n14;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n47;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
xnor (out,n0,n397);
nand (n0,n1,n396);
nand (n1,n2,n17);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
xor (n6,n7,n12);
and (n7,n8,n9);
wire s0n9,s1n9,notn9;
or (n9,s0n9,s1n9);
not(notn9,n4);
and (s0n9,notn9,n10);
and (s1n9,n4,n11);
and (n12,n13,n14);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n4);
and (s0n14,notn14,n15);
and (s1n14,n4,n16);
nand (n17,n18,n3);
nand (n18,n19,n395);
or (n19,n20,n226);
not (n20,n21);
or (n21,n22,n225);
and (n22,n23,n182);
or (n23,n24,n181);
and (n24,n25,n150);
xor (n25,n26,n117);
or (n26,n27,n116);
and (n27,n28,n91);
xor (n28,n29,n60);
nand (n29,n30,n55);
or (n30,n31,n40);
not (n31,n32);
nand (n32,n33,n38);
or (n33,n34,n13);
not (n34,n35);
wire s0n35,s1n35,notn35;
or (n35,s0n35,s1n35);
not(notn35,n4);
and (s0n35,notn35,n36);
and (s1n35,n4,n37);
or (n38,n35,n39);
not (n39,n13);
nand (n40,n41,n52);
nor (n41,n42,n50);
and (n42,n43,n47);
not (n43,n44);
wire s0n44,s1n44,notn44;
or (n44,s0n44,s1n44);
not(notn44,n4);
and (s0n44,notn44,n45);
and (s1n44,n4,n46);
wire s0n47,s1n47,notn47;
or (n47,s0n47,s1n47);
not(notn47,n4);
and (s0n47,notn47,n48);
and (s1n47,n4,n49);
and (n50,n44,n51);
not (n51,n47);
nand (n52,n53,n54);
or (n53,n43,n35);
nand (n54,n35,n43);
or (n55,n41,n56);
nor (n56,n57,n58);
and (n57,n8,n34);
and (n58,n59,n35);
not (n59,n8);
nand (n60,n61,n85);
or (n61,n62,n72);
not (n62,n63);
nand (n63,n64,n70);
or (n64,n65,n68);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n4);
and (s0n65,notn65,n66);
and (s1n65,n4,n67);
not (n68,n69);
or (n70,n71,n69);
not (n71,n65);
not (n72,n73);
and (n73,n74,n81);
nand (n74,n75,n80);
or (n75,n76,n65);
not (n76,n77);
wire s0n77,s1n77,notn77;
or (n77,s0n77,s1n77);
not(notn77,n4);
and (s0n77,notn77,n78);
and (s1n77,n4,n79);
nand (n80,n65,n76);
not (n81,n82);
nand (n82,n83,n84);
or (n83,n76,n14);
nand (n84,n14,n76);
nand (n85,n82,n86);
nor (n86,n87,n89);
and (n87,n88,n65);
and (n89,n90,n71);
not (n90,n88);
nand (n91,n92,n110);
or (n92,n93,n105);
nand (n93,n94,n102);
not (n94,n95);
nand (n95,n96,n101);
or (n96,n97,n65);
not (n97,n98);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n4);
and (s0n98,notn98,n99);
and (s1n98,n4,n100);
nand (n101,n65,n97);
nand (n102,n103,n104);
or (n103,n97,n47);
nand (n104,n47,n97);
nor (n105,n106,n108);
and (n106,n51,n107);
and (n108,n47,n109);
not (n109,n107);
or (n110,n94,n111);
nor (n111,n112,n114);
and (n112,n51,n113);
and (n114,n47,n115);
not (n115,n113);
and (n116,n29,n60);
xor (n117,n118,n144);
xor (n118,n119,n127);
and (n119,n120,n13);
not (n120,n121);
nand (n121,n35,n122);
not (n122,n123);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n4);
and (s0n123,notn123,1'b0);
and (s1n123,n4,n125);
and (n125,n126,n37);
nand (n127,n128,n137);
or (n128,n129,n132);
not (n129,n130);
nor (n130,n131,n9);
not (n131,n14);
nor (n132,n133,n136);
and (n133,n134,n14);
not (n134,n135);
and (n136,n135,n131);
or (n137,n138,n143);
nor (n138,n139,n141);
and (n139,n131,n140);
and (n141,n14,n142);
not (n142,n140);
not (n143,n9);
nand (n144,n145,n146);
or (n145,n40,n56);
or (n146,n41,n147);
nor (n147,n148,n149);
and (n148,n107,n34);
and (n149,n109,n35);
xor (n150,n151,n167);
xor (n151,n152,n161);
nand (n152,n153,n155);
or (n153,n72,n154);
not (n154,n86);
or (n155,n81,n156);
nor (n156,n157,n159);
and (n157,n71,n158);
and (n159,n65,n160);
not (n160,n158);
nand (n161,n162,n163);
or (n162,n93,n111);
or (n163,n94,n164);
nor (n164,n165,n166);
and (n165,n51,n69);
and (n166,n47,n68);
and (n167,n168,n173);
nor (n168,n169,n34);
nor (n169,n170,n172);
and (n170,n51,n171);
nand (n171,n44,n13);
and (n172,n43,n39);
nand (n173,n174,n179);
or (n174,n175,n129);
not (n175,n176);
nor (n176,n177,n178);
and (n177,n158,n14);
and (n178,n160,n131);
nand (n179,n180,n9);
not (n180,n132);
and (n181,n26,n117);
xor (n182,n183,n208);
xor (n183,n184,n205);
xor (n184,n185,n197);
xor (n185,n186,n193);
nand (n186,n187,n188);
or (n187,n147,n40);
nand (n188,n189,n192);
nor (n189,n190,n191);
and (n190,n113,n35);
and (n191,n115,n34);
not (n192,n41);
nor (n193,n121,n194);
nor (n194,n195,n196);
and (n195,n123,n59);
and (n196,n122,n8);
nand (n197,n198,n199);
or (n198,n129,n138);
or (n199,n200,n143);
nor (n200,n201,n203);
and (n201,n131,n202);
and (n203,n14,n204);
not (n204,n202);
or (n205,n206,n207);
and (n206,n151,n167);
and (n207,n152,n161);
xor (n208,n209,n222);
xor (n209,n210,n216);
nand (n210,n211,n212);
or (n211,n93,n164);
or (n212,n94,n213);
nor (n213,n214,n215);
and (n214,n51,n88);
and (n215,n47,n90);
nand (n216,n217,n218);
or (n217,n72,n156);
or (n218,n219,n81);
nor (n219,n220,n221);
and (n220,n71,n135);
and (n221,n65,n134);
or (n222,n223,n224);
and (n223,n118,n144);
and (n224,n119,n127);
nor (n225,n23,n182);
not (n226,n227);
nand (n227,n228,n394);
or (n228,n229,n389);
nor (n229,n230,n387);
and (n230,n231,n376);
or (n231,n232,n375);
and (n232,n233,n291);
xor (n233,n234,n274);
or (n234,n235,n273);
and (n235,n236,n258);
xor (n236,n237,n247);
nand (n237,n238,n243);
or (n238,n239,n72);
not (n239,n240);
nor (n240,n241,n242);
and (n241,n109,n71);
and (n242,n107,n65);
nand (n243,n82,n244);
nor (n244,n245,n246);
and (n245,n113,n65);
and (n246,n71,n115);
nand (n247,n248,n253);
or (n248,n249,n94);
not (n249,n250);
nor (n250,n251,n252);
and (n251,n8,n47);
and (n252,n59,n51);
nand (n253,n254,n255);
not (n254,n93);
nand (n255,n256,n257);
or (n256,n51,n13);
or (n257,n47,n39);
xor (n258,n259,n264);
and (n259,n260,n47);
nand (n260,n261,n263);
or (n261,n65,n262);
and (n262,n13,n98);
or (n263,n98,n13);
nand (n264,n265,n269);
or (n265,n129,n266);
nor (n266,n267,n268);
and (n267,n131,n69);
and (n268,n14,n68);
or (n269,n270,n143);
nor (n270,n271,n272);
and (n271,n88,n131);
and (n272,n90,n14);
and (n273,n237,n247);
xor (n274,n275,n280);
xor (n275,n276,n279);
nand (n276,n277,n278);
or (n277,n249,n93);
or (n278,n94,n105);
and (n279,n259,n264);
xor (n280,n281,n287);
xor (n281,n282,n283);
and (n282,n192,n13);
nand (n283,n284,n285);
or (n284,n143,n175);
nand (n285,n286,n130);
not (n286,n270);
nand (n287,n288,n290);
or (n288,n289,n72);
not (n289,n244);
nand (n290,n82,n63);
or (n291,n292,n374);
and (n292,n293,n314);
xor (n293,n294,n313);
or (n294,n295,n312);
and (n295,n296,n305);
xor (n296,n297,n298);
and (n297,n95,n13);
nand (n298,n299,n304);
or (n299,n300,n72);
not (n300,n301);
nor (n301,n302,n303);
and (n302,n8,n65);
and (n303,n59,n71);
nand (n304,n240,n82);
nand (n305,n306,n311);
or (n306,n129,n307);
not (n307,n308);
nor (n308,n309,n310);
and (n309,n115,n131);
and (n310,n113,n14);
or (n311,n266,n143);
and (n312,n297,n298);
xor (n313,n236,n258);
or (n314,n315,n373);
and (n315,n316,n372);
xor (n316,n317,n331);
nor (n317,n318,n326);
not (n318,n319);
nand (n319,n320,n325);
or (n320,n321,n129);
not (n321,n322);
nand (n322,n323,n324);
or (n323,n109,n14);
nand (n324,n14,n109);
nand (n325,n308,n9);
nand (n326,n327,n65);
nand (n327,n328,n330);
or (n328,n14,n329);
and (n329,n13,n77);
or (n330,n77,n13);
nand (n331,n332,n370);
or (n332,n333,n356);
not (n333,n334);
nand (n334,n335,n355);
or (n335,n336,n345);
nor (n336,n337,n344);
nand (n337,n338,n343);
or (n338,n339,n129);
not (n339,n340);
nand (n340,n341,n342);
or (n341,n59,n14);
nand (n342,n14,n59);
nand (n343,n322,n9);
nor (n344,n81,n39);
nand (n345,n346,n353);
nand (n346,n347,n352);
or (n347,n348,n129);
not (n348,n349);
nand (n349,n350,n351);
or (n350,n131,n13);
or (n351,n14,n39);
nand (n352,n340,n9);
nor (n353,n354,n131);
and (n354,n13,n9);
nand (n355,n337,n344);
not (n356,n357);
nand (n357,n358,n366);
not (n358,n359);
nand (n359,n360,n365);
or (n360,n361,n72);
not (n361,n362);
nand (n362,n363,n364);
or (n363,n71,n13);
or (n364,n65,n39);
nand (n365,n82,n301);
nor (n366,n367,n369);
and (n367,n318,n368);
not (n368,n326);
and (n369,n319,n326);
nand (n370,n371,n359);
not (n371,n366);
xor (n372,n296,n305);
and (n373,n317,n331);
and (n374,n294,n313);
and (n375,n234,n274);
or (n376,n377,n384);
xor (n377,n378,n383);
xor (n378,n379,n380);
xor (n379,n168,n173);
or (n380,n381,n382);
and (n381,n281,n287);
and (n382,n282,n283);
xor (n383,n28,n91);
or (n384,n385,n386);
and (n385,n275,n280);
and (n386,n276,n279);
not (n387,n388);
nand (n388,n377,n384);
nor (n389,n390,n391);
xor (n390,n25,n150);
or (n391,n392,n393);
and (n392,n378,n383);
and (n393,n379,n380);
nand (n394,n390,n391);
or (n395,n227,n21);
and (n397,n396,n398);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n4);
and (s0n398,notn398,n399);
and (s1n398,n4,n6);
xor (n399,n400,n605);
xor (n400,n401,n603);
xor (n401,n402,n602);
xor (n402,n403,n593);
xor (n403,n404,n592);
xor (n404,n405,n577);
xor (n405,n406,n576);
xor (n406,n407,n556);
xor (n407,n408,n555);
xor (n408,n409,n529);
xor (n409,n410,n528);
xor (n410,n411,n499);
xor (n411,n412,n498);
xor (n412,n413,n460);
xor (n413,n414,n459);
xor (n414,n415,n418);
xor (n415,n416,n417);
and (n416,n202,n9);
and (n417,n140,n14);
or (n418,n419,n422);
and (n419,n420,n421);
and (n420,n140,n9);
and (n421,n135,n14);
and (n422,n423,n424);
xor (n423,n420,n421);
or (n424,n425,n427);
and (n425,n426,n177);
and (n426,n135,n9);
and (n427,n428,n429);
xor (n428,n426,n177);
or (n429,n430,n433);
and (n430,n431,n432);
and (n431,n158,n9);
and (n432,n88,n14);
and (n433,n434,n435);
xor (n434,n431,n432);
or (n435,n436,n439);
and (n436,n437,n438);
and (n437,n88,n9);
and (n438,n69,n14);
and (n439,n440,n441);
xor (n440,n437,n438);
or (n441,n442,n444);
and (n442,n443,n310);
and (n443,n69,n9);
and (n444,n445,n446);
xor (n445,n443,n310);
or (n446,n447,n450);
and (n447,n448,n449);
and (n448,n113,n9);
and (n449,n107,n14);
and (n450,n451,n452);
xor (n451,n448,n449);
or (n452,n453,n456);
and (n453,n454,n455);
and (n454,n107,n9);
and (n455,n8,n14);
and (n456,n457,n458);
xor (n457,n454,n455);
and (n458,n7,n12);
and (n459,n135,n77);
or (n460,n461,n464);
and (n461,n462,n463);
xor (n462,n423,n424);
and (n463,n158,n77);
and (n464,n465,n466);
xor (n465,n462,n463);
or (n466,n467,n470);
and (n467,n468,n469);
xor (n468,n428,n429);
and (n469,n88,n77);
and (n470,n471,n472);
xor (n471,n468,n469);
or (n472,n473,n476);
and (n473,n474,n475);
xor (n474,n434,n435);
and (n475,n69,n77);
and (n476,n477,n478);
xor (n477,n474,n475);
or (n478,n479,n482);
and (n479,n480,n481);
xor (n480,n440,n441);
and (n481,n113,n77);
and (n482,n483,n484);
xor (n483,n480,n481);
or (n484,n485,n488);
and (n485,n486,n487);
xor (n486,n445,n446);
and (n487,n107,n77);
and (n488,n489,n490);
xor (n489,n486,n487);
or (n490,n491,n494);
and (n491,n492,n493);
xor (n492,n451,n452);
and (n493,n8,n77);
and (n494,n495,n496);
xor (n495,n492,n493);
and (n496,n497,n329);
xor (n497,n457,n458);
and (n498,n158,n65);
or (n499,n500,n502);
and (n500,n501,n87);
xor (n501,n465,n466);
and (n502,n503,n504);
xor (n503,n501,n87);
or (n504,n505,n508);
and (n505,n506,n507);
xor (n506,n471,n472);
and (n507,n69,n65);
and (n508,n509,n510);
xor (n509,n506,n507);
or (n510,n511,n513);
and (n511,n512,n245);
xor (n512,n477,n478);
and (n513,n514,n515);
xor (n514,n512,n245);
or (n515,n516,n518);
and (n516,n517,n242);
xor (n517,n483,n484);
and (n518,n519,n520);
xor (n519,n517,n242);
or (n520,n521,n523);
and (n521,n522,n302);
xor (n522,n489,n490);
and (n523,n524,n525);
xor (n524,n522,n302);
and (n525,n526,n527);
xor (n526,n495,n496);
and (n527,n13,n65);
and (n528,n88,n98);
or (n529,n530,n533);
and (n530,n531,n532);
xor (n531,n503,n504);
and (n532,n69,n98);
and (n533,n534,n535);
xor (n534,n531,n532);
or (n535,n536,n539);
and (n536,n537,n538);
xor (n537,n509,n510);
and (n538,n113,n98);
and (n539,n540,n541);
xor (n540,n537,n538);
or (n541,n542,n545);
and (n542,n543,n544);
xor (n543,n514,n515);
and (n544,n107,n98);
and (n545,n546,n547);
xor (n546,n543,n544);
or (n547,n548,n551);
and (n548,n549,n550);
xor (n549,n519,n520);
and (n550,n8,n98);
and (n551,n552,n553);
xor (n552,n549,n550);
and (n553,n554,n262);
xor (n554,n524,n525);
and (n555,n69,n47);
or (n556,n557,n560);
and (n557,n558,n559);
xor (n558,n534,n535);
and (n559,n113,n47);
and (n560,n561,n562);
xor (n561,n558,n559);
or (n562,n563,n566);
and (n563,n564,n565);
xor (n564,n540,n541);
and (n565,n107,n47);
and (n566,n567,n568);
xor (n567,n564,n565);
or (n568,n569,n571);
and (n569,n570,n251);
xor (n570,n546,n547);
and (n571,n572,n573);
xor (n572,n570,n251);
and (n573,n574,n575);
xor (n574,n552,n553);
and (n575,n13,n47);
and (n576,n113,n44);
or (n577,n578,n581);
and (n578,n579,n580);
xor (n579,n561,n562);
and (n580,n107,n44);
and (n581,n582,n583);
xor (n582,n579,n580);
or (n583,n584,n587);
and (n584,n585,n586);
xor (n585,n567,n568);
and (n586,n8,n44);
and (n587,n588,n589);
xor (n588,n585,n586);
and (n589,n590,n591);
xor (n590,n572,n573);
not (n591,n171);
and (n592,n107,n35);
or (n593,n594,n597);
and (n594,n595,n596);
xor (n595,n582,n583);
and (n596,n8,n35);
and (n597,n598,n599);
xor (n598,n595,n596);
and (n599,n600,n601);
xor (n600,n588,n589);
and (n601,n13,n35);
and (n602,n8,n123);
and (n603,n604,n605);
xor (n604,n598,n599);
and (n605,n13,n123);
endmodule
