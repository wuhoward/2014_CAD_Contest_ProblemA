module top (out,n21,n25,n29,n32,n39,n41,n48,n49,n58
        ,n65,n67,n73,n79,n85,n94,n96,n103,n110,n120
        ,n126,n135,n146,n147,n151,n156,n178,n184,n203,n220
        ,n234,n285,n363,n424,n503,n1661,n1662,n1665);
output out;
input n21;
input n25;
input n29;
input n32;
input n39;
input n41;
input n48;
input n49;
input n58;
input n65;
input n67;
input n73;
input n79;
input n85;
input n94;
input n96;
input n103;
input n110;
input n120;
input n126;
input n135;
input n146;
input n147;
input n151;
input n156;
input n178;
input n184;
input n203;
input n220;
input n234;
input n285;
input n363;
input n424;
input n503;
input n1661;
input n1662;
input n1665;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1663;
wire n1664;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
xor (out,n0,n1666);
nand (n0,n1,n1663);
or (n1,n2,n1659);
not (n2,n3);
nor (n3,n4,n1657);
and (n4,n5,n1597);
nand (n5,n6,n1078);
nor (n6,n7,n1064);
and (n7,n8,n739);
and (n8,n9,n604);
nor (n9,n10,n515);
nor (n10,n11,n435);
xor (n11,n12,n343);
xor (n12,n13,n188);
or (n13,n14,n187);
and (n14,n15,n160);
xor (n15,n16,n88);
xor (n16,n17,n60);
xor (n17,n18,n33);
nand (n18,n19,n31);
or (n19,n20,n22);
not (n20,n21);
not (n22,n23);
nor (n23,n24,n26);
not (n24,n25);
nand (n26,n27,n30);
or (n27,n28,n25);
not (n28,n29);
nand (n30,n25,n28);
nand (n31,n26,n32);
nand (n33,n34,n54);
or (n34,n35,n43);
not (n35,n36);
nor (n36,n37,n42);
and (n37,n38,n40);
not (n38,n39);
not (n40,n41);
and (n42,n39,n41);
nand (n43,n44,n51);
not (n44,n45);
nand (n45,n46,n50);
or (n46,n47,n49);
not (n47,n48);
nand (n50,n49,n47);
nand (n51,n52,n53);
nand (n52,n47,n41);
nand (n53,n48,n40);
nand (n54,n45,n55);
nor (n55,n56,n59);
and (n56,n57,n40);
not (n57,n58);
and (n59,n58,n41);
nand (n60,n61,n81);
or (n61,n62,n75);
nand (n62,n63,n69);
nand (n63,n64,n68);
or (n64,n65,n66);
not (n66,n67);
nand (n68,n66,n65);
not (n69,n70);
nand (n70,n71,n74);
or (n71,n72,n65);
not (n72,n73);
nand (n74,n65,n72);
not (n75,n76);
nor (n76,n77,n80);
and (n77,n78,n66);
not (n78,n79);
and (n80,n79,n67);
or (n81,n69,n82);
not (n82,n83);
nor (n83,n84,n86);
and (n84,n85,n67);
and (n86,n87,n66);
not (n87,n85);
xor (n88,n89,n137);
xor (n89,n90,n114);
nand (n90,n91,n106);
or (n91,n92,n99);
nor (n92,n93,n97);
and (n93,n94,n95);
not (n95,n96);
and (n97,n98,n96);
not (n98,n94);
nand (n99,n100,n105);
nor (n100,n101,n104);
and (n101,n102,n41);
not (n102,n103);
and (n104,n103,n40);
xor (n105,n102,n98);
nand (n106,n107,n113);
not (n107,n108);
nor (n108,n109,n111);
and (n109,n98,n110);
and (n111,n112,n94);
not (n112,n110);
not (n113,n100);
nand (n114,n115,n131);
or (n115,n116,n122);
not (n116,n117);
nor (n117,n118,n121);
and (n118,n119,n28);
not (n119,n120);
and (n121,n120,n29);
nand (n122,n123,n128);
not (n123,n124);
nand (n124,n125,n127);
or (n125,n98,n126);
nand (n127,n98,n126);
nand (n128,n129,n130);
or (n129,n126,n28);
nand (n130,n28,n126);
nand (n131,n124,n132);
nand (n132,n133,n136);
or (n133,n29,n134);
not (n134,n135);
or (n136,n28,n135);
not (n137,n138);
nor (n138,n139,n159);
and (n139,n140,n153);
not (n140,n141);
nand (n141,n142,n149);
not (n142,n143);
nand (n143,n144,n148);
or (n144,n145,n147);
not (n145,n146);
nand (n148,n145,n147);
nand (n149,n150,n152);
or (n150,n151,n145);
nand (n152,n145,n151);
nor (n153,n154,n158);
and (n154,n155,n157);
not (n155,n156);
not (n157,n151);
and (n158,n156,n151);
nor (n159,n142,n157);
or (n160,n161,n186);
and (n161,n162,n171);
xor (n162,n163,n138);
nand (n163,n164,n170);
or (n164,n165,n122);
not (n165,n166);
nor (n166,n167,n169);
and (n167,n168,n28);
not (n168,n32);
and (n169,n32,n29);
nand (n170,n124,n117);
nand (n171,n172,n147);
nor (n172,n173,n180);
and (n173,n174,n175);
not (n174,n62);
nor (n175,n176,n179);
and (n176,n177,n66);
not (n177,n178);
and (n179,n178,n67);
and (n180,n70,n181);
nor (n181,n182,n185);
and (n182,n183,n66);
not (n183,n184);
and (n185,n184,n67);
and (n186,n163,n138);
and (n187,n16,n88);
xor (n188,n189,n297);
xor (n189,n190,n248);
xor (n190,n191,n245);
xor (n191,n192,n210);
not (n192,n193);
nand (n193,n194,n209);
or (n194,n195,n199);
not (n195,n196);
nor (n196,n197,n198);
and (n197,n156,n73);
and (n198,n155,n72);
not (n199,n200);
nor (n200,n201,n205);
nand (n201,n202,n204);
or (n202,n157,n203);
nand (n204,n203,n157);
nor (n205,n206,n208);
and (n206,n207,n73);
not (n207,n203);
and (n208,n203,n72);
nand (n209,n201,n73);
or (n210,n211,n244);
and (n211,n212,n223);
xor (n212,n213,n215);
nand (n213,n214,n151);
or (n214,n143,n140);
nand (n215,n216,n222);
or (n216,n217,n199);
not (n217,n218);
nand (n218,n219,n221);
or (n219,n220,n72);
nand (n221,n72,n220);
nand (n222,n196,n201);
nand (n223,n224,n240);
or (n224,n225,n230);
not (n225,n226);
nand (n226,n227,n228);
or (n227,n49,n177);
or (n228,n229,n178);
not (n229,n49);
not (n230,n231);
nor (n231,n232,n237);
nor (n232,n233,n235);
and (n233,n234,n229);
and (n235,n49,n236);
not (n236,n234);
nand (n237,n238,n239);
or (n238,n66,n234);
nand (n239,n234,n66);
nand (n240,n237,n241);
nor (n241,n242,n243);
and (n242,n183,n229);
and (n243,n184,n49);
and (n244,n213,n215);
or (n245,n246,n247);
and (n246,n17,n60);
and (n247,n18,n33);
or (n248,n249,n296);
and (n249,n250,n295);
xor (n250,n251,n272);
or (n251,n252,n271);
and (n252,n253,n265);
xor (n253,n254,n261);
nand (n254,n255,n260);
or (n255,n256,n43);
not (n256,n257);
nand (n257,n258,n259);
or (n258,n110,n40);
nand (n259,n40,n110);
nand (n260,n36,n45);
nand (n261,n262,n264);
or (n262,n263,n62);
not (n263,n181);
nand (n264,n70,n76);
nand (n265,n266,n270);
or (n266,n99,n267);
nor (n267,n268,n269);
and (n268,n135,n98);
and (n269,n94,n134);
or (n270,n92,n100);
and (n271,n254,n261);
or (n272,n273,n294);
and (n273,n274,n287);
xor (n274,n275,n282);
nand (n275,n276,n281);
or (n276,n277,n199);
not (n277,n278);
nor (n278,n279,n280);
and (n279,n87,n72);
and (n280,n85,n73);
nand (n281,n218,n201);
nand (n282,n283,n286);
or (n283,n284,n22);
not (n284,n285);
nand (n286,n26,n21);
nand (n287,n288,n293);
or (n288,n289,n230);
not (n289,n290);
nor (n290,n291,n292);
and (n291,n57,n229);
and (n292,n58,n49);
nand (n293,n237,n226);
and (n294,n275,n282);
xor (n295,n212,n223);
and (n296,n251,n272);
xor (n297,n298,n340);
xor (n298,n299,n316);
xor (n299,n300,n313);
xor (n300,n301,n308);
nand (n301,n302,n304);
or (n302,n303,n230);
not (n303,n241);
nand (n304,n237,n305);
nor (n305,n306,n307);
and (n306,n78,n229);
and (n307,n79,n49);
nand (n308,n309,n311);
or (n309,n310,n122);
not (n310,n132);
nand (n311,n124,n312);
xnor (n312,n95,n29);
nand (n313,n314,n315);
or (n314,n168,n22);
nand (n315,n26,n120);
xor (n316,n317,n332);
xor (n317,n318,n325);
nand (n318,n319,n320);
or (n319,n82,n62);
nand (n320,n70,n321);
nor (n321,n322,n324);
and (n322,n323,n66);
not (n323,n220);
and (n324,n220,n67);
nand (n325,n326,n328);
or (n326,n327,n43);
not (n327,n55);
or (n328,n44,n329);
nor (n329,n330,n331);
and (n330,n177,n41);
and (n331,n178,n40);
nand (n332,n333,n338);
or (n333,n334,n100);
not (n334,n335);
nand (n335,n336,n337);
or (n336,n38,n94);
or (n337,n39,n98);
nand (n338,n107,n339);
not (n339,n99);
or (n340,n341,n342);
and (n341,n89,n137);
and (n342,n90,n114);
or (n343,n344,n434);
and (n344,n345,n399);
xor (n345,n346,n347);
xor (n346,n250,n295);
or (n347,n348,n398);
and (n348,n349,n397);
xor (n349,n350,n374);
or (n350,n351,n373);
and (n351,n352,n365);
xor (n352,n353,n360);
nand (n353,n354,n359);
or (n354,n355,n122);
not (n355,n356);
nor (n356,n357,n358);
and (n357,n20,n28);
and (n358,n21,n29);
nand (n359,n166,n124);
nand (n360,n361,n364);
or (n361,n362,n22);
not (n362,n363);
nand (n364,n26,n285);
nand (n365,n366,n368);
or (n366,n367,n142);
not (n367,n153);
or (n368,n141,n369);
not (n369,n370);
or (n370,n371,n372);
and (n371,n323,n151);
and (n372,n220,n157);
and (n373,n353,n360);
or (n374,n375,n396);
and (n375,n376,n390);
xor (n376,n377,n384);
nand (n377,n378,n383);
or (n378,n379,n230);
not (n379,n380);
nor (n380,n381,n382);
and (n381,n38,n229);
and (n382,n39,n49);
nand (n383,n237,n290);
nand (n384,n385,n389);
or (n385,n386,n199);
nor (n386,n387,n388);
and (n387,n78,n73);
and (n388,n79,n72);
nand (n389,n278,n201);
nand (n390,n391,n395);
or (n391,n43,n392);
nor (n392,n393,n394);
and (n393,n40,n96);
and (n394,n41,n95);
or (n395,n44,n256);
and (n396,n377,n384);
xor (n397,n253,n265);
and (n398,n350,n374);
or (n399,n400,n433);
and (n400,n401,n404);
xor (n401,n402,n403);
xor (n402,n274,n287);
xor (n403,n162,n171);
and (n404,n405,n427);
or (n405,n406,n426);
and (n406,n407,n421);
xor (n407,n408,n414);
nand (n408,n409,n413);
or (n409,n410,n62);
nor (n410,n411,n412);
and (n411,n57,n67);
and (n412,n58,n66);
nand (n413,n175,n70);
nand (n414,n415,n420);
or (n415,n416,n122);
not (n416,n417);
nand (n417,n418,n419);
or (n418,n29,n284);
or (n419,n28,n285);
nand (n420,n124,n356);
nand (n421,n422,n425);
or (n422,n423,n22);
not (n423,n424);
nand (n425,n26,n363);
and (n426,n408,n414);
nand (n427,n428,n432);
or (n428,n99,n429);
nor (n429,n430,n431);
and (n430,n98,n120);
and (n431,n94,n119);
or (n432,n100,n267);
and (n433,n402,n403);
and (n434,n346,n347);
or (n435,n436,n514);
and (n436,n437,n440);
xor (n437,n438,n439);
xor (n438,n15,n160);
xor (n439,n345,n399);
or (n440,n441,n513);
and (n441,n442,n477);
xor (n442,n443,n444);
xor (n443,n349,n397);
or (n444,n445,n476);
and (n445,n446,n474);
xor (n446,n447,n473);
or (n447,n448,n472);
and (n448,n449,n464);
xor (n449,n450,n457);
nand (n450,n451,n456);
or (n451,n452,n141);
not (n452,n453);
nor (n453,n454,n455);
and (n454,n87,n157);
and (n455,n85,n151);
nand (n456,n143,n370);
nand (n457,n458,n463);
or (n458,n459,n230);
not (n459,n460);
nand (n460,n461,n462);
or (n461,n49,n112);
or (n462,n229,n110);
nand (n463,n237,n380);
nand (n464,n465,n470);
or (n465,n199,n466);
not (n466,n467);
nor (n467,n468,n469);
and (n468,n72,n183);
and (n469,n184,n73);
or (n470,n386,n471);
not (n471,n201);
and (n472,n450,n457);
xor (n473,n376,n390);
nand (n474,n475,n171);
or (n475,n147,n172);
and (n476,n447,n473);
or (n477,n478,n512);
and (n478,n479,n511);
xor (n479,n480,n481);
xor (n480,n352,n365);
or (n481,n482,n510);
and (n482,n483,n499);
xor (n483,n484,n492);
nand (n484,n485,n490);
or (n485,n486,n43);
not (n486,n487);
nor (n487,n488,n489);
and (n488,n134,n40);
and (n489,n135,n41);
nand (n490,n491,n45);
not (n491,n392);
nand (n492,n493,n498);
or (n493,n494,n99);
not (n494,n495);
nand (n495,n496,n497);
or (n496,n94,n168);
or (n497,n98,n32);
or (n498,n100,n429);
nand (n499,n500,n509);
or (n500,n501,n504);
nand (n501,n502,n147);
not (n502,n503);
not (n504,n505);
nor (n505,n506,n508);
and (n506,n155,n507);
not (n507,n147);
and (n508,n156,n147);
or (n509,n507,n502);
and (n510,n484,n492);
xor (n511,n405,n427);
and (n512,n480,n481);
and (n513,n443,n444);
and (n514,n438,n439);
nor (n515,n516,n517);
xor (n516,n437,n440);
or (n517,n518,n603);
and (n518,n519,n602);
xor (n519,n520,n521);
xor (n520,n401,n404);
or (n521,n522,n601);
and (n522,n523,n600);
xor (n523,n524,n593);
or (n524,n525,n592);
and (n525,n526,n568);
xor (n526,n527,n545);
or (n527,n528,n544);
and (n528,n529,n537);
xor (n529,n530,n531);
and (n530,n26,n424);
nand (n531,n532,n533);
or (n532,n502,n504);
or (n533,n534,n501);
nor (n534,n535,n536);
and (n535,n507,n220);
and (n536,n147,n323);
nand (n537,n538,n543);
or (n538,n141,n539);
not (n539,n540);
nor (n540,n541,n542);
and (n541,n78,n157);
and (n542,n79,n151);
nand (n543,n143,n453);
and (n544,n530,n531);
or (n545,n546,n567);
and (n546,n547,n561);
xor (n547,n548,n555);
nand (n548,n549,n554);
or (n549,n550,n199);
not (n550,n551);
nand (n551,n552,n553);
or (n552,n73,n177);
or (n553,n72,n178);
nand (n554,n467,n201);
nand (n555,n556,n560);
or (n556,n557,n43);
nor (n557,n558,n559);
and (n558,n119,n41);
and (n559,n120,n40);
nand (n560,n487,n45);
nand (n561,n562,n563);
or (n562,n494,n100);
or (n563,n99,n564);
nor (n564,n565,n566);
and (n565,n21,n98);
and (n566,n94,n20);
and (n567,n548,n555);
or (n568,n569,n591);
and (n569,n570,n584);
xor (n570,n571,n578);
nand (n571,n572,n577);
or (n572,n573,n122);
not (n573,n574);
nand (n574,n575,n576);
or (n575,n29,n362);
or (n576,n28,n363);
nand (n577,n417,n124);
nand (n578,n579,n583);
or (n579,n62,n580);
nor (n580,n581,n582);
and (n581,n38,n67);
and (n582,n39,n66);
or (n583,n69,n410);
nand (n584,n585,n589);
or (n585,n230,n586);
nor (n586,n587,n588);
and (n587,n95,n49);
and (n588,n96,n229);
or (n589,n590,n459);
not (n590,n237);
and (n591,n571,n578);
and (n592,n527,n545);
or (n593,n594,n599);
and (n594,n595,n598);
xor (n595,n596,n597);
xor (n596,n407,n421);
xor (n597,n449,n464);
xor (n598,n483,n499);
and (n599,n596,n597);
xor (n600,n446,n474);
and (n601,n524,n593);
xor (n602,n442,n477);
and (n603,n520,n521);
nor (n604,n605,n677);
nor (n605,n606,n674);
xor (n606,n607,n671);
xor (n607,n608,n654);
xor (n608,n609,n637);
xor (n609,n610,n613);
or (n610,n611,n612);
and (n611,n300,n313);
and (n612,n301,n308);
xor (n613,n614,n629);
xor (n614,n615,n622);
nand (n615,n616,n617);
or (n616,n334,n99);
nand (n617,n618,n113);
not (n618,n619);
nor (n619,n620,n621);
and (n620,n58,n98);
and (n621,n94,n57);
nand (n622,n623,n625);
or (n623,n624,n230);
not (n624,n305);
or (n625,n590,n626);
nor (n626,n627,n628);
and (n627,n87,n49);
and (n628,n85,n229);
nand (n629,n630,n632);
or (n630,n122,n631);
not (n631,n312);
or (n632,n123,n633);
not (n633,n634);
nor (n634,n635,n636);
and (n635,n112,n28);
and (n636,n110,n29);
xor (n637,n638,n648);
xor (n638,n639,n641);
nand (n639,n640,n73);
or (n640,n201,n200);
nand (n641,n642,n644);
or (n642,n62,n643);
not (n643,n321);
or (n644,n69,n645);
nor (n645,n646,n647);
and (n646,n66,n156);
and (n647,n67,n155);
nand (n648,n649,n650);
or (n649,n43,n329);
or (n650,n44,n651);
nor (n651,n652,n653);
and (n652,n40,n184);
and (n653,n41,n183);
xor (n654,n655,n668);
xor (n655,n656,n665);
xor (n656,n657,n662);
xor (n657,n658,n193);
nand (n658,n659,n660);
or (n659,n22,n119);
or (n660,n661,n134);
not (n661,n26);
or (n662,n663,n664);
and (n663,n317,n332);
and (n664,n318,n325);
or (n665,n666,n667);
and (n666,n191,n245);
and (n667,n192,n210);
or (n668,n669,n670);
and (n669,n298,n340);
and (n670,n299,n316);
or (n671,n672,n673);
and (n672,n189,n297);
and (n673,n190,n248);
or (n674,n675,n676);
and (n675,n12,n343);
and (n676,n13,n188);
nor (n677,n678,n736);
xor (n678,n679,n733);
xor (n679,n680,n707);
xor (n680,n681,n688);
xor (n681,n682,n685);
or (n682,n683,n684);
and (n683,n614,n629);
and (n684,n615,n622);
or (n685,n686,n687);
and (n686,n638,n648);
and (n687,n639,n641);
xor (n688,n689,n704);
xor (n689,n690,n696);
nand (n690,n691,n692);
or (n691,n99,n619);
or (n692,n693,n100);
nor (n693,n694,n695);
and (n694,n178,n98);
and (n695,n94,n177);
nand (n696,n697,n702);
or (n697,n698,n123);
not (n698,n699);
nor (n699,n700,n701);
and (n700,n38,n28);
and (n701,n39,n29);
nand (n702,n703,n634);
not (n703,n122);
nand (n704,n705,n706);
or (n705,n62,n645);
or (n706,n69,n66);
xor (n707,n708,n730);
xor (n708,n709,n727);
xor (n709,n710,n720);
xor (n710,n711,n714);
nand (n711,n712,n713);
or (n712,n22,n134);
or (n713,n661,n95);
nand (n714,n715,n716);
or (n715,n651,n43);
or (n716,n44,n717);
nor (n717,n718,n719);
and (n718,n40,n79);
and (n719,n41,n78);
not (n720,n721);
nand (n721,n722,n723);
or (n722,n230,n626);
or (n723,n590,n724);
nor (n724,n725,n726);
and (n725,n323,n49);
and (n726,n220,n229);
or (n727,n728,n729);
and (n728,n657,n662);
and (n729,n658,n193);
or (n730,n731,n732);
and (n731,n609,n637);
and (n732,n610,n613);
or (n733,n734,n735);
and (n734,n655,n668);
and (n735,n656,n665);
or (n736,n737,n738);
and (n737,n607,n671);
and (n738,n608,n654);
nand (n739,n740,n1058);
or (n740,n741,n1040);
not (n741,n742);
nor (n742,n743,n1039);
and (n743,n744,n980);
nand (n744,n745,n888);
xor (n745,n746,n875);
xor (n746,n747,n748);
xor (n747,n595,n598);
or (n748,n749,n874);
and (n749,n750,n845);
xor (n750,n751,n798);
or (n751,n752,n797);
and (n752,n753,n773);
xor (n753,n754,n760);
nand (n754,n755,n759);
or (n755,n99,n756);
nor (n756,n757,n758);
and (n757,n98,n285);
and (n758,n94,n284);
or (n759,n100,n564);
xor (n760,n761,n767);
nor (n761,n762,n28);
nor (n762,n763,n765);
and (n763,n764,n98);
nand (n764,n424,n126);
and (n765,n423,n766);
not (n766,n126);
nand (n767,n768,n772);
or (n768,n769,n501);
nor (n769,n770,n771);
and (n770,n87,n147);
and (n771,n85,n507);
or (n772,n534,n502);
or (n773,n774,n796);
and (n774,n775,n785);
xor (n775,n776,n777);
nor (n776,n123,n423);
nand (n777,n778,n783);
or (n778,n501,n779);
not (n779,n780);
nor (n780,n781,n782);
and (n781,n78,n507);
and (n782,n79,n147);
nand (n783,n784,n503);
not (n784,n769);
nand (n785,n786,n791);
or (n786,n141,n787);
not (n787,n788);
nand (n788,n789,n790);
or (n789,n151,n177);
or (n790,n157,n178);
or (n791,n142,n792);
not (n792,n793);
nand (n793,n794,n795);
or (n794,n151,n183);
or (n795,n157,n184);
and (n796,n776,n777);
and (n797,n754,n760);
xor (n798,n799,n822);
xor (n799,n800,n801);
and (n800,n761,n767);
or (n801,n802,n821);
and (n802,n803,n814);
xor (n803,n804,n807);
nand (n804,n805,n806);
or (n805,n792,n141);
nand (n806,n143,n540);
nand (n807,n808,n813);
or (n808,n809,n122);
not (n809,n810);
nand (n810,n811,n812);
or (n811,n28,n424);
or (n812,n29,n423);
nand (n813,n574,n124);
nand (n814,n815,n820);
or (n815,n62,n816);
not (n816,n817);
nor (n817,n818,n819);
and (n818,n112,n66);
and (n819,n110,n67);
or (n820,n69,n580);
and (n821,n804,n807);
or (n822,n823,n844);
and (n823,n824,n838);
xor (n824,n825,n832);
nand (n825,n826,n831);
or (n826,n827,n230);
not (n827,n828);
nor (n828,n829,n830);
and (n829,n134,n229);
and (n830,n135,n49);
or (n831,n586,n590);
nand (n832,n833,n837);
or (n833,n834,n199);
nor (n834,n835,n836);
and (n835,n72,n58);
and (n836,n73,n57);
nand (n837,n201,n551);
nand (n838,n839,n843);
or (n839,n43,n840);
nor (n840,n841,n842);
and (n841,n40,n32);
and (n842,n41,n168);
or (n843,n44,n557);
and (n844,n825,n832);
or (n845,n846,n873);
and (n846,n847,n872);
xor (n847,n848,n871);
or (n848,n849,n870);
and (n849,n850,n864);
xor (n850,n851,n858);
nand (n851,n852,n857);
or (n852,n853,n62);
not (n853,n854);
nand (n854,n855,n856);
or (n855,n67,n95);
or (n856,n66,n96);
nand (n857,n70,n817);
nand (n858,n859,n863);
or (n859,n230,n860);
nor (n860,n861,n862);
and (n861,n229,n120);
and (n862,n49,n119);
nand (n863,n237,n828);
nand (n864,n865,n869);
or (n865,n199,n866);
nor (n866,n867,n868);
and (n867,n72,n39);
and (n868,n73,n38);
or (n869,n834,n471);
and (n870,n851,n858);
xor (n871,n824,n838);
xor (n872,n803,n814);
and (n873,n848,n871);
and (n874,n751,n798);
xor (n875,n876,n881);
xor (n876,n877,n880);
or (n877,n878,n879);
and (n878,n799,n822);
and (n879,n800,n801);
xor (n880,n526,n568);
or (n881,n882,n887);
and (n882,n883,n886);
xor (n883,n884,n885);
xor (n884,n547,n561);
xor (n885,n529,n537);
xor (n886,n570,n584);
and (n887,n884,n885);
or (n888,n889,n979);
and (n889,n890,n978);
xor (n890,n891,n892);
xor (n891,n883,n886);
or (n892,n893,n977);
and (n893,n894,n925);
xor (n894,n895,n924);
or (n895,n896,n923);
and (n896,n897,n911);
xor (n897,n898,n905);
nand (n898,n899,n903);
or (n899,n900,n43);
nor (n900,n901,n902);
and (n901,n20,n41);
and (n902,n21,n40);
nand (n903,n904,n45);
not (n904,n840);
nand (n905,n906,n910);
or (n906,n907,n99);
nor (n907,n908,n909);
and (n908,n98,n363);
and (n909,n94,n362);
or (n910,n100,n756);
and (n911,n912,n917);
nor (n912,n913,n98);
nor (n913,n914,n916);
and (n914,n915,n40);
nand (n915,n424,n103);
and (n916,n423,n102);
nand (n917,n918,n919);
or (n918,n502,n779);
or (n919,n920,n501);
nor (n920,n921,n922);
and (n921,n183,n147);
and (n922,n184,n507);
and (n923,n898,n905);
xor (n924,n753,n773);
or (n925,n926,n976);
and (n926,n927,n975);
xor (n927,n928,n953);
or (n928,n929,n952);
and (n929,n930,n945);
xor (n930,n931,n938);
nand (n931,n932,n937);
or (n932,n933,n141);
not (n933,n934);
nor (n934,n935,n936);
and (n935,n57,n157);
and (n936,n58,n151);
nand (n937,n788,n143);
nand (n938,n939,n944);
or (n939,n940,n62);
not (n940,n941);
nand (n941,n942,n943);
or (n942,n67,n134);
or (n943,n66,n135);
nand (n944,n70,n854);
nand (n945,n946,n951);
or (n946,n230,n947);
not (n947,n948);
nand (n948,n949,n950);
or (n949,n49,n168);
or (n950,n229,n32);
or (n951,n590,n860);
and (n952,n931,n938);
or (n953,n954,n974);
and (n954,n955,n968);
xor (n955,n956,n962);
nand (n956,n957,n961);
or (n957,n199,n958);
nor (n958,n959,n960);
and (n959,n72,n110);
and (n960,n73,n112);
or (n961,n866,n471);
nand (n962,n963,n967);
or (n963,n43,n964);
nor (n964,n965,n966);
and (n965,n40,n285);
and (n966,n41,n284);
or (n967,n900,n44);
nand (n968,n969,n973);
or (n969,n99,n970);
nor (n970,n971,n972);
and (n971,n423,n94);
and (n972,n424,n98);
or (n973,n907,n100);
and (n974,n956,n962);
xor (n975,n775,n785);
and (n976,n928,n953);
and (n977,n895,n924);
xor (n978,n750,n845);
and (n979,n891,n892);
nand (n980,n981,n982);
xor (n981,n890,n978);
or (n982,n983,n1038);
and (n983,n984,n1037);
xor (n984,n985,n986);
xor (n985,n847,n872);
or (n986,n987,n1036);
and (n987,n988,n991);
xor (n988,n989,n990);
xor (n989,n850,n864);
xor (n990,n897,n911);
or (n991,n992,n1035);
and (n992,n993,n1013);
xor (n993,n994,n995);
xor (n994,n912,n917);
or (n995,n996,n1012);
and (n996,n997,n1006);
xor (n997,n998,n999);
and (n998,n113,n424);
nand (n999,n1000,n1005);
or (n1000,n1001,n141);
not (n1001,n1002);
nand (n1002,n1003,n1004);
or (n1003,n151,n38);
or (n1004,n157,n39);
nand (n1005,n143,n934);
nand (n1006,n1007,n1008);
or (n1007,n940,n69);
or (n1008,n62,n1009);
nor (n1009,n1010,n1011);
and (n1010,n119,n67);
and (n1011,n120,n66);
and (n1012,n998,n999);
or (n1013,n1014,n1034);
and (n1014,n1015,n1028);
xor (n1015,n1016,n1022);
nand (n1016,n1017,n1021);
or (n1017,n1018,n230);
nor (n1018,n1019,n1020);
and (n1019,n20,n49);
and (n1020,n21,n229);
nand (n1021,n948,n237);
nand (n1022,n1023,n1027);
or (n1023,n1024,n501);
nor (n1024,n1025,n1026);
and (n1025,n507,n178);
and (n1026,n147,n177);
or (n1027,n920,n502);
nand (n1028,n1029,n1033);
or (n1029,n1030,n43);
nor (n1030,n1031,n1032);
and (n1031,n40,n363);
and (n1032,n41,n362);
or (n1033,n964,n44);
and (n1034,n1016,n1022);
and (n1035,n994,n995);
and (n1036,n989,n990);
xor (n1037,n894,n925);
and (n1038,n985,n986);
nor (n1039,n745,n888);
not (n1040,n1041);
nor (n1041,n1042,n1053);
nor (n1042,n1043,n1044);
xor (n1043,n519,n602);
or (n1044,n1045,n1052);
and (n1045,n1046,n1051);
xor (n1046,n1047,n1048);
xor (n1047,n479,n511);
or (n1048,n1049,n1050);
and (n1049,n876,n881);
and (n1050,n877,n880);
xor (n1051,n523,n600);
and (n1052,n1047,n1048);
nor (n1053,n1054,n1055);
xor (n1054,n1046,n1051);
or (n1055,n1056,n1057);
and (n1056,n746,n875);
and (n1057,n747,n748);
nor (n1058,n1059,n1063);
and (n1059,n1060,n1061);
not (n1060,n1042);
not (n1061,n1062);
nand (n1062,n1054,n1055);
and (n1063,n1043,n1044);
nand (n1064,n1065,n1072);
or (n1065,n1066,n1067);
not (n1066,n604);
not (n1067,n1068);
nor (n1068,n1069,n10);
and (n1069,n1070,n1071);
nand (n1070,n435,n11);
nand (n1071,n516,n517);
nor (n1072,n1073,n1077);
and (n1073,n1074,n1075);
not (n1074,n677);
not (n1075,n1076);
nand (n1076,n606,n674);
and (n1077,n678,n736);
nand (n1078,n8,n1079,n1082);
and (n1079,n1041,n1080);
nor (n1080,n1039,n1081);
nor (n1081,n981,n982);
nand (n1082,n1083,n1584);
or (n1083,n1084,n1520);
not (n1084,n1085);
nand (n1085,n1086,n1509,n1519);
nand (n1086,n1087,n1265,n1369);
nand (n1087,n1088,n1229);
not (n1088,n1089);
xor (n1089,n1090,n1188);
xor (n1090,n1091,n1126);
xor (n1091,n1092,n1108);
xor (n1092,n1093,n1099);
nand (n1093,n1094,n1098);
or (n1094,n43,n1095);
nor (n1095,n1096,n1097);
and (n1096,n423,n41);
and (n1097,n40,n424);
or (n1098,n44,n1030);
nand (n1099,n1100,n1104);
or (n1100,n199,n1101);
nor (n1101,n1102,n1103);
and (n1102,n72,n135);
and (n1103,n73,n134);
or (n1104,n1105,n471);
nor (n1105,n1106,n1107);
and (n1106,n72,n96);
and (n1107,n73,n95);
nand (n1108,n1109,n1125);
or (n1109,n1110,n1117);
not (n1110,n1111);
nand (n1111,n1112,n41);
nand (n1112,n1113,n1114);
or (n1113,n424,n48);
nand (n1114,n1115,n229);
not (n1115,n1116);
and (n1116,n424,n48);
not (n1117,n1118);
nand (n1118,n1119,n1124);
or (n1119,n1120,n141);
not (n1120,n1121);
nand (n1121,n1122,n1123);
or (n1122,n151,n112);
or (n1123,n157,n110);
nand (n1124,n143,n1002);
or (n1125,n1118,n1111);
xor (n1126,n1127,n1177);
xor (n1127,n1128,n1149);
or (n1128,n1129,n1148);
and (n1129,n1130,n1138);
xor (n1130,n1131,n1132);
and (n1131,n45,n424);
nand (n1132,n1133,n1137);
or (n1133,n1134,n141);
nor (n1134,n1135,n1136);
and (n1135,n95,n151);
and (n1136,n96,n157);
nand (n1137,n143,n1121);
nand (n1138,n1139,n1144);
or (n1139,n62,n1140);
not (n1140,n1141);
nor (n1141,n1142,n1143);
and (n1142,n20,n66);
and (n1143,n21,n67);
or (n1144,n69,n1145);
nor (n1145,n1146,n1147);
and (n1146,n32,n66);
and (n1147,n168,n67);
and (n1148,n1131,n1132);
or (n1149,n1150,n1176);
and (n1150,n1151,n1170);
xor (n1151,n1152,n1161);
nand (n1152,n1153,n1157);
or (n1153,n230,n1154);
nor (n1154,n1155,n1156);
and (n1155,n362,n49);
and (n1156,n363,n229);
or (n1157,n590,n1158);
nor (n1158,n1159,n1160);
and (n1159,n285,n229);
and (n1160,n284,n49);
nand (n1161,n1162,n1166);
or (n1162,n1163,n501);
nor (n1163,n1164,n1165);
and (n1164,n507,n39);
and (n1165,n147,n38);
or (n1166,n1167,n502);
nor (n1167,n1168,n1169);
and (n1168,n507,n58);
and (n1169,n147,n57);
nand (n1170,n1171,n1175);
or (n1171,n199,n1172);
nor (n1172,n1173,n1174);
and (n1173,n72,n120);
and (n1174,n73,n119);
or (n1175,n1101,n471);
and (n1176,n1152,n1161);
xor (n1177,n1178,n1185);
xor (n1178,n1179,n1182);
nand (n1179,n1180,n1181);
or (n1180,n62,n1145);
or (n1181,n1009,n69);
nand (n1182,n1183,n1184);
or (n1183,n230,n1158);
or (n1184,n590,n1018);
nand (n1185,n1186,n1187);
or (n1186,n1167,n501);
or (n1187,n1024,n502);
or (n1188,n1189,n1228);
and (n1189,n1190,n1227);
xor (n1190,n1191,n1204);
and (n1191,n1192,n1198);
and (n1192,n1193,n49);
nand (n1193,n1194,n1195);
or (n1194,n424,n234);
nand (n1195,n1196,n66);
not (n1196,n1197);
and (n1197,n424,n234);
nand (n1198,n1199,n1203);
or (n1199,n141,n1200);
nor (n1200,n1201,n1202);
and (n1201,n157,n135);
and (n1202,n151,n134);
or (n1203,n142,n1134);
or (n1204,n1205,n1226);
and (n1205,n1206,n1220);
xor (n1206,n1207,n1214);
nand (n1207,n1208,n1213);
or (n1208,n1209,n62);
not (n1209,n1210);
nor (n1210,n1211,n1212);
and (n1211,n285,n67);
and (n1212,n284,n66);
nand (n1213,n70,n1141);
nand (n1214,n1215,n1219);
or (n1215,n230,n1216);
nor (n1216,n1217,n1218);
and (n1217,n49,n423);
and (n1218,n229,n424);
or (n1219,n590,n1154);
nand (n1220,n1221,n1225);
or (n1221,n501,n1222);
nor (n1222,n1223,n1224);
and (n1223,n507,n110);
and (n1224,n147,n112);
or (n1225,n1163,n502);
and (n1226,n1207,n1214);
xor (n1227,n1130,n1138);
and (n1228,n1191,n1204);
not (n1229,n1230);
or (n1230,n1231,n1264);
and (n1231,n1232,n1263);
xor (n1232,n1233,n1234);
xor (n1233,n1151,n1170);
or (n1234,n1235,n1262);
and (n1235,n1236,n1244);
xor (n1236,n1237,n1243);
nand (n1237,n1238,n1242);
or (n1238,n199,n1239);
nor (n1239,n1240,n1241);
and (n1240,n72,n32);
and (n1241,n73,n168);
or (n1242,n1172,n471);
xor (n1243,n1192,n1198);
or (n1244,n1245,n1261);
and (n1245,n1246,n1254);
xor (n1246,n1247,n1248);
and (n1247,n237,n424);
nand (n1248,n1249,n1253);
or (n1249,n1250,n501);
nor (n1250,n1251,n1252);
and (n1251,n507,n96);
and (n1252,n147,n95);
or (n1253,n1222,n502);
nand (n1254,n1255,n1260);
or (n1255,n62,n1256);
not (n1256,n1257);
nand (n1257,n1258,n1259);
or (n1258,n67,n362);
or (n1259,n66,n363);
or (n1260,n69,n1209);
and (n1261,n1247,n1248);
and (n1262,n1237,n1243);
xor (n1263,n1190,n1227);
and (n1264,n1233,n1234);
nor (n1265,n1266,n1306);
not (n1266,n1267);
or (n1267,n1268,n1269);
xor (n1268,n1232,n1263);
or (n1269,n1270,n1305);
and (n1270,n1271,n1304);
xor (n1271,n1272,n1273);
xor (n1272,n1206,n1220);
or (n1273,n1274,n1303);
and (n1274,n1275,n1288);
xor (n1275,n1276,n1282);
nand (n1276,n1277,n1281);
or (n1277,n141,n1278);
nor (n1278,n1279,n1280);
and (n1279,n157,n120);
and (n1280,n151,n119);
or (n1281,n142,n1200);
nand (n1282,n1283,n1287);
or (n1283,n199,n1284);
nor (n1284,n1285,n1286);
and (n1285,n72,n21);
and (n1286,n73,n20);
or (n1287,n1239,n471);
and (n1288,n1289,n1296);
nor (n1289,n1290,n66);
nor (n1290,n1291,n1294);
and (n1291,n1292,n72);
not (n1292,n1293);
and (n1293,n424,n65);
and (n1294,n423,n1295);
not (n1295,n65);
nand (n1296,n1297,n1302);
or (n1297,n501,n1298);
not (n1298,n1299);
nor (n1299,n1300,n1301);
and (n1300,n135,n147);
and (n1301,n134,n507);
or (n1302,n1250,n502);
and (n1303,n1276,n1282);
xor (n1304,n1236,n1244);
and (n1305,n1272,n1273);
nand (n1306,n1307,n1363);
not (n1307,n1308);
nor (n1308,n1309,n1338);
xor (n1309,n1310,n1337);
xor (n1310,n1311,n1336);
or (n1311,n1312,n1335);
and (n1312,n1313,n1329);
xor (n1313,n1314,n1321);
nand (n1314,n1315,n1320);
or (n1315,n1316,n62);
not (n1316,n1317);
nand (n1317,n1318,n1319);
or (n1318,n66,n424);
or (n1319,n67,n423);
nand (n1320,n70,n1257);
nand (n1321,n1322,n1327);
or (n1322,n1323,n141);
not (n1323,n1324);
nand (n1324,n1325,n1326);
or (n1325,n151,n168);
or (n1326,n157,n32);
nand (n1327,n1328,n143);
not (n1328,n1278);
nand (n1329,n1330,n1334);
or (n1330,n199,n1331);
nor (n1331,n1332,n1333);
and (n1332,n72,n285);
and (n1333,n73,n284);
or (n1334,n1284,n471);
and (n1335,n1314,n1321);
xor (n1336,n1246,n1254);
xor (n1337,n1275,n1288);
or (n1338,n1339,n1362);
and (n1339,n1340,n1361);
xor (n1340,n1341,n1342);
xor (n1341,n1289,n1296);
or (n1342,n1343,n1360);
and (n1343,n1344,n1353);
xor (n1344,n1345,n1346);
and (n1345,n70,n424);
nand (n1346,n1347,n1348);
or (n1347,n502,n1298);
or (n1348,n1349,n501);
not (n1349,n1350);
nand (n1350,n1351,n1352);
or (n1351,n120,n507);
nand (n1352,n507,n120);
nand (n1353,n1354,n1359);
or (n1354,n1355,n141);
not (n1355,n1356);
nand (n1356,n1357,n1358);
or (n1357,n151,n20);
or (n1358,n157,n21);
nand (n1359,n143,n1324);
and (n1360,n1345,n1346);
xor (n1361,n1313,n1329);
and (n1362,n1341,n1342);
not (n1363,n1364);
nor (n1364,n1365,n1366);
xor (n1365,n1271,n1304);
or (n1366,n1367,n1368);
and (n1367,n1310,n1337);
and (n1368,n1311,n1336);
or (n1369,n1370,n1508);
and (n1370,n1371,n1398);
xor (n1371,n1372,n1397);
or (n1372,n1373,n1396);
and (n1373,n1374,n1395);
xor (n1374,n1375,n1381);
nand (n1375,n1376,n1380);
or (n1376,n199,n1377);
nor (n1377,n1378,n1379);
and (n1378,n72,n363);
and (n1379,n73,n362);
or (n1380,n1331,n471);
nor (n1381,n1382,n1390);
not (n1382,n1383);
nand (n1383,n1384,n1389);
or (n1384,n501,n1385);
not (n1385,n1386);
nor (n1386,n1387,n1388);
and (n1387,n32,n147);
and (n1388,n168,n507);
nand (n1389,n1350,n503);
nand (n1390,n1391,n73);
nand (n1391,n1392,n1394);
or (n1392,n1393,n151);
and (n1393,n424,n203);
or (n1394,n424,n203);
xor (n1395,n1344,n1353);
and (n1396,n1375,n1381);
xor (n1397,n1340,n1361);
or (n1398,n1399,n1507);
and (n1399,n1400,n1424);
xor (n1400,n1401,n1423);
or (n1401,n1402,n1422);
and (n1402,n1403,n1418);
xor (n1403,n1404,n1411);
nand (n1404,n1405,n1410);
or (n1405,n1406,n141);
not (n1406,n1407);
nor (n1407,n1408,n1409);
and (n1408,n284,n157);
and (n1409,n285,n151);
nand (n1410,n143,n1356);
nand (n1411,n1412,n1417);
or (n1412,n1413,n199);
not (n1413,n1414);
nand (n1414,n1415,n1416);
or (n1415,n72,n424);
or (n1416,n423,n73);
or (n1417,n1377,n471);
nand (n1418,n1419,n1421);
or (n1419,n1420,n1382);
not (n1420,n1390);
or (n1421,n1383,n1390);
and (n1422,n1404,n1411);
xor (n1423,n1374,n1395);
or (n1424,n1425,n1506);
and (n1425,n1426,n1447);
xor (n1426,n1427,n1446);
or (n1427,n1428,n1445);
and (n1428,n1429,n1438);
xor (n1429,n1430,n1431);
and (n1430,n201,n424);
nand (n1431,n1432,n1437);
or (n1432,n1433,n141);
not (n1433,n1434);
nor (n1434,n1435,n1436);
and (n1435,n362,n157);
and (n1436,n363,n151);
nand (n1437,n143,n1407);
nand (n1438,n1439,n1440);
or (n1439,n502,n1385);
or (n1440,n501,n1441);
not (n1441,n1442);
nor (n1442,n1443,n1444);
and (n1443,n20,n507);
and (n1444,n21,n147);
and (n1445,n1430,n1431);
xor (n1446,n1403,n1418);
nand (n1447,n1448,n1505);
or (n1448,n1449,n1465);
nor (n1449,n1450,n1451);
xor (n1450,n1429,n1438);
and (n1451,n1452,n1459);
nand (n1452,n1453,n1454);
nand (n1453,n1442,n503);
nand (n1454,n1455,n1458);
nor (n1455,n1456,n1457);
and (n1456,n284,n507);
and (n1457,n285,n147);
not (n1458,n501);
not (n1459,n1460);
nand (n1460,n1461,n151);
nand (n1461,n1462,n1464);
or (n1462,n1463,n147);
and (n1463,n424,n146);
or (n1464,n424,n146);
nor (n1465,n1466,n1504);
and (n1466,n1467,n1478);
nand (n1467,n1468,n1472);
nor (n1468,n1469,n1471);
and (n1469,n1470,n1459);
not (n1470,n1452);
and (n1471,n1452,n1460);
nor (n1472,n1473,n1474);
and (n1473,n143,n1434);
and (n1474,n140,n1475);
nand (n1475,n1476,n1477);
or (n1476,n157,n424);
or (n1477,n423,n151);
nand (n1478,n1479,n1502);
or (n1479,n1480,n1494);
not (n1480,n1481);
and (n1481,n1482,n1492);
nand (n1482,n1483,n1488);
or (n1483,n502,n1484);
not (n1484,n1485);
nor (n1485,n1486,n1487);
and (n1486,n362,n507);
and (n1487,n363,n147);
nand (n1488,n1489,n1458);
nand (n1489,n1490,n1491);
or (n1490,n507,n424);
or (n1491,n147,n423);
nor (n1492,n1493,n507);
and (n1493,n424,n503);
not (n1494,n1495);
nand (n1495,n1496,n1501);
not (n1496,n1497);
nand (n1497,n1498,n1500);
or (n1498,n502,n1499);
not (n1499,n1455);
nand (n1500,n1485,n1458);
nand (n1501,n143,n424);
nand (n1502,n1503,n1497);
not (n1503,n1501);
nor (n1504,n1468,n1472);
nand (n1505,n1450,n1451);
and (n1506,n1427,n1446);
and (n1507,n1401,n1423);
and (n1508,n1372,n1397);
nand (n1509,n1510,n1087);
or (n1510,n1511,n1513);
not (n1511,n1512);
nand (n1512,n1268,n1269);
not (n1513,n1514);
nand (n1514,n1267,n1515);
nand (n1515,n1516,n1518);
or (n1516,n1364,n1517);
nand (n1517,n1309,n1338);
nand (n1518,n1365,n1366);
nand (n1519,n1089,n1230);
not (n1520,n1521);
nor (n1521,n1522,n1547);
nor (n1522,n1523,n1524);
xor (n1523,n984,n1037);
or (n1524,n1525,n1546);
and (n1525,n1526,n1529);
xor (n1526,n1527,n1528);
xor (n1527,n927,n975);
xor (n1528,n988,n991);
or (n1529,n1530,n1545);
and (n1530,n1531,n1534);
xor (n1531,n1532,n1533);
xor (n1532,n955,n968);
xor (n1533,n930,n945);
or (n1534,n1535,n1544);
and (n1535,n1536,n1541);
xor (n1536,n1537,n1540);
nand (n1537,n1538,n1539);
or (n1538,n199,n1105);
or (n1539,n958,n471);
and (n1540,n1118,n1110);
or (n1541,n1542,n1543);
and (n1542,n1178,n1185);
and (n1543,n1179,n1182);
and (n1544,n1537,n1540);
and (n1545,n1532,n1533);
and (n1546,n1527,n1528);
nand (n1547,n1548,n1577);
nor (n1548,n1549,n1572);
nor (n1549,n1550,n1563);
xor (n1550,n1551,n1562);
xor (n1551,n1552,n1553);
xor (n1552,n993,n1013);
or (n1553,n1554,n1561);
and (n1554,n1555,n1558);
xor (n1555,n1556,n1557);
xor (n1556,n1015,n1028);
xor (n1557,n997,n1006);
or (n1558,n1559,n1560);
and (n1559,n1092,n1108);
and (n1560,n1093,n1099);
and (n1561,n1556,n1557);
xor (n1562,n1531,n1534);
or (n1563,n1564,n1571);
and (n1564,n1565,n1570);
xor (n1565,n1566,n1567);
xor (n1566,n1536,n1541);
or (n1567,n1568,n1569);
and (n1568,n1127,n1177);
and (n1569,n1128,n1149);
xor (n1570,n1555,n1558);
and (n1571,n1566,n1567);
nor (n1572,n1573,n1576);
or (n1573,n1574,n1575);
and (n1574,n1090,n1188);
and (n1575,n1091,n1126);
xor (n1576,n1565,n1570);
nand (n1577,n1578,n1580);
not (n1578,n1579);
xor (n1579,n1526,n1529);
not (n1580,n1581);
or (n1581,n1582,n1583);
and (n1582,n1551,n1562);
and (n1583,n1552,n1553);
nor (n1584,n1585,n1596);
and (n1585,n1586,n1587);
not (n1586,n1522);
nand (n1587,n1588,n1595);
or (n1588,n1589,n1590);
not (n1589,n1577);
not (n1590,n1591);
nand (n1591,n1592,n1594);
or (n1592,n1549,n1593);
nand (n1593,n1573,n1576);
nand (n1594,n1550,n1563);
nand (n1595,n1579,n1581);
and (n1596,n1523,n1524);
not (n1597,n1598);
nand (n1598,n1599,n1656);
not (n1599,n1600);
nor (n1600,n1601,n1604);
or (n1601,n1602,n1603);
and (n1602,n679,n733);
and (n1603,n680,n707);
xor (n1604,n1605,n1653);
xor (n1605,n1606,n1609);
or (n1606,n1607,n1608);
and (n1607,n681,n688);
and (n1608,n682,n685);
xor (n1609,n1610,n1631);
xor (n1610,n1611,n1628);
xor (n1611,n1612,n1622);
xor (n1612,n1613,n1615);
nand (n1613,n1614,n67);
or (n1614,n174,n70);
nand (n1615,n1616,n1617);
or (n1616,n724,n230);
nand (n1617,n1618,n237);
not (n1618,n1619);
nor (n1619,n1620,n1621);
and (n1620,n229,n156);
and (n1621,n49,n155);
nand (n1622,n1623,n1624);
or (n1623,n693,n99);
or (n1624,n100,n1625);
nor (n1625,n1626,n1627);
and (n1626,n98,n184);
and (n1627,n94,n183);
or (n1628,n1629,n1630);
and (n1629,n710,n720);
and (n1630,n711,n714);
xor (n1631,n1632,n1636);
xor (n1632,n721,n1633);
or (n1633,n1634,n1635);
and (n1634,n689,n704);
and (n1635,n690,n696);
xor (n1636,n1637,n1650);
xor (n1637,n1638,n1644);
nand (n1638,n1639,n1640);
or (n1639,n698,n122);
nand (n1640,n124,n1641);
nor (n1641,n1642,n1643);
and (n1642,n57,n28);
and (n1643,n58,n29);
nand (n1644,n1645,n1646);
or (n1645,n717,n43);
or (n1646,n44,n1647);
nor (n1647,n1648,n1649);
and (n1648,n87,n41);
and (n1649,n85,n40);
nand (n1650,n1651,n1652);
or (n1651,n95,n22);
or (n1652,n661,n112);
or (n1653,n1654,n1655);
and (n1654,n708,n730);
and (n1655,n709,n727);
nand (n1656,n1601,n1604);
and (n1657,n1658,n1598);
not (n1658,n5);
nand (n1659,n1660,n1662);
not (n1660,n1661);
nand (n1663,n1664,n1665);
nor (n1664,n1662,n1661);
wire s0n1666,s1n1666,notn1666;
or (n1666,s0n1666,s1n1666);
not(notn1666,n1661);
and (s0n1666,notn1666,n1667);
and (s1n1666,n1661,1'b0);
wire s0n1667,s1n1667,notn1667;
or (n1667,s0n1667,s1n1667);
not(notn1667,n1662);
and (s0n1667,notn1667,n1665);
and (s1n1667,n1662,n1668);
xor (n1668,n1669,n2912);
xor (n1669,n1670,n2911);
xor (n1670,n1671,n2864);
xor (n1671,n1672,n701);
xor (n1672,n1673,n2807);
xor (n1673,n1674,n2806);
xor (n1674,n1675,n2743);
xor (n1675,n1676,n2742);
xor (n1676,n1677,n2673);
xor (n1677,n1678,n2672);
xor (n1678,n1679,n2600);
xor (n1679,n1680,n2599);
xor (n1680,n1681,n2519);
xor (n1681,n1682,n2518);
xor (n1682,n1683,n2436);
xor (n1683,n1684,n2435);
xor (n1684,n1685,n2343);
xor (n1685,n1686,n2342);
or (n1686,n1687,n2255);
and (n1687,n1688,n2254);
or (n1688,n1689,n2160);
and (n1689,n1690,n2159);
or (n1690,n1691,n2066);
and (n1691,n1692,n197);
or (n1692,n1693,n1972);
and (n1693,n1694,n1971);
or (n1694,n1695,n1881);
and (n1695,n1696,n158);
or (n1696,n1697,n1787);
and (n1697,n1698,n1786);
and (n1698,n508,n1699);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
and (n1701,n156,n503);
and (n1702,n220,n147);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
or (n1705,n1706,n1709);
and (n1706,n1707,n1708);
and (n1707,n220,n503);
and (n1708,n85,n147);
and (n1709,n1710,n1711);
xor (n1710,n1707,n1708);
or (n1711,n1712,n1714);
and (n1712,n1713,n782);
and (n1713,n85,n503);
and (n1714,n1715,n1716);
xor (n1715,n1713,n782);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
and (n1718,n79,n503);
and (n1719,n184,n147);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
and (n1724,n184,n503);
and (n1725,n178,n147);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
or (n1728,n1729,n1732);
and (n1729,n1730,n1731);
and (n1730,n178,n503);
and (n1731,n58,n147);
and (n1732,n1733,n1734);
xor (n1733,n1730,n1731);
or (n1734,n1735,n1738);
and (n1735,n1736,n1737);
and (n1736,n58,n503);
and (n1737,n39,n147);
and (n1738,n1739,n1740);
xor (n1739,n1736,n1737);
or (n1740,n1741,n1744);
and (n1741,n1742,n1743);
and (n1742,n39,n503);
and (n1743,n110,n147);
and (n1744,n1745,n1746);
xor (n1745,n1742,n1743);
or (n1746,n1747,n1750);
and (n1747,n1748,n1749);
and (n1748,n110,n503);
and (n1749,n96,n147);
and (n1750,n1751,n1752);
xor (n1751,n1748,n1749);
or (n1752,n1753,n1755);
and (n1753,n1754,n1300);
and (n1754,n96,n503);
and (n1755,n1756,n1757);
xor (n1756,n1754,n1300);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
and (n1759,n135,n503);
and (n1760,n120,n147);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1766);
and (n1764,n1765,n1387);
and (n1765,n120,n503);
and (n1766,n1767,n1768);
xor (n1767,n1765,n1387);
or (n1768,n1769,n1771);
and (n1769,n1770,n1444);
and (n1770,n32,n503);
and (n1771,n1772,n1773);
xor (n1772,n1770,n1444);
or (n1773,n1774,n1776);
and (n1774,n1775,n1457);
and (n1775,n21,n503);
and (n1776,n1777,n1778);
xor (n1777,n1775,n1457);
or (n1778,n1779,n1781);
and (n1779,n1780,n1487);
and (n1780,n285,n503);
and (n1781,n1782,n1783);
xor (n1782,n1780,n1487);
and (n1783,n1784,n1785);
and (n1784,n363,n503);
and (n1785,n424,n147);
and (n1786,n156,n146);
and (n1787,n1788,n1789);
xor (n1788,n1698,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n508,n1699);
and (n1792,n220,n146);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1704,n1705);
and (n1798,n85,n146);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1710,n1711);
and (n1804,n79,n146);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1715,n1716);
and (n1810,n184,n146);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1721,n1722);
and (n1816,n178,n146);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1727,n1728);
and (n1822,n58,n146);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
xor (n1827,n1733,n1734);
and (n1828,n39,n146);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
or (n1831,n1832,n1835);
and (n1832,n1833,n1834);
xor (n1833,n1739,n1740);
and (n1834,n110,n146);
and (n1835,n1836,n1837);
xor (n1836,n1833,n1834);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
xor (n1839,n1745,n1746);
and (n1840,n96,n146);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
or (n1843,n1844,n1847);
and (n1844,n1845,n1846);
xor (n1845,n1751,n1752);
and (n1846,n135,n146);
and (n1847,n1848,n1849);
xor (n1848,n1845,n1846);
or (n1849,n1850,n1853);
and (n1850,n1851,n1852);
xor (n1851,n1756,n1757);
and (n1852,n120,n146);
and (n1853,n1854,n1855);
xor (n1854,n1851,n1852);
or (n1855,n1856,n1859);
and (n1856,n1857,n1858);
xor (n1857,n1762,n1763);
and (n1858,n32,n146);
and (n1859,n1860,n1861);
xor (n1860,n1857,n1858);
or (n1861,n1862,n1865);
and (n1862,n1863,n1864);
xor (n1863,n1767,n1768);
and (n1864,n21,n146);
and (n1865,n1866,n1867);
xor (n1866,n1863,n1864);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
xor (n1869,n1772,n1773);
and (n1870,n285,n146);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
or (n1873,n1874,n1877);
and (n1874,n1875,n1876);
xor (n1875,n1777,n1778);
and (n1876,n363,n146);
and (n1877,n1878,n1879);
xor (n1878,n1875,n1876);
and (n1879,n1880,n1463);
xor (n1880,n1782,n1783);
and (n1881,n1882,n1883);
xor (n1882,n1696,n158);
or (n1883,n1884,n1887);
and (n1884,n1885,n1886);
xor (n1885,n1788,n1789);
and (n1886,n220,n151);
and (n1887,n1888,n1889);
xor (n1888,n1885,n1886);
or (n1889,n1890,n1892);
and (n1890,n1891,n455);
xor (n1891,n1794,n1795);
and (n1892,n1893,n1894);
xor (n1893,n1891,n455);
or (n1894,n1895,n1897);
and (n1895,n1896,n542);
xor (n1896,n1800,n1801);
and (n1897,n1898,n1899);
xor (n1898,n1896,n542);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1806,n1807);
and (n1902,n184,n151);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1812,n1813);
and (n1908,n178,n151);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
or (n1911,n1912,n1914);
and (n1912,n1913,n936);
xor (n1913,n1818,n1819);
and (n1914,n1915,n1916);
xor (n1915,n1913,n936);
or (n1916,n1917,n1920);
and (n1917,n1918,n1919);
xor (n1918,n1824,n1825);
and (n1919,n39,n151);
and (n1920,n1921,n1922);
xor (n1921,n1918,n1919);
or (n1922,n1923,n1926);
and (n1923,n1924,n1925);
xor (n1924,n1830,n1831);
and (n1925,n110,n151);
and (n1926,n1927,n1928);
xor (n1927,n1924,n1925);
or (n1928,n1929,n1932);
and (n1929,n1930,n1931);
xor (n1930,n1836,n1837);
and (n1931,n96,n151);
and (n1932,n1933,n1934);
xor (n1933,n1930,n1931);
or (n1934,n1935,n1938);
and (n1935,n1936,n1937);
xor (n1936,n1842,n1843);
and (n1937,n135,n151);
and (n1938,n1939,n1940);
xor (n1939,n1936,n1937);
or (n1940,n1941,n1944);
and (n1941,n1942,n1943);
xor (n1942,n1848,n1849);
and (n1943,n120,n151);
and (n1944,n1945,n1946);
xor (n1945,n1942,n1943);
or (n1946,n1947,n1950);
and (n1947,n1948,n1949);
xor (n1948,n1854,n1855);
and (n1949,n32,n151);
and (n1950,n1951,n1952);
xor (n1951,n1948,n1949);
or (n1952,n1953,n1956);
and (n1953,n1954,n1955);
xor (n1954,n1860,n1861);
and (n1955,n21,n151);
and (n1956,n1957,n1958);
xor (n1957,n1954,n1955);
or (n1958,n1959,n1961);
and (n1959,n1960,n1409);
xor (n1960,n1866,n1867);
and (n1961,n1962,n1963);
xor (n1962,n1960,n1409);
or (n1963,n1964,n1966);
and (n1964,n1965,n1436);
xor (n1965,n1872,n1873);
and (n1966,n1967,n1968);
xor (n1967,n1965,n1436);
and (n1968,n1969,n1970);
xor (n1969,n1878,n1879);
and (n1970,n424,n151);
and (n1971,n156,n203);
and (n1972,n1973,n1974);
xor (n1973,n1694,n1971);
or (n1974,n1975,n1978);
and (n1975,n1976,n1977);
xor (n1976,n1882,n1883);
and (n1977,n220,n203);
and (n1978,n1979,n1980);
xor (n1979,n1976,n1977);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
xor (n1982,n1888,n1889);
and (n1983,n85,n203);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1893,n1894);
and (n1989,n79,n203);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1996);
and (n1993,n1994,n1995);
xor (n1994,n1898,n1899);
and (n1995,n184,n203);
and (n1996,n1997,n1998);
xor (n1997,n1994,n1995);
or (n1998,n1999,n2002);
and (n1999,n2000,n2001);
xor (n2000,n1904,n1905);
and (n2001,n178,n203);
and (n2002,n2003,n2004);
xor (n2003,n2000,n2001);
or (n2004,n2005,n2008);
and (n2005,n2006,n2007);
xor (n2006,n1910,n1911);
and (n2007,n58,n203);
and (n2008,n2009,n2010);
xor (n2009,n2006,n2007);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1915,n1916);
and (n2013,n39,n203);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
or (n2016,n2017,n2020);
and (n2017,n2018,n2019);
xor (n2018,n1921,n1922);
and (n2019,n110,n203);
and (n2020,n2021,n2022);
xor (n2021,n2018,n2019);
or (n2022,n2023,n2026);
and (n2023,n2024,n2025);
xor (n2024,n1927,n1928);
and (n2025,n96,n203);
and (n2026,n2027,n2028);
xor (n2027,n2024,n2025);
or (n2028,n2029,n2032);
and (n2029,n2030,n2031);
xor (n2030,n1933,n1934);
and (n2031,n135,n203);
and (n2032,n2033,n2034);
xor (n2033,n2030,n2031);
or (n2034,n2035,n2038);
and (n2035,n2036,n2037);
xor (n2036,n1939,n1940);
and (n2037,n120,n203);
and (n2038,n2039,n2040);
xor (n2039,n2036,n2037);
or (n2040,n2041,n2044);
and (n2041,n2042,n2043);
xor (n2042,n1945,n1946);
and (n2043,n32,n203);
and (n2044,n2045,n2046);
xor (n2045,n2042,n2043);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1951,n1952);
and (n2049,n21,n203);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
or (n2052,n2053,n2056);
and (n2053,n2054,n2055);
xor (n2054,n1957,n1958);
and (n2055,n285,n203);
and (n2056,n2057,n2058);
xor (n2057,n2054,n2055);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n1962,n1963);
and (n2061,n363,n203);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
and (n2064,n2065,n1393);
xor (n2065,n1967,n1968);
and (n2066,n2067,n2068);
xor (n2067,n1692,n197);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n1973,n1974);
and (n2071,n220,n73);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2077);
and (n2075,n2076,n280);
xor (n2076,n1979,n1980);
and (n2077,n2078,n2079);
xor (n2078,n2076,n280);
or (n2079,n2080,n2083);
and (n2080,n2081,n2082);
xor (n2081,n1985,n1986);
and (n2082,n79,n73);
and (n2083,n2084,n2085);
xor (n2084,n2081,n2082);
or (n2085,n2086,n2088);
and (n2086,n2087,n469);
xor (n2087,n1991,n1992);
and (n2088,n2089,n2090);
xor (n2089,n2087,n469);
or (n2090,n2091,n2094);
and (n2091,n2092,n2093);
xor (n2092,n1997,n1998);
and (n2093,n178,n73);
and (n2094,n2095,n2096);
xor (n2095,n2092,n2093);
or (n2096,n2097,n2100);
and (n2097,n2098,n2099);
xor (n2098,n2003,n2004);
and (n2099,n58,n73);
and (n2100,n2101,n2102);
xor (n2101,n2098,n2099);
or (n2102,n2103,n2106);
and (n2103,n2104,n2105);
xor (n2104,n2009,n2010);
and (n2105,n39,n73);
and (n2106,n2107,n2108);
xor (n2107,n2104,n2105);
or (n2108,n2109,n2112);
and (n2109,n2110,n2111);
xor (n2110,n2015,n2016);
and (n2111,n110,n73);
and (n2112,n2113,n2114);
xor (n2113,n2110,n2111);
or (n2114,n2115,n2118);
and (n2115,n2116,n2117);
xor (n2116,n2021,n2022);
and (n2117,n96,n73);
and (n2118,n2119,n2120);
xor (n2119,n2116,n2117);
or (n2120,n2121,n2124);
and (n2121,n2122,n2123);
xor (n2122,n2027,n2028);
and (n2123,n135,n73);
and (n2124,n2125,n2126);
xor (n2125,n2122,n2123);
or (n2126,n2127,n2130);
and (n2127,n2128,n2129);
xor (n2128,n2033,n2034);
and (n2129,n120,n73);
and (n2130,n2131,n2132);
xor (n2131,n2128,n2129);
or (n2132,n2133,n2136);
and (n2133,n2134,n2135);
xor (n2134,n2039,n2040);
and (n2135,n32,n73);
and (n2136,n2137,n2138);
xor (n2137,n2134,n2135);
or (n2138,n2139,n2142);
and (n2139,n2140,n2141);
xor (n2140,n2045,n2046);
and (n2141,n21,n73);
and (n2142,n2143,n2144);
xor (n2143,n2140,n2141);
or (n2144,n2145,n2148);
and (n2145,n2146,n2147);
xor (n2146,n2051,n2052);
and (n2147,n285,n73);
and (n2148,n2149,n2150);
xor (n2149,n2146,n2147);
or (n2150,n2151,n2154);
and (n2151,n2152,n2153);
xor (n2152,n2057,n2058);
and (n2153,n363,n73);
and (n2154,n2155,n2156);
xor (n2155,n2152,n2153);
and (n2156,n2157,n2158);
xor (n2157,n2063,n2064);
and (n2158,n424,n73);
and (n2159,n156,n65);
and (n2160,n2161,n2162);
xor (n2161,n1690,n2159);
or (n2162,n2163,n2166);
and (n2163,n2164,n2165);
xor (n2164,n2067,n2068);
and (n2165,n220,n65);
and (n2166,n2167,n2168);
xor (n2167,n2164,n2165);
or (n2168,n2169,n2172);
and (n2169,n2170,n2171);
xor (n2170,n2073,n2074);
and (n2171,n85,n65);
and (n2172,n2173,n2174);
xor (n2173,n2170,n2171);
or (n2174,n2175,n2178);
and (n2175,n2176,n2177);
xor (n2176,n2078,n2079);
and (n2177,n79,n65);
and (n2178,n2179,n2180);
xor (n2179,n2176,n2177);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2084,n2085);
and (n2183,n184,n65);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2089,n2090);
and (n2189,n178,n65);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2095,n2096);
and (n2195,n58,n65);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2101,n2102);
and (n2201,n39,n65);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2107,n2108);
and (n2207,n110,n65);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2113,n2114);
and (n2213,n96,n65);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2119,n2120);
and (n2219,n135,n65);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2125,n2126);
and (n2225,n120,n65);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2131,n2132);
and (n2231,n32,n65);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2137,n2138);
and (n2237,n21,n65);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
or (n2240,n2241,n2244);
and (n2241,n2242,n2243);
xor (n2242,n2143,n2144);
and (n2243,n285,n65);
and (n2244,n2245,n2246);
xor (n2245,n2242,n2243);
or (n2246,n2247,n2250);
and (n2247,n2248,n2249);
xor (n2248,n2149,n2150);
and (n2249,n363,n65);
and (n2250,n2251,n2252);
xor (n2251,n2248,n2249);
and (n2252,n2253,n1293);
xor (n2253,n2155,n2156);
and (n2254,n156,n67);
and (n2255,n2256,n2257);
xor (n2256,n1688,n2254);
or (n2257,n2258,n2260);
and (n2258,n2259,n324);
xor (n2259,n2161,n2162);
and (n2260,n2261,n2262);
xor (n2261,n2259,n324);
or (n2262,n2263,n2265);
and (n2263,n2264,n84);
xor (n2264,n2167,n2168);
and (n2265,n2266,n2267);
xor (n2266,n2264,n84);
or (n2267,n2268,n2270);
and (n2268,n2269,n80);
xor (n2269,n2173,n2174);
and (n2270,n2271,n2272);
xor (n2271,n2269,n80);
or (n2272,n2273,n2275);
and (n2273,n2274,n185);
xor (n2274,n2179,n2180);
and (n2275,n2276,n2277);
xor (n2276,n2274,n185);
or (n2277,n2278,n2280);
and (n2278,n2279,n179);
xor (n2279,n2185,n2186);
and (n2280,n2281,n2282);
xor (n2281,n2279,n179);
or (n2282,n2283,n2286);
and (n2283,n2284,n2285);
xor (n2284,n2191,n2192);
and (n2285,n58,n67);
and (n2286,n2287,n2288);
xor (n2287,n2284,n2285);
or (n2288,n2289,n2292);
and (n2289,n2290,n2291);
xor (n2290,n2197,n2198);
and (n2291,n39,n67);
and (n2292,n2293,n2294);
xor (n2293,n2290,n2291);
or (n2294,n2295,n2297);
and (n2295,n2296,n819);
xor (n2296,n2203,n2204);
and (n2297,n2298,n2299);
xor (n2298,n2296,n819);
or (n2299,n2300,n2303);
and (n2300,n2301,n2302);
xor (n2301,n2209,n2210);
and (n2302,n96,n67);
and (n2303,n2304,n2305);
xor (n2304,n2301,n2302);
or (n2305,n2306,n2309);
and (n2306,n2307,n2308);
xor (n2307,n2215,n2216);
and (n2308,n135,n67);
and (n2309,n2310,n2311);
xor (n2310,n2307,n2308);
or (n2311,n2312,n2315);
and (n2312,n2313,n2314);
xor (n2313,n2221,n2222);
and (n2314,n120,n67);
and (n2315,n2316,n2317);
xor (n2316,n2313,n2314);
or (n2317,n2318,n2321);
and (n2318,n2319,n2320);
xor (n2319,n2227,n2228);
and (n2320,n32,n67);
and (n2321,n2322,n2323);
xor (n2322,n2319,n2320);
or (n2323,n2324,n2326);
and (n2324,n2325,n1143);
xor (n2325,n2233,n2234);
and (n2326,n2327,n2328);
xor (n2327,n2325,n1143);
or (n2328,n2329,n2331);
and (n2329,n2330,n1211);
xor (n2330,n2239,n2240);
and (n2331,n2332,n2333);
xor (n2332,n2330,n1211);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2245,n2246);
and (n2336,n363,n67);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
and (n2339,n2340,n2341);
xor (n2340,n2251,n2252);
and (n2341,n424,n67);
and (n2342,n156,n234);
or (n2343,n2344,n2347);
and (n2344,n2345,n2346);
xor (n2345,n2256,n2257);
and (n2346,n220,n234);
and (n2347,n2348,n2349);
xor (n2348,n2345,n2346);
or (n2349,n2350,n2353);
and (n2350,n2351,n2352);
xor (n2351,n2261,n2262);
and (n2352,n85,n234);
and (n2353,n2354,n2355);
xor (n2354,n2351,n2352);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2266,n2267);
and (n2358,n79,n234);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2271,n2272);
and (n2364,n184,n234);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2276,n2277);
and (n2370,n178,n234);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2281,n2282);
and (n2376,n58,n234);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2287,n2288);
and (n2382,n39,n234);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2293,n2294);
and (n2388,n110,n234);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2298,n2299);
and (n2394,n96,n234);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2304,n2305);
and (n2400,n135,n234);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
or (n2403,n2404,n2407);
and (n2404,n2405,n2406);
xor (n2405,n2310,n2311);
and (n2406,n120,n234);
and (n2407,n2408,n2409);
xor (n2408,n2405,n2406);
or (n2409,n2410,n2413);
and (n2410,n2411,n2412);
xor (n2411,n2316,n2317);
and (n2412,n32,n234);
and (n2413,n2414,n2415);
xor (n2414,n2411,n2412);
or (n2415,n2416,n2419);
and (n2416,n2417,n2418);
xor (n2417,n2322,n2323);
and (n2418,n21,n234);
and (n2419,n2420,n2421);
xor (n2420,n2417,n2418);
or (n2421,n2422,n2425);
and (n2422,n2423,n2424);
xor (n2423,n2327,n2328);
and (n2424,n285,n234);
and (n2425,n2426,n2427);
xor (n2426,n2423,n2424);
or (n2427,n2428,n2431);
and (n2428,n2429,n2430);
xor (n2429,n2332,n2333);
and (n2430,n363,n234);
and (n2431,n2432,n2433);
xor (n2432,n2429,n2430);
and (n2433,n2434,n1197);
xor (n2434,n2338,n2339);
and (n2435,n220,n49);
or (n2436,n2437,n2440);
and (n2437,n2438,n2439);
xor (n2438,n2348,n2349);
and (n2439,n85,n49);
and (n2440,n2441,n2442);
xor (n2441,n2438,n2439);
or (n2442,n2443,n2445);
and (n2443,n2444,n307);
xor (n2444,n2354,n2355);
and (n2445,n2446,n2447);
xor (n2446,n2444,n307);
or (n2447,n2448,n2450);
and (n2448,n2449,n243);
xor (n2449,n2360,n2361);
and (n2450,n2451,n2452);
xor (n2451,n2449,n243);
or (n2452,n2453,n2456);
and (n2453,n2454,n2455);
xor (n2454,n2366,n2367);
and (n2455,n178,n49);
and (n2456,n2457,n2458);
xor (n2457,n2454,n2455);
or (n2458,n2459,n2461);
and (n2459,n2460,n292);
xor (n2460,n2372,n2373);
and (n2461,n2462,n2463);
xor (n2462,n2460,n292);
or (n2463,n2464,n2466);
and (n2464,n2465,n382);
xor (n2465,n2378,n2379);
and (n2466,n2467,n2468);
xor (n2467,n2465,n382);
or (n2468,n2469,n2472);
and (n2469,n2470,n2471);
xor (n2470,n2384,n2385);
and (n2471,n110,n49);
and (n2472,n2473,n2474);
xor (n2473,n2470,n2471);
or (n2474,n2475,n2478);
and (n2475,n2476,n2477);
xor (n2476,n2390,n2391);
and (n2477,n96,n49);
and (n2478,n2479,n2480);
xor (n2479,n2476,n2477);
or (n2480,n2481,n2483);
and (n2481,n2482,n830);
xor (n2482,n2396,n2397);
and (n2483,n2484,n2485);
xor (n2484,n2482,n830);
or (n2485,n2486,n2489);
and (n2486,n2487,n2488);
xor (n2487,n2402,n2403);
and (n2488,n120,n49);
and (n2489,n2490,n2491);
xor (n2490,n2487,n2488);
or (n2491,n2492,n2495);
and (n2492,n2493,n2494);
xor (n2493,n2408,n2409);
and (n2494,n32,n49);
and (n2495,n2496,n2497);
xor (n2496,n2493,n2494);
or (n2497,n2498,n2501);
and (n2498,n2499,n2500);
xor (n2499,n2414,n2415);
and (n2500,n21,n49);
and (n2501,n2502,n2503);
xor (n2502,n2499,n2500);
or (n2503,n2504,n2507);
and (n2504,n2505,n2506);
xor (n2505,n2420,n2421);
and (n2506,n285,n49);
and (n2507,n2508,n2509);
xor (n2508,n2505,n2506);
or (n2509,n2510,n2513);
and (n2510,n2511,n2512);
xor (n2511,n2426,n2427);
and (n2512,n363,n49);
and (n2513,n2514,n2515);
xor (n2514,n2511,n2512);
and (n2515,n2516,n2517);
xor (n2516,n2432,n2433);
and (n2517,n424,n49);
and (n2518,n85,n48);
or (n2519,n2520,n2523);
and (n2520,n2521,n2522);
xor (n2521,n2441,n2442);
and (n2522,n79,n48);
and (n2523,n2524,n2525);
xor (n2524,n2521,n2522);
or (n2525,n2526,n2529);
and (n2526,n2527,n2528);
xor (n2527,n2446,n2447);
and (n2528,n184,n48);
and (n2529,n2530,n2531);
xor (n2530,n2527,n2528);
or (n2531,n2532,n2535);
and (n2532,n2533,n2534);
xor (n2533,n2451,n2452);
and (n2534,n178,n48);
and (n2535,n2536,n2537);
xor (n2536,n2533,n2534);
or (n2537,n2538,n2541);
and (n2538,n2539,n2540);
xor (n2539,n2457,n2458);
and (n2540,n58,n48);
and (n2541,n2542,n2543);
xor (n2542,n2539,n2540);
or (n2543,n2544,n2547);
and (n2544,n2545,n2546);
xor (n2545,n2462,n2463);
and (n2546,n39,n48);
and (n2547,n2548,n2549);
xor (n2548,n2545,n2546);
or (n2549,n2550,n2553);
and (n2550,n2551,n2552);
xor (n2551,n2467,n2468);
and (n2552,n110,n48);
and (n2553,n2554,n2555);
xor (n2554,n2551,n2552);
or (n2555,n2556,n2559);
and (n2556,n2557,n2558);
xor (n2557,n2473,n2474);
and (n2558,n96,n48);
and (n2559,n2560,n2561);
xor (n2560,n2557,n2558);
or (n2561,n2562,n2565);
and (n2562,n2563,n2564);
xor (n2563,n2479,n2480);
and (n2564,n135,n48);
and (n2565,n2566,n2567);
xor (n2566,n2563,n2564);
or (n2567,n2568,n2571);
and (n2568,n2569,n2570);
xor (n2569,n2484,n2485);
and (n2570,n120,n48);
and (n2571,n2572,n2573);
xor (n2572,n2569,n2570);
or (n2573,n2574,n2577);
and (n2574,n2575,n2576);
xor (n2575,n2490,n2491);
and (n2576,n32,n48);
and (n2577,n2578,n2579);
xor (n2578,n2575,n2576);
or (n2579,n2580,n2583);
and (n2580,n2581,n2582);
xor (n2581,n2496,n2497);
and (n2582,n21,n48);
and (n2583,n2584,n2585);
xor (n2584,n2581,n2582);
or (n2585,n2586,n2589);
and (n2586,n2587,n2588);
xor (n2587,n2502,n2503);
and (n2588,n285,n48);
and (n2589,n2590,n2591);
xor (n2590,n2587,n2588);
or (n2591,n2592,n2595);
and (n2592,n2593,n2594);
xor (n2593,n2508,n2509);
and (n2594,n363,n48);
and (n2595,n2596,n2597);
xor (n2596,n2593,n2594);
and (n2597,n2598,n1116);
xor (n2598,n2514,n2515);
and (n2599,n79,n41);
or (n2600,n2601,n2604);
and (n2601,n2602,n2603);
xor (n2602,n2524,n2525);
and (n2603,n184,n41);
and (n2604,n2605,n2606);
xor (n2605,n2602,n2603);
or (n2606,n2607,n2610);
and (n2607,n2608,n2609);
xor (n2608,n2530,n2531);
and (n2609,n178,n41);
and (n2610,n2611,n2612);
xor (n2611,n2608,n2609);
or (n2612,n2613,n2615);
and (n2613,n2614,n59);
xor (n2614,n2536,n2537);
and (n2615,n2616,n2617);
xor (n2616,n2614,n59);
or (n2617,n2618,n2620);
and (n2618,n2619,n42);
xor (n2619,n2542,n2543);
and (n2620,n2621,n2622);
xor (n2621,n2619,n42);
or (n2622,n2623,n2626);
and (n2623,n2624,n2625);
xor (n2624,n2548,n2549);
and (n2625,n110,n41);
and (n2626,n2627,n2628);
xor (n2627,n2624,n2625);
or (n2628,n2629,n2632);
and (n2629,n2630,n2631);
xor (n2630,n2554,n2555);
and (n2631,n96,n41);
and (n2632,n2633,n2634);
xor (n2633,n2630,n2631);
or (n2634,n2635,n2637);
and (n2635,n2636,n489);
xor (n2636,n2560,n2561);
and (n2637,n2638,n2639);
xor (n2638,n2636,n489);
or (n2639,n2640,n2643);
and (n2640,n2641,n2642);
xor (n2641,n2566,n2567);
and (n2642,n120,n41);
and (n2643,n2644,n2645);
xor (n2644,n2641,n2642);
or (n2645,n2646,n2649);
and (n2646,n2647,n2648);
xor (n2647,n2572,n2573);
and (n2648,n32,n41);
and (n2649,n2650,n2651);
xor (n2650,n2647,n2648);
or (n2651,n2652,n2655);
and (n2652,n2653,n2654);
xor (n2653,n2578,n2579);
and (n2654,n21,n41);
and (n2655,n2656,n2657);
xor (n2656,n2653,n2654);
or (n2657,n2658,n2661);
and (n2658,n2659,n2660);
xor (n2659,n2584,n2585);
and (n2660,n285,n41);
and (n2661,n2662,n2663);
xor (n2662,n2659,n2660);
or (n2663,n2664,n2667);
and (n2664,n2665,n2666);
xor (n2665,n2590,n2591);
and (n2666,n363,n41);
and (n2667,n2668,n2669);
xor (n2668,n2665,n2666);
and (n2669,n2670,n2671);
xor (n2670,n2596,n2597);
and (n2671,n424,n41);
and (n2672,n184,n103);
or (n2673,n2674,n2677);
and (n2674,n2675,n2676);
xor (n2675,n2605,n2606);
and (n2676,n178,n103);
and (n2677,n2678,n2679);
xor (n2678,n2675,n2676);
or (n2679,n2680,n2683);
and (n2680,n2681,n2682);
xor (n2681,n2611,n2612);
and (n2682,n58,n103);
and (n2683,n2684,n2685);
xor (n2684,n2681,n2682);
or (n2685,n2686,n2689);
and (n2686,n2687,n2688);
xor (n2687,n2616,n2617);
and (n2688,n39,n103);
and (n2689,n2690,n2691);
xor (n2690,n2687,n2688);
or (n2691,n2692,n2695);
and (n2692,n2693,n2694);
xor (n2693,n2621,n2622);
and (n2694,n110,n103);
and (n2695,n2696,n2697);
xor (n2696,n2693,n2694);
or (n2697,n2698,n2701);
and (n2698,n2699,n2700);
xor (n2699,n2627,n2628);
and (n2700,n96,n103);
and (n2701,n2702,n2703);
xor (n2702,n2699,n2700);
or (n2703,n2704,n2707);
and (n2704,n2705,n2706);
xor (n2705,n2633,n2634);
and (n2706,n135,n103);
and (n2707,n2708,n2709);
xor (n2708,n2705,n2706);
or (n2709,n2710,n2713);
and (n2710,n2711,n2712);
xor (n2711,n2638,n2639);
and (n2712,n120,n103);
and (n2713,n2714,n2715);
xor (n2714,n2711,n2712);
or (n2715,n2716,n2719);
and (n2716,n2717,n2718);
xor (n2717,n2644,n2645);
and (n2718,n32,n103);
and (n2719,n2720,n2721);
xor (n2720,n2717,n2718);
or (n2721,n2722,n2725);
and (n2722,n2723,n2724);
xor (n2723,n2650,n2651);
and (n2724,n21,n103);
and (n2725,n2726,n2727);
xor (n2726,n2723,n2724);
or (n2727,n2728,n2731);
and (n2728,n2729,n2730);
xor (n2729,n2656,n2657);
and (n2730,n285,n103);
and (n2731,n2732,n2733);
xor (n2732,n2729,n2730);
or (n2733,n2734,n2737);
and (n2734,n2735,n2736);
xor (n2735,n2662,n2663);
and (n2736,n363,n103);
and (n2737,n2738,n2739);
xor (n2738,n2735,n2736);
and (n2739,n2740,n2741);
xor (n2740,n2668,n2669);
not (n2741,n915);
and (n2742,n178,n94);
or (n2743,n2744,n2747);
and (n2744,n2745,n2746);
xor (n2745,n2678,n2679);
and (n2746,n58,n94);
and (n2747,n2748,n2749);
xor (n2748,n2745,n2746);
or (n2749,n2750,n2753);
and (n2750,n2751,n2752);
xor (n2751,n2684,n2685);
and (n2752,n39,n94);
and (n2753,n2754,n2755);
xor (n2754,n2751,n2752);
or (n2755,n2756,n2759);
and (n2756,n2757,n2758);
xor (n2757,n2690,n2691);
and (n2758,n110,n94);
and (n2759,n2760,n2761);
xor (n2760,n2757,n2758);
or (n2761,n2762,n2765);
and (n2762,n2763,n2764);
xor (n2763,n2696,n2697);
and (n2764,n96,n94);
and (n2765,n2766,n2767);
xor (n2766,n2763,n2764);
or (n2767,n2768,n2771);
and (n2768,n2769,n2770);
xor (n2769,n2702,n2703);
and (n2770,n135,n94);
and (n2771,n2772,n2773);
xor (n2772,n2769,n2770);
or (n2773,n2774,n2777);
and (n2774,n2775,n2776);
xor (n2775,n2708,n2709);
and (n2776,n120,n94);
and (n2777,n2778,n2779);
xor (n2778,n2775,n2776);
or (n2779,n2780,n2783);
and (n2780,n2781,n2782);
xor (n2781,n2714,n2715);
and (n2782,n32,n94);
and (n2783,n2784,n2785);
xor (n2784,n2781,n2782);
or (n2785,n2786,n2789);
and (n2786,n2787,n2788);
xor (n2787,n2720,n2721);
and (n2788,n21,n94);
and (n2789,n2790,n2791);
xor (n2790,n2787,n2788);
or (n2791,n2792,n2795);
and (n2792,n2793,n2794);
xor (n2793,n2726,n2727);
and (n2794,n285,n94);
and (n2795,n2796,n2797);
xor (n2796,n2793,n2794);
or (n2797,n2798,n2801);
and (n2798,n2799,n2800);
xor (n2799,n2732,n2733);
and (n2800,n363,n94);
and (n2801,n2802,n2803);
xor (n2802,n2799,n2800);
and (n2803,n2804,n2805);
xor (n2804,n2738,n2739);
and (n2805,n424,n94);
and (n2806,n58,n126);
or (n2807,n2808,n2811);
and (n2808,n2809,n2810);
xor (n2809,n2748,n2749);
and (n2810,n39,n126);
and (n2811,n2812,n2813);
xor (n2812,n2809,n2810);
or (n2813,n2814,n2817);
and (n2814,n2815,n2816);
xor (n2815,n2754,n2755);
and (n2816,n110,n126);
and (n2817,n2818,n2819);
xor (n2818,n2815,n2816);
or (n2819,n2820,n2823);
and (n2820,n2821,n2822);
xor (n2821,n2760,n2761);
and (n2822,n96,n126);
and (n2823,n2824,n2825);
xor (n2824,n2821,n2822);
or (n2825,n2826,n2829);
and (n2826,n2827,n2828);
xor (n2827,n2766,n2767);
and (n2828,n135,n126);
and (n2829,n2830,n2831);
xor (n2830,n2827,n2828);
or (n2831,n2832,n2835);
and (n2832,n2833,n2834);
xor (n2833,n2772,n2773);
and (n2834,n120,n126);
and (n2835,n2836,n2837);
xor (n2836,n2833,n2834);
or (n2837,n2838,n2841);
and (n2838,n2839,n2840);
xor (n2839,n2778,n2779);
and (n2840,n32,n126);
and (n2841,n2842,n2843);
xor (n2842,n2839,n2840);
or (n2843,n2844,n2847);
and (n2844,n2845,n2846);
xor (n2845,n2784,n2785);
and (n2846,n21,n126);
and (n2847,n2848,n2849);
xor (n2848,n2845,n2846);
or (n2849,n2850,n2853);
and (n2850,n2851,n2852);
xor (n2851,n2790,n2791);
and (n2852,n285,n126);
and (n2853,n2854,n2855);
xor (n2854,n2851,n2852);
or (n2855,n2856,n2859);
and (n2856,n2857,n2858);
xor (n2857,n2796,n2797);
and (n2858,n363,n126);
and (n2859,n2860,n2861);
xor (n2860,n2857,n2858);
and (n2861,n2862,n2863);
xor (n2862,n2802,n2803);
not (n2863,n764);
or (n2864,n2865,n2867);
and (n2865,n2866,n636);
xor (n2866,n2812,n2813);
and (n2867,n2868,n2869);
xor (n2868,n2866,n636);
or (n2869,n2870,n2873);
and (n2870,n2871,n2872);
xor (n2871,n2818,n2819);
and (n2872,n96,n29);
and (n2873,n2874,n2875);
xor (n2874,n2871,n2872);
or (n2875,n2876,n2879);
and (n2876,n2877,n2878);
xor (n2877,n2824,n2825);
and (n2878,n135,n29);
and (n2879,n2880,n2881);
xor (n2880,n2877,n2878);
or (n2881,n2882,n2884);
and (n2882,n2883,n121);
xor (n2883,n2830,n2831);
and (n2884,n2885,n2886);
xor (n2885,n2883,n121);
or (n2886,n2887,n2889);
and (n2887,n2888,n169);
xor (n2888,n2836,n2837);
and (n2889,n2890,n2891);
xor (n2890,n2888,n169);
or (n2891,n2892,n2894);
and (n2892,n2893,n358);
xor (n2893,n2842,n2843);
and (n2894,n2895,n2896);
xor (n2895,n2893,n358);
or (n2896,n2897,n2900);
and (n2897,n2898,n2899);
xor (n2898,n2848,n2849);
and (n2899,n285,n29);
and (n2900,n2901,n2902);
xor (n2901,n2898,n2899);
or (n2902,n2903,n2906);
and (n2903,n2904,n2905);
xor (n2904,n2854,n2855);
and (n2905,n363,n29);
and (n2906,n2907,n2908);
xor (n2907,n2904,n2905);
and (n2908,n2909,n2910);
xor (n2909,n2860,n2861);
and (n2910,n424,n29);
and (n2911,n110,n25);
or (n2912,n2913,n2916);
and (n2913,n2914,n2915);
xor (n2914,n2868,n2869);
and (n2915,n96,n25);
and (n2916,n2917,n2918);
xor (n2917,n2914,n2915);
or (n2918,n2919,n2922);
and (n2919,n2920,n2921);
xor (n2920,n2874,n2875);
and (n2921,n135,n25);
and (n2922,n2923,n2924);
xor (n2923,n2920,n2921);
or (n2924,n2925,n2928);
and (n2925,n2926,n2927);
xor (n2926,n2880,n2881);
and (n2927,n120,n25);
and (n2928,n2929,n2930);
xor (n2929,n2926,n2927);
or (n2930,n2931,n2934);
and (n2931,n2932,n2933);
xor (n2932,n2885,n2886);
and (n2933,n32,n25);
and (n2934,n2935,n2936);
xor (n2935,n2932,n2933);
or (n2936,n2937,n2940);
and (n2937,n2938,n2939);
xor (n2938,n2890,n2891);
and (n2939,n21,n25);
and (n2940,n2941,n2942);
xor (n2941,n2938,n2939);
or (n2942,n2943,n2946);
and (n2943,n2944,n2945);
xor (n2944,n2895,n2896);
and (n2945,n285,n25);
and (n2946,n2947,n2948);
xor (n2947,n2944,n2945);
or (n2948,n2949,n2952);
and (n2949,n2950,n2951);
xor (n2950,n2901,n2902);
and (n2951,n363,n25);
and (n2952,n2953,n2954);
xor (n2953,n2950,n2951);
and (n2954,n2955,n2956);
xor (n2955,n2907,n2908);
and (n2956,n424,n25);
endmodule
