module top (out,n3,n6,n7,n27,n29,n35,n41,n47,n54
        ,n56,n64,n65,n73,n77,n81,n86,n96,n102,n103
        ,n111,n123,n133,n142,n143,n149,n157,n167,n172,n182
        ,n190,n251,n252,n281,n373,n436,n497,n584);
output out;
input n3;
input n6;
input n7;
input n27;
input n29;
input n35;
input n41;
input n47;
input n54;
input n56;
input n64;
input n65;
input n73;
input n77;
input n81;
input n86;
input n96;
input n102;
input n103;
input n111;
input n123;
input n133;
input n142;
input n143;
input n149;
input n157;
input n167;
input n172;
input n182;
input n190;
input n251;
input n252;
input n281;
input n373;
input n436;
input n497;
input n584;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
xor (out,n0,n1542);
nand (n0,n1,n8);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nor (n5,n6,n7);
nand (n8,n9,n1539);
nand (n9,n10,n1538);
or (n10,n11,n510);
nand (n11,n12,n509);
not (n12,n13);
nor (n13,n14,n387);
xor (n14,n15,n329);
xor (n15,n16,n196);
xor (n16,n17,n135);
xor (n17,n18,n88);
or (n18,n19,n87);
and (n19,n20,n74);
xor (n20,n21,n49);
nand (n21,n22,n43);
or (n22,n23,n31);
not (n23,n24);
nor (n24,n25,n30);
and (n25,n26,n28);
not (n26,n27);
not (n28,n29);
and (n30,n27,n29);
not (n31,n32);
nor (n32,n33,n38);
nor (n33,n34,n36);
and (n34,n35,n28);
and (n36,n29,n37);
not (n37,n35);
nand (n38,n39,n42);
or (n39,n40,n35);
not (n40,n41);
nand (n42,n35,n40);
nand (n43,n38,n44);
nor (n44,n45,n48);
and (n45,n46,n28);
not (n46,n47);
and (n48,n47,n29);
nand (n49,n50,n70);
or (n50,n51,n59);
not (n51,n52);
nand (n52,n53,n57);
or (n53,n54,n55);
not (n55,n56);
or (n57,n58,n56);
not (n58,n54);
nand (n59,n60,n67);
not (n60,n61);
nand (n61,n62,n66);
or (n62,n63,n65);
not (n63,n64);
nand (n66,n63,n65);
nand (n67,n68,n69);
or (n68,n65,n58);
nand (n69,n58,n65);
nand (n70,n61,n71);
xnor (n71,n72,n54);
not (n72,n73);
nand (n74,n75,n85);
or (n75,n76,n78);
not (n76,n77);
not (n78,n79);
nor (n79,n80,n82);
not (n80,n81);
nand (n82,n83,n84);
or (n83,n58,n81);
nand (n84,n81,n58);
nand (n85,n82,n86);
and (n87,n21,n49);
xor (n88,n89,n125);
xor (n89,n90,n115);
nand (n90,n91,n107);
or (n91,n92,n98);
not (n92,n93);
nand (n93,n94,n97);
or (n94,n95,n64);
not (n95,n96);
or (n97,n96,n63);
nand (n98,n99,n106);
nor (n99,n100,n104);
and (n100,n101,n103);
not (n101,n102);
and (n104,n102,n105);
not (n105,n103);
xor (n106,n101,n63);
nand (n107,n108,n114);
not (n108,n109);
nor (n109,n110,n112);
and (n110,n111,n63);
and (n112,n64,n113);
not (n113,n111);
not (n114,n99);
nand (n115,n116,n118);
or (n116,n117,n31);
not (n117,n44);
or (n118,n119,n120);
not (n119,n38);
nor (n120,n121,n124);
and (n121,n122,n29);
not (n122,n123);
and (n124,n123,n28);
nand (n125,n126,n128);
or (n126,n59,n127);
not (n127,n71);
or (n128,n60,n129);
not (n129,n130);
nor (n130,n131,n134);
and (n131,n132,n58);
not (n132,n133);
and (n134,n133,n54);
xor (n135,n136,n175);
xor (n136,n137,n152);
nand (n137,n138,n149);
or (n138,n139,n145);
nand (n139,n140,n144);
or (n140,n141,n143);
not (n141,n142);
nand (n144,n143,n141);
nor (n145,n139,n146);
nor (n146,n147,n150);
and (n147,n148,n149);
not (n148,n143);
and (n150,n143,n151);
not (n151,n149);
nand (n152,n153,n169);
or (n153,n154,n163);
nand (n154,n155,n159);
nand (n155,n156,n158);
or (n156,n157,n40);
nand (n158,n40,n157);
not (n159,n160);
nand (n160,n161,n162);
or (n161,n151,n157);
nand (n162,n157,n151);
not (n163,n164);
nor (n164,n165,n168);
and (n165,n166,n40);
not (n166,n167);
and (n168,n167,n41);
or (n169,n159,n170);
nor (n170,n171,n173);
and (n171,n40,n172);
and (n173,n41,n174);
not (n174,n172);
nand (n175,n176,n192);
or (n176,n177,n187);
nand (n177,n178,n184);
not (n178,n179);
nand (n179,n180,n183);
or (n180,n181,n29);
not (n181,n182);
nand (n183,n29,n181);
nand (n184,n185,n186);
nand (n185,n181,n103);
nand (n186,n182,n105);
nor (n187,n188,n191);
and (n188,n189,n103);
not (n189,n190);
and (n191,n190,n105);
or (n192,n178,n193);
nor (n193,n194,n195);
and (n194,n105,n27);
and (n195,n103,n26);
xor (n196,n197,n299);
xor (n197,n198,n239);
xor (n198,n199,n213);
xor (n199,n200,n205);
nand (n200,n201,n203);
or (n201,n78,n202);
not (n202,n86);
or (n203,n204,n55);
not (n204,n82);
nand (n205,n206,n212);
or (n206,n207,n211);
not (n207,n208);
nor (n208,n209,n210);
and (n209,n172,n149);
and (n210,n174,n151);
not (n211,n145);
nand (n212,n139,n149);
or (n213,n214,n238);
and (n214,n215,n230);
xor (n215,n216,n223);
nand (n216,n217,n222);
or (n217,n218,n154);
not (n218,n219);
nor (n219,n220,n221);
and (n220,n123,n41);
and (n221,n122,n40);
nand (n222,n160,n164);
nand (n223,n224,n229);
or (n224,n225,n177);
not (n225,n226);
nor (n226,n227,n228);
and (n227,n113,n105);
and (n228,n111,n103);
or (n229,n178,n187);
nand (n230,n231,n232);
or (n231,n92,n99);
nand (n232,n233,n237);
not (n233,n234);
nor (n234,n235,n236);
and (n235,n63,n133);
and (n236,n132,n64);
not (n237,n98);
and (n238,n216,n223);
or (n239,n240,n298);
and (n240,n241,n275);
xor (n241,n242,n243);
not (n242,n205);
or (n243,n244,n274);
and (n244,n245,n267);
xor (n245,n246,n260);
nand (n246,n247,n142);
or (n247,n248,n254);
nand (n248,n249,n253);
or (n249,n250,n252);
not (n250,n251);
nand (n253,n250,n252);
not (n254,n255);
nand (n255,n256,n257);
not (n256,n248);
nand (n257,n258,n259);
or (n258,n142,n250);
nand (n259,n250,n142);
nand (n260,n261,n266);
or (n261,n262,n211);
not (n262,n263);
nand (n263,n264,n265);
or (n264,n167,n151);
nand (n265,n151,n167);
nand (n266,n208,n139);
nand (n267,n268,n273);
or (n268,n269,n31);
not (n269,n270);
nand (n270,n271,n272);
or (n271,n29,n189);
or (n272,n28,n190);
nand (n273,n38,n24);
and (n274,n246,n260);
or (n275,n276,n297);
and (n276,n277,n290);
xor (n277,n278,n283);
nand (n278,n279,n282);
or (n279,n280,n78);
not (n280,n281);
nand (n282,n82,n77);
nand (n283,n284,n289);
or (n284,n285,n177);
not (n285,n286);
nor (n286,n287,n288);
and (n287,n95,n105);
and (n288,n96,n103);
nand (n289,n179,n226);
nand (n290,n291,n296);
or (n291,n154,n292);
not (n292,n293);
nor (n293,n294,n295);
and (n294,n46,n40);
and (n295,n47,n41);
or (n296,n159,n218);
and (n297,n278,n283);
and (n298,n242,n243);
or (n299,n300,n328);
and (n300,n301,n304);
xor (n301,n302,n303);
xor (n302,n20,n74);
xor (n303,n215,n230);
or (n304,n305,n327);
and (n305,n306,n320);
xor (n306,n307,n313);
nand (n307,n308,n312);
or (n308,n309,n98);
nor (n309,n310,n311);
and (n310,n64,n72);
and (n311,n63,n73);
nand (n312,n233,n114);
nand (n313,n314,n319);
or (n314,n315,n59);
not (n315,n316);
nor (n316,n317,n318);
and (n317,n202,n58);
and (n318,n86,n54);
nand (n319,n61,n52);
not (n320,n321);
nor (n321,n322,n326);
and (n322,n254,n323);
nor (n323,n324,n325);
and (n324,n174,n141);
and (n325,n172,n142);
nor (n326,n256,n141);
and (n327,n307,n313);
and (n328,n302,n303);
or (n329,n330,n386);
and (n330,n331,n385);
xor (n331,n332,n333);
xor (n332,n241,n275);
or (n333,n334,n384);
and (n334,n335,n383);
xor (n335,n336,n360);
or (n336,n337,n359);
and (n337,n338,n353);
xor (n338,n339,n346);
nand (n339,n340,n345);
or (n340,n341,n177);
not (n341,n342);
nand (n342,n343,n344);
or (n343,n133,n105);
nand (n344,n105,n133);
nand (n345,n286,n179);
nand (n346,n347,n352);
or (n347,n348,n154);
not (n348,n349);
nor (n349,n350,n351);
and (n350,n26,n40);
and (n351,n27,n41);
nand (n352,n160,n293);
nand (n353,n354,n358);
or (n354,n98,n355);
nor (n355,n356,n357);
and (n356,n56,n63);
and (n357,n64,n55);
or (n358,n309,n99);
and (n359,n339,n346);
or (n360,n361,n382);
and (n361,n362,n375);
xor (n362,n363,n370);
nand (n363,n364,n369);
or (n364,n365,n211);
not (n365,n366);
nor (n366,n367,n368);
and (n367,n122,n151);
and (n368,n123,n149);
nand (n369,n263,n139);
nand (n370,n371,n374);
or (n371,n372,n78);
not (n372,n373);
nand (n374,n82,n281);
nand (n375,n376,n381);
or (n376,n377,n31);
not (n377,n378);
nor (n378,n379,n380);
and (n379,n113,n28);
and (n380,n111,n29);
nand (n381,n38,n270);
and (n382,n363,n370);
xor (n383,n245,n267);
and (n384,n336,n360);
xor (n385,n301,n304);
and (n386,n332,n333);
or (n387,n388,n508);
and (n388,n389,n416);
xor (n389,n390,n415);
or (n390,n391,n414);
and (n391,n392,n395);
xor (n392,n393,n394);
xor (n393,n277,n290);
xor (n394,n306,n320);
or (n395,n396,n413);
and (n396,n397,n405);
xor (n397,n398,n321);
nand (n398,n399,n404);
or (n399,n400,n59);
not (n400,n401);
nor (n401,n402,n403);
and (n402,n76,n58);
and (n403,n77,n54);
nand (n404,n61,n316);
nand (n405,n406,n252);
nor (n406,n407,n412);
and (n407,n408,n409);
not (n408,n154);
nor (n409,n410,n411);
and (n410,n189,n40);
and (n411,n190,n41);
and (n412,n160,n349);
and (n413,n398,n321);
and (n414,n393,n394);
xor (n415,n331,n385);
or (n416,n417,n507);
and (n417,n418,n472);
xor (n418,n419,n420);
xor (n419,n335,n383);
or (n420,n421,n471);
and (n421,n422,n470);
xor (n422,n423,n447);
or (n423,n424,n446);
and (n424,n425,n438);
xor (n425,n426,n433);
nand (n426,n427,n432);
or (n427,n428,n59);
not (n428,n429);
nor (n429,n430,n431);
and (n430,n280,n58);
and (n431,n281,n54);
nand (n432,n401,n61);
nand (n433,n434,n437);
or (n434,n435,n78);
not (n435,n436);
nand (n437,n82,n373);
nand (n438,n439,n441);
or (n439,n440,n256);
not (n440,n323);
or (n441,n255,n442);
not (n442,n443);
or (n443,n444,n445);
and (n444,n166,n142);
and (n445,n167,n141);
and (n446,n426,n433);
or (n447,n448,n469);
and (n448,n449,n463);
xor (n449,n450,n457);
nand (n450,n451,n456);
or (n451,n452,n31);
not (n452,n453);
nor (n453,n454,n455);
and (n454,n95,n28);
and (n455,n96,n29);
nand (n456,n38,n378);
nand (n457,n458,n462);
or (n458,n459,n211);
nor (n459,n460,n461);
and (n460,n46,n149);
and (n461,n47,n151);
nand (n462,n366,n139);
nand (n463,n464,n468);
or (n464,n177,n465);
nor (n465,n466,n467);
and (n466,n105,n73);
and (n467,n103,n72);
or (n468,n178,n341);
and (n469,n450,n457);
xor (n470,n338,n353);
and (n471,n423,n447);
or (n472,n473,n506);
and (n473,n474,n477);
xor (n474,n475,n476);
xor (n475,n362,n375);
xor (n476,n397,n405);
and (n477,n478,n500);
or (n478,n479,n499);
and (n479,n480,n494);
xor (n480,n481,n487);
nand (n481,n482,n486);
or (n482,n483,n154);
nor (n483,n484,n485);
and (n484,n113,n41);
and (n485,n111,n40);
nand (n486,n409,n160);
nand (n487,n488,n493);
or (n488,n489,n59);
not (n489,n490);
nand (n490,n491,n492);
or (n491,n54,n372);
or (n492,n58,n373);
nand (n493,n61,n429);
nand (n494,n495,n498);
or (n495,n496,n78);
not (n496,n497);
nand (n498,n82,n436);
and (n499,n481,n487);
nand (n500,n501,n505);
or (n501,n98,n502);
nor (n502,n503,n504);
and (n503,n63,n86);
and (n504,n64,n202);
or (n505,n99,n355);
and (n506,n475,n476);
and (n507,n419,n420);
and (n508,n390,n415);
nand (n509,n14,n387);
nand (n510,n511,n1533);
or (n511,n512,n684);
not (n512,n513);
nor (n513,n514,n596);
nor (n514,n515,n516);
xor (n515,n389,n416);
or (n516,n517,n595);
and (n517,n518,n521);
xor (n518,n519,n520);
xor (n519,n392,n395);
xor (n520,n418,n472);
or (n521,n522,n594);
and (n522,n523,n558);
xor (n523,n524,n525);
xor (n524,n422,n470);
or (n525,n526,n557);
and (n526,n527,n555);
xor (n527,n528,n554);
or (n528,n529,n553);
and (n529,n530,n545);
xor (n530,n531,n538);
nand (n531,n532,n537);
or (n532,n533,n255);
not (n533,n534);
nor (n534,n535,n536);
and (n535,n122,n141);
and (n536,n123,n142);
nand (n537,n248,n443);
nand (n538,n539,n544);
or (n539,n540,n31);
not (n540,n541);
nand (n541,n542,n543);
or (n542,n29,n132);
or (n543,n28,n133);
nand (n544,n38,n453);
nand (n545,n546,n551);
or (n546,n211,n547);
not (n547,n548);
nor (n548,n549,n550);
and (n549,n151,n26);
and (n550,n27,n149);
or (n551,n459,n552);
not (n552,n139);
and (n553,n531,n538);
xor (n554,n449,n463);
nand (n555,n556,n405);
or (n556,n252,n406);
and (n557,n528,n554);
or (n558,n559,n593);
and (n559,n560,n592);
xor (n560,n561,n562);
xor (n561,n425,n438);
or (n562,n563,n591);
and (n563,n564,n580);
xor (n564,n565,n573);
nand (n565,n566,n571);
or (n566,n567,n177);
not (n567,n568);
nor (n568,n569,n570);
and (n569,n55,n105);
and (n570,n56,n103);
nand (n571,n572,n179);
not (n572,n465);
nand (n573,n574,n579);
or (n574,n575,n98);
not (n575,n576);
nand (n576,n577,n578);
or (n577,n64,n76);
or (n578,n63,n77);
or (n579,n99,n502);
nand (n580,n581,n590);
or (n581,n582,n585);
nand (n582,n583,n252);
not (n583,n584);
not (n585,n586);
nor (n586,n587,n589);
and (n587,n174,n588);
not (n588,n252);
and (n589,n172,n252);
or (n590,n588,n583);
and (n591,n565,n573);
xor (n592,n478,n500);
and (n593,n561,n562);
and (n594,n524,n525);
and (n595,n519,n520);
nor (n596,n597,n598);
xor (n597,n518,n521);
or (n598,n599,n683);
and (n599,n600,n682);
xor (n600,n601,n602);
xor (n601,n474,n477);
or (n602,n603,n681);
and (n603,n604,n680);
xor (n604,n605,n673);
or (n605,n606,n672);
and (n606,n607,n649);
xor (n607,n608,n626);
or (n608,n609,n625);
and (n609,n610,n618);
xor (n610,n611,n612);
and (n611,n82,n497);
nand (n612,n613,n614);
or (n613,n583,n585);
or (n614,n615,n582);
nor (n615,n616,n617);
and (n616,n588,n167);
and (n617,n252,n166);
nand (n618,n619,n624);
or (n619,n255,n620);
not (n620,n621);
nor (n621,n622,n623);
and (n622,n46,n141);
and (n623,n47,n142);
nand (n624,n248,n534);
and (n625,n611,n612);
or (n626,n627,n648);
and (n627,n628,n642);
xor (n628,n629,n636);
nand (n629,n630,n635);
or (n630,n631,n211);
not (n631,n632);
nand (n632,n633,n634);
or (n633,n149,n189);
or (n634,n151,n190);
nand (n635,n548,n139);
nand (n636,n637,n641);
or (n637,n638,n177);
nor (n638,n639,n640);
and (n639,n202,n103);
and (n640,n86,n105);
nand (n641,n568,n179);
nand (n642,n643,n644);
or (n643,n575,n99);
or (n644,n98,n645);
nor (n645,n646,n647);
and (n646,n281,n63);
and (n647,n64,n280);
and (n648,n629,n636);
or (n649,n650,n671);
and (n650,n651,n665);
xor (n651,n652,n659);
nand (n652,n653,n658);
or (n653,n654,n59);
not (n654,n655);
nand (n655,n656,n657);
or (n656,n54,n435);
or (n657,n58,n436);
nand (n658,n490,n61);
nand (n659,n660,n664);
or (n660,n154,n661);
nor (n661,n662,n663);
and (n662,n95,n41);
and (n663,n96,n40);
or (n664,n159,n483);
nand (n665,n666,n670);
or (n666,n31,n667);
nor (n667,n668,n669);
and (n668,n72,n29);
and (n669,n73,n28);
or (n670,n119,n540);
and (n671,n652,n659);
and (n672,n608,n626);
or (n673,n674,n679);
and (n674,n675,n678);
xor (n675,n676,n677);
xor (n676,n480,n494);
xor (n677,n530,n545);
xor (n678,n564,n580);
and (n679,n676,n677);
xor (n680,n527,n555);
and (n681,n605,n673);
xor (n682,n523,n558);
and (n683,n601,n602);
not (n684,n685);
nand (n685,n686,n1518);
or (n686,n687,n1448);
not (n687,n688);
nand (n688,n689,n1435);
or (n689,n690,n1141);
not (n690,n691);
nand (n691,n692,n1130,n1140);
nand (n692,n693,n886,n990);
nand (n693,n694,n850);
not (n694,n695);
xor (n695,n696,n809);
xor (n696,n697,n738);
xor (n697,n698,n717);
xor (n698,n699,n708);
nand (n699,n700,n704);
or (n700,n177,n701);
nor (n701,n702,n703);
and (n702,n496,n103);
and (n703,n105,n497);
or (n704,n178,n705);
nor (n705,n706,n707);
and (n706,n105,n436);
and (n707,n103,n435);
nand (n708,n709,n713);
or (n709,n211,n710);
nor (n710,n711,n712);
and (n711,n151,n56);
and (n712,n149,n55);
or (n713,n714,n552);
nor (n714,n715,n716);
and (n715,n151,n73);
and (n716,n149,n72);
nand (n717,n718,n737);
or (n718,n719,n726);
not (n719,n720);
nand (n720,n721,n103);
nand (n721,n722,n723);
or (n722,n497,n182);
nand (n723,n724,n28);
not (n724,n725);
and (n725,n497,n182);
not (n726,n727);
nand (n727,n728,n733);
or (n728,n729,n255);
not (n729,n730);
nand (n730,n731,n732);
or (n731,n142,n132);
or (n732,n141,n133);
nand (n733,n248,n734);
nand (n734,n735,n736);
or (n735,n142,n95);
or (n736,n141,n96);
or (n737,n727,n720);
xor (n738,n739,n789);
xor (n739,n740,n761);
or (n740,n741,n760);
and (n741,n742,n750);
xor (n742,n743,n744);
and (n743,n179,n497);
nand (n744,n745,n749);
or (n745,n746,n255);
nor (n746,n747,n748);
and (n747,n72,n142);
and (n748,n73,n141);
nand (n749,n248,n730);
nand (n750,n751,n756);
or (n751,n154,n752);
not (n752,n753);
nor (n753,n754,n755);
and (n754,n280,n40);
and (n755,n281,n41);
or (n756,n159,n757);
nor (n757,n758,n759);
and (n758,n77,n40);
and (n759,n76,n41);
and (n760,n743,n744);
or (n761,n762,n788);
and (n762,n763,n782);
xor (n763,n764,n773);
nand (n764,n765,n769);
or (n765,n31,n766);
nor (n766,n767,n768);
and (n767,n435,n29);
and (n768,n436,n28);
or (n769,n119,n770);
nor (n770,n771,n772);
and (n771,n373,n28);
and (n772,n372,n29);
nand (n773,n774,n778);
or (n774,n775,n582);
nor (n775,n776,n777);
and (n776,n588,n96);
and (n777,n252,n95);
or (n778,n779,n583);
nor (n779,n780,n781);
and (n780,n588,n111);
and (n781,n252,n113);
nand (n782,n783,n787);
or (n783,n211,n784);
nor (n784,n785,n786);
and (n785,n151,n86);
and (n786,n149,n202);
or (n787,n710,n552);
and (n788,n764,n773);
xor (n789,n790,n803);
xor (n790,n791,n797);
nand (n791,n792,n793);
or (n792,n154,n757);
or (n793,n794,n159);
nor (n794,n795,n796);
and (n795,n202,n41);
and (n796,n86,n40);
nand (n797,n798,n799);
or (n798,n31,n770);
or (n799,n119,n800);
nor (n800,n801,n802);
and (n801,n280,n29);
and (n802,n281,n28);
nand (n803,n804,n805);
or (n804,n779,n582);
or (n805,n806,n583);
nor (n806,n807,n808);
and (n807,n588,n190);
and (n808,n252,n189);
or (n809,n810,n849);
and (n810,n811,n848);
xor (n811,n812,n825);
and (n812,n813,n819);
and (n813,n814,n29);
nand (n814,n815,n816);
or (n815,n497,n35);
nand (n816,n817,n40);
not (n817,n818);
and (n818,n497,n35);
nand (n819,n820,n824);
or (n820,n255,n821);
nor (n821,n822,n823);
and (n822,n141,n56);
and (n823,n142,n55);
or (n824,n256,n746);
or (n825,n826,n847);
and (n826,n827,n841);
xor (n827,n828,n835);
nand (n828,n829,n834);
or (n829,n830,n154);
not (n830,n831);
nor (n831,n832,n833);
and (n832,n373,n41);
and (n833,n372,n40);
nand (n834,n160,n753);
nand (n835,n836,n840);
or (n836,n31,n837);
nor (n837,n838,n839);
and (n838,n29,n496);
and (n839,n28,n497);
or (n840,n119,n766);
nand (n841,n842,n846);
or (n842,n582,n843);
nor (n843,n844,n845);
and (n844,n588,n133);
and (n845,n252,n132);
or (n846,n775,n583);
and (n847,n828,n835);
xor (n848,n742,n750);
and (n849,n812,n825);
not (n850,n851);
or (n851,n852,n885);
and (n852,n853,n884);
xor (n853,n854,n855);
xor (n854,n763,n782);
or (n855,n856,n883);
and (n856,n857,n865);
xor (n857,n858,n864);
nand (n858,n859,n863);
or (n859,n211,n860);
nor (n860,n861,n862);
and (n861,n151,n77);
and (n862,n149,n76);
or (n863,n784,n552);
xor (n864,n813,n819);
or (n865,n866,n882);
and (n866,n867,n875);
xor (n867,n868,n869);
and (n868,n38,n497);
nand (n869,n870,n874);
or (n870,n871,n582);
nor (n871,n872,n873);
and (n872,n588,n73);
and (n873,n252,n72);
or (n874,n843,n583);
nand (n875,n876,n881);
or (n876,n154,n877);
not (n877,n878);
nand (n878,n879,n880);
or (n879,n41,n435);
or (n880,n40,n436);
or (n881,n159,n830);
and (n882,n868,n869);
and (n883,n858,n864);
xor (n884,n811,n848);
and (n885,n854,n855);
nor (n886,n887,n927);
not (n887,n888);
or (n888,n889,n890);
xor (n889,n853,n884);
or (n890,n891,n926);
and (n891,n892,n925);
xor (n892,n893,n894);
xor (n893,n827,n841);
or (n894,n895,n924);
and (n895,n896,n909);
xor (n896,n897,n903);
nand (n897,n898,n902);
or (n898,n255,n899);
nor (n899,n900,n901);
and (n900,n141,n86);
and (n901,n142,n202);
or (n902,n256,n821);
nand (n903,n904,n908);
or (n904,n211,n905);
nor (n905,n906,n907);
and (n906,n151,n281);
and (n907,n149,n280);
or (n908,n860,n552);
and (n909,n910,n917);
nor (n910,n911,n40);
nor (n911,n912,n915);
and (n912,n913,n151);
not (n913,n914);
and (n914,n497,n157);
and (n915,n496,n916);
not (n916,n157);
nand (n917,n918,n923);
or (n918,n582,n919);
not (n919,n920);
nor (n920,n921,n922);
and (n921,n56,n252);
and (n922,n55,n588);
or (n923,n871,n583);
and (n924,n897,n903);
xor (n925,n857,n865);
and (n926,n893,n894);
nand (n927,n928,n984);
not (n928,n929);
nor (n929,n930,n959);
xor (n930,n931,n958);
xor (n931,n932,n957);
or (n932,n933,n956);
and (n933,n934,n950);
xor (n934,n935,n942);
nand (n935,n936,n941);
or (n936,n937,n154);
not (n937,n938);
nand (n938,n939,n940);
or (n939,n40,n497);
or (n940,n41,n496);
nand (n941,n160,n878);
nand (n942,n943,n948);
or (n943,n944,n255);
not (n944,n945);
nand (n945,n946,n947);
or (n946,n142,n76);
or (n947,n141,n77);
nand (n948,n949,n248);
not (n949,n899);
nand (n950,n951,n955);
or (n951,n211,n952);
nor (n952,n953,n954);
and (n953,n151,n373);
and (n954,n149,n372);
or (n955,n905,n552);
and (n956,n935,n942);
xor (n957,n867,n875);
xor (n958,n896,n909);
or (n959,n960,n983);
and (n960,n961,n982);
xor (n961,n962,n963);
xor (n962,n910,n917);
or (n963,n964,n981);
and (n964,n965,n974);
xor (n965,n966,n967);
and (n966,n160,n497);
nand (n967,n968,n969);
or (n968,n583,n919);
or (n969,n970,n582);
not (n970,n971);
nand (n971,n972,n973);
or (n972,n86,n588);
nand (n973,n588,n86);
nand (n974,n975,n980);
or (n975,n976,n255);
not (n976,n977);
nand (n977,n978,n979);
or (n978,n142,n280);
or (n979,n141,n281);
nand (n980,n248,n945);
and (n981,n966,n967);
xor (n982,n934,n950);
and (n983,n962,n963);
not (n984,n985);
nor (n985,n986,n987);
xor (n986,n892,n925);
or (n987,n988,n989);
and (n988,n931,n958);
and (n989,n932,n957);
or (n990,n991,n1129);
and (n991,n992,n1019);
xor (n992,n993,n1018);
or (n993,n994,n1017);
and (n994,n995,n1016);
xor (n995,n996,n1002);
nand (n996,n997,n1001);
or (n997,n211,n998);
nor (n998,n999,n1000);
and (n999,n151,n436);
and (n1000,n149,n435);
or (n1001,n952,n552);
nor (n1002,n1003,n1011);
not (n1003,n1004);
nand (n1004,n1005,n1010);
or (n1005,n582,n1006);
not (n1006,n1007);
nor (n1007,n1008,n1009);
and (n1008,n77,n252);
and (n1009,n76,n588);
nand (n1010,n971,n584);
nand (n1011,n1012,n149);
nand (n1012,n1013,n1015);
or (n1013,n1014,n142);
and (n1014,n497,n143);
or (n1015,n497,n143);
xor (n1016,n965,n974);
and (n1017,n996,n1002);
xor (n1018,n961,n982);
or (n1019,n1020,n1128);
and (n1020,n1021,n1045);
xor (n1021,n1022,n1044);
or (n1022,n1023,n1043);
and (n1023,n1024,n1039);
xor (n1024,n1025,n1032);
nand (n1025,n1026,n1031);
or (n1026,n1027,n255);
not (n1027,n1028);
nor (n1028,n1029,n1030);
and (n1029,n372,n141);
and (n1030,n373,n142);
nand (n1031,n248,n977);
nand (n1032,n1033,n1038);
or (n1033,n1034,n211);
not (n1034,n1035);
nand (n1035,n1036,n1037);
or (n1036,n151,n497);
or (n1037,n496,n149);
or (n1038,n998,n552);
nand (n1039,n1040,n1042);
or (n1040,n1041,n1003);
not (n1041,n1011);
or (n1042,n1004,n1011);
and (n1043,n1025,n1032);
xor (n1044,n995,n1016);
or (n1045,n1046,n1127);
and (n1046,n1047,n1068);
xor (n1047,n1048,n1067);
or (n1048,n1049,n1066);
and (n1049,n1050,n1059);
xor (n1050,n1051,n1052);
and (n1051,n139,n497);
nand (n1052,n1053,n1058);
or (n1053,n1054,n255);
not (n1054,n1055);
nor (n1055,n1056,n1057);
and (n1056,n435,n141);
and (n1057,n436,n142);
nand (n1058,n248,n1028);
nand (n1059,n1060,n1061);
or (n1060,n583,n1006);
or (n1061,n582,n1062);
not (n1062,n1063);
nor (n1063,n1064,n1065);
and (n1064,n280,n588);
and (n1065,n281,n252);
and (n1066,n1051,n1052);
xor (n1067,n1024,n1039);
nand (n1068,n1069,n1126);
or (n1069,n1070,n1086);
nor (n1070,n1071,n1072);
xor (n1071,n1050,n1059);
and (n1072,n1073,n1080);
nand (n1073,n1074,n1075);
nand (n1074,n1063,n584);
nand (n1075,n1076,n1079);
nor (n1076,n1077,n1078);
and (n1077,n372,n588);
and (n1078,n373,n252);
not (n1079,n582);
not (n1080,n1081);
nand (n1081,n1082,n142);
nand (n1082,n1083,n1085);
or (n1083,n1084,n252);
and (n1084,n497,n251);
or (n1085,n497,n251);
nor (n1086,n1087,n1125);
and (n1087,n1088,n1099);
nand (n1088,n1089,n1093);
nor (n1089,n1090,n1092);
and (n1090,n1091,n1080);
not (n1091,n1073);
and (n1092,n1073,n1081);
nor (n1093,n1094,n1095);
and (n1094,n248,n1055);
and (n1095,n254,n1096);
nand (n1096,n1097,n1098);
or (n1097,n141,n497);
or (n1098,n496,n142);
nand (n1099,n1100,n1123);
or (n1100,n1101,n1115);
not (n1101,n1102);
and (n1102,n1103,n1113);
nand (n1103,n1104,n1109);
or (n1104,n583,n1105);
not (n1105,n1106);
nor (n1106,n1107,n1108);
and (n1107,n435,n588);
and (n1108,n436,n252);
nand (n1109,n1110,n1079);
nand (n1110,n1111,n1112);
or (n1111,n588,n497);
or (n1112,n252,n496);
nor (n1113,n1114,n588);
and (n1114,n497,n584);
not (n1115,n1116);
nand (n1116,n1117,n1122);
not (n1117,n1118);
nand (n1118,n1119,n1121);
or (n1119,n583,n1120);
not (n1120,n1076);
nand (n1121,n1106,n1079);
nand (n1122,n248,n497);
nand (n1123,n1124,n1118);
not (n1124,n1122);
nor (n1125,n1089,n1093);
nand (n1126,n1071,n1072);
and (n1127,n1048,n1067);
and (n1128,n1022,n1044);
and (n1129,n993,n1018);
nand (n1130,n1131,n693);
or (n1131,n1132,n1134);
not (n1132,n1133);
nand (n1133,n889,n890);
not (n1134,n1135);
nand (n1135,n888,n1136);
nand (n1136,n1137,n1139);
or (n1137,n985,n1138);
nand (n1138,n930,n959);
nand (n1139,n986,n987);
nand (n1140,n695,n851);
not (n1141,n1142);
nor (n1142,n1143,n1398);
nor (n1143,n1144,n1375);
xor (n1144,n1145,n1297);
xor (n1145,n1146,n1215);
xor (n1146,n1147,n1195);
xor (n1147,n1148,n1180);
or (n1148,n1149,n1179);
and (n1149,n1150,n1170);
xor (n1150,n1151,n1161);
nand (n1151,n1152,n1157);
or (n1152,n1153,n154);
not (n1153,n1154);
nand (n1154,n1155,n1156);
or (n1155,n41,n72);
or (n1156,n40,n73);
nand (n1157,n160,n1158);
nor (n1158,n1159,n1160);
and (n1159,n132,n40);
and (n1160,n133,n41);
nand (n1161,n1162,n1166);
or (n1162,n31,n1163);
nor (n1163,n1164,n1165);
and (n1164,n28,n86);
and (n1165,n29,n202);
nand (n1166,n38,n1167);
nor (n1167,n1168,n1169);
and (n1168,n55,n28);
and (n1169,n56,n29);
nand (n1170,n1171,n1175);
or (n1171,n211,n1172);
nor (n1172,n1173,n1174);
and (n1173,n151,n96);
and (n1174,n149,n95);
or (n1175,n1176,n552);
nor (n1176,n1177,n1178);
and (n1177,n151,n111);
and (n1178,n149,n113);
and (n1179,n1151,n1161);
xor (n1180,n1181,n1189);
xor (n1181,n1182,n1186);
nand (n1182,n1183,n1185);
or (n1183,n1184,n31);
not (n1184,n1167);
or (n1185,n667,n119);
nand (n1186,n1187,n1188);
or (n1187,n1176,n211);
nand (n1188,n139,n632);
nand (n1189,n1190,n1194);
or (n1190,n177,n1191);
nor (n1191,n1192,n1193);
and (n1192,n105,n77);
and (n1193,n103,n76);
or (n1194,n178,n638);
xor (n1195,n1196,n1211);
xor (n1196,n1197,n1204);
nand (n1197,n1198,n1203);
or (n1198,n1199,n255);
not (n1199,n1200);
nand (n1200,n1201,n1202);
or (n1201,n142,n26);
or (n1202,n141,n27);
nand (n1203,n248,n621);
nand (n1204,n1205,n1210);
or (n1205,n1206,n59);
not (n1206,n1207);
nand (n1207,n1208,n1209);
or (n1208,n58,n497);
or (n1209,n54,n496);
nand (n1210,n655,n61);
nand (n1211,n1212,n1214);
or (n1212,n154,n1213);
not (n1213,n1158);
or (n1214,n159,n661);
or (n1215,n1216,n1296);
and (n1216,n1217,n1253);
xor (n1217,n1218,n1219);
xor (n1218,n1150,n1170);
xor (n1219,n1220,n1237);
xor (n1220,n1221,n1228);
nand (n1221,n1222,n1226);
or (n1222,n1223,n177);
nor (n1223,n1224,n1225);
and (n1224,n280,n103);
and (n1225,n281,n105);
nand (n1226,n1227,n179);
not (n1227,n1191);
nand (n1228,n1229,n1233);
or (n1229,n1230,n98);
nor (n1230,n1231,n1232);
and (n1231,n63,n436);
and (n1232,n64,n435);
or (n1233,n99,n1234);
nor (n1234,n1235,n1236);
and (n1235,n63,n373);
and (n1236,n64,n372);
and (n1237,n1238,n1243);
nor (n1238,n1239,n63);
nor (n1239,n1240,n1242);
and (n1240,n1241,n105);
nand (n1241,n497,n102);
and (n1242,n496,n101);
nand (n1243,n1244,n1249);
or (n1244,n583,n1245);
not (n1245,n1246);
nor (n1246,n1247,n1248);
and (n1247,n46,n588);
and (n1248,n47,n252);
or (n1249,n1250,n582);
nor (n1250,n1251,n1252);
and (n1251,n26,n252);
and (n1252,n27,n588);
or (n1253,n1254,n1295);
and (n1254,n1255,n1276);
xor (n1255,n1256,n1257);
xor (n1256,n1238,n1243);
or (n1257,n1258,n1275);
and (n1258,n1259,n1268);
xor (n1259,n1260,n1261);
and (n1260,n114,n497);
nand (n1261,n1262,n1264);
or (n1262,n1263,n255);
not (n1263,n734);
nand (n1264,n248,n1265);
nor (n1265,n1266,n1267);
and (n1266,n113,n141);
and (n1267,n111,n142);
nand (n1268,n1269,n1274);
or (n1269,n1270,n159);
not (n1270,n1271);
nand (n1271,n1272,n1273);
or (n1272,n41,n55);
or (n1273,n40,n56);
or (n1274,n154,n794);
and (n1275,n1260,n1261);
or (n1276,n1277,n1294);
and (n1277,n1278,n1288);
xor (n1278,n1279,n1285);
nand (n1279,n1280,n1281);
or (n1280,n800,n31);
nand (n1281,n1282,n38);
nand (n1282,n1283,n1284);
or (n1283,n29,n76);
or (n1284,n28,n77);
nand (n1285,n1286,n1287);
or (n1286,n806,n582);
or (n1287,n1250,n583);
nand (n1288,n1289,n1290);
or (n1289,n705,n177);
or (n1290,n1291,n178);
nor (n1291,n1292,n1293);
and (n1292,n105,n373);
and (n1293,n103,n372);
and (n1294,n1279,n1285);
and (n1295,n1256,n1257);
and (n1296,n1218,n1219);
xor (n1297,n1298,n1336);
xor (n1298,n1299,n1302);
or (n1299,n1300,n1301);
and (n1300,n1220,n1237);
and (n1301,n1221,n1228);
xor (n1302,n1303,n1320);
xor (n1303,n1304,n1307);
nand (n1304,n1305,n1306);
or (n1305,n98,n1234);
or (n1306,n99,n645);
xor (n1307,n1308,n1314);
nor (n1308,n1309,n58);
nor (n1309,n1310,n1312);
and (n1310,n1311,n63);
nand (n1311,n497,n65);
and (n1312,n496,n1313);
not (n1313,n65);
nand (n1314,n1315,n1319);
or (n1315,n1316,n582);
nor (n1316,n1317,n1318);
and (n1317,n122,n252);
and (n1318,n123,n588);
or (n1319,n615,n583);
or (n1320,n1321,n1335);
and (n1321,n1322,n1328);
xor (n1322,n1323,n1324);
nor (n1323,n60,n496);
nand (n1324,n1325,n1326);
or (n1325,n582,n1245);
nand (n1326,n1327,n584);
not (n1327,n1316);
nand (n1328,n1329,n1334);
or (n1329,n255,n1330);
not (n1330,n1331);
nand (n1331,n1332,n1333);
or (n1332,n142,n189);
or (n1333,n141,n190);
or (n1334,n256,n1199);
and (n1335,n1323,n1324);
or (n1336,n1337,n1374);
and (n1337,n1338,n1373);
xor (n1338,n1339,n1354);
or (n1339,n1340,n1353);
and (n1340,n1341,n1349);
xor (n1341,n1342,n1346);
nand (n1342,n1343,n1345);
or (n1343,n1344,n255);
not (n1344,n1265);
nand (n1345,n1331,n248);
nand (n1346,n1347,n1348);
or (n1347,n1270,n154);
nand (n1348,n160,n1154);
nand (n1349,n1350,n1352);
or (n1350,n31,n1351);
not (n1351,n1282);
or (n1352,n119,n1163);
and (n1353,n1342,n1346);
or (n1354,n1355,n1372);
and (n1355,n1356,n1366);
xor (n1356,n1357,n1363);
nand (n1357,n1358,n1362);
or (n1358,n211,n1359);
nor (n1359,n1360,n1361);
and (n1360,n151,n133);
and (n1361,n149,n132);
or (n1362,n1172,n552);
nand (n1363,n1364,n1365);
or (n1364,n177,n1291);
or (n1365,n1223,n178);
nand (n1366,n1367,n1371);
or (n1367,n98,n1368);
nor (n1368,n1369,n1370);
and (n1369,n496,n64);
and (n1370,n497,n63);
or (n1371,n1230,n99);
and (n1372,n1357,n1363);
xor (n1373,n1322,n1328);
and (n1374,n1339,n1354);
or (n1375,n1376,n1397);
and (n1376,n1377,n1380);
xor (n1377,n1378,n1379);
xor (n1378,n1338,n1373);
xor (n1379,n1217,n1253);
or (n1380,n1381,n1396);
and (n1381,n1382,n1385);
xor (n1382,n1383,n1384);
xor (n1383,n1356,n1366);
xor (n1384,n1341,n1349);
or (n1385,n1386,n1395);
and (n1386,n1387,n1392);
xor (n1387,n1388,n1391);
nand (n1388,n1389,n1390);
or (n1389,n211,n714);
or (n1390,n1359,n552);
and (n1391,n727,n719);
or (n1392,n1393,n1394);
and (n1393,n790,n803);
and (n1394,n791,n797);
and (n1395,n1388,n1391);
and (n1396,n1383,n1384);
and (n1397,n1378,n1379);
nand (n1398,n1399,n1428);
nor (n1399,n1400,n1423);
nor (n1400,n1401,n1414);
xor (n1401,n1402,n1413);
xor (n1402,n1403,n1404);
xor (n1403,n1255,n1276);
or (n1404,n1405,n1412);
and (n1405,n1406,n1409);
xor (n1406,n1407,n1408);
xor (n1407,n1278,n1288);
xor (n1408,n1259,n1268);
or (n1409,n1410,n1411);
and (n1410,n698,n717);
and (n1411,n699,n708);
and (n1412,n1407,n1408);
xor (n1413,n1382,n1385);
or (n1414,n1415,n1422);
and (n1415,n1416,n1421);
xor (n1416,n1417,n1418);
xor (n1417,n1387,n1392);
or (n1418,n1419,n1420);
and (n1419,n739,n789);
and (n1420,n740,n761);
xor (n1421,n1406,n1409);
and (n1422,n1417,n1418);
nor (n1423,n1424,n1427);
or (n1424,n1425,n1426);
and (n1425,n696,n809);
and (n1426,n697,n738);
xor (n1427,n1416,n1421);
nand (n1428,n1429,n1431);
not (n1429,n1430);
xor (n1430,n1377,n1380);
not (n1431,n1432);
or (n1432,n1433,n1434);
and (n1433,n1402,n1413);
and (n1434,n1403,n1404);
nor (n1435,n1436,n1447);
and (n1436,n1437,n1438);
not (n1437,n1143);
nand (n1438,n1439,n1446);
or (n1439,n1440,n1441);
not (n1440,n1428);
not (n1441,n1442);
nand (n1442,n1443,n1445);
or (n1443,n1400,n1444);
nand (n1444,n1424,n1427);
nand (n1445,n1401,n1414);
nand (n1446,n1430,n1432);
and (n1447,n1144,n1375);
not (n1448,n1449);
and (n1449,n1450,n1501);
nor (n1450,n1451,n1482);
nor (n1451,n1452,n1453);
xor (n1452,n600,n682);
or (n1453,n1454,n1481);
and (n1454,n1455,n1480);
xor (n1455,n1456,n1457);
xor (n1456,n560,n592);
or (n1457,n1458,n1479);
and (n1458,n1459,n1472);
xor (n1459,n1460,n1471);
or (n1460,n1461,n1470);
and (n1461,n1462,n1467);
xor (n1462,n1463,n1464);
and (n1463,n1308,n1314);
or (n1464,n1465,n1466);
and (n1465,n1196,n1211);
and (n1466,n1197,n1204);
or (n1467,n1468,n1469);
and (n1468,n1181,n1189);
and (n1469,n1182,n1186);
and (n1470,n1463,n1464);
xor (n1471,n607,n649);
or (n1472,n1473,n1478);
and (n1473,n1474,n1477);
xor (n1474,n1475,n1476);
xor (n1475,n628,n642);
xor (n1476,n610,n618);
xor (n1477,n651,n665);
and (n1478,n1475,n1476);
and (n1479,n1460,n1471);
xor (n1480,n604,n680);
and (n1481,n1456,n1457);
nor (n1482,n1483,n1484);
xor (n1483,n1455,n1480);
or (n1484,n1485,n1500);
and (n1485,n1486,n1499);
xor (n1486,n1487,n1488);
xor (n1487,n675,n678);
or (n1488,n1489,n1498);
and (n1489,n1490,n1495);
xor (n1490,n1491,n1494);
or (n1491,n1492,n1493);
and (n1492,n1303,n1320);
and (n1493,n1304,n1307);
xor (n1494,n1462,n1467);
or (n1495,n1496,n1497);
and (n1496,n1147,n1195);
and (n1497,n1148,n1180);
and (n1498,n1491,n1494);
xor (n1499,n1459,n1472);
and (n1500,n1487,n1488);
nor (n1501,n1502,n1513);
nor (n1502,n1503,n1504);
xor (n1503,n1486,n1499);
or (n1504,n1505,n1512);
and (n1505,n1506,n1511);
xor (n1506,n1507,n1508);
xor (n1507,n1474,n1477);
or (n1508,n1509,n1510);
and (n1509,n1298,n1336);
and (n1510,n1299,n1302);
xor (n1511,n1490,n1495);
and (n1512,n1507,n1508);
nor (n1513,n1514,n1515);
xor (n1514,n1506,n1511);
or (n1515,n1516,n1517);
and (n1516,n1145,n1297);
and (n1517,n1146,n1215);
not (n1518,n1519);
nand (n1519,n1520,n1527);
or (n1520,n1521,n1526);
not (n1521,n1522);
nor (n1522,n1523,n1502);
and (n1523,n1524,n1525);
nand (n1524,n1503,n1504);
nand (n1525,n1514,n1515);
not (n1526,n1450);
nor (n1527,n1528,n1532);
and (n1528,n1529,n1530);
not (n1529,n1451);
not (n1530,n1531);
nand (n1531,n1483,n1484);
and (n1532,n1452,n1453);
not (n1533,n1534);
nor (n1534,n1535,n514);
and (n1535,n1536,n1537);
nand (n1536,n516,n515);
nand (n1537,n597,n598);
nand (n1538,n510,n11);
not (n1539,n1540);
nand (n1540,n1541,n6);
not (n1541,n7);
wire s0n1542,s1n1542,notn1542;
or (n1542,s0n1542,s1n1542);
not(notn1542,n7);
and (s0n1542,notn1542,n1543);
and (s1n1542,n7,1'b0);
wire s0n1543,s1n1543,notn1543;
or (n1543,s0n1543,s1n1543);
not(notn1543,n6);
and (s0n1543,notn1543,n3);
and (s1n1543,n6,n1544);
xor (n1544,n1545,n2684);
xor (n1545,n1546,n2683);
xor (n1546,n1547,n2647);
xor (n1547,n1548,n2646);
xor (n1548,n1549,n2601);
xor (n1549,n1550,n2600);
xor (n1550,n1551,n2549);
xor (n1551,n1552,n2548);
xor (n1552,n1553,n2491);
xor (n1553,n1554,n2490);
xor (n1554,n1555,n2430);
xor (n1555,n1556,n2429);
xor (n1556,n1557,n2361);
xor (n1557,n1558,n2360);
xor (n1558,n1559,n2289);
xor (n1559,n1560,n48);
xor (n1560,n1561,n2209);
xor (n1561,n1562,n2208);
xor (n1562,n1563,n2128);
xor (n1563,n1564,n168);
xor (n1564,n1565,n2036);
xor (n1565,n1566,n2035);
or (n1566,n1567,n1942);
and (n1567,n1568,n209);
or (n1568,n1569,n1848);
and (n1569,n1570,n1847);
or (n1570,n1571,n1757);
and (n1571,n1572,n325);
or (n1572,n1573,n1663);
and (n1573,n1574,n1662);
and (n1574,n589,n1575);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
and (n1577,n172,n584);
and (n1578,n167,n252);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
and (n1583,n167,n584);
and (n1584,n123,n252);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1590);
and (n1588,n1589,n1248);
and (n1589,n123,n584);
and (n1590,n1591,n1592);
xor (n1591,n1589,n1248);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
and (n1594,n47,n584);
and (n1595,n27,n252);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
and (n1600,n27,n584);
and (n1601,n190,n252);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
and (n1606,n190,n584);
and (n1607,n111,n252);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
and (n1612,n111,n584);
and (n1613,n96,n252);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
and (n1618,n96,n584);
and (n1619,n133,n252);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
and (n1624,n133,n584);
and (n1625,n73,n252);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1631);
and (n1629,n1630,n921);
and (n1630,n73,n584);
and (n1631,n1632,n1633);
xor (n1632,n1630,n921);
or (n1633,n1634,n1637);
and (n1634,n1635,n1636);
and (n1635,n56,n584);
and (n1636,n86,n252);
and (n1637,n1638,n1639);
xor (n1638,n1635,n1636);
or (n1639,n1640,n1642);
and (n1640,n1641,n1008);
and (n1641,n86,n584);
and (n1642,n1643,n1644);
xor (n1643,n1641,n1008);
or (n1644,n1645,n1647);
and (n1645,n1646,n1065);
and (n1646,n77,n584);
and (n1647,n1648,n1649);
xor (n1648,n1646,n1065);
or (n1649,n1650,n1652);
and (n1650,n1651,n1078);
and (n1651,n281,n584);
and (n1652,n1653,n1654);
xor (n1653,n1651,n1078);
or (n1654,n1655,n1657);
and (n1655,n1656,n1108);
and (n1656,n373,n584);
and (n1657,n1658,n1659);
xor (n1658,n1656,n1108);
and (n1659,n1660,n1661);
and (n1660,n436,n584);
and (n1661,n497,n252);
and (n1662,n172,n251);
and (n1663,n1664,n1665);
xor (n1664,n1574,n1662);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n589,n1575);
and (n1668,n167,n251);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1580,n1581);
and (n1674,n123,n251);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1586,n1587);
and (n1680,n47,n251);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1591,n1592);
and (n1686,n27,n251);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
or (n1689,n1690,n1693);
and (n1690,n1691,n1692);
xor (n1691,n1597,n1598);
and (n1692,n190,n251);
and (n1693,n1694,n1695);
xor (n1694,n1691,n1692);
or (n1695,n1696,n1699);
and (n1696,n1697,n1698);
xor (n1697,n1603,n1604);
and (n1698,n111,n251);
and (n1699,n1700,n1701);
xor (n1700,n1697,n1698);
or (n1701,n1702,n1705);
and (n1702,n1703,n1704);
xor (n1703,n1609,n1610);
and (n1704,n96,n251);
and (n1705,n1706,n1707);
xor (n1706,n1703,n1704);
or (n1707,n1708,n1711);
and (n1708,n1709,n1710);
xor (n1709,n1615,n1616);
and (n1710,n133,n251);
and (n1711,n1712,n1713);
xor (n1712,n1709,n1710);
or (n1713,n1714,n1717);
and (n1714,n1715,n1716);
xor (n1715,n1621,n1622);
and (n1716,n73,n251);
and (n1717,n1718,n1719);
xor (n1718,n1715,n1716);
or (n1719,n1720,n1723);
and (n1720,n1721,n1722);
xor (n1721,n1627,n1628);
and (n1722,n56,n251);
and (n1723,n1724,n1725);
xor (n1724,n1721,n1722);
or (n1725,n1726,n1729);
and (n1726,n1727,n1728);
xor (n1727,n1632,n1633);
and (n1728,n86,n251);
and (n1729,n1730,n1731);
xor (n1730,n1727,n1728);
or (n1731,n1732,n1735);
and (n1732,n1733,n1734);
xor (n1733,n1638,n1639);
and (n1734,n77,n251);
and (n1735,n1736,n1737);
xor (n1736,n1733,n1734);
or (n1737,n1738,n1741);
and (n1738,n1739,n1740);
xor (n1739,n1643,n1644);
and (n1740,n281,n251);
and (n1741,n1742,n1743);
xor (n1742,n1739,n1740);
or (n1743,n1744,n1747);
and (n1744,n1745,n1746);
xor (n1745,n1648,n1649);
and (n1746,n373,n251);
and (n1747,n1748,n1749);
xor (n1748,n1745,n1746);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
xor (n1751,n1653,n1654);
and (n1752,n436,n251);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
and (n1755,n1756,n1084);
xor (n1756,n1658,n1659);
and (n1757,n1758,n1759);
xor (n1758,n1572,n325);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1664,n1665);
and (n1762,n167,n142);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
or (n1765,n1766,n1768);
and (n1766,n1767,n536);
xor (n1767,n1670,n1671);
and (n1768,n1769,n1770);
xor (n1769,n1767,n536);
or (n1770,n1771,n1773);
and (n1771,n1772,n623);
xor (n1772,n1676,n1677);
and (n1773,n1774,n1775);
xor (n1774,n1772,n623);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1682,n1683);
and (n1778,n27,n142);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1688,n1689);
and (n1784,n190,n142);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1790);
and (n1788,n1789,n1267);
xor (n1789,n1694,n1695);
and (n1790,n1791,n1792);
xor (n1791,n1789,n1267);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1700,n1701);
and (n1795,n96,n142);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1706,n1707);
and (n1801,n133,n142);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1712,n1713);
and (n1807,n73,n142);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1718,n1719);
and (n1813,n56,n142);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1724,n1725);
and (n1819,n86,n142);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
or (n1822,n1823,n1826);
and (n1823,n1824,n1825);
xor (n1824,n1730,n1731);
and (n1825,n77,n142);
and (n1826,n1827,n1828);
xor (n1827,n1824,n1825);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1736,n1737);
and (n1831,n281,n142);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1837);
and (n1835,n1836,n1030);
xor (n1836,n1742,n1743);
and (n1837,n1838,n1839);
xor (n1838,n1836,n1030);
or (n1839,n1840,n1842);
and (n1840,n1841,n1057);
xor (n1841,n1748,n1749);
and (n1842,n1843,n1844);
xor (n1843,n1841,n1057);
and (n1844,n1845,n1846);
xor (n1845,n1754,n1755);
and (n1846,n497,n142);
and (n1847,n172,n143);
and (n1848,n1849,n1850);
xor (n1849,n1570,n1847);
or (n1850,n1851,n1854);
and (n1851,n1852,n1853);
xor (n1852,n1758,n1759);
and (n1853,n167,n143);
and (n1854,n1855,n1856);
xor (n1855,n1852,n1853);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n1764,n1765);
and (n1859,n123,n143);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1769,n1770);
and (n1865,n47,n143);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
or (n1868,n1869,n1872);
and (n1869,n1870,n1871);
xor (n1870,n1774,n1775);
and (n1871,n27,n143);
and (n1872,n1873,n1874);
xor (n1873,n1870,n1871);
or (n1874,n1875,n1878);
and (n1875,n1876,n1877);
xor (n1876,n1780,n1781);
and (n1877,n190,n143);
and (n1878,n1879,n1880);
xor (n1879,n1876,n1877);
or (n1880,n1881,n1884);
and (n1881,n1882,n1883);
xor (n1882,n1786,n1787);
and (n1883,n111,n143);
and (n1884,n1885,n1886);
xor (n1885,n1882,n1883);
or (n1886,n1887,n1890);
and (n1887,n1888,n1889);
xor (n1888,n1791,n1792);
and (n1889,n96,n143);
and (n1890,n1891,n1892);
xor (n1891,n1888,n1889);
or (n1892,n1893,n1896);
and (n1893,n1894,n1895);
xor (n1894,n1797,n1798);
and (n1895,n133,n143);
and (n1896,n1897,n1898);
xor (n1897,n1894,n1895);
or (n1898,n1899,n1902);
and (n1899,n1900,n1901);
xor (n1900,n1803,n1804);
and (n1901,n73,n143);
and (n1902,n1903,n1904);
xor (n1903,n1900,n1901);
or (n1904,n1905,n1908);
and (n1905,n1906,n1907);
xor (n1906,n1809,n1810);
and (n1907,n56,n143);
and (n1908,n1909,n1910);
xor (n1909,n1906,n1907);
or (n1910,n1911,n1914);
and (n1911,n1912,n1913);
xor (n1912,n1815,n1816);
and (n1913,n86,n143);
and (n1914,n1915,n1916);
xor (n1915,n1912,n1913);
or (n1916,n1917,n1920);
and (n1917,n1918,n1919);
xor (n1918,n1821,n1822);
and (n1919,n77,n143);
and (n1920,n1921,n1922);
xor (n1921,n1918,n1919);
or (n1922,n1923,n1926);
and (n1923,n1924,n1925);
xor (n1924,n1827,n1828);
and (n1925,n281,n143);
and (n1926,n1927,n1928);
xor (n1927,n1924,n1925);
or (n1928,n1929,n1932);
and (n1929,n1930,n1931);
xor (n1930,n1833,n1834);
and (n1931,n373,n143);
and (n1932,n1933,n1934);
xor (n1933,n1930,n1931);
or (n1934,n1935,n1938);
and (n1935,n1936,n1937);
xor (n1936,n1838,n1839);
and (n1937,n436,n143);
and (n1938,n1939,n1940);
xor (n1939,n1936,n1937);
and (n1940,n1941,n1014);
xor (n1941,n1843,n1844);
and (n1942,n1943,n1944);
xor (n1943,n1568,n209);
or (n1944,n1945,n1948);
and (n1945,n1946,n1947);
xor (n1946,n1849,n1850);
and (n1947,n167,n149);
and (n1948,n1949,n1950);
xor (n1949,n1946,n1947);
or (n1950,n1951,n1953);
and (n1951,n1952,n368);
xor (n1952,n1855,n1856);
and (n1953,n1954,n1955);
xor (n1954,n1952,n368);
or (n1955,n1956,n1959);
and (n1956,n1957,n1958);
xor (n1957,n1861,n1862);
and (n1958,n47,n149);
and (n1959,n1960,n1961);
xor (n1960,n1957,n1958);
or (n1961,n1962,n1964);
and (n1962,n1963,n550);
xor (n1963,n1867,n1868);
and (n1964,n1965,n1966);
xor (n1965,n1963,n550);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
xor (n1968,n1873,n1874);
and (n1969,n190,n149);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
xor (n1974,n1879,n1880);
and (n1975,n111,n149);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
xor (n1980,n1885,n1886);
and (n1981,n96,n149);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
xor (n1986,n1891,n1892);
and (n1987,n133,n149);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
or (n1990,n1991,n1994);
and (n1991,n1992,n1993);
xor (n1992,n1897,n1898);
and (n1993,n73,n149);
and (n1994,n1995,n1996);
xor (n1995,n1992,n1993);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
xor (n1998,n1903,n1904);
and (n1999,n56,n149);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2006);
and (n2003,n2004,n2005);
xor (n2004,n1909,n1910);
and (n2005,n86,n149);
and (n2006,n2007,n2008);
xor (n2007,n2004,n2005);
or (n2008,n2009,n2012);
and (n2009,n2010,n2011);
xor (n2010,n1915,n1916);
and (n2011,n77,n149);
and (n2012,n2013,n2014);
xor (n2013,n2010,n2011);
or (n2014,n2015,n2018);
and (n2015,n2016,n2017);
xor (n2016,n1921,n1922);
and (n2017,n281,n149);
and (n2018,n2019,n2020);
xor (n2019,n2016,n2017);
or (n2020,n2021,n2024);
and (n2021,n2022,n2023);
xor (n2022,n1927,n1928);
and (n2023,n373,n149);
and (n2024,n2025,n2026);
xor (n2025,n2022,n2023);
or (n2026,n2027,n2030);
and (n2027,n2028,n2029);
xor (n2028,n1933,n1934);
and (n2029,n436,n149);
and (n2030,n2031,n2032);
xor (n2031,n2028,n2029);
and (n2032,n2033,n2034);
xor (n2033,n1939,n1940);
and (n2034,n497,n149);
and (n2035,n172,n157);
or (n2036,n2037,n2040);
and (n2037,n2038,n2039);
xor (n2038,n1943,n1944);
and (n2039,n167,n157);
and (n2040,n2041,n2042);
xor (n2041,n2038,n2039);
or (n2042,n2043,n2046);
and (n2043,n2044,n2045);
xor (n2044,n1949,n1950);
and (n2045,n123,n157);
and (n2046,n2047,n2048);
xor (n2047,n2044,n2045);
or (n2048,n2049,n2052);
and (n2049,n2050,n2051);
xor (n2050,n1954,n1955);
and (n2051,n47,n157);
and (n2052,n2053,n2054);
xor (n2053,n2050,n2051);
or (n2054,n2055,n2058);
and (n2055,n2056,n2057);
xor (n2056,n1960,n1961);
and (n2057,n27,n157);
and (n2058,n2059,n2060);
xor (n2059,n2056,n2057);
or (n2060,n2061,n2064);
and (n2061,n2062,n2063);
xor (n2062,n1965,n1966);
and (n2063,n190,n157);
and (n2064,n2065,n2066);
xor (n2065,n2062,n2063);
or (n2066,n2067,n2070);
and (n2067,n2068,n2069);
xor (n2068,n1971,n1972);
and (n2069,n111,n157);
and (n2070,n2071,n2072);
xor (n2071,n2068,n2069);
or (n2072,n2073,n2076);
and (n2073,n2074,n2075);
xor (n2074,n1977,n1978);
and (n2075,n96,n157);
and (n2076,n2077,n2078);
xor (n2077,n2074,n2075);
or (n2078,n2079,n2082);
and (n2079,n2080,n2081);
xor (n2080,n1983,n1984);
and (n2081,n133,n157);
and (n2082,n2083,n2084);
xor (n2083,n2080,n2081);
or (n2084,n2085,n2088);
and (n2085,n2086,n2087);
xor (n2086,n1989,n1990);
and (n2087,n73,n157);
and (n2088,n2089,n2090);
xor (n2089,n2086,n2087);
or (n2090,n2091,n2094);
and (n2091,n2092,n2093);
xor (n2092,n1995,n1996);
and (n2093,n56,n157);
and (n2094,n2095,n2096);
xor (n2095,n2092,n2093);
or (n2096,n2097,n2100);
and (n2097,n2098,n2099);
xor (n2098,n2001,n2002);
and (n2099,n86,n157);
and (n2100,n2101,n2102);
xor (n2101,n2098,n2099);
or (n2102,n2103,n2106);
and (n2103,n2104,n2105);
xor (n2104,n2007,n2008);
and (n2105,n77,n157);
and (n2106,n2107,n2108);
xor (n2107,n2104,n2105);
or (n2108,n2109,n2112);
and (n2109,n2110,n2111);
xor (n2110,n2013,n2014);
and (n2111,n281,n157);
and (n2112,n2113,n2114);
xor (n2113,n2110,n2111);
or (n2114,n2115,n2118);
and (n2115,n2116,n2117);
xor (n2116,n2019,n2020);
and (n2117,n373,n157);
and (n2118,n2119,n2120);
xor (n2119,n2116,n2117);
or (n2120,n2121,n2124);
and (n2121,n2122,n2123);
xor (n2122,n2025,n2026);
and (n2123,n436,n157);
and (n2124,n2125,n2126);
xor (n2125,n2122,n2123);
and (n2126,n2127,n914);
xor (n2127,n2031,n2032);
or (n2128,n2129,n2131);
and (n2129,n2130,n220);
xor (n2130,n2041,n2042);
and (n2131,n2132,n2133);
xor (n2132,n2130,n220);
or (n2133,n2134,n2136);
and (n2134,n2135,n295);
xor (n2135,n2047,n2048);
and (n2136,n2137,n2138);
xor (n2137,n2135,n295);
or (n2138,n2139,n2141);
and (n2139,n2140,n351);
xor (n2140,n2053,n2054);
and (n2141,n2142,n2143);
xor (n2142,n2140,n351);
or (n2143,n2144,n2146);
and (n2144,n2145,n411);
xor (n2145,n2059,n2060);
and (n2146,n2147,n2148);
xor (n2147,n2145,n411);
or (n2148,n2149,n2152);
and (n2149,n2150,n2151);
xor (n2150,n2065,n2066);
and (n2151,n111,n41);
and (n2152,n2153,n2154);
xor (n2153,n2150,n2151);
or (n2154,n2155,n2158);
and (n2155,n2156,n2157);
xor (n2156,n2071,n2072);
and (n2157,n96,n41);
and (n2158,n2159,n2160);
xor (n2159,n2156,n2157);
or (n2160,n2161,n2163);
and (n2161,n2162,n1160);
xor (n2162,n2077,n2078);
and (n2163,n2164,n2165);
xor (n2164,n2162,n1160);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2083,n2084);
and (n2168,n73,n41);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2089,n2090);
and (n2174,n56,n41);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
or (n2177,n2178,n2181);
and (n2178,n2179,n2180);
xor (n2179,n2095,n2096);
and (n2180,n86,n41);
and (n2181,n2182,n2183);
xor (n2182,n2179,n2180);
or (n2183,n2184,n2187);
and (n2184,n2185,n2186);
xor (n2185,n2101,n2102);
and (n2186,n77,n41);
and (n2187,n2188,n2189);
xor (n2188,n2185,n2186);
or (n2189,n2190,n2192);
and (n2190,n2191,n755);
xor (n2191,n2107,n2108);
and (n2192,n2193,n2194);
xor (n2193,n2191,n755);
or (n2194,n2195,n2197);
and (n2195,n2196,n832);
xor (n2196,n2113,n2114);
and (n2197,n2198,n2199);
xor (n2198,n2196,n832);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2119,n2120);
and (n2202,n436,n41);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
and (n2205,n2206,n2207);
xor (n2206,n2125,n2126);
and (n2207,n497,n41);
and (n2208,n123,n35);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2132,n2133);
and (n2212,n47,n35);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
or (n2215,n2216,n2219);
and (n2216,n2217,n2218);
xor (n2217,n2137,n2138);
and (n2218,n27,n35);
and (n2219,n2220,n2221);
xor (n2220,n2217,n2218);
or (n2221,n2222,n2225);
and (n2222,n2223,n2224);
xor (n2223,n2142,n2143);
and (n2224,n190,n35);
and (n2225,n2226,n2227);
xor (n2226,n2223,n2224);
or (n2227,n2228,n2231);
and (n2228,n2229,n2230);
xor (n2229,n2147,n2148);
and (n2230,n111,n35);
and (n2231,n2232,n2233);
xor (n2232,n2229,n2230);
or (n2233,n2234,n2237);
and (n2234,n2235,n2236);
xor (n2235,n2153,n2154);
and (n2236,n96,n35);
and (n2237,n2238,n2239);
xor (n2238,n2235,n2236);
or (n2239,n2240,n2243);
and (n2240,n2241,n2242);
xor (n2241,n2159,n2160);
and (n2242,n133,n35);
and (n2243,n2244,n2245);
xor (n2244,n2241,n2242);
or (n2245,n2246,n2249);
and (n2246,n2247,n2248);
xor (n2247,n2164,n2165);
and (n2248,n73,n35);
and (n2249,n2250,n2251);
xor (n2250,n2247,n2248);
or (n2251,n2252,n2255);
and (n2252,n2253,n2254);
xor (n2253,n2170,n2171);
and (n2254,n56,n35);
and (n2255,n2256,n2257);
xor (n2256,n2253,n2254);
or (n2257,n2258,n2261);
and (n2258,n2259,n2260);
xor (n2259,n2176,n2177);
and (n2260,n86,n35);
and (n2261,n2262,n2263);
xor (n2262,n2259,n2260);
or (n2263,n2264,n2267);
and (n2264,n2265,n2266);
xor (n2265,n2182,n2183);
and (n2266,n77,n35);
and (n2267,n2268,n2269);
xor (n2268,n2265,n2266);
or (n2269,n2270,n2273);
and (n2270,n2271,n2272);
xor (n2271,n2188,n2189);
and (n2272,n281,n35);
and (n2273,n2274,n2275);
xor (n2274,n2271,n2272);
or (n2275,n2276,n2279);
and (n2276,n2277,n2278);
xor (n2277,n2193,n2194);
and (n2278,n373,n35);
and (n2279,n2280,n2281);
xor (n2280,n2277,n2278);
or (n2281,n2282,n2285);
and (n2282,n2283,n2284);
xor (n2283,n2198,n2199);
and (n2284,n436,n35);
and (n2285,n2286,n2287);
xor (n2286,n2283,n2284);
and (n2287,n2288,n818);
xor (n2288,n2204,n2205);
or (n2289,n2290,n2292);
and (n2290,n2291,n30);
xor (n2291,n2214,n2215);
and (n2292,n2293,n2294);
xor (n2293,n2291,n30);
or (n2294,n2295,n2298);
and (n2295,n2296,n2297);
xor (n2296,n2220,n2221);
and (n2297,n190,n29);
and (n2298,n2299,n2300);
xor (n2299,n2296,n2297);
or (n2300,n2301,n2303);
and (n2301,n2302,n380);
xor (n2302,n2226,n2227);
and (n2303,n2304,n2305);
xor (n2304,n2302,n380);
or (n2305,n2306,n2308);
and (n2306,n2307,n455);
xor (n2307,n2232,n2233);
and (n2308,n2309,n2310);
xor (n2309,n2307,n455);
or (n2310,n2311,n2314);
and (n2311,n2312,n2313);
xor (n2312,n2238,n2239);
and (n2313,n133,n29);
and (n2314,n2315,n2316);
xor (n2315,n2312,n2313);
or (n2316,n2317,n2320);
and (n2317,n2318,n2319);
xor (n2318,n2244,n2245);
and (n2319,n73,n29);
and (n2320,n2321,n2322);
xor (n2321,n2318,n2319);
or (n2322,n2323,n2325);
and (n2323,n2324,n1169);
xor (n2324,n2250,n2251);
and (n2325,n2326,n2327);
xor (n2326,n2324,n1169);
or (n2327,n2328,n2331);
and (n2328,n2329,n2330);
xor (n2329,n2256,n2257);
and (n2330,n86,n29);
and (n2331,n2332,n2333);
xor (n2332,n2329,n2330);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2262,n2263);
and (n2336,n77,n29);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
or (n2339,n2340,n2343);
and (n2340,n2341,n2342);
xor (n2341,n2268,n2269);
and (n2342,n281,n29);
and (n2343,n2344,n2345);
xor (n2344,n2341,n2342);
or (n2345,n2346,n2349);
and (n2346,n2347,n2348);
xor (n2347,n2274,n2275);
and (n2348,n373,n29);
and (n2349,n2350,n2351);
xor (n2350,n2347,n2348);
or (n2351,n2352,n2355);
and (n2352,n2353,n2354);
xor (n2353,n2280,n2281);
and (n2354,n436,n29);
and (n2355,n2356,n2357);
xor (n2356,n2353,n2354);
and (n2357,n2358,n2359);
xor (n2358,n2286,n2287);
and (n2359,n497,n29);
and (n2360,n27,n182);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2293,n2294);
and (n2364,n190,n182);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2299,n2300);
and (n2370,n111,n182);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2304,n2305);
and (n2376,n96,n182);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2309,n2310);
and (n2382,n133,n182);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2315,n2316);
and (n2388,n73,n182);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2321,n2322);
and (n2394,n56,n182);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2326,n2327);
and (n2400,n86,n182);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
or (n2403,n2404,n2407);
and (n2404,n2405,n2406);
xor (n2405,n2332,n2333);
and (n2406,n77,n182);
and (n2407,n2408,n2409);
xor (n2408,n2405,n2406);
or (n2409,n2410,n2413);
and (n2410,n2411,n2412);
xor (n2411,n2338,n2339);
and (n2412,n281,n182);
and (n2413,n2414,n2415);
xor (n2414,n2411,n2412);
or (n2415,n2416,n2419);
and (n2416,n2417,n2418);
xor (n2417,n2344,n2345);
and (n2418,n373,n182);
and (n2419,n2420,n2421);
xor (n2420,n2417,n2418);
or (n2421,n2422,n2425);
and (n2422,n2423,n2424);
xor (n2423,n2350,n2351);
and (n2424,n436,n182);
and (n2425,n2426,n2427);
xor (n2426,n2423,n2424);
and (n2427,n2428,n725);
xor (n2428,n2356,n2357);
and (n2429,n190,n103);
or (n2430,n2431,n2433);
and (n2431,n2432,n228);
xor (n2432,n2366,n2367);
and (n2433,n2434,n2435);
xor (n2434,n2432,n228);
or (n2435,n2436,n2438);
and (n2436,n2437,n288);
xor (n2437,n2372,n2373);
and (n2438,n2439,n2440);
xor (n2439,n2437,n288);
or (n2440,n2441,n2444);
and (n2441,n2442,n2443);
xor (n2442,n2378,n2379);
and (n2443,n133,n103);
and (n2444,n2445,n2446);
xor (n2445,n2442,n2443);
or (n2446,n2447,n2450);
and (n2447,n2448,n2449);
xor (n2448,n2384,n2385);
and (n2449,n73,n103);
and (n2450,n2451,n2452);
xor (n2451,n2448,n2449);
or (n2452,n2453,n2455);
and (n2453,n2454,n570);
xor (n2454,n2390,n2391);
and (n2455,n2456,n2457);
xor (n2456,n2454,n570);
or (n2457,n2458,n2461);
and (n2458,n2459,n2460);
xor (n2459,n2396,n2397);
and (n2460,n86,n103);
and (n2461,n2462,n2463);
xor (n2462,n2459,n2460);
or (n2463,n2464,n2467);
and (n2464,n2465,n2466);
xor (n2465,n2402,n2403);
and (n2466,n77,n103);
and (n2467,n2468,n2469);
xor (n2468,n2465,n2466);
or (n2469,n2470,n2473);
and (n2470,n2471,n2472);
xor (n2471,n2408,n2409);
and (n2472,n281,n103);
and (n2473,n2474,n2475);
xor (n2474,n2471,n2472);
or (n2475,n2476,n2479);
and (n2476,n2477,n2478);
xor (n2477,n2414,n2415);
and (n2478,n373,n103);
and (n2479,n2480,n2481);
xor (n2480,n2477,n2478);
or (n2481,n2482,n2485);
and (n2482,n2483,n2484);
xor (n2483,n2420,n2421);
and (n2484,n436,n103);
and (n2485,n2486,n2487);
xor (n2486,n2483,n2484);
and (n2487,n2488,n2489);
xor (n2488,n2426,n2427);
and (n2489,n497,n103);
and (n2490,n111,n102);
or (n2491,n2492,n2495);
and (n2492,n2493,n2494);
xor (n2493,n2434,n2435);
and (n2494,n96,n102);
and (n2495,n2496,n2497);
xor (n2496,n2493,n2494);
or (n2497,n2498,n2501);
and (n2498,n2499,n2500);
xor (n2499,n2439,n2440);
and (n2500,n133,n102);
and (n2501,n2502,n2503);
xor (n2502,n2499,n2500);
or (n2503,n2504,n2507);
and (n2504,n2505,n2506);
xor (n2505,n2445,n2446);
and (n2506,n73,n102);
and (n2507,n2508,n2509);
xor (n2508,n2505,n2506);
or (n2509,n2510,n2513);
and (n2510,n2511,n2512);
xor (n2511,n2451,n2452);
and (n2512,n56,n102);
and (n2513,n2514,n2515);
xor (n2514,n2511,n2512);
or (n2515,n2516,n2519);
and (n2516,n2517,n2518);
xor (n2517,n2456,n2457);
and (n2518,n86,n102);
and (n2519,n2520,n2521);
xor (n2520,n2517,n2518);
or (n2521,n2522,n2525);
and (n2522,n2523,n2524);
xor (n2523,n2462,n2463);
and (n2524,n77,n102);
and (n2525,n2526,n2527);
xor (n2526,n2523,n2524);
or (n2527,n2528,n2531);
and (n2528,n2529,n2530);
xor (n2529,n2468,n2469);
and (n2530,n281,n102);
and (n2531,n2532,n2533);
xor (n2532,n2529,n2530);
or (n2533,n2534,n2537);
and (n2534,n2535,n2536);
xor (n2535,n2474,n2475);
and (n2536,n373,n102);
and (n2537,n2538,n2539);
xor (n2538,n2535,n2536);
or (n2539,n2540,n2543);
and (n2540,n2541,n2542);
xor (n2541,n2480,n2481);
and (n2542,n436,n102);
and (n2543,n2544,n2545);
xor (n2544,n2541,n2542);
and (n2545,n2546,n2547);
xor (n2546,n2486,n2487);
not (n2547,n1241);
and (n2548,n96,n64);
or (n2549,n2550,n2553);
and (n2550,n2551,n2552);
xor (n2551,n2496,n2497);
and (n2552,n133,n64);
and (n2553,n2554,n2555);
xor (n2554,n2551,n2552);
or (n2555,n2556,n2559);
and (n2556,n2557,n2558);
xor (n2557,n2502,n2503);
and (n2558,n73,n64);
and (n2559,n2560,n2561);
xor (n2560,n2557,n2558);
or (n2561,n2562,n2565);
and (n2562,n2563,n2564);
xor (n2563,n2508,n2509);
and (n2564,n56,n64);
and (n2565,n2566,n2567);
xor (n2566,n2563,n2564);
or (n2567,n2568,n2571);
and (n2568,n2569,n2570);
xor (n2569,n2514,n2515);
and (n2570,n86,n64);
and (n2571,n2572,n2573);
xor (n2572,n2569,n2570);
or (n2573,n2574,n2577);
and (n2574,n2575,n2576);
xor (n2575,n2520,n2521);
and (n2576,n77,n64);
and (n2577,n2578,n2579);
xor (n2578,n2575,n2576);
or (n2579,n2580,n2583);
and (n2580,n2581,n2582);
xor (n2581,n2526,n2527);
and (n2582,n281,n64);
and (n2583,n2584,n2585);
xor (n2584,n2581,n2582);
or (n2585,n2586,n2589);
and (n2586,n2587,n2588);
xor (n2587,n2532,n2533);
and (n2588,n373,n64);
and (n2589,n2590,n2591);
xor (n2590,n2587,n2588);
or (n2591,n2592,n2595);
and (n2592,n2593,n2594);
xor (n2593,n2538,n2539);
and (n2594,n436,n64);
and (n2595,n2596,n2597);
xor (n2596,n2593,n2594);
and (n2597,n2598,n2599);
xor (n2598,n2544,n2545);
and (n2599,n497,n64);
and (n2600,n133,n65);
or (n2601,n2602,n2605);
and (n2602,n2603,n2604);
xor (n2603,n2554,n2555);
and (n2604,n73,n65);
and (n2605,n2606,n2607);
xor (n2606,n2603,n2604);
or (n2607,n2608,n2611);
and (n2608,n2609,n2610);
xor (n2609,n2560,n2561);
and (n2610,n56,n65);
and (n2611,n2612,n2613);
xor (n2612,n2609,n2610);
or (n2613,n2614,n2617);
and (n2614,n2615,n2616);
xor (n2615,n2566,n2567);
and (n2616,n86,n65);
and (n2617,n2618,n2619);
xor (n2618,n2615,n2616);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
xor (n2621,n2572,n2573);
and (n2622,n77,n65);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
xor (n2627,n2578,n2579);
and (n2628,n281,n65);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
xor (n2633,n2584,n2585);
and (n2634,n373,n65);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
xor (n2639,n2590,n2591);
and (n2640,n436,n65);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
and (n2643,n2644,n2645);
xor (n2644,n2596,n2597);
not (n2645,n1311);
and (n2646,n73,n54);
or (n2647,n2648,n2651);
and (n2648,n2649,n2650);
xor (n2649,n2606,n2607);
and (n2650,n56,n54);
and (n2651,n2652,n2653);
xor (n2652,n2649,n2650);
or (n2653,n2654,n2656);
and (n2654,n2655,n318);
xor (n2655,n2612,n2613);
and (n2656,n2657,n2658);
xor (n2657,n2655,n318);
or (n2658,n2659,n2661);
and (n2659,n2660,n403);
xor (n2660,n2618,n2619);
and (n2661,n2662,n2663);
xor (n2662,n2660,n403);
or (n2663,n2664,n2666);
and (n2664,n2665,n431);
xor (n2665,n2624,n2625);
and (n2666,n2667,n2668);
xor (n2667,n2665,n431);
or (n2668,n2669,n2672);
and (n2669,n2670,n2671);
xor (n2670,n2630,n2631);
and (n2671,n373,n54);
and (n2672,n2673,n2674);
xor (n2673,n2670,n2671);
or (n2674,n2675,n2678);
and (n2675,n2676,n2677);
xor (n2676,n2636,n2637);
and (n2677,n436,n54);
and (n2678,n2679,n2680);
xor (n2679,n2676,n2677);
and (n2680,n2681,n2682);
xor (n2681,n2642,n2643);
and (n2682,n497,n54);
and (n2683,n56,n81);
or (n2684,n2685,n2688);
and (n2685,n2686,n2687);
xor (n2686,n2652,n2653);
and (n2687,n86,n81);
and (n2688,n2689,n2690);
xor (n2689,n2686,n2687);
or (n2690,n2691,n2694);
and (n2691,n2692,n2693);
xor (n2692,n2657,n2658);
and (n2693,n77,n81);
and (n2694,n2695,n2696);
xor (n2695,n2692,n2693);
or (n2696,n2697,n2700);
and (n2697,n2698,n2699);
xor (n2698,n2662,n2663);
and (n2699,n281,n81);
and (n2700,n2701,n2702);
xor (n2701,n2698,n2699);
or (n2702,n2703,n2706);
and (n2703,n2704,n2705);
xor (n2704,n2667,n2668);
and (n2705,n373,n81);
and (n2706,n2707,n2708);
xor (n2707,n2704,n2705);
or (n2708,n2709,n2712);
and (n2709,n2710,n2711);
xor (n2710,n2673,n2674);
and (n2711,n436,n81);
and (n2712,n2713,n2714);
xor (n2713,n2710,n2711);
and (n2714,n2715,n2716);
xor (n2715,n2679,n2680);
and (n2716,n497,n81);
endmodule
