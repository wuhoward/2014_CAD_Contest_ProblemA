module top (out,n21,n22,n25,n29,n31,n35,n42,n50,n52
        ,n57,n64,n71,n84,n90,n92,n103,n110,n112,n119
        ,n125,n139,n140,n149,n154,n165,n174,n183,n188,n192
        ,n209,n214,n221,n250,n285,n286,n294,n295,n306,n314
        ,n322,n329,n340,n350,n363,n458,n465);
output out;
input n21;
input n22;
input n25;
input n29;
input n31;
input n35;
input n42;
input n50;
input n52;
input n57;
input n64;
input n71;
input n84;
input n90;
input n92;
input n103;
input n110;
input n112;
input n119;
input n125;
input n139;
input n140;
input n149;
input n154;
input n165;
input n174;
input n183;
input n188;
input n192;
input n209;
input n214;
input n221;
input n250;
input n285;
input n286;
input n294;
input n295;
input n306;
input n314;
input n322;
input n329;
input n340;
input n350;
input n363;
input n458;
input n465;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
xor (out,n0,n1749);
nand (n0,n1,n1748);
or (n1,n2,n700);
not (n2,n3);
nor (n3,n4,n699);
not (n4,n5);
nand (n5,n6,n609);
xor (n6,n7,n596);
xor (n7,n8,n380);
xor (n8,n9,n269);
xor (n9,n10,n200);
or (n10,n11,n199);
and (n11,n12,n158);
xor (n12,n13,n75);
or (n13,n14,n74);
and (n14,n15,n44);
xor (n15,n16,n26);
and (n16,n17,n25);
not (n17,n18);
and (n18,n19,n23);
nand (n19,n20,n22);
not (n20,n21);
nand (n23,n24,n21);
not (n24,n22);
nand (n26,n27,n38);
or (n27,n28,n32);
nand (n28,n29,n30);
not (n30,n31);
nor (n32,n33,n36);
and (n33,n34,n35);
not (n34,n29);
and (n36,n29,n37);
not (n37,n35);
or (n38,n39,n30);
nor (n39,n40,n43);
and (n40,n41,n29);
not (n41,n42);
and (n43,n42,n34);
nand (n44,n45,n66);
or (n45,n46,n60);
not (n46,n47);
nor (n47,n48,n54);
nand (n48,n49,n53);
or (n49,n50,n51);
not (n51,n52);
nand (n53,n50,n51);
nor (n54,n55,n58);
and (n55,n50,n56);
not (n56,n57);
and (n58,n57,n59);
not (n59,n50);
not (n60,n61);
nor (n61,n62,n65);
and (n62,n63,n56);
not (n63,n64);
and (n65,n64,n57);
or (n66,n67,n68);
not (n67,n48);
not (n68,n69);
nor (n69,n70,n72);
and (n70,n71,n57);
and (n72,n73,n56);
not (n73,n71);
and (n74,n16,n26);
or (n75,n76,n157);
and (n76,n77,n133);
xor (n77,n78,n105);
nand (n78,n79,n98);
or (n79,n80,n86);
not (n80,n81);
nand (n81,n82,n85);
or (n82,n22,n83);
not (n83,n84);
or (n85,n24,n84);
not (n86,n87);
nor (n87,n88,n94);
nand (n88,n89,n93);
or (n89,n90,n91);
not (n91,n92);
nand (n93,n90,n91);
nor (n94,n95,n96);
and (n95,n24,n90);
and (n96,n22,n97);
not (n97,n90);
or (n98,n99,n100);
not (n99,n88);
nor (n100,n101,n104);
and (n101,n102,n22);
not (n102,n103);
and (n104,n103,n24);
nand (n105,n106,n121);
or (n106,n107,n115);
not (n107,n108);
nand (n108,n109,n113);
or (n109,n110,n111);
not (n111,n112);
or (n113,n114,n112);
not (n114,n110);
not (n115,n116);
nand (n116,n117,n120);
or (n117,n57,n118);
not (n118,n119);
nand (n120,n57,n118);
nand (n121,n122,n128);
not (n122,n123);
nor (n123,n124,n126);
and (n124,n114,n125);
and (n126,n110,n127);
not (n127,n125);
not (n128,n129);
nand (n129,n115,n130);
nand (n130,n131,n132);
or (n131,n110,n118);
nand (n132,n110,n118);
nand (n133,n134,n151);
or (n134,n135,n146);
nand (n135,n136,n143);
nor (n136,n137,n141);
and (n137,n138,n140);
not (n138,n139);
and (n141,n142,n139);
not (n142,n140);
nand (n143,n144,n145);
or (n144,n139,n51);
nand (n145,n139,n51);
nor (n146,n147,n150);
and (n147,n148,n52);
not (n148,n149);
and (n150,n149,n51);
or (n151,n136,n152);
nor (n152,n153,n155);
and (n153,n51,n154);
and (n155,n52,n156);
not (n156,n154);
and (n157,n78,n105);
xor (n158,n159,n177);
xor (n159,n160,n168);
nand (n160,n161,n162);
or (n161,n28,n39);
or (n162,n163,n30);
nor (n163,n164,n166);
and (n164,n34,n165);
and (n166,n29,n167);
not (n167,n165);
nand (n168,n169,n170);
or (n169,n135,n152);
nand (n170,n171,n172);
not (n171,n136);
nor (n172,n173,n175);
and (n173,n174,n52);
and (n175,n176,n51);
not (n176,n174);
nand (n177,n178,n195);
or (n178,n179,n190);
nand (n179,n180,n185);
nor (n180,n181,n184);
and (n181,n110,n182);
not (n182,n183);
and (n184,n114,n183);
nand (n185,n186,n189);
or (n186,n183,n187);
not (n187,n188);
nand (n189,n187,n183);
nor (n190,n191,n193);
and (n191,n187,n192);
and (n193,n188,n194);
not (n194,n192);
or (n195,n180,n196);
nor (n196,n197,n198);
and (n197,n187,n125);
and (n198,n188,n127);
and (n199,n13,n75);
xor (n200,n201,n234);
xor (n201,n202,n231);
and (n202,n203,n210);
and (n203,n204,n209);
nand (n204,n205,n206);
or (n205,n25,n21);
nand (n206,n207,n24);
not (n207,n208);
and (n208,n25,n21);
nand (n210,n211,n227);
or (n211,n212,n217);
nor (n212,n213,n215);
and (n213,n142,n214);
and (n215,n140,n216);
not (n216,n214);
not (n217,n218);
nor (n218,n219,n223);
nand (n219,n220,n222);
or (n220,n221,n34);
nand (n222,n34,n221);
nor (n223,n224,n225);
and (n224,n142,n221);
and (n225,n140,n226);
not (n226,n221);
nand (n227,n219,n228);
nor (n228,n229,n230);
and (n229,n35,n140);
and (n230,n37,n142);
or (n231,n232,n233);
and (n232,n159,n177);
and (n233,n160,n168);
or (n234,n235,n268);
and (n235,n236,n252);
xor (n236,n237,n244);
nand (n237,n238,n239);
or (n238,n107,n129);
nand (n239,n240,n116);
not (n240,n241);
nor (n241,n242,n243);
and (n242,n63,n110);
and (n243,n64,n114);
nand (n244,n245,n246);
or (n245,n86,n100);
nand (n246,n88,n247);
nor (n247,n248,n251);
and (n248,n249,n24);
not (n249,n250);
and (n251,n250,n22);
nand (n252,n253,n264);
or (n253,n254,n260);
not (n254,n255);
nor (n255,n17,n256);
nor (n256,n257,n258);
and (n257,n20,n209);
and (n258,n21,n259);
not (n259,n209);
nor (n260,n261,n263);
and (n261,n262,n209);
not (n262,n25);
and (n263,n259,n25);
or (n264,n18,n265);
nor (n265,n266,n267);
and (n266,n259,n84);
and (n267,n209,n83);
and (n268,n237,n244);
or (n269,n270,n379);
and (n270,n271,n333);
xor (n271,n272,n332);
xor (n272,n273,n308);
xor (n273,n274,n280);
nand (n274,n275,n276);
or (n275,n68,n46);
nand (n276,n48,n277);
nor (n277,n278,n279);
and (n278,n149,n57);
and (n279,n148,n56);
nand (n280,n281,n302);
or (n281,n282,n289);
nor (n282,n283,n287);
and (n283,n284,n286);
not (n284,n285);
and (n287,n285,n288);
not (n288,n286);
nand (n289,n290,n297);
not (n290,n291);
nand (n291,n292,n296);
or (n292,n293,n295);
not (n293,n294);
nand (n296,n293,n295);
not (n297,n298);
nor (n298,n299,n301);
and (n299,n300,n286);
not (n300,n295);
and (n301,n295,n288);
nand (n302,n291,n303);
nand (n303,n304,n307);
or (n304,n286,n305);
not (n305,n306);
or (n307,n288,n306);
nand (n308,n309,n325);
or (n309,n310,n320);
not (n310,n311);
nor (n311,n312,n317);
nor (n312,n313,n315);
and (n313,n91,n314);
and (n315,n92,n316);
not (n316,n314);
nor (n317,n318,n319);
and (n318,n314,n286);
and (n319,n316,n288);
nor (n320,n321,n323);
and (n321,n91,n322);
and (n323,n92,n324);
not (n324,n322);
or (n325,n326,n327);
not (n326,n317);
nor (n327,n328,n330);
and (n328,n91,n329);
and (n330,n92,n331);
not (n331,n329);
xor (n332,n236,n252);
or (n333,n334,n378);
and (n334,n335,n366);
xor (n335,n336,n344);
nand (n336,n337,n343);
or (n337,n179,n338);
nor (n338,n339,n341);
and (n339,n187,n340);
and (n341,n188,n342);
not (n342,n340);
or (n343,n180,n190);
nand (n344,n345,n359);
or (n345,n346,n356);
not (n346,n347);
nor (n347,n348,n352);
nand (n348,n349,n351);
or (n349,n350,n187);
nand (n351,n350,n187);
nor (n352,n353,n354);
and (n353,n293,n350);
and (n354,n294,n355);
not (n355,n350);
nor (n356,n357,n358);
and (n357,n306,n293);
and (n358,n294,n305);
or (n359,n360,n361);
not (n360,n348);
nor (n361,n362,n364);
and (n362,n293,n363);
and (n364,n294,n365);
not (n365,n363);
and (n366,n367,n372);
nor (n367,n368,n24);
nor (n368,n369,n371);
and (n369,n370,n91);
nand (n370,n25,n90);
and (n371,n262,n97);
nand (n372,n373,n377);
or (n373,n28,n374);
nor (n374,n375,n376);
and (n375,n34,n214);
and (n376,n29,n216);
or (n377,n32,n30);
and (n378,n336,n344);
and (n379,n272,n332);
xor (n380,n381,n515);
xor (n381,n382,n433);
xor (n382,n383,n411);
xor (n383,n384,n387);
or (n384,n385,n386);
and (n385,n273,n308);
and (n386,n274,n280);
xor (n387,n388,n402);
xor (n388,n389,n396);
nand (n389,n390,n392);
or (n390,n391,n135);
not (n391,n172);
nand (n392,n171,n393);
nor (n393,n394,n395);
and (n394,n214,n52);
and (n395,n216,n51);
nand (n396,n397,n398);
or (n397,n179,n196);
or (n398,n399,n180);
nor (n399,n400,n401);
and (n400,n187,n112);
and (n401,n188,n111);
nand (n402,n403,n407);
or (n403,n346,n404);
nor (n404,n405,n406);
and (n405,n293,n340);
and (n406,n294,n342);
or (n407,n360,n408);
nor (n408,n409,n410);
and (n409,n293,n192);
and (n410,n294,n194);
xor (n411,n412,n426);
xor (n412,n413,n420);
nand (n413,n414,n416);
or (n414,n415,n289);
not (n415,n303);
nand (n416,n417,n291);
nor (n417,n418,n419);
and (n418,n363,n286);
and (n419,n365,n288);
nand (n420,n421,n422);
or (n421,n310,n327);
or (n422,n326,n423);
nor (n423,n424,n425);
and (n424,n91,n285);
and (n425,n92,n284);
nand (n426,n427,n428);
or (n427,n129,n241);
or (n428,n115,n429);
not (n429,n430);
nand (n430,n431,n432);
or (n431,n110,n73);
or (n432,n114,n71);
xor (n433,n434,n483);
xor (n434,n435,n460);
xor (n435,n436,n452);
xor (n436,n437,n444);
nand (n437,n438,n440);
or (n438,n439,n86);
not (n439,n247);
nand (n440,n441,n88);
nor (n441,n442,n443);
and (n442,n324,n24);
and (n443,n322,n22);
nand (n444,n445,n450);
or (n445,n446,n18);
not (n446,n447);
nand (n447,n448,n449);
or (n448,n209,n102);
or (n449,n259,n103);
nand (n450,n451,n255);
not (n451,n265);
nand (n452,n453,n454);
or (n453,n28,n163);
or (n454,n455,n30);
nor (n455,n456,n459);
and (n456,n457,n29);
not (n457,n458);
and (n459,n458,n34);
xor (n460,n461,n476);
xor (n461,n462,n468);
nor (n462,n463,n262);
nor (n463,n464,n466);
and (n464,n259,n465);
and (n466,n209,n467);
not (n467,n465);
nand (n468,n469,n471);
or (n469,n470,n217);
not (n470,n228);
nand (n471,n472,n219);
not (n472,n473);
nor (n473,n474,n475);
and (n474,n41,n140);
and (n475,n42,n142);
nand (n476,n477,n479);
or (n477,n478,n46);
not (n478,n277);
nand (n479,n48,n480);
nand (n480,n481,n482);
or (n481,n57,n156);
or (n482,n56,n154);
or (n483,n484,n514);
and (n484,n485,n490);
xor (n485,n486,n489);
nand (n486,n487,n488);
or (n487,n346,n361);
or (n488,n360,n404);
xor (n489,n203,n210);
or (n490,n491,n513);
and (n491,n492,n506);
xor (n492,n493,n500);
nand (n493,n494,n499);
or (n494,n495,n289);
not (n495,n496);
nor (n496,n497,n498);
and (n497,n331,n288);
and (n498,n329,n286);
or (n499,n290,n282);
nand (n500,n501,n505);
or (n501,n310,n502);
nor (n502,n503,n504);
and (n503,n91,n250);
and (n504,n92,n249);
or (n505,n326,n320);
nand (n506,n507,n511);
or (n507,n217,n508);
nor (n508,n509,n510);
and (n509,n142,n174);
and (n510,n140,n176);
or (n511,n512,n212);
not (n512,n219);
and (n513,n493,n500);
and (n514,n486,n489);
or (n515,n516,n595);
and (n516,n517,n594);
xor (n517,n518,n593);
or (n518,n519,n592);
and (n519,n520,n568);
xor (n520,n521,n544);
or (n521,n522,n543);
and (n522,n523,n537);
xor (n523,n524,n531);
nand (n524,n525,n530);
or (n525,n526,n46);
not (n526,n527);
nor (n527,n528,n529);
and (n528,n112,n57);
and (n529,n111,n56);
nand (n530,n61,n48);
nand (n531,n532,n536);
or (n532,n533,n289);
nor (n533,n534,n535);
and (n534,n322,n288);
and (n535,n324,n286);
nand (n536,n496,n291);
nand (n537,n538,n542);
or (n538,n310,n539);
nor (n539,n540,n541);
and (n540,n91,n103);
and (n541,n92,n102);
or (n542,n502,n326);
and (n543,n524,n531);
or (n544,n545,n567);
and (n545,n546,n561);
xor (n546,n547,n555);
nand (n547,n548,n553);
or (n548,n549,n135);
not (n549,n550);
nand (n550,n551,n552);
or (n551,n52,n73);
or (n552,n51,n71);
nand (n553,n554,n171);
not (n554,n146);
nand (n555,n556,n560);
or (n556,n179,n557);
nor (n557,n558,n559);
and (n558,n363,n187);
and (n559,n188,n365);
or (n560,n338,n180);
nand (n561,n562,n566);
or (n562,n346,n563);
nor (n563,n564,n565);
and (n564,n285,n293);
and (n565,n294,n284);
or (n566,n360,n356);
and (n567,n547,n555);
or (n568,n569,n591);
and (n569,n570,n584);
xor (n570,n571,n578);
nand (n571,n572,n576);
or (n572,n573,n217);
nor (n573,n574,n575);
and (n574,n154,n142);
and (n575,n156,n140);
nand (n576,n577,n219);
not (n577,n508);
nand (n578,n579,n580);
or (n579,n80,n99);
or (n580,n86,n581);
nor (n581,n582,n583);
and (n582,n22,n262);
and (n583,n24,n25);
nand (n584,n585,n590);
or (n585,n129,n586);
not (n586,n587);
nor (n587,n588,n589);
and (n588,n194,n114);
and (n589,n192,n110);
or (n590,n115,n123);
and (n591,n571,n578);
and (n592,n521,n544);
xor (n593,n485,n490);
xor (n594,n12,n158);
and (n595,n518,n593);
or (n596,n597,n608);
and (n597,n598,n607);
xor (n598,n599,n606);
or (n599,n600,n605);
and (n600,n601,n604);
xor (n601,n602,n603);
xor (n602,n15,n44);
xor (n603,n492,n506);
xor (n604,n77,n133);
and (n605,n602,n603);
xor (n606,n271,n333);
xor (n607,n517,n594);
and (n608,n599,n606);
or (n609,n610,n698);
and (n610,n611,n691);
xor (n611,n612,n690);
or (n612,n613,n689);
and (n613,n614,n660);
xor (n614,n615,n616);
xor (n615,n335,n366);
or (n616,n617,n659);
and (n617,n618,n637);
xor (n618,n619,n620);
xor (n619,n367,n372);
or (n620,n621,n636);
and (n621,n622,n630);
xor (n622,n623,n624);
and (n623,n88,n25);
nand (n624,n625,n629);
or (n625,n28,n626);
nor (n626,n627,n628);
and (n627,n34,n174);
and (n628,n29,n176);
or (n629,n374,n30);
nand (n630,n631,n635);
or (n631,n46,n632);
nor (n632,n633,n634);
and (n633,n56,n125);
and (n634,n57,n127);
or (n635,n67,n526);
and (n636,n623,n624);
or (n637,n638,n658);
and (n638,n639,n652);
xor (n639,n640,n646);
nand (n640,n641,n645);
or (n641,n289,n642);
nor (n642,n643,n644);
and (n643,n288,n250);
and (n644,n286,n249);
or (n645,n290,n533);
nand (n646,n647,n651);
or (n647,n310,n648);
nor (n648,n649,n650);
and (n649,n91,n84);
and (n650,n92,n83);
or (n651,n326,n539);
nand (n652,n653,n657);
or (n653,n217,n654);
nor (n654,n655,n656);
and (n655,n142,n149);
and (n656,n140,n148);
or (n657,n512,n573);
and (n658,n640,n646);
and (n659,n619,n620);
or (n660,n661,n688);
and (n661,n662,n687);
xor (n662,n663,n686);
or (n663,n664,n685);
and (n664,n665,n679);
xor (n665,n666,n673);
nand (n666,n667,n672);
or (n667,n668,n129);
not (n668,n669);
nand (n669,n670,n671);
or (n670,n110,n342);
or (n671,n114,n340);
nand (n672,n116,n587);
nand (n673,n674,n678);
or (n674,n675,n135);
nor (n675,n676,n677);
and (n676,n51,n64);
and (n677,n52,n63);
nand (n678,n171,n550);
nand (n679,n680,n684);
or (n680,n179,n681);
nor (n681,n682,n683);
and (n682,n187,n306);
and (n683,n188,n305);
or (n684,n180,n557);
and (n685,n666,n673);
xor (n686,n546,n561);
xor (n687,n523,n537);
and (n688,n663,n686);
and (n689,n615,n616);
xor (n690,n598,n607);
or (n691,n692,n697);
and (n692,n693,n696);
xor (n693,n694,n695);
xor (n694,n520,n568);
xor (n695,n601,n604);
xor (n696,n614,n660);
and (n697,n694,n695);
and (n698,n612,n690);
nor (n699,n6,n609);
not (n700,n701);
and (n701,n702,n1743);
nand (n702,n703,n1724);
nand (n703,n704,n1710);
or (n704,n705,n1480);
not (n705,n706);
nand (n706,n707,n1470,n1479);
nand (n707,n708,n1162,n1379);
or (n708,n709,n1161);
and (n709,n710,n903);
xor (n710,n711,n834);
or (n711,n712,n833);
and (n712,n713,n794);
xor (n713,n714,n743);
xor (n714,n715,n734);
xor (n715,n716,n725);
nand (n716,n717,n721);
or (n717,n129,n718);
nor (n718,n719,n720);
and (n719,n114,n84);
and (n720,n110,n83);
or (n721,n115,n722);
nor (n722,n723,n724);
and (n723,n114,n103);
and (n724,n110,n102);
nand (n725,n726,n730);
or (n726,n727,n28);
nor (n727,n728,n729);
and (n728,n34,n340);
and (n729,n29,n342);
or (n730,n731,n30);
nor (n731,n732,n733);
and (n732,n34,n192);
and (n733,n29,n194);
nand (n734,n735,n739);
or (n735,n135,n736);
nor (n736,n737,n738);
and (n737,n51,n329);
and (n738,n52,n331);
or (n739,n136,n740);
nor (n740,n741,n742);
and (n741,n51,n285);
and (n742,n52,n284);
or (n743,n744,n793);
and (n744,n745,n768);
xor (n745,n746,n752);
nand (n746,n747,n751);
or (n747,n135,n748);
nor (n748,n749,n750);
and (n749,n51,n322);
and (n750,n52,n324);
or (n751,n136,n736);
xor (n752,n753,n759);
and (n753,n754,n110);
nand (n754,n755,n756);
or (n755,n25,n119);
nand (n756,n757,n56);
not (n757,n758);
and (n758,n25,n119);
nand (n759,n760,n764);
or (n760,n217,n761);
nor (n761,n762,n763);
and (n762,n142,n285);
and (n763,n140,n284);
or (n764,n512,n765);
nor (n765,n766,n767);
and (n766,n142,n306);
and (n767,n140,n305);
or (n768,n769,n792);
and (n769,n770,n781);
xor (n770,n771,n772);
and (n771,n116,n25);
nand (n772,n773,n777);
or (n773,n28,n774);
nor (n774,n775,n776);
and (n775,n34,n306);
and (n776,n29,n305);
or (n777,n778,n30);
nor (n778,n779,n780);
and (n779,n34,n363);
and (n780,n29,n365);
nand (n781,n782,n787);
or (n782,n783,n46);
not (n783,n784);
nor (n784,n785,n786);
and (n785,n84,n57);
and (n786,n83,n56);
nand (n787,n788,n48);
not (n788,n789);
nor (n789,n790,n791);
and (n790,n56,n103);
and (n791,n57,n102);
and (n792,n771,n772);
and (n793,n746,n752);
xor (n794,n795,n818);
xor (n795,n796,n797);
and (n796,n753,n759);
or (n797,n798,n817);
and (n798,n799,n814);
xor (n799,n800,n806);
nand (n800,n801,n802);
or (n801,n46,n789);
or (n802,n67,n803);
nor (n803,n804,n805);
and (n804,n56,n250);
and (n805,n57,n249);
nand (n806,n807,n812);
or (n807,n808,n129);
not (n808,n809);
nand (n809,n810,n811);
or (n810,n114,n25);
or (n811,n262,n110);
nand (n812,n813,n116);
not (n813,n718);
nand (n814,n815,n816);
or (n815,n28,n778);
or (n816,n727,n30);
and (n817,n800,n806);
xor (n818,n819,n827);
xor (n819,n820,n821);
nor (n820,n180,n262);
nand (n821,n822,n823);
or (n822,n217,n765);
or (n823,n512,n824);
nor (n824,n825,n826);
and (n825,n142,n363);
and (n826,n140,n365);
nand (n827,n828,n829);
or (n828,n46,n803);
or (n829,n67,n830);
nor (n830,n831,n832);
and (n831,n56,n322);
and (n832,n57,n324);
and (n833,n714,n743);
xor (n834,n835,n900);
xor (n835,n836,n871);
xor (n836,n837,n853);
xor (n837,n838,n847);
nand (n838,n839,n843);
or (n839,n179,n840);
nor (n840,n841,n842);
and (n841,n262,n188);
and (n842,n187,n25);
or (n843,n180,n844);
nor (n844,n845,n846);
and (n845,n187,n84);
and (n846,n188,n83);
nand (n847,n848,n849);
or (n848,n135,n740);
or (n849,n136,n850);
nor (n850,n851,n852);
and (n851,n51,n306);
and (n852,n52,n305);
nand (n853,n854,n870);
or (n854,n855,n862);
not (n855,n856);
nand (n856,n857,n188);
nand (n857,n858,n859);
or (n858,n25,n183);
nand (n859,n860,n114);
not (n860,n861);
and (n861,n25,n183);
not (n862,n863);
nand (n863,n864,n865);
or (n864,n217,n824);
or (n865,n512,n866);
not (n866,n867);
nand (n867,n868,n869);
or (n868,n140,n342);
or (n869,n142,n340);
or (n870,n863,n856);
xor (n871,n872,n879);
xor (n872,n873,n876);
or (n873,n874,n875);
and (n874,n819,n827);
and (n875,n820,n821);
or (n876,n877,n878);
and (n877,n715,n734);
and (n878,n716,n725);
xor (n879,n880,n893);
xor (n880,n881,n887);
nand (n881,n882,n883);
or (n882,n46,n830);
or (n883,n67,n884);
nor (n884,n885,n886);
and (n885,n56,n329);
and (n886,n57,n331);
nand (n887,n888,n889);
or (n888,n129,n722);
or (n889,n115,n890);
nor (n890,n891,n892);
and (n891,n114,n250);
and (n892,n110,n249);
nand (n893,n894,n899);
or (n894,n30,n895);
not (n895,n896);
nor (n896,n897,n898);
and (n897,n125,n29);
and (n898,n127,n34);
or (n899,n731,n28);
or (n900,n901,n902);
and (n901,n795,n818);
and (n902,n796,n797);
or (n903,n904,n1160);
and (n904,n905,n945);
xor (n905,n906,n944);
or (n906,n907,n943);
and (n907,n908,n942);
xor (n908,n909,n910);
xor (n909,n799,n814);
or (n910,n911,n941);
and (n911,n912,n927);
xor (n912,n913,n919);
nand (n913,n914,n918);
or (n914,n217,n915);
nor (n915,n916,n917);
and (n916,n331,n140);
and (n917,n329,n142);
or (n918,n512,n761);
nand (n919,n920,n925);
or (n920,n921,n135);
not (n921,n922);
nand (n922,n923,n924);
or (n923,n52,n249);
or (n924,n51,n250);
nand (n925,n926,n171);
not (n926,n748);
and (n927,n928,n934);
nor (n928,n929,n56);
nor (n929,n930,n933);
and (n930,n931,n51);
not (n931,n932);
and (n932,n25,n50);
and (n933,n262,n59);
nand (n934,n935,n940);
or (n935,n28,n936);
not (n936,n937);
nor (n937,n938,n939);
and (n938,n284,n34);
and (n939,n285,n29);
or (n940,n774,n30);
and (n941,n913,n919);
xor (n942,n745,n768);
and (n943,n909,n910);
xor (n944,n713,n794);
or (n945,n946,n1159);
and (n946,n947,n981);
xor (n947,n948,n980);
or (n948,n949,n979);
and (n949,n950,n978);
xor (n950,n951,n977);
or (n951,n952,n976);
and (n952,n953,n969);
xor (n953,n954,n961);
nand (n954,n955,n960);
or (n955,n956,n46);
not (n956,n957);
nand (n957,n958,n959);
or (n958,n56,n25);
or (n959,n262,n57);
nand (n960,n48,n784);
nand (n961,n962,n967);
or (n962,n963,n217);
not (n963,n964);
nor (n964,n965,n966);
and (n965,n324,n142);
and (n966,n322,n140);
nand (n967,n968,n219);
not (n968,n915);
nand (n969,n970,n975);
or (n970,n971,n135);
not (n971,n972);
nor (n972,n973,n974);
and (n973,n103,n52);
and (n974,n102,n51);
nand (n975,n171,n922);
and (n976,n954,n961);
xor (n977,n770,n781);
xor (n978,n912,n927);
and (n979,n951,n977);
xor (n980,n908,n942);
nand (n981,n982,n1158);
or (n982,n983,n1013);
not (n983,n984);
nand (n984,n985,n987);
not (n985,n986);
xor (n986,n950,n978);
not (n987,n988);
or (n988,n989,n1012);
and (n989,n990,n1011);
xor (n990,n991,n992);
xor (n991,n928,n934);
or (n992,n993,n1010);
and (n993,n994,n1003);
xor (n994,n995,n996);
and (n995,n48,n25);
nand (n996,n997,n1002);
or (n997,n28,n998);
not (n998,n999);
nor (n999,n1000,n1001);
and (n1000,n329,n29);
and (n1001,n331,n34);
nand (n1002,n937,n31);
nand (n1003,n1004,n1009);
or (n1004,n1005,n217);
not (n1005,n1006);
nor (n1006,n1007,n1008);
and (n1007,n249,n142);
and (n1008,n250,n140);
nand (n1009,n219,n964);
and (n1010,n995,n996);
xor (n1011,n953,n969);
and (n1012,n991,n992);
not (n1013,n1014);
nand (n1014,n1015,n1157);
or (n1015,n1016,n1047);
not (n1016,n1017);
nand (n1017,n1018,n1020);
not (n1018,n1019);
xor (n1019,n990,n1011);
not (n1020,n1021);
or (n1021,n1022,n1046);
and (n1022,n1023,n1045);
xor (n1023,n1024,n1031);
nand (n1024,n1025,n1030);
or (n1025,n1026,n135);
not (n1026,n1027);
nor (n1027,n1028,n1029);
and (n1028,n84,n52);
and (n1029,n83,n51);
nand (n1030,n171,n972);
and (n1031,n1032,n1037);
and (n1032,n1033,n52);
nand (n1033,n1034,n1036);
or (n1034,n1035,n140);
and (n1035,n25,n139);
or (n1036,n25,n139);
nand (n1037,n1038,n1039);
or (n1038,n30,n998);
nand (n1039,n1040,n1044);
not (n1040,n1041);
nor (n1041,n1042,n1043);
and (n1042,n322,n34);
and (n1043,n324,n29);
not (n1044,n28);
xor (n1045,n994,n1003);
and (n1046,n1024,n1031);
not (n1047,n1048);
nand (n1048,n1049,n1156);
or (n1049,n1050,n1074);
not (n1050,n1051);
nand (n1051,n1052,n1054);
not (n1052,n1053);
xor (n1053,n1023,n1045);
not (n1054,n1055);
or (n1055,n1056,n1073);
and (n1056,n1057,n1072);
xor (n1057,n1058,n1065);
nand (n1058,n1059,n1064);
or (n1059,n1060,n217);
not (n1060,n1061);
nor (n1061,n1062,n1063);
and (n1062,n102,n142);
and (n1063,n103,n140);
nand (n1064,n219,n1006);
nand (n1065,n1066,n1071);
or (n1066,n1067,n135);
not (n1067,n1068);
nand (n1068,n1069,n1070);
or (n1069,n51,n25);
or (n1070,n52,n262);
nand (n1071,n171,n1027);
xor (n1072,n1032,n1037);
and (n1073,n1058,n1065);
not (n1074,n1075);
nand (n1075,n1076,n1155);
or (n1076,n1077,n1101);
not (n1077,n1078);
nand (n1078,n1079,n1081);
not (n1079,n1080);
xor (n1080,n1057,n1072);
not (n1081,n1082);
or (n1082,n1083,n1100);
and (n1083,n1084,n1093);
xor (n1084,n1085,n1086);
and (n1085,n171,n25);
nand (n1086,n1087,n1092);
or (n1087,n1088,n217);
not (n1088,n1089);
nor (n1089,n1090,n1091);
and (n1090,n84,n140);
and (n1091,n83,n142);
nand (n1092,n219,n1061);
nand (n1093,n1094,n1099);
or (n1094,n28,n1095);
not (n1095,n1096);
nor (n1096,n1097,n1098);
and (n1097,n249,n34);
and (n1098,n250,n29);
or (n1099,n1041,n30);
and (n1100,n1085,n1086);
not (n1101,n1102);
nand (n1102,n1103,n1154);
or (n1103,n1104,n1120);
nor (n1104,n1105,n1106);
xor (n1105,n1084,n1093);
and (n1106,n1107,n1113);
nor (n1107,n1108,n142);
nor (n1108,n1109,n1110);
and (n1109,n226,n262);
and (n1110,n1111,n34);
not (n1111,n1112);
and (n1112,n25,n221);
nand (n1113,n1114,n1115);
or (n1114,n30,n1095);
nand (n1115,n1116,n1044);
not (n1116,n1117);
nor (n1117,n1118,n1119);
and (n1118,n34,n103);
and (n1119,n29,n102);
not (n1120,n1121);
or (n1121,n1122,n1153);
and (n1122,n1123,n1132);
xor (n1123,n1124,n1131);
nand (n1124,n1125,n1130);
or (n1125,n1126,n217);
not (n1126,n1127);
nand (n1127,n1128,n1129);
or (n1128,n142,n25);
or (n1129,n140,n262);
nand (n1130,n219,n1089);
xor (n1131,n1107,n1113);
or (n1132,n1133,n1152);
and (n1133,n1134,n1142);
xor (n1134,n1135,n1136);
nor (n1135,n512,n262);
nand (n1136,n1137,n1141);
or (n1137,n1138,n28);
nor (n1138,n1139,n1140);
and (n1139,n34,n84);
and (n1140,n29,n83);
or (n1141,n1117,n30);
nor (n1142,n1143,n1150);
nor (n1143,n1144,n1146);
and (n1144,n1145,n31);
not (n1145,n1138);
nor (n1146,n1147,n28);
nor (n1147,n1148,n1149);
and (n1148,n25,n34);
and (n1149,n262,n29);
or (n1150,n1151,n34);
and (n1151,n25,n31);
and (n1152,n1135,n1136);
and (n1153,n1124,n1131);
nand (n1154,n1105,n1106);
nand (n1155,n1080,n1082);
nand (n1156,n1053,n1055);
nand (n1157,n1019,n1021);
nand (n1158,n986,n988);
and (n1159,n948,n980);
and (n1160,n906,n944);
and (n1161,n711,n834);
nor (n1162,n1163,n1361);
not (n1163,n1164);
or (n1164,n1165,n1346);
xor (n1165,n1166,n1329);
xor (n1166,n1167,n1251);
xor (n1167,n1168,n1233);
xor (n1168,n1169,n1201);
or (n1169,n1170,n1200);
and (n1170,n1171,n1191);
xor (n1171,n1172,n1181);
nand (n1172,n1173,n1177);
or (n1173,n217,n1174);
nor (n1174,n1175,n1176);
and (n1175,n142,n192);
and (n1176,n140,n194);
or (n1177,n512,n1178);
nor (n1178,n1179,n1180);
and (n1179,n142,n125);
and (n1180,n140,n127);
nand (n1181,n1182,n1186);
or (n1182,n46,n1183);
nor (n1183,n1184,n1185);
and (n1184,n56,n285);
and (n1185,n57,n284);
or (n1186,n67,n1187);
not (n1187,n1188);
nor (n1188,n1189,n1190);
and (n1189,n306,n57);
and (n1190,n305,n56);
nand (n1191,n1192,n1196);
or (n1192,n129,n1193);
nor (n1193,n1194,n1195);
and (n1194,n114,n322);
and (n1195,n110,n324);
or (n1196,n115,n1197);
nor (n1197,n1198,n1199);
and (n1198,n114,n329);
and (n1199,n110,n331);
and (n1200,n1172,n1181);
or (n1201,n1202,n1232);
and (n1202,n1203,n1222);
xor (n1203,n1204,n1213);
nand (n1204,n1205,n1209);
or (n1205,n135,n1206);
nor (n1206,n1207,n1208);
and (n1207,n51,n363);
and (n1208,n52,n365);
or (n1209,n136,n1210);
nor (n1210,n1211,n1212);
and (n1211,n51,n340);
and (n1212,n52,n342);
nand (n1213,n1214,n1218);
or (n1214,n179,n1215);
nor (n1215,n1216,n1217);
and (n1216,n187,n103);
and (n1217,n188,n102);
or (n1218,n180,n1219);
nor (n1219,n1220,n1221);
and (n1220,n187,n250);
and (n1221,n188,n249);
nand (n1222,n1223,n1228);
or (n1223,n1224,n360);
not (n1224,n1225);
nand (n1225,n1226,n1227);
or (n1226,n83,n294);
or (n1227,n293,n84);
or (n1228,n346,n1229);
nor (n1229,n1230,n1231);
and (n1230,n262,n294);
and (n1231,n25,n293);
and (n1232,n1204,n1213);
xor (n1233,n1234,n1245);
xor (n1234,n1235,n1236);
nor (n1235,n290,n262);
nand (n1236,n1237,n1241);
or (n1237,n28,n1238);
nor (n1238,n1239,n1240);
and (n1239,n34,n64);
and (n1240,n29,n63);
or (n1241,n1242,n30);
nor (n1242,n1243,n1244);
and (n1243,n34,n71);
and (n1244,n29,n73);
nand (n1245,n1246,n1247);
or (n1246,n217,n1178);
or (n1247,n512,n1248);
nor (n1248,n1249,n1250);
and (n1249,n142,n112);
and (n1250,n140,n111);
xor (n1251,n1252,n1300);
xor (n1252,n1253,n1274);
xor (n1253,n1254,n1268);
xor (n1254,n1255,n1262);
nand (n1255,n1256,n1257);
or (n1256,n1187,n46);
nand (n1257,n1258,n48);
not (n1258,n1259);
nor (n1259,n1260,n1261);
and (n1260,n56,n363);
and (n1261,n57,n365);
nand (n1262,n1263,n1264);
or (n1263,n129,n1197);
or (n1264,n115,n1265);
nor (n1265,n1266,n1267);
and (n1266,n284,n110);
and (n1267,n285,n114);
nand (n1268,n1269,n1270);
or (n1269,n135,n1210);
or (n1270,n136,n1271);
nor (n1271,n1272,n1273);
and (n1272,n51,n192);
and (n1273,n52,n194);
xor (n1274,n1275,n1288);
xor (n1275,n1276,n1282);
nand (n1276,n1277,n1278);
or (n1277,n179,n1219);
or (n1278,n180,n1279);
nor (n1279,n1280,n1281);
and (n1280,n187,n322);
and (n1281,n188,n324);
nand (n1282,n1283,n1284);
or (n1283,n1224,n346);
or (n1284,n360,n1285);
nor (n1285,n1286,n1287);
and (n1286,n293,n103);
and (n1287,n294,n102);
and (n1288,n1289,n1294);
nor (n1289,n1290,n293);
nor (n1290,n1291,n1293);
and (n1291,n1292,n187);
nand (n1292,n25,n350);
and (n1293,n262,n355);
nand (n1294,n1295,n1299);
or (n1295,n1296,n28);
nor (n1296,n1297,n1298);
and (n1297,n34,n112);
and (n1298,n29,n111);
or (n1299,n1238,n30);
or (n1300,n1301,n1328);
and (n1301,n1302,n1315);
xor (n1302,n1303,n1304);
xor (n1303,n1289,n1294);
or (n1304,n1305,n1314);
and (n1305,n1306,n1311);
xor (n1306,n1307,n1308);
nor (n1307,n360,n262);
nand (n1308,n1309,n1310);
or (n1309,n866,n217);
or (n1310,n512,n1174);
nand (n1311,n1312,n1313);
or (n1312,n46,n884);
or (n1313,n67,n1183);
and (n1314,n1307,n1308);
or (n1315,n1316,n1327);
and (n1316,n1317,n1324);
xor (n1317,n1318,n1321);
nand (n1318,n1319,n1320);
or (n1319,n129,n890);
or (n1320,n115,n1193);
nand (n1321,n1322,n1323);
or (n1322,n28,n895);
or (n1323,n1296,n30);
nand (n1324,n1325,n1326);
or (n1325,n179,n844);
or (n1326,n180,n1215);
and (n1327,n1318,n1321);
and (n1328,n1303,n1304);
or (n1329,n1330,n1345);
and (n1330,n1331,n1334);
xor (n1331,n1332,n1333);
xor (n1332,n1203,n1222);
xor (n1333,n1171,n1191);
or (n1334,n1335,n1344);
and (n1335,n1336,n1341);
xor (n1336,n1337,n1340);
nand (n1337,n1338,n1339);
or (n1338,n135,n850);
or (n1339,n136,n1206);
nor (n1340,n862,n856);
or (n1341,n1342,n1343);
and (n1342,n880,n893);
and (n1343,n881,n887);
and (n1344,n1337,n1340);
and (n1345,n1332,n1333);
or (n1346,n1347,n1360);
and (n1347,n1348,n1359);
xor (n1348,n1349,n1350);
xor (n1349,n1302,n1315);
or (n1350,n1351,n1358);
and (n1351,n1352,n1355);
xor (n1352,n1353,n1354);
xor (n1353,n1317,n1324);
xor (n1354,n1306,n1311);
or (n1355,n1356,n1357);
and (n1356,n837,n853);
and (n1357,n838,n847);
and (n1358,n1353,n1354);
xor (n1359,n1331,n1334);
and (n1360,n1349,n1350);
nand (n1361,n1362,n1374);
not (n1362,n1363);
nor (n1363,n1364,n1365);
xor (n1364,n1348,n1359);
or (n1365,n1366,n1373);
and (n1366,n1367,n1372);
xor (n1367,n1368,n1369);
xor (n1368,n1336,n1341);
or (n1369,n1370,n1371);
and (n1370,n872,n879);
and (n1371,n873,n876);
xor (n1372,n1352,n1355);
and (n1373,n1368,n1369);
or (n1374,n1375,n1378);
or (n1375,n1376,n1377);
and (n1376,n835,n900);
and (n1377,n836,n871);
xor (n1378,n1367,n1372);
or (n1379,n1380,n1467);
xor (n1380,n1381,n1436);
xor (n1381,n1382,n1433);
xor (n1382,n1383,n1409);
xor (n1383,n1384,n1387);
or (n1384,n1385,n1386);
and (n1385,n1254,n1268);
and (n1386,n1255,n1262);
xor (n1387,n1388,n1403);
xor (n1388,n1389,n1396);
nand (n1389,n1390,n1391);
or (n1390,n1265,n129);
nand (n1391,n1392,n116);
not (n1392,n1393);
nor (n1393,n1394,n1395);
and (n1394,n306,n114);
and (n1395,n110,n305);
nand (n1396,n1397,n1398);
or (n1397,n1271,n135);
nand (n1398,n1399,n171);
not (n1399,n1400);
nor (n1400,n1401,n1402);
and (n1401,n51,n125);
and (n1402,n52,n127);
nand (n1403,n1404,n1405);
or (n1404,n179,n1279);
or (n1405,n180,n1406);
nor (n1406,n1407,n1408);
and (n1407,n187,n329);
and (n1408,n188,n331);
xor (n1409,n1410,n1427);
xor (n1410,n1411,n1418);
nand (n1411,n1412,n1416);
or (n1412,n1413,n512);
nor (n1413,n1414,n1415);
and (n1414,n142,n64);
and (n1415,n140,n63);
nand (n1416,n1417,n218);
not (n1417,n1248);
nand (n1418,n1419,n1423);
or (n1419,n289,n1420);
nor (n1420,n1421,n1422);
and (n1421,n286,n262);
and (n1422,n288,n25);
or (n1423,n290,n1424);
nor (n1424,n1425,n1426);
and (n1425,n288,n84);
and (n1426,n286,n83);
nand (n1427,n1428,n1429);
or (n1428,n46,n1259);
or (n1429,n67,n1430);
nor (n1430,n1431,n1432);
and (n1431,n56,n340);
and (n1432,n57,n342);
or (n1433,n1434,n1435);
and (n1434,n1252,n1300);
and (n1435,n1253,n1274);
xor (n1436,n1437,n1464);
xor (n1437,n1438,n1441);
or (n1438,n1439,n1440);
and (n1439,n1275,n1288);
and (n1440,n1276,n1282);
xor (n1441,n1442,n1461);
xor (n1442,n1443,n1449);
nand (n1443,n1444,n1445);
or (n1444,n346,n1285);
or (n1445,n360,n1446);
nor (n1446,n1447,n1448);
and (n1447,n293,n250);
and (n1448,n294,n249);
xor (n1449,n1450,n1455);
nor (n1450,n1451,n288);
nor (n1451,n1452,n1454);
and (n1452,n1453,n293);
nand (n1453,n25,n295);
and (n1454,n262,n300);
nand (n1455,n1456,n1457);
or (n1456,n28,n1242);
or (n1457,n1458,n30);
nor (n1458,n1459,n1460);
and (n1459,n34,n149);
and (n1460,n29,n148);
or (n1461,n1462,n1463);
and (n1462,n1234,n1245);
and (n1463,n1235,n1236);
or (n1464,n1465,n1466);
and (n1465,n1168,n1233);
and (n1466,n1169,n1201);
or (n1467,n1468,n1469);
and (n1468,n1166,n1329);
and (n1469,n1167,n1251);
nand (n1470,n1471,n1379);
nand (n1471,n1472,n1478);
or (n1472,n1163,n1473);
not (n1473,n1474);
nand (n1474,n1475,n1477);
or (n1475,n1363,n1476);
nand (n1476,n1375,n1378);
nand (n1477,n1364,n1365);
nand (n1478,n1165,n1346);
nand (n1479,n1380,n1467);
not (n1480,n1481);
and (n1481,n1482,n1671,n1704);
not (n1482,n1483);
nor (n1483,n1484,n1642);
xor (n1484,n1485,n1627);
xor (n1485,n1486,n1535);
xor (n1486,n1487,n1534);
xor (n1487,n1488,n1489);
xor (n1488,n570,n584);
or (n1489,n1490,n1533);
and (n1490,n1491,n1510);
xor (n1491,n1492,n1498);
nand (n1492,n1493,n1497);
or (n1493,n346,n1494);
nor (n1494,n1495,n1496);
and (n1495,n293,n329);
and (n1496,n294,n331);
or (n1497,n360,n563);
and (n1498,n1499,n1504);
nor (n1499,n1500,n91);
nor (n1500,n1501,n1503);
and (n1501,n1502,n288);
nand (n1502,n25,n314);
and (n1503,n262,n316);
nand (n1504,n1505,n1509);
or (n1505,n28,n1506);
nor (n1506,n1507,n1508);
and (n1507,n34,n154);
and (n1508,n29,n156);
or (n1509,n626,n30);
or (n1510,n1511,n1532);
and (n1511,n1512,n1526);
xor (n1512,n1513,n1520);
nand (n1513,n1514,n1518);
or (n1514,n1515,n46);
nor (n1515,n1516,n1517);
and (n1516,n56,n192);
and (n1517,n57,n194);
nand (n1518,n1519,n48);
not (n1519,n632);
nand (n1520,n1521,n1525);
or (n1521,n289,n1522);
nor (n1522,n1523,n1524);
and (n1523,n288,n103);
and (n1524,n286,n102);
or (n1525,n290,n642);
nand (n1526,n1527,n1531);
or (n1527,n310,n1528);
nor (n1528,n1529,n1530);
and (n1529,n262,n92);
and (n1530,n91,n25);
or (n1531,n326,n648);
and (n1532,n1513,n1520);
and (n1533,n1492,n1498);
xor (n1534,n618,n637);
or (n1535,n1536,n1626);
and (n1536,n1537,n1619);
xor (n1537,n1538,n1594);
or (n1538,n1539,n1593);
and (n1539,n1540,n1577);
xor (n1540,n1541,n1555);
or (n1541,n1542,n1554);
and (n1542,n1543,n1548);
xor (n1543,n1544,n1545);
and (n1544,n317,n25);
nand (n1545,n1546,n1547);
or (n1546,n28,n1458);
or (n1547,n1506,n30);
nand (n1548,n1549,n1550);
or (n1549,n217,n1413);
or (n1550,n512,n1551);
nor (n1551,n1552,n1553);
and (n1552,n142,n71);
and (n1553,n140,n73);
and (n1554,n1544,n1545);
or (n1555,n1556,n1576);
and (n1556,n1557,n1570);
xor (n1557,n1558,n1564);
nand (n1558,n1559,n1560);
or (n1559,n135,n1400);
or (n1560,n136,n1561);
nor (n1561,n1562,n1563);
and (n1562,n51,n112);
and (n1563,n52,n111);
nand (n1564,n1565,n1566);
or (n1565,n179,n1406);
or (n1566,n180,n1567);
nor (n1567,n1568,n1569);
and (n1568,n187,n285);
and (n1569,n188,n284);
nand (n1570,n1571,n1572);
or (n1571,n346,n1446);
or (n1572,n360,n1573);
nor (n1573,n1574,n1575);
and (n1574,n293,n322);
and (n1575,n294,n324);
and (n1576,n1558,n1564);
or (n1577,n1578,n1592);
and (n1578,n1579,n1586);
xor (n1579,n1580,n1583);
nand (n1580,n1581,n1582);
or (n1581,n289,n1424);
or (n1582,n290,n1522);
nand (n1583,n1584,n1585);
or (n1584,n46,n1430);
or (n1585,n67,n1515);
nand (n1586,n1587,n1588);
or (n1587,n129,n1393);
or (n1588,n115,n1589);
nor (n1589,n1590,n1591);
and (n1590,n114,n363);
and (n1591,n110,n365);
and (n1592,n1580,n1583);
and (n1593,n1541,n1555);
or (n1594,n1595,n1618);
and (n1595,n1596,n1609);
xor (n1596,n1597,n1598);
xor (n1597,n1512,n1526);
xor (n1598,n1599,n1606);
xor (n1599,n1600,n1603);
nand (n1600,n1601,n1602);
or (n1601,n217,n1551);
or (n1602,n512,n654);
nand (n1603,n1604,n1605);
or (n1604,n129,n1589);
or (n1605,n115,n668);
nand (n1606,n1607,n1608);
or (n1607,n135,n1561);
or (n1608,n136,n675);
xor (n1609,n1610,n1617);
xor (n1610,n1611,n1614);
nand (n1611,n1612,n1613);
or (n1612,n179,n1567);
or (n1613,n180,n681);
nand (n1614,n1615,n1616);
or (n1615,n346,n1573);
or (n1616,n360,n1494);
xor (n1617,n1499,n1504);
and (n1618,n1597,n1598);
xor (n1619,n1620,n1625);
xor (n1620,n1621,n1624);
or (n1621,n1622,n1623);
and (n1622,n1599,n1606);
and (n1623,n1600,n1603);
xor (n1624,n665,n679);
xor (n1625,n622,n630);
and (n1626,n1538,n1594);
xor (n1627,n1628,n1633);
xor (n1628,n1629,n1632);
or (n1629,n1630,n1631);
and (n1630,n1620,n1625);
and (n1631,n1621,n1624);
xor (n1632,n662,n687);
or (n1633,n1634,n1641);
and (n1634,n1635,n1640);
xor (n1635,n1636,n1637);
xor (n1636,n639,n652);
or (n1637,n1638,n1639);
and (n1638,n1610,n1617);
and (n1639,n1611,n1614);
xor (n1640,n1491,n1510);
and (n1641,n1636,n1637);
or (n1642,n1643,n1670);
and (n1643,n1644,n1669);
xor (n1644,n1645,n1646);
xor (n1645,n1635,n1640);
or (n1646,n1647,n1668);
and (n1647,n1648,n1661);
xor (n1648,n1649,n1660);
or (n1649,n1650,n1659);
and (n1650,n1651,n1656);
xor (n1651,n1652,n1653);
and (n1652,n1450,n1455);
or (n1653,n1654,n1655);
and (n1654,n1410,n1427);
and (n1655,n1411,n1418);
or (n1656,n1657,n1658);
and (n1657,n1388,n1403);
and (n1658,n1389,n1396);
and (n1659,n1652,n1653);
xor (n1660,n1540,n1577);
or (n1661,n1662,n1667);
and (n1662,n1663,n1666);
xor (n1663,n1664,n1665);
xor (n1664,n1557,n1570);
xor (n1665,n1543,n1548);
xor (n1666,n1579,n1586);
and (n1667,n1664,n1665);
and (n1668,n1649,n1660);
xor (n1669,n1537,n1619);
and (n1670,n1645,n1646);
and (n1671,n1672,n1699);
nand (n1672,n1673,n1689);
not (n1673,n1674);
xor (n1674,n1675,n1688);
xor (n1675,n1676,n1677);
xor (n1676,n1596,n1609);
or (n1677,n1678,n1687);
and (n1678,n1679,n1684);
xor (n1679,n1680,n1683);
or (n1680,n1681,n1682);
and (n1681,n1442,n1461);
and (n1682,n1443,n1449);
xor (n1683,n1651,n1656);
or (n1684,n1685,n1686);
and (n1685,n1383,n1409);
and (n1686,n1384,n1387);
and (n1687,n1680,n1683);
xor (n1688,n1648,n1661);
not (n1689,n1690);
or (n1690,n1691,n1698);
and (n1691,n1692,n1697);
xor (n1692,n1693,n1694);
xor (n1693,n1663,n1666);
or (n1694,n1695,n1696);
and (n1695,n1437,n1464);
and (n1696,n1438,n1441);
xor (n1697,n1679,n1684);
and (n1698,n1693,n1694);
or (n1699,n1700,n1703);
or (n1700,n1701,n1702);
and (n1701,n1381,n1436);
and (n1702,n1382,n1433);
xor (n1703,n1692,n1697);
not (n1704,n1705);
nor (n1705,n1706,n1707);
xor (n1706,n1644,n1669);
or (n1707,n1708,n1709);
and (n1708,n1675,n1688);
and (n1709,n1676,n1677);
not (n1710,n1711);
nand (n1711,n1712,n1723);
or (n1712,n1713,n1483);
nor (n1713,n1714,n1722);
and (n1714,n1715,n1704);
not (n1715,n1716);
nand (n1716,n1717,n1672);
or (n1717,n1718,n1720);
not (n1718,n1719);
nand (n1719,n1703,n1700);
not (n1720,n1721);
nand (n1721,n1674,n1690);
and (n1722,n1706,n1707);
nand (n1723,n1484,n1642);
nor (n1724,n1725,n1738);
nor (n1725,n1726,n1727);
xor (n1726,n611,n691);
or (n1727,n1728,n1737);
and (n1728,n1729,n1736);
xor (n1729,n1730,n1733);
or (n1730,n1731,n1732);
and (n1731,n1487,n1534);
and (n1732,n1488,n1489);
or (n1733,n1734,n1735);
and (n1734,n1628,n1633);
and (n1735,n1629,n1632);
xor (n1736,n693,n696);
and (n1737,n1730,n1733);
nor (n1738,n1739,n1740);
xor (n1739,n1729,n1736);
or (n1740,n1741,n1742);
and (n1741,n1485,n1627);
and (n1742,n1486,n1535);
not (n1743,n1744);
nand (n1744,n1745,n1747);
or (n1745,n1725,n1746);
nand (n1746,n1739,n1740);
nand (n1747,n1726,n1727);
or (n1748,n701,n3);
xor (n1749,n1750,n3110);
xor (n1750,n1751,n3107);
xor (n1751,n1752,n3106);
xor (n1752,n1753,n3098);
xor (n1753,n1754,n3097);
xor (n1754,n1755,n3082);
xor (n1755,n1756,n251);
xor (n1756,n1757,n3061);
xor (n1757,n1758,n3060);
xor (n1758,n1759,n3033);
xor (n1759,n1760,n3032);
xor (n1760,n1761,n2999);
xor (n1761,n1762,n2998);
xor (n1762,n1763,n2960);
xor (n1763,n1764,n2959);
xor (n1764,n1765,n2914);
xor (n1765,n1766,n2913);
xor (n1766,n1767,n2862);
xor (n1767,n1768,n2861);
xor (n1768,n1769,n2804);
xor (n1769,n1770,n2803);
xor (n1770,n1771,n2740);
xor (n1771,n1772,n2739);
xor (n1772,n1773,n2671);
xor (n1773,n1774,n2670);
xor (n1774,n1775,n2596);
xor (n1775,n1776,n2595);
xor (n1776,n1777,n2515);
xor (n1777,n1778,n2514);
xor (n1778,n1779,n2432);
xor (n1779,n1780,n278);
xor (n1780,n1781,n2340);
xor (n1781,n1782,n2339);
xor (n1782,n1783,n2242);
xor (n1783,n1784,n173);
xor (n1784,n1785,n2138);
xor (n1785,n1786,n2137);
xor (n1786,n1787,n2030);
xor (n1787,n1788,n229);
xor (n1788,n1789,n1914);
xor (n1789,n1790,n1913);
xor (n1790,n1791,n1794);
xor (n1791,n1792,n1793);
and (n1792,n458,n31);
and (n1793,n165,n29);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
and (n1796,n165,n31);
and (n1797,n42,n29);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
and (n1802,n42,n31);
and (n1803,n35,n29);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
and (n1808,n35,n31);
and (n1809,n214,n29);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
and (n1814,n214,n31);
and (n1815,n174,n29);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
and (n1820,n174,n31);
and (n1821,n154,n29);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
and (n1826,n154,n31);
and (n1827,n149,n29);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
and (n1832,n149,n31);
and (n1833,n71,n29);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
and (n1838,n71,n31);
and (n1839,n64,n29);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
and (n1844,n64,n31);
and (n1845,n112,n29);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1851);
and (n1849,n1850,n897);
and (n1850,n112,n31);
and (n1851,n1852,n1853);
xor (n1852,n1850,n897);
or (n1853,n1854,n1857);
and (n1854,n1855,n1856);
and (n1855,n125,n31);
and (n1856,n192,n29);
and (n1857,n1858,n1859);
xor (n1858,n1855,n1856);
or (n1859,n1860,n1863);
and (n1860,n1861,n1862);
and (n1861,n192,n31);
and (n1862,n340,n29);
and (n1863,n1864,n1865);
xor (n1864,n1861,n1862);
or (n1865,n1866,n1869);
and (n1866,n1867,n1868);
and (n1867,n340,n31);
and (n1868,n363,n29);
and (n1869,n1870,n1871);
xor (n1870,n1867,n1868);
or (n1871,n1872,n1875);
and (n1872,n1873,n1874);
and (n1873,n363,n31);
and (n1874,n306,n29);
and (n1875,n1876,n1877);
xor (n1876,n1873,n1874);
or (n1877,n1878,n1880);
and (n1878,n1879,n939);
and (n1879,n306,n31);
and (n1880,n1881,n1882);
xor (n1881,n1879,n939);
or (n1882,n1883,n1885);
and (n1883,n1884,n1000);
and (n1884,n285,n31);
and (n1885,n1886,n1887);
xor (n1886,n1884,n1000);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
and (n1889,n329,n31);
and (n1890,n322,n29);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
or (n1893,n1894,n1896);
and (n1894,n1895,n1098);
and (n1895,n322,n31);
and (n1896,n1897,n1898);
xor (n1897,n1895,n1098);
or (n1898,n1899,n1902);
and (n1899,n1900,n1901);
and (n1900,n250,n31);
and (n1901,n103,n29);
and (n1902,n1903,n1904);
xor (n1903,n1900,n1901);
or (n1904,n1905,n1908);
and (n1905,n1906,n1907);
and (n1906,n103,n31);
and (n1907,n84,n29);
and (n1908,n1909,n1910);
xor (n1909,n1906,n1907);
and (n1910,n1911,n1912);
and (n1911,n84,n31);
and (n1912,n25,n29);
and (n1913,n42,n221);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1799,n1800);
and (n1917,n35,n221);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
or (n1920,n1921,n1924);
and (n1921,n1922,n1923);
xor (n1922,n1805,n1806);
and (n1923,n214,n221);
and (n1924,n1925,n1926);
xor (n1925,n1922,n1923);
or (n1926,n1927,n1930);
and (n1927,n1928,n1929);
xor (n1928,n1811,n1812);
and (n1929,n174,n221);
and (n1930,n1931,n1932);
xor (n1931,n1928,n1929);
or (n1932,n1933,n1936);
and (n1933,n1934,n1935);
xor (n1934,n1817,n1818);
and (n1935,n154,n221);
and (n1936,n1937,n1938);
xor (n1937,n1934,n1935);
or (n1938,n1939,n1942);
and (n1939,n1940,n1941);
xor (n1940,n1823,n1824);
and (n1941,n149,n221);
and (n1942,n1943,n1944);
xor (n1943,n1940,n1941);
or (n1944,n1945,n1948);
and (n1945,n1946,n1947);
xor (n1946,n1829,n1830);
and (n1947,n71,n221);
and (n1948,n1949,n1950);
xor (n1949,n1946,n1947);
or (n1950,n1951,n1954);
and (n1951,n1952,n1953);
xor (n1952,n1835,n1836);
and (n1953,n64,n221);
and (n1954,n1955,n1956);
xor (n1955,n1952,n1953);
or (n1956,n1957,n1960);
and (n1957,n1958,n1959);
xor (n1958,n1841,n1842);
and (n1959,n112,n221);
and (n1960,n1961,n1962);
xor (n1961,n1958,n1959);
or (n1962,n1963,n1966);
and (n1963,n1964,n1965);
xor (n1964,n1847,n1848);
and (n1965,n125,n221);
and (n1966,n1967,n1968);
xor (n1967,n1964,n1965);
or (n1968,n1969,n1972);
and (n1969,n1970,n1971);
xor (n1970,n1852,n1853);
and (n1971,n192,n221);
and (n1972,n1973,n1974);
xor (n1973,n1970,n1971);
or (n1974,n1975,n1978);
and (n1975,n1976,n1977);
xor (n1976,n1858,n1859);
and (n1977,n340,n221);
and (n1978,n1979,n1980);
xor (n1979,n1976,n1977);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
xor (n1982,n1864,n1865);
and (n1983,n363,n221);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1870,n1871);
and (n1989,n306,n221);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1996);
and (n1993,n1994,n1995);
xor (n1994,n1876,n1877);
and (n1995,n285,n221);
and (n1996,n1997,n1998);
xor (n1997,n1994,n1995);
or (n1998,n1999,n2002);
and (n1999,n2000,n2001);
xor (n2000,n1881,n1882);
and (n2001,n329,n221);
and (n2002,n2003,n2004);
xor (n2003,n2000,n2001);
or (n2004,n2005,n2008);
and (n2005,n2006,n2007);
xor (n2006,n1886,n1887);
and (n2007,n322,n221);
and (n2008,n2009,n2010);
xor (n2009,n2006,n2007);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1892,n1893);
and (n2013,n250,n221);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
or (n2016,n2017,n2020);
and (n2017,n2018,n2019);
xor (n2018,n1897,n1898);
and (n2019,n103,n221);
and (n2020,n2021,n2022);
xor (n2021,n2018,n2019);
or (n2022,n2023,n2026);
and (n2023,n2024,n2025);
xor (n2024,n1903,n1904);
and (n2025,n84,n221);
and (n2026,n2027,n2028);
xor (n2027,n2024,n2025);
and (n2028,n2029,n1112);
xor (n2029,n1909,n1910);
or (n2030,n2031,n2034);
and (n2031,n2032,n2033);
xor (n2032,n1919,n1920);
and (n2033,n214,n140);
and (n2034,n2035,n2036);
xor (n2035,n2032,n2033);
or (n2036,n2037,n2040);
and (n2037,n2038,n2039);
xor (n2038,n1925,n1926);
and (n2039,n174,n140);
and (n2040,n2041,n2042);
xor (n2041,n2038,n2039);
or (n2042,n2043,n2046);
and (n2043,n2044,n2045);
xor (n2044,n1931,n1932);
and (n2045,n154,n140);
and (n2046,n2047,n2048);
xor (n2047,n2044,n2045);
or (n2048,n2049,n2052);
and (n2049,n2050,n2051);
xor (n2050,n1937,n1938);
and (n2051,n149,n140);
and (n2052,n2053,n2054);
xor (n2053,n2050,n2051);
or (n2054,n2055,n2058);
and (n2055,n2056,n2057);
xor (n2056,n1943,n1944);
and (n2057,n71,n140);
and (n2058,n2059,n2060);
xor (n2059,n2056,n2057);
or (n2060,n2061,n2064);
and (n2061,n2062,n2063);
xor (n2062,n1949,n1950);
and (n2063,n64,n140);
and (n2064,n2065,n2066);
xor (n2065,n2062,n2063);
or (n2066,n2067,n2070);
and (n2067,n2068,n2069);
xor (n2068,n1955,n1956);
and (n2069,n112,n140);
and (n2070,n2071,n2072);
xor (n2071,n2068,n2069);
or (n2072,n2073,n2076);
and (n2073,n2074,n2075);
xor (n2074,n1961,n1962);
and (n2075,n125,n140);
and (n2076,n2077,n2078);
xor (n2077,n2074,n2075);
or (n2078,n2079,n2082);
and (n2079,n2080,n2081);
xor (n2080,n1967,n1968);
and (n2081,n192,n140);
and (n2082,n2083,n2084);
xor (n2083,n2080,n2081);
or (n2084,n2085,n2088);
and (n2085,n2086,n2087);
xor (n2086,n1973,n1974);
and (n2087,n340,n140);
and (n2088,n2089,n2090);
xor (n2089,n2086,n2087);
or (n2090,n2091,n2094);
and (n2091,n2092,n2093);
xor (n2092,n1979,n1980);
and (n2093,n363,n140);
and (n2094,n2095,n2096);
xor (n2095,n2092,n2093);
or (n2096,n2097,n2100);
and (n2097,n2098,n2099);
xor (n2098,n1985,n1986);
and (n2099,n306,n140);
and (n2100,n2101,n2102);
xor (n2101,n2098,n2099);
or (n2102,n2103,n2106);
and (n2103,n2104,n2105);
xor (n2104,n1991,n1992);
and (n2105,n285,n140);
and (n2106,n2107,n2108);
xor (n2107,n2104,n2105);
or (n2108,n2109,n2112);
and (n2109,n2110,n2111);
xor (n2110,n1997,n1998);
and (n2111,n329,n140);
and (n2112,n2113,n2114);
xor (n2113,n2110,n2111);
or (n2114,n2115,n2117);
and (n2115,n2116,n966);
xor (n2116,n2003,n2004);
and (n2117,n2118,n2119);
xor (n2118,n2116,n966);
or (n2119,n2120,n2122);
and (n2120,n2121,n1008);
xor (n2121,n2009,n2010);
and (n2122,n2123,n2124);
xor (n2123,n2121,n1008);
or (n2124,n2125,n2127);
and (n2125,n2126,n1063);
xor (n2126,n2015,n2016);
and (n2127,n2128,n2129);
xor (n2128,n2126,n1063);
or (n2129,n2130,n2132);
and (n2130,n2131,n1090);
xor (n2131,n2021,n2022);
and (n2132,n2133,n2134);
xor (n2133,n2131,n1090);
and (n2134,n2135,n2136);
xor (n2135,n2027,n2028);
and (n2136,n25,n140);
and (n2137,n214,n139);
or (n2138,n2139,n2142);
and (n2139,n2140,n2141);
xor (n2140,n2035,n2036);
and (n2141,n174,n139);
and (n2142,n2143,n2144);
xor (n2143,n2140,n2141);
or (n2144,n2145,n2148);
and (n2145,n2146,n2147);
xor (n2146,n2041,n2042);
and (n2147,n154,n139);
and (n2148,n2149,n2150);
xor (n2149,n2146,n2147);
or (n2150,n2151,n2154);
and (n2151,n2152,n2153);
xor (n2152,n2047,n2048);
and (n2153,n149,n139);
and (n2154,n2155,n2156);
xor (n2155,n2152,n2153);
or (n2156,n2157,n2160);
and (n2157,n2158,n2159);
xor (n2158,n2053,n2054);
and (n2159,n71,n139);
and (n2160,n2161,n2162);
xor (n2161,n2158,n2159);
or (n2162,n2163,n2166);
and (n2163,n2164,n2165);
xor (n2164,n2059,n2060);
and (n2165,n64,n139);
and (n2166,n2167,n2168);
xor (n2167,n2164,n2165);
or (n2168,n2169,n2172);
and (n2169,n2170,n2171);
xor (n2170,n2065,n2066);
and (n2171,n112,n139);
and (n2172,n2173,n2174);
xor (n2173,n2170,n2171);
or (n2174,n2175,n2178);
and (n2175,n2176,n2177);
xor (n2176,n2071,n2072);
and (n2177,n125,n139);
and (n2178,n2179,n2180);
xor (n2179,n2176,n2177);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2077,n2078);
and (n2183,n192,n139);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2083,n2084);
and (n2189,n340,n139);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2089,n2090);
and (n2195,n363,n139);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2095,n2096);
and (n2201,n306,n139);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2101,n2102);
and (n2207,n285,n139);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2107,n2108);
and (n2213,n329,n139);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2113,n2114);
and (n2219,n322,n139);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2118,n2119);
and (n2225,n250,n139);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2123,n2124);
and (n2231,n103,n139);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2128,n2129);
and (n2237,n84,n139);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
and (n2240,n2241,n1035);
xor (n2241,n2133,n2134);
or (n2242,n2243,n2246);
and (n2243,n2244,n2245);
xor (n2244,n2143,n2144);
and (n2245,n154,n52);
and (n2246,n2247,n2248);
xor (n2247,n2244,n2245);
or (n2248,n2249,n2252);
and (n2249,n2250,n2251);
xor (n2250,n2149,n2150);
and (n2251,n149,n52);
and (n2252,n2253,n2254);
xor (n2253,n2250,n2251);
or (n2254,n2255,n2258);
and (n2255,n2256,n2257);
xor (n2256,n2155,n2156);
and (n2257,n71,n52);
and (n2258,n2259,n2260);
xor (n2259,n2256,n2257);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2161,n2162);
and (n2263,n64,n52);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2167,n2168);
and (n2269,n112,n52);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2173,n2174);
and (n2275,n125,n52);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2282);
and (n2279,n2280,n2281);
xor (n2280,n2179,n2180);
and (n2281,n192,n52);
and (n2282,n2283,n2284);
xor (n2283,n2280,n2281);
or (n2284,n2285,n2288);
and (n2285,n2286,n2287);
xor (n2286,n2185,n2186);
and (n2287,n340,n52);
and (n2288,n2289,n2290);
xor (n2289,n2286,n2287);
or (n2290,n2291,n2294);
and (n2291,n2292,n2293);
xor (n2292,n2191,n2192);
and (n2293,n363,n52);
and (n2294,n2295,n2296);
xor (n2295,n2292,n2293);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2197,n2198);
and (n2299,n306,n52);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
or (n2302,n2303,n2306);
and (n2303,n2304,n2305);
xor (n2304,n2203,n2204);
and (n2305,n285,n52);
and (n2306,n2307,n2308);
xor (n2307,n2304,n2305);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2209,n2210);
and (n2311,n329,n52);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2215,n2216);
and (n2317,n322,n52);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
or (n2320,n2321,n2324);
and (n2321,n2322,n2323);
xor (n2322,n2221,n2222);
and (n2323,n250,n52);
and (n2324,n2325,n2326);
xor (n2325,n2322,n2323);
or (n2326,n2327,n2329);
and (n2327,n2328,n973);
xor (n2328,n2227,n2228);
and (n2329,n2330,n2331);
xor (n2330,n2328,n973);
or (n2331,n2332,n2334);
and (n2332,n2333,n1028);
xor (n2333,n2233,n2234);
and (n2334,n2335,n2336);
xor (n2335,n2333,n1028);
and (n2336,n2337,n2338);
xor (n2337,n2239,n2240);
and (n2338,n25,n52);
and (n2339,n154,n50);
or (n2340,n2341,n2344);
and (n2341,n2342,n2343);
xor (n2342,n2247,n2248);
and (n2343,n149,n50);
and (n2344,n2345,n2346);
xor (n2345,n2342,n2343);
or (n2346,n2347,n2350);
and (n2347,n2348,n2349);
xor (n2348,n2253,n2254);
and (n2349,n71,n50);
and (n2350,n2351,n2352);
xor (n2351,n2348,n2349);
or (n2352,n2353,n2356);
and (n2353,n2354,n2355);
xor (n2354,n2259,n2260);
and (n2355,n64,n50);
and (n2356,n2357,n2358);
xor (n2357,n2354,n2355);
or (n2358,n2359,n2362);
and (n2359,n2360,n2361);
xor (n2360,n2265,n2266);
and (n2361,n112,n50);
and (n2362,n2363,n2364);
xor (n2363,n2360,n2361);
or (n2364,n2365,n2368);
and (n2365,n2366,n2367);
xor (n2366,n2271,n2272);
and (n2367,n125,n50);
and (n2368,n2369,n2370);
xor (n2369,n2366,n2367);
or (n2370,n2371,n2374);
and (n2371,n2372,n2373);
xor (n2372,n2277,n2278);
and (n2373,n192,n50);
and (n2374,n2375,n2376);
xor (n2375,n2372,n2373);
or (n2376,n2377,n2380);
and (n2377,n2378,n2379);
xor (n2378,n2283,n2284);
and (n2379,n340,n50);
and (n2380,n2381,n2382);
xor (n2381,n2378,n2379);
or (n2382,n2383,n2386);
and (n2383,n2384,n2385);
xor (n2384,n2289,n2290);
and (n2385,n363,n50);
and (n2386,n2387,n2388);
xor (n2387,n2384,n2385);
or (n2388,n2389,n2392);
and (n2389,n2390,n2391);
xor (n2390,n2295,n2296);
and (n2391,n306,n50);
and (n2392,n2393,n2394);
xor (n2393,n2390,n2391);
or (n2394,n2395,n2398);
and (n2395,n2396,n2397);
xor (n2396,n2301,n2302);
and (n2397,n285,n50);
and (n2398,n2399,n2400);
xor (n2399,n2396,n2397);
or (n2400,n2401,n2404);
and (n2401,n2402,n2403);
xor (n2402,n2307,n2308);
and (n2403,n329,n50);
and (n2404,n2405,n2406);
xor (n2405,n2402,n2403);
or (n2406,n2407,n2410);
and (n2407,n2408,n2409);
xor (n2408,n2313,n2314);
and (n2409,n322,n50);
and (n2410,n2411,n2412);
xor (n2411,n2408,n2409);
or (n2412,n2413,n2416);
and (n2413,n2414,n2415);
xor (n2414,n2319,n2320);
and (n2415,n250,n50);
and (n2416,n2417,n2418);
xor (n2417,n2414,n2415);
or (n2418,n2419,n2422);
and (n2419,n2420,n2421);
xor (n2420,n2325,n2326);
and (n2421,n103,n50);
and (n2422,n2423,n2424);
xor (n2423,n2420,n2421);
or (n2424,n2425,n2428);
and (n2425,n2426,n2427);
xor (n2426,n2330,n2331);
and (n2427,n84,n50);
and (n2428,n2429,n2430);
xor (n2429,n2426,n2427);
and (n2430,n2431,n932);
xor (n2431,n2335,n2336);
or (n2432,n2433,n2435);
and (n2433,n2434,n70);
xor (n2434,n2345,n2346);
and (n2435,n2436,n2437);
xor (n2436,n2434,n70);
or (n2437,n2438,n2440);
and (n2438,n2439,n65);
xor (n2439,n2351,n2352);
and (n2440,n2441,n2442);
xor (n2441,n2439,n65);
or (n2442,n2443,n2445);
and (n2443,n2444,n528);
xor (n2444,n2357,n2358);
and (n2445,n2446,n2447);
xor (n2446,n2444,n528);
or (n2447,n2448,n2451);
and (n2448,n2449,n2450);
xor (n2449,n2363,n2364);
and (n2450,n125,n57);
and (n2451,n2452,n2453);
xor (n2452,n2449,n2450);
or (n2453,n2454,n2457);
and (n2454,n2455,n2456);
xor (n2455,n2369,n2370);
and (n2456,n192,n57);
and (n2457,n2458,n2459);
xor (n2458,n2455,n2456);
or (n2459,n2460,n2463);
and (n2460,n2461,n2462);
xor (n2461,n2375,n2376);
and (n2462,n340,n57);
and (n2463,n2464,n2465);
xor (n2464,n2461,n2462);
or (n2465,n2466,n2469);
and (n2466,n2467,n2468);
xor (n2467,n2381,n2382);
and (n2468,n363,n57);
and (n2469,n2470,n2471);
xor (n2470,n2467,n2468);
or (n2471,n2472,n2474);
and (n2472,n2473,n1189);
xor (n2473,n2387,n2388);
and (n2474,n2475,n2476);
xor (n2475,n2473,n1189);
or (n2476,n2477,n2480);
and (n2477,n2478,n2479);
xor (n2478,n2393,n2394);
and (n2479,n285,n57);
and (n2480,n2481,n2482);
xor (n2481,n2478,n2479);
or (n2482,n2483,n2486);
and (n2483,n2484,n2485);
xor (n2484,n2399,n2400);
and (n2485,n329,n57);
and (n2486,n2487,n2488);
xor (n2487,n2484,n2485);
or (n2488,n2489,n2492);
and (n2489,n2490,n2491);
xor (n2490,n2405,n2406);
and (n2491,n322,n57);
and (n2492,n2493,n2494);
xor (n2493,n2490,n2491);
or (n2494,n2495,n2498);
and (n2495,n2496,n2497);
xor (n2496,n2411,n2412);
and (n2497,n250,n57);
and (n2498,n2499,n2500);
xor (n2499,n2496,n2497);
or (n2500,n2501,n2504);
and (n2501,n2502,n2503);
xor (n2502,n2417,n2418);
and (n2503,n103,n57);
and (n2504,n2505,n2506);
xor (n2505,n2502,n2503);
or (n2506,n2507,n2509);
and (n2507,n2508,n785);
xor (n2508,n2423,n2424);
and (n2509,n2510,n2511);
xor (n2510,n2508,n785);
and (n2511,n2512,n2513);
xor (n2512,n2429,n2430);
and (n2513,n25,n57);
and (n2514,n71,n119);
or (n2515,n2516,n2519);
and (n2516,n2517,n2518);
xor (n2517,n2436,n2437);
and (n2518,n64,n119);
and (n2519,n2520,n2521);
xor (n2520,n2517,n2518);
or (n2521,n2522,n2525);
and (n2522,n2523,n2524);
xor (n2523,n2441,n2442);
and (n2524,n112,n119);
and (n2525,n2526,n2527);
xor (n2526,n2523,n2524);
or (n2527,n2528,n2531);
and (n2528,n2529,n2530);
xor (n2529,n2446,n2447);
and (n2530,n125,n119);
and (n2531,n2532,n2533);
xor (n2532,n2529,n2530);
or (n2533,n2534,n2537);
and (n2534,n2535,n2536);
xor (n2535,n2452,n2453);
and (n2536,n192,n119);
and (n2537,n2538,n2539);
xor (n2538,n2535,n2536);
or (n2539,n2540,n2543);
and (n2540,n2541,n2542);
xor (n2541,n2458,n2459);
and (n2542,n340,n119);
and (n2543,n2544,n2545);
xor (n2544,n2541,n2542);
or (n2545,n2546,n2549);
and (n2546,n2547,n2548);
xor (n2547,n2464,n2465);
and (n2548,n363,n119);
and (n2549,n2550,n2551);
xor (n2550,n2547,n2548);
or (n2551,n2552,n2555);
and (n2552,n2553,n2554);
xor (n2553,n2470,n2471);
and (n2554,n306,n119);
and (n2555,n2556,n2557);
xor (n2556,n2553,n2554);
or (n2557,n2558,n2561);
and (n2558,n2559,n2560);
xor (n2559,n2475,n2476);
and (n2560,n285,n119);
and (n2561,n2562,n2563);
xor (n2562,n2559,n2560);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2481,n2482);
and (n2566,n329,n119);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2487,n2488);
and (n2572,n322,n119);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
or (n2575,n2576,n2579);
and (n2576,n2577,n2578);
xor (n2577,n2493,n2494);
and (n2578,n250,n119);
and (n2579,n2580,n2581);
xor (n2580,n2577,n2578);
or (n2581,n2582,n2585);
and (n2582,n2583,n2584);
xor (n2583,n2499,n2500);
and (n2584,n103,n119);
and (n2585,n2586,n2587);
xor (n2586,n2583,n2584);
or (n2587,n2588,n2591);
and (n2588,n2589,n2590);
xor (n2589,n2505,n2506);
and (n2590,n84,n119);
and (n2591,n2592,n2593);
xor (n2592,n2589,n2590);
and (n2593,n2594,n758);
xor (n2594,n2510,n2511);
and (n2595,n64,n110);
or (n2596,n2597,n2600);
and (n2597,n2598,n2599);
xor (n2598,n2520,n2521);
and (n2599,n112,n110);
and (n2600,n2601,n2602);
xor (n2601,n2598,n2599);
or (n2602,n2603,n2606);
and (n2603,n2604,n2605);
xor (n2604,n2526,n2527);
and (n2605,n125,n110);
and (n2606,n2607,n2608);
xor (n2607,n2604,n2605);
or (n2608,n2609,n2611);
and (n2609,n2610,n589);
xor (n2610,n2532,n2533);
and (n2611,n2612,n2613);
xor (n2612,n2610,n589);
or (n2613,n2614,n2617);
and (n2614,n2615,n2616);
xor (n2615,n2538,n2539);
and (n2616,n340,n110);
and (n2617,n2618,n2619);
xor (n2618,n2615,n2616);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
xor (n2621,n2544,n2545);
and (n2622,n363,n110);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
xor (n2627,n2550,n2551);
and (n2628,n306,n110);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
xor (n2633,n2556,n2557);
and (n2634,n285,n110);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
xor (n2639,n2562,n2563);
and (n2640,n329,n110);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
or (n2643,n2644,n2647);
and (n2644,n2645,n2646);
xor (n2645,n2568,n2569);
and (n2646,n322,n110);
and (n2647,n2648,n2649);
xor (n2648,n2645,n2646);
or (n2649,n2650,n2653);
and (n2650,n2651,n2652);
xor (n2651,n2574,n2575);
and (n2652,n250,n110);
and (n2653,n2654,n2655);
xor (n2654,n2651,n2652);
or (n2655,n2656,n2659);
and (n2656,n2657,n2658);
xor (n2657,n2580,n2581);
and (n2658,n103,n110);
and (n2659,n2660,n2661);
xor (n2660,n2657,n2658);
or (n2661,n2662,n2665);
and (n2662,n2663,n2664);
xor (n2663,n2586,n2587);
and (n2664,n84,n110);
and (n2665,n2666,n2667);
xor (n2666,n2663,n2664);
and (n2667,n2668,n2669);
xor (n2668,n2592,n2593);
and (n2669,n25,n110);
and (n2670,n112,n183);
or (n2671,n2672,n2675);
and (n2672,n2673,n2674);
xor (n2673,n2601,n2602);
and (n2674,n125,n183);
and (n2675,n2676,n2677);
xor (n2676,n2673,n2674);
or (n2677,n2678,n2681);
and (n2678,n2679,n2680);
xor (n2679,n2607,n2608);
and (n2680,n192,n183);
and (n2681,n2682,n2683);
xor (n2682,n2679,n2680);
or (n2683,n2684,n2687);
and (n2684,n2685,n2686);
xor (n2685,n2612,n2613);
and (n2686,n340,n183);
and (n2687,n2688,n2689);
xor (n2688,n2685,n2686);
or (n2689,n2690,n2693);
and (n2690,n2691,n2692);
xor (n2691,n2618,n2619);
and (n2692,n363,n183);
and (n2693,n2694,n2695);
xor (n2694,n2691,n2692);
or (n2695,n2696,n2699);
and (n2696,n2697,n2698);
xor (n2697,n2624,n2625);
and (n2698,n306,n183);
and (n2699,n2700,n2701);
xor (n2700,n2697,n2698);
or (n2701,n2702,n2705);
and (n2702,n2703,n2704);
xor (n2703,n2630,n2631);
and (n2704,n285,n183);
and (n2705,n2706,n2707);
xor (n2706,n2703,n2704);
or (n2707,n2708,n2711);
and (n2708,n2709,n2710);
xor (n2709,n2636,n2637);
and (n2710,n329,n183);
and (n2711,n2712,n2713);
xor (n2712,n2709,n2710);
or (n2713,n2714,n2717);
and (n2714,n2715,n2716);
xor (n2715,n2642,n2643);
and (n2716,n322,n183);
and (n2717,n2718,n2719);
xor (n2718,n2715,n2716);
or (n2719,n2720,n2723);
and (n2720,n2721,n2722);
xor (n2721,n2648,n2649);
and (n2722,n250,n183);
and (n2723,n2724,n2725);
xor (n2724,n2721,n2722);
or (n2725,n2726,n2729);
and (n2726,n2727,n2728);
xor (n2727,n2654,n2655);
and (n2728,n103,n183);
and (n2729,n2730,n2731);
xor (n2730,n2727,n2728);
or (n2731,n2732,n2735);
and (n2732,n2733,n2734);
xor (n2733,n2660,n2661);
and (n2734,n84,n183);
and (n2735,n2736,n2737);
xor (n2736,n2733,n2734);
and (n2737,n2738,n861);
xor (n2738,n2666,n2667);
and (n2739,n125,n188);
or (n2740,n2741,n2744);
and (n2741,n2742,n2743);
xor (n2742,n2676,n2677);
and (n2743,n192,n188);
and (n2744,n2745,n2746);
xor (n2745,n2742,n2743);
or (n2746,n2747,n2750);
and (n2747,n2748,n2749);
xor (n2748,n2682,n2683);
and (n2749,n340,n188);
and (n2750,n2751,n2752);
xor (n2751,n2748,n2749);
or (n2752,n2753,n2756);
and (n2753,n2754,n2755);
xor (n2754,n2688,n2689);
and (n2755,n363,n188);
and (n2756,n2757,n2758);
xor (n2757,n2754,n2755);
or (n2758,n2759,n2762);
and (n2759,n2760,n2761);
xor (n2760,n2694,n2695);
and (n2761,n306,n188);
and (n2762,n2763,n2764);
xor (n2763,n2760,n2761);
or (n2764,n2765,n2768);
and (n2765,n2766,n2767);
xor (n2766,n2700,n2701);
and (n2767,n285,n188);
and (n2768,n2769,n2770);
xor (n2769,n2766,n2767);
or (n2770,n2771,n2774);
and (n2771,n2772,n2773);
xor (n2772,n2706,n2707);
and (n2773,n329,n188);
and (n2774,n2775,n2776);
xor (n2775,n2772,n2773);
or (n2776,n2777,n2780);
and (n2777,n2778,n2779);
xor (n2778,n2712,n2713);
and (n2779,n322,n188);
and (n2780,n2781,n2782);
xor (n2781,n2778,n2779);
or (n2782,n2783,n2786);
and (n2783,n2784,n2785);
xor (n2784,n2718,n2719);
and (n2785,n250,n188);
and (n2786,n2787,n2788);
xor (n2787,n2784,n2785);
or (n2788,n2789,n2792);
and (n2789,n2790,n2791);
xor (n2790,n2724,n2725);
and (n2791,n103,n188);
and (n2792,n2793,n2794);
xor (n2793,n2790,n2791);
or (n2794,n2795,n2798);
and (n2795,n2796,n2797);
xor (n2796,n2730,n2731);
and (n2797,n84,n188);
and (n2798,n2799,n2800);
xor (n2799,n2796,n2797);
and (n2800,n2801,n2802);
xor (n2801,n2736,n2737);
and (n2802,n25,n188);
and (n2803,n192,n350);
or (n2804,n2805,n2808);
and (n2805,n2806,n2807);
xor (n2806,n2745,n2746);
and (n2807,n340,n350);
and (n2808,n2809,n2810);
xor (n2809,n2806,n2807);
or (n2810,n2811,n2814);
and (n2811,n2812,n2813);
xor (n2812,n2751,n2752);
and (n2813,n363,n350);
and (n2814,n2815,n2816);
xor (n2815,n2812,n2813);
or (n2816,n2817,n2820);
and (n2817,n2818,n2819);
xor (n2818,n2757,n2758);
and (n2819,n306,n350);
and (n2820,n2821,n2822);
xor (n2821,n2818,n2819);
or (n2822,n2823,n2826);
and (n2823,n2824,n2825);
xor (n2824,n2763,n2764);
and (n2825,n285,n350);
and (n2826,n2827,n2828);
xor (n2827,n2824,n2825);
or (n2828,n2829,n2832);
and (n2829,n2830,n2831);
xor (n2830,n2769,n2770);
and (n2831,n329,n350);
and (n2832,n2833,n2834);
xor (n2833,n2830,n2831);
or (n2834,n2835,n2838);
and (n2835,n2836,n2837);
xor (n2836,n2775,n2776);
and (n2837,n322,n350);
and (n2838,n2839,n2840);
xor (n2839,n2836,n2837);
or (n2840,n2841,n2844);
and (n2841,n2842,n2843);
xor (n2842,n2781,n2782);
and (n2843,n250,n350);
and (n2844,n2845,n2846);
xor (n2845,n2842,n2843);
or (n2846,n2847,n2850);
and (n2847,n2848,n2849);
xor (n2848,n2787,n2788);
and (n2849,n103,n350);
and (n2850,n2851,n2852);
xor (n2851,n2848,n2849);
or (n2852,n2853,n2856);
and (n2853,n2854,n2855);
xor (n2854,n2793,n2794);
and (n2855,n84,n350);
and (n2856,n2857,n2858);
xor (n2857,n2854,n2855);
and (n2858,n2859,n2860);
xor (n2859,n2799,n2800);
not (n2860,n1292);
and (n2861,n340,n294);
or (n2862,n2863,n2866);
and (n2863,n2864,n2865);
xor (n2864,n2809,n2810);
and (n2865,n363,n294);
and (n2866,n2867,n2868);
xor (n2867,n2864,n2865);
or (n2868,n2869,n2872);
and (n2869,n2870,n2871);
xor (n2870,n2815,n2816);
and (n2871,n306,n294);
and (n2872,n2873,n2874);
xor (n2873,n2870,n2871);
or (n2874,n2875,n2878);
and (n2875,n2876,n2877);
xor (n2876,n2821,n2822);
and (n2877,n285,n294);
and (n2878,n2879,n2880);
xor (n2879,n2876,n2877);
or (n2880,n2881,n2884);
and (n2881,n2882,n2883);
xor (n2882,n2827,n2828);
and (n2883,n329,n294);
and (n2884,n2885,n2886);
xor (n2885,n2882,n2883);
or (n2886,n2887,n2890);
and (n2887,n2888,n2889);
xor (n2888,n2833,n2834);
and (n2889,n322,n294);
and (n2890,n2891,n2892);
xor (n2891,n2888,n2889);
or (n2892,n2893,n2896);
and (n2893,n2894,n2895);
xor (n2894,n2839,n2840);
and (n2895,n250,n294);
and (n2896,n2897,n2898);
xor (n2897,n2894,n2895);
or (n2898,n2899,n2902);
and (n2899,n2900,n2901);
xor (n2900,n2845,n2846);
and (n2901,n103,n294);
and (n2902,n2903,n2904);
xor (n2903,n2900,n2901);
or (n2904,n2905,n2908);
and (n2905,n2906,n2907);
xor (n2906,n2851,n2852);
and (n2907,n84,n294);
and (n2908,n2909,n2910);
xor (n2909,n2906,n2907);
and (n2910,n2911,n2912);
xor (n2911,n2857,n2858);
and (n2912,n25,n294);
and (n2913,n363,n295);
or (n2914,n2915,n2918);
and (n2915,n2916,n2917);
xor (n2916,n2867,n2868);
and (n2917,n306,n295);
and (n2918,n2919,n2920);
xor (n2919,n2916,n2917);
or (n2920,n2921,n2924);
and (n2921,n2922,n2923);
xor (n2922,n2873,n2874);
and (n2923,n285,n295);
and (n2924,n2925,n2926);
xor (n2925,n2922,n2923);
or (n2926,n2927,n2930);
and (n2927,n2928,n2929);
xor (n2928,n2879,n2880);
and (n2929,n329,n295);
and (n2930,n2931,n2932);
xor (n2931,n2928,n2929);
or (n2932,n2933,n2936);
and (n2933,n2934,n2935);
xor (n2934,n2885,n2886);
and (n2935,n322,n295);
and (n2936,n2937,n2938);
xor (n2937,n2934,n2935);
or (n2938,n2939,n2942);
and (n2939,n2940,n2941);
xor (n2940,n2891,n2892);
and (n2941,n250,n295);
and (n2942,n2943,n2944);
xor (n2943,n2940,n2941);
or (n2944,n2945,n2948);
and (n2945,n2946,n2947);
xor (n2946,n2897,n2898);
and (n2947,n103,n295);
and (n2948,n2949,n2950);
xor (n2949,n2946,n2947);
or (n2950,n2951,n2954);
and (n2951,n2952,n2953);
xor (n2952,n2903,n2904);
and (n2953,n84,n295);
and (n2954,n2955,n2956);
xor (n2955,n2952,n2953);
and (n2956,n2957,n2958);
xor (n2957,n2909,n2910);
not (n2958,n1453);
and (n2959,n306,n286);
or (n2960,n2961,n2964);
and (n2961,n2962,n2963);
xor (n2962,n2919,n2920);
and (n2963,n285,n286);
and (n2964,n2965,n2966);
xor (n2965,n2962,n2963);
or (n2966,n2967,n2969);
and (n2967,n2968,n498);
xor (n2968,n2925,n2926);
and (n2969,n2970,n2971);
xor (n2970,n2968,n498);
or (n2971,n2972,n2975);
and (n2972,n2973,n2974);
xor (n2973,n2931,n2932);
and (n2974,n322,n286);
and (n2975,n2976,n2977);
xor (n2976,n2973,n2974);
or (n2977,n2978,n2981);
and (n2978,n2979,n2980);
xor (n2979,n2937,n2938);
and (n2980,n250,n286);
and (n2981,n2982,n2983);
xor (n2982,n2979,n2980);
or (n2983,n2984,n2987);
and (n2984,n2985,n2986);
xor (n2985,n2943,n2944);
and (n2986,n103,n286);
and (n2987,n2988,n2989);
xor (n2988,n2985,n2986);
or (n2989,n2990,n2993);
and (n2990,n2991,n2992);
xor (n2991,n2949,n2950);
and (n2992,n84,n286);
and (n2993,n2994,n2995);
xor (n2994,n2991,n2992);
and (n2995,n2996,n2997);
xor (n2996,n2955,n2956);
and (n2997,n25,n286);
and (n2998,n285,n314);
or (n2999,n3000,n3003);
and (n3000,n3001,n3002);
xor (n3001,n2965,n2966);
and (n3002,n329,n314);
and (n3003,n3004,n3005);
xor (n3004,n3001,n3002);
or (n3005,n3006,n3009);
and (n3006,n3007,n3008);
xor (n3007,n2970,n2971);
and (n3008,n322,n314);
and (n3009,n3010,n3011);
xor (n3010,n3007,n3008);
or (n3011,n3012,n3015);
and (n3012,n3013,n3014);
xor (n3013,n2976,n2977);
and (n3014,n250,n314);
and (n3015,n3016,n3017);
xor (n3016,n3013,n3014);
or (n3017,n3018,n3021);
and (n3018,n3019,n3020);
xor (n3019,n2982,n2983);
and (n3020,n103,n314);
and (n3021,n3022,n3023);
xor (n3022,n3019,n3020);
or (n3023,n3024,n3027);
and (n3024,n3025,n3026);
xor (n3025,n2988,n2989);
and (n3026,n84,n314);
and (n3027,n3028,n3029);
xor (n3028,n3025,n3026);
and (n3029,n3030,n3031);
xor (n3030,n2994,n2995);
not (n3031,n1502);
and (n3032,n329,n92);
or (n3033,n3034,n3037);
and (n3034,n3035,n3036);
xor (n3035,n3004,n3005);
and (n3036,n322,n92);
and (n3037,n3038,n3039);
xor (n3038,n3035,n3036);
or (n3039,n3040,n3043);
and (n3040,n3041,n3042);
xor (n3041,n3010,n3011);
and (n3042,n250,n92);
and (n3043,n3044,n3045);
xor (n3044,n3041,n3042);
or (n3045,n3046,n3049);
and (n3046,n3047,n3048);
xor (n3047,n3016,n3017);
and (n3048,n103,n92);
and (n3049,n3050,n3051);
xor (n3050,n3047,n3048);
or (n3051,n3052,n3055);
and (n3052,n3053,n3054);
xor (n3053,n3022,n3023);
and (n3054,n84,n92);
and (n3055,n3056,n3057);
xor (n3056,n3053,n3054);
and (n3057,n3058,n3059);
xor (n3058,n3028,n3029);
and (n3059,n25,n92);
and (n3060,n322,n90);
or (n3061,n3062,n3065);
and (n3062,n3063,n3064);
xor (n3063,n3038,n3039);
and (n3064,n250,n90);
and (n3065,n3066,n3067);
xor (n3066,n3063,n3064);
or (n3067,n3068,n3071);
and (n3068,n3069,n3070);
xor (n3069,n3044,n3045);
and (n3070,n103,n90);
and (n3071,n3072,n3073);
xor (n3072,n3069,n3070);
or (n3073,n3074,n3077);
and (n3074,n3075,n3076);
xor (n3075,n3050,n3051);
and (n3076,n84,n90);
and (n3077,n3078,n3079);
xor (n3078,n3075,n3076);
and (n3079,n3080,n3081);
xor (n3080,n3056,n3057);
not (n3081,n370);
or (n3082,n3083,n3086);
and (n3083,n3084,n3085);
xor (n3084,n3066,n3067);
and (n3085,n103,n22);
and (n3086,n3087,n3088);
xor (n3087,n3084,n3085);
or (n3088,n3089,n3092);
and (n3089,n3090,n3091);
xor (n3090,n3072,n3073);
and (n3091,n84,n22);
and (n3092,n3093,n3094);
xor (n3093,n3090,n3091);
and (n3094,n3095,n3096);
xor (n3095,n3078,n3079);
and (n3096,n25,n22);
and (n3097,n103,n21);
or (n3098,n3099,n3102);
and (n3099,n3100,n3101);
xor (n3100,n3087,n3088);
and (n3101,n84,n21);
and (n3102,n3103,n3104);
xor (n3103,n3100,n3101);
and (n3104,n3105,n208);
xor (n3105,n3093,n3094);
and (n3106,n84,n209);
and (n3107,n3108,n3109);
xor (n3108,n3103,n3104);
and (n3109,n25,n209);
not (n3110,n3111);
nand (n3111,n25,n465);
endmodule
