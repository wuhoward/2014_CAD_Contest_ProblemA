module top (out,n20,n21,n25,n27,n29,n30,n31,n34,n35
        ,n36,n42,n43,n44,n52,n53,n57,n59,n61,n62
        ,n65,n67,n69,n71,n72,n73,n74,n75,n76,n77
        ,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87
        ,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97
        ,n98,n99,n106,n107,n108,n119,n120,n121,n127,n128
        ,n129,n138,n139,n140,n147,n148,n149,n160,n161,n162
        ,n166,n167,n168,n176,n177,n178,n190,n191,n192,n201
        ,n202,n203,n209,n210,n211,n220,n221,n222,n226,n227
        ,n228,n236,n237,n238,n242,n243,n244,n254,n255,n256
        ,n267,n268,n269,n278,n279,n280,n283,n284,n285,n293
        ,n294,n295,n312,n313,n314,n325,n326,n327,n334,n335
        ,n336,n346,n347,n348,n357,n358,n359,n366,n367,n368
        ,n375,n376,n377,n386,n387,n388,n396,n397,n398,n405
        ,n406,n407,n1241,n1242,n1246,n1248,n1250,n1253,n1254,n1258
        ,n1260,n1262,n1263,n1266,n1268,n1270,n1272,n1273,n1274,n1275
        ,n1276,n1277,n1278,n1279,n1280,n1281,n1282,n1283,n1284,n1285
        ,n1286,n1287,n1288,n1289,n1290,n1291,n1292,n1293,n1294,n1295
        ,n1296,n1297,n1298,n1299,n1300,n1303,n1304,n1307,n1308,n1309);
output out;
input n20;
input n21;
input n25;
input n27;
input n29;
input n30;
input n31;
input n34;
input n35;
input n36;
input n42;
input n43;
input n44;
input n52;
input n53;
input n57;
input n59;
input n61;
input n62;
input n65;
input n67;
input n69;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n81;
input n82;
input n83;
input n84;
input n85;
input n86;
input n87;
input n88;
input n89;
input n90;
input n91;
input n92;
input n93;
input n94;
input n95;
input n96;
input n97;
input n98;
input n99;
input n106;
input n107;
input n108;
input n119;
input n120;
input n121;
input n127;
input n128;
input n129;
input n138;
input n139;
input n140;
input n147;
input n148;
input n149;
input n160;
input n161;
input n162;
input n166;
input n167;
input n168;
input n176;
input n177;
input n178;
input n190;
input n191;
input n192;
input n201;
input n202;
input n203;
input n209;
input n210;
input n211;
input n220;
input n221;
input n222;
input n226;
input n227;
input n228;
input n236;
input n237;
input n238;
input n242;
input n243;
input n244;
input n254;
input n255;
input n256;
input n267;
input n268;
input n269;
input n278;
input n279;
input n280;
input n283;
input n284;
input n285;
input n293;
input n294;
input n295;
input n312;
input n313;
input n314;
input n325;
input n326;
input n327;
input n334;
input n335;
input n336;
input n346;
input n347;
input n348;
input n357;
input n358;
input n359;
input n366;
input n367;
input n368;
input n375;
input n376;
input n377;
input n386;
input n387;
input n388;
input n396;
input n397;
input n398;
input n405;
input n406;
input n407;
input n1241;
input n1242;
input n1246;
input n1248;
input n1250;
input n1253;
input n1254;
input n1258;
input n1260;
input n1262;
input n1263;
input n1266;
input n1268;
input n1270;
input n1272;
input n1273;
input n1274;
input n1275;
input n1276;
input n1277;
input n1278;
input n1279;
input n1280;
input n1281;
input n1282;
input n1283;
input n1284;
input n1285;
input n1286;
input n1287;
input n1288;
input n1289;
input n1290;
input n1291;
input n1292;
input n1293;
input n1294;
input n1295;
input n1296;
input n1297;
input n1298;
input n1299;
input n1300;
input n1303;
input n1304;
input n1307;
input n1308;
input n1309;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n32;
wire n33;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n58;
wire n60;
wire n63;
wire n64;
wire n66;
wire n68;
wire n70;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n163;
wire n164;
wire n165;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n223;
wire n224;
wire n225;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n239;
wire n240;
wire n241;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n281;
wire n282;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1243;
wire n1244;
wire n1245;
wire n1247;
wire n1249;
wire n1251;
wire n1252;
wire n1255;
wire n1256;
wire n1257;
wire n1259;
wire n1261;
wire n1264;
wire n1265;
wire n1267;
wire n1269;
wire n1271;
wire n1301;
wire n1302;
wire n1305;
wire n1306;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
xnor (out,n0,n1314);
nand (n0,n1,n1232);
nand (n1,n2,n1231);
or (n2,n3,n699);
nand (n3,n4,n698);
nand (n4,n5,n635);
not (n5,n6);
xor (n6,n7,n588);
xor (n7,n8,n411);
xor (n8,n9,n302);
xor (n9,n10,n194);
xor (n10,n11,n152);
xor (n11,n12,n110);
nand (n12,n13,n101);
or (n13,n14,n47);
not (n14,n15);
nor (n15,n16,n37);
not (n16,n17);
xnor (n17,n18,n32);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n31);
and (s0n18,notn18,n19);
and (s1n18,n31,n30);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,n20);
and (s1n19,n22,n21);
and (n22,n23,n28);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
not (n28,n29);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n31);
and (s0n32,notn32,n33);
and (s1n32,n31,n36);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n22);
and (s0n33,notn33,n34);
and (s1n33,n22,n35);
nor (n37,n38,n45);
and (n38,n39,n40);
not (n39,n32);
wire s0n40,s1n40,notn40;
or (n40,s0n40,s1n40);
not(notn40,n31);
and (s0n40,notn40,n41);
and (s1n40,n31,n44);
wire s0n41,s1n41,notn41;
or (n41,s0n41,s1n41);
not(notn41,n22);
and (s0n41,notn41,n42);
and (s1n41,n22,n43);
and (n45,n32,n46);
not (n46,n40);
not (n47,n48);
nand (n48,n49,n100);
or (n49,n46,n50);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n63);
and (s0n50,notn50,n51);
and (s1n50,n63,n62);
wire s0n51,s1n51,notn51;
or (n51,s0n51,s1n51);
not(notn51,n54);
and (s0n51,notn51,n52);
and (s1n51,n54,n53);
and (n54,n55,n60);
and (n55,n56,n58);
not (n56,n57);
not (n58,n59);
not (n60,n61);
and (n63,n64,n66);
not (n64,n65);
or (n66,n67,n68);
and (n68,n69,n70);
or (n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99);
nand (n100,n50,n46);
nand (n101,n102,n16);
nand (n102,n103,n109);
or (n103,n46,n104);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n63);
and (s0n104,notn104,n105);
and (s1n104,n63,n108);
wire s0n105,s1n105,notn105;
or (n105,s0n105,s1n105);
not(notn105,n54);
and (s0n105,notn105,n106);
and (s1n105,n54,n107);
nand (n109,n104,n46);
nand (n110,n111,n142);
or (n111,n112,n132);
not (n112,n113);
and (n113,n114,n123);
nand (n114,n115,n122);
or (n115,n116,n18);
not (n116,n117);
wire s0n117,s1n117,notn117;
or (n117,s0n117,s1n117);
not(notn117,n31);
and (s0n117,notn117,n118);
and (s1n117,n31,n121);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n22);
and (s0n118,notn118,n119);
and (s1n118,n22,n120);
nand (n122,n18,n116);
nor (n123,n124,n130);
and (n124,n125,n116);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n31);
and (s0n125,notn125,n126);
and (s1n125,n31,n129);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n22);
and (s0n126,notn126,n127);
and (s1n126,n22,n128);
and (n130,n131,n117);
not (n131,n125);
not (n132,n133);
nand (n133,n134,n141);
or (n134,n135,n136);
not (n135,n18);
wire s0n136,s1n136,notn136;
or (n136,s0n136,s1n136);
not(notn136,n63);
and (s0n136,notn136,n137);
and (s1n136,n63,n140);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n54);
and (s0n137,notn137,n138);
and (s1n137,n54,n139);
nand (n141,n136,n135);
nand (n142,n143,n151);
nand (n143,n144,n150);
or (n144,n135,n145);
wire s0n145,s1n145,notn145;
or (n145,s0n145,s1n145);
not(notn145,n63);
and (s0n145,notn145,n146);
and (s1n145,n63,n149);
wire s0n146,s1n146,notn146;
or (n146,s0n146,s1n146);
not(notn146,n54);
and (s0n146,notn146,n147);
and (s1n146,n54,n148);
nand (n150,n145,n135);
not (n151,n123);
nand (n152,n153,n180);
or (n153,n154,n170);
not (n154,n155);
nor (n155,n156,n169);
and (n156,n157,n163);
not (n157,n158);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n31);
and (s0n158,notn158,n159);
and (s1n158,n31,n162);
wire s0n159,s1n159,notn159;
or (n159,s0n159,s1n159);
not(notn159,n22);
and (s0n159,notn159,n160);
and (s1n159,n22,n161);
not (n163,n164);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n63);
and (s0n164,notn164,n165);
and (s1n164,n63,n168);
wire s0n165,s1n165,notn165;
or (n165,s0n165,s1n165);
not(notn165,n54);
and (s0n165,notn165,n166);
and (s1n165,n54,n167);
and (n169,n164,n158);
not (n170,n171);
nand (n171,n172,n179);
or (n172,n173,n40);
not (n173,n174);
wire s0n174,s1n174,notn174;
or (n174,s0n174,s1n174);
not(notn174,n31);
and (s0n174,notn174,n175);
and (s1n174,n31,n178);
wire s0n175,s1n175,notn175;
or (n175,s0n175,s1n175);
not(notn175,n22);
and (s0n175,notn175,n176);
and (s1n175,n22,n177);
nand (n179,n173,n40);
or (n180,n181,n185);
nand (n181,n170,n182);
nor (n182,n183,n184);
and (n183,n174,n158);
and (n184,n173,n157);
nor (n185,n186,n193);
and (n186,n158,n187);
not (n187,n188);
wire s0n188,s1n188,notn188;
or (n188,s0n188,s1n188);
not(notn188,n63);
and (s0n188,notn188,n189);
and (s1n188,n63,n192);
wire s0n189,s1n189,notn189;
or (n189,s0n189,s1n189);
not(notn189,n54);
and (s0n189,notn189,n190);
and (s1n189,n54,n191);
and (n193,n157,n188);
xor (n194,n195,n259);
xor (n195,n196,n212);
nor (n196,n197,n206);
nor (n197,n198,n204);
and (n198,n199,n157);
wire s0n199,s1n199,notn199;
or (n199,s0n199,s1n199);
not(notn199,n31);
and (s0n199,notn199,n200);
and (s1n199,n31,n203);
wire s0n200,s1n200,notn200;
or (n200,s0n200,s1n200);
not(notn200,n22);
and (s0n200,notn200,n201);
and (s1n200,n22,n202);
and (n204,n205,n158);
not (n205,n199);
not (n206,n207);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n63);
and (s0n207,notn207,n208);
and (s1n207,n63,n211);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n54);
and (s0n208,notn208,n209);
and (s1n208,n54,n210);
nand (n212,n213,n249);
or (n213,n214,n230);
not (n214,n215);
nor (n215,n216,n229);
and (n216,n217,n223);
not (n217,n218);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n31);
and (s0n218,notn218,n219);
and (s1n218,n31,n222);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n22);
and (s0n219,notn219,n220);
and (s1n219,n22,n221);
not (n223,n224);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n63);
and (s0n224,notn224,n225);
and (s1n224,n63,n228);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n54);
and (s0n225,notn225,n226);
and (s1n225,n54,n227);
and (n229,n224,n218);
nand (n230,n231,n246);
not (n231,n232);
nand (n232,n233,n245);
or (n233,n234,n239);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n31);
and (s0n234,notn234,n235);
and (s1n234,n31,n238);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n22);
and (s0n235,notn235,n236);
and (s1n235,n22,n237);
not (n239,n240);
wire s0n240,s1n240,notn240;
or (n240,s0n240,s1n240);
not(notn240,n31);
and (s0n240,notn240,n241);
and (s1n240,n31,n244);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n22);
and (s0n241,notn241,n242);
and (s1n241,n22,n243);
nand (n245,n239,n234);
nand (n246,n247,n248);
or (n247,n239,n218);
nand (n248,n218,n239);
nand (n249,n250,n232);
nor (n250,n251,n257);
and (n251,n252,n218);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n63);
and (s0n252,notn252,n253);
and (s1n252,n63,n256);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n54);
and (s0n253,notn253,n254);
and (s1n253,n54,n255);
and (n257,n217,n258);
not (n258,n252);
nand (n259,n260,n287);
or (n260,n261,n272);
not (n261,n262);
nand (n262,n263,n270);
or (n263,n264,n234);
not (n264,n265);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n63);
and (s0n265,notn265,n266);
and (s1n265,n63,n269);
wire s0n266,s1n266,notn266;
or (n266,s0n266,s1n266);
not(notn266,n54);
and (s0n266,notn266,n267);
and (s1n266,n54,n268);
or (n270,n265,n271);
not (n271,n234);
not (n272,n273);
nand (n273,n274,n286);
or (n274,n275,n281);
not (n275,n276);
wire s0n276,s1n276,notn276;
or (n276,s0n276,s1n276);
not(notn276,n31);
and (s0n276,notn276,n277);
and (s1n276,n31,n280);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n22);
and (s0n277,notn277,n278);
and (s1n277,n22,n279);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n31);
and (s0n281,notn281,n282);
and (s1n281,n31,n285);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n22);
and (s0n282,notn282,n283);
and (s1n282,n22,n284);
nand (n286,n281,n275);
nand (n287,n288,n297);
nor (n288,n289,n296);
and (n289,n271,n290);
not (n290,n291);
wire s0n291,s1n291,notn291;
or (n291,s0n291,s1n291);
not(notn291,n63);
and (s0n291,notn291,n292);
and (s1n291,n63,n295);
wire s0n292,s1n292,notn292;
or (n292,s0n292,s1n292);
not(notn292,n54);
and (s0n292,notn292,n293);
and (s1n292,n54,n294);
and (n296,n291,n234);
nor (n297,n273,n298);
not (n298,n299);
nand (n299,n300,n301);
or (n300,n234,n275);
nand (n301,n275,n234);
xor (n302,n303,n380);
xor (n303,n304,n338);
nand (n304,n305,n329);
or (n305,n306,n320);
not (n306,n307);
nor (n307,n308,n317);
nor (n308,n309,n315);
and (n309,n131,n310);
wire s0n310,s1n310,notn310;
or (n310,s0n310,s1n310);
not(notn310,n31);
and (s0n310,notn310,n311);
and (s1n310,n31,n314);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n22);
and (s0n311,notn311,n312);
and (s1n311,n22,n313);
and (n315,n125,n316);
not (n316,n310);
nand (n317,n318,n319);
or (n318,n316,n218);
nand (n319,n218,n316);
not (n320,n321);
nand (n321,n322,n328);
or (n322,n131,n323);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n63);
and (s0n323,notn323,n324);
and (s1n323,n63,n327);
wire s0n324,s1n324,notn324;
or (n324,s0n324,s1n324);
not(notn324,n54);
and (s0n324,notn324,n325);
and (s1n324,n54,n326);
nand (n328,n323,n131);
nand (n329,n330,n317);
nand (n330,n331,n337);
or (n331,n131,n332);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n63);
and (s0n332,notn332,n333);
and (s1n332,n63,n336);
wire s0n333,s1n333,notn333;
or (n333,s0n333,s1n333);
not(notn333,n54);
and (s0n333,notn333,n334);
and (s1n333,n54,n335);
nand (n337,n332,n131);
nand (n338,n339,n370);
or (n339,n340,n351);
not (n340,n341);
nand (n341,n342,n349);
or (n342,n281,n343);
not (n343,n344);
wire s0n344,s1n344,notn344;
or (n344,s0n344,s1n344);
not(notn344,n63);
and (s0n344,notn344,n345);
and (s1n344,n63,n348);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n54);
and (s0n345,notn345,n346);
and (s1n345,n54,n347);
or (n349,n344,n350);
not (n350,n281);
not (n351,n352);
nor (n352,n353,n362);
nor (n353,n354,n360);
and (n354,n350,n355);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n31);
and (s0n355,notn355,n356);
and (s1n355,n31,n359);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n22);
and (s0n356,notn356,n357);
and (s1n356,n22,n358);
and (n360,n281,n361);
not (n361,n355);
nand (n362,n363,n369);
or (n363,n364,n361);
wire s0n364,s1n364,notn364;
or (n364,s0n364,s1n364);
not(notn364,n31);
and (s0n364,notn364,n365);
and (s1n364,n31,n368);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n22);
and (s0n365,notn365,n366);
and (s1n365,n22,n367);
nand (n369,n361,n364);
nand (n370,n362,n371);
nor (n371,n372,n378);
and (n372,n373,n281);
wire s0n373,s1n373,notn373;
or (n373,s0n373,s1n373);
not(notn373,n63);
and (s0n373,notn373,n374);
and (s1n373,n63,n377);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n54);
and (s0n374,notn374,n375);
and (s1n374,n54,n376);
and (n378,n350,n379);
not (n379,n373);
nand (n380,n381,n400);
or (n381,n382,n390);
not (n382,n383);
nor (n383,n384,n389);
wire s0n384,s1n384,notn384;
or (n384,s0n384,s1n384);
not(notn384,n31);
and (s0n384,notn384,n385);
and (s1n384,n31,n388);
wire s0n385,s1n385,notn385;
or (n385,s0n385,s1n385);
not(notn385,n22);
and (s0n385,notn385,n386);
and (s1n385,n22,n387);
not (n389,n364);
not (n390,n391);
nand (n391,n392,n399);
or (n392,n364,n393);
not (n393,n394);
wire s0n394,s1n394,notn394;
or (n394,s0n394,s1n394);
not(notn394,n63);
and (s0n394,notn394,n395);
and (s1n394,n63,n398);
wire s0n395,s1n395,notn395;
or (n395,s0n395,s1n395);
not(notn395,n54);
and (s0n395,notn395,n396);
and (s1n395,n54,n397);
nand (n399,n393,n364);
or (n400,n401,n410);
nor (n401,n402,n408);
and (n402,n403,n389);
wire s0n403,s1n403,notn403;
or (n403,s0n403,s1n403);
not(notn403,n63);
and (s0n403,notn403,n404);
and (s1n403,n63,n407);
wire s0n404,s1n404,notn404;
or (n404,s0n404,s1n404);
not(notn404,n54);
and (s0n404,notn404,n405);
and (s1n404,n54,n406);
and (n408,n409,n364);
not (n409,n403);
not (n410,n384);
or (n411,n412,n587);
and (n412,n413,n516);
xor (n413,n414,n456);
or (n414,n415,n455);
and (n415,n416,n437);
xor (n416,n417,n427);
nand (n417,n418,n423);
or (n418,n419,n14);
not (n419,n420);
nand (n420,n421,n422);
or (n421,n46,n188);
nand (n422,n188,n46);
nand (n423,n424,n16);
nand (n424,n425,n426);
or (n425,n46,n164);
nand (n426,n164,n46);
nand (n427,n428,n433);
or (n428,n429,n351);
not (n429,n430);
nand (n430,n431,n432);
or (n431,n281,n290);
nand (n432,n281,n290);
nand (n433,n362,n434);
nor (n434,n435,n436);
and (n435,n350,n264);
and (n436,n265,n281);
and (n437,n438,n444);
nor (n438,n439,n46);
and (n439,n440,n443);
nand (n440,n441,n135);
not (n441,n442);
and (n442,n207,n32);
nand (n443,n206,n39);
nand (n444,n445,n450);
or (n445,n446,n230);
not (n446,n447);
nand (n447,n448,n449);
or (n448,n217,n145);
nand (n449,n145,n217);
nand (n450,n451,n232);
nand (n451,n452,n454);
or (n452,n218,n453);
not (n453,n323);
nand (n454,n453,n218);
and (n455,n417,n427);
xor (n456,n457,n480);
xor (n457,n458,n466);
nand (n458,n459,n464);
or (n459,n181,n460);
not (n460,n461);
nor (n461,n462,n463);
and (n462,n157,n206);
and (n463,n207,n158);
nand (n464,n465,n171);
not (n465,n185);
xor (n466,n467,n473);
nor (n467,n468,n157);
and (n468,n469,n472);
nand (n469,n470,n46);
not (n470,n471);
and (n471,n207,n174);
nand (n472,n206,n173);
nand (n473,n474,n479);
or (n474,n475,n230);
not (n475,n476);
nand (n476,n477,n478);
or (n477,n217,n332);
nand (n478,n332,n217);
nand (n479,n215,n232);
or (n480,n481,n515);
and (n481,n482,n504);
xor (n482,n483,n494);
nand (n483,n484,n490);
or (n484,n485,n489);
not (n485,n486);
nand (n486,n487,n488);
or (n487,n234,n223);
nand (n488,n223,n234);
not (n489,n297);
nand (n490,n491,n273);
nand (n491,n492,n493);
or (n492,n234,n258);
nand (n493,n258,n234);
nand (n494,n495,n500);
or (n495,n306,n496);
not (n496,n497);
nand (n497,n498,n499);
or (n498,n131,n136);
nand (n499,n136,n131);
nand (n500,n501,n317);
nand (n501,n502,n503);
or (n502,n131,n145);
nand (n503,n145,n131);
nand (n504,n505,n510);
or (n505,n123,n506);
not (n506,n507);
nand (n507,n508,n509);
or (n508,n135,n104);
nand (n509,n104,n135);
nand (n510,n113,n511);
nor (n511,n512,n513);
and (n512,n18,n50);
and (n513,n135,n514);
not (n514,n50);
and (n515,n483,n494);
or (n516,n517,n586);
and (n517,n518,n572);
xor (n518,n519,n544);
or (n519,n520,n543);
and (n520,n521,n536);
xor (n521,n522,n529);
nand (n522,n523,n528);
or (n523,n524,n112);
not (n524,n525);
nand (n525,n526,n527);
or (n526,n135,n164);
nand (n527,n164,n135);
nand (n528,n511,n151);
nand (n529,n530,n535);
or (n530,n531,n14);
not (n531,n532);
nand (n532,n533,n534);
or (n533,n46,n207);
nand (n534,n207,n46);
nand (n535,n420,n16);
nand (n536,n537,n542);
or (n537,n538,n351);
not (n538,n539);
nand (n539,n540,n541);
or (n540,n281,n258);
nand (n541,n258,n281);
nand (n542,n430,n362);
and (n543,n522,n529);
or (n544,n545,n571);
and (n545,n546,n564);
xor (n546,n547,n557);
nand (n547,n548,n553);
or (n548,n549,n382);
not (n549,n550);
nand (n550,n551,n552);
or (n551,n389,n265);
nand (n552,n265,n389);
nand (n553,n554,n384);
nand (n554,n555,n556);
or (n555,n364,n343);
nand (n556,n343,n364);
nand (n557,n558,n563);
or (n558,n559,n489);
not (n559,n560);
nand (n560,n561,n562);
or (n561,n271,n332);
nand (n562,n332,n271);
nand (n563,n273,n486);
nand (n564,n565,n570);
or (n565,n306,n566);
not (n566,n567);
nand (n567,n568,n569);
or (n568,n131,n104);
nand (n569,n104,n131);
nand (n570,n497,n317);
and (n571,n547,n557);
xor (n572,n573,n579);
xor (n573,n574,n575);
and (n574,n171,n207);
nand (n575,n576,n578);
or (n576,n577,n230);
not (n577,n451);
nand (n578,n476,n232);
nand (n579,n580,n582);
or (n580,n581,n382);
not (n581,n554);
nand (n582,n583,n384);
nand (n583,n584,n585);
or (n584,n364,n379);
nand (n585,n379,n364);
and (n586,n519,n544);
and (n587,n414,n456);
xor (n588,n589,n626);
xor (n589,n590,n593);
or (n590,n591,n592);
and (n591,n457,n480);
and (n592,n458,n466);
xor (n593,n594,n610);
xor (n594,n595,n596);
and (n595,n467,n473);
or (n596,n597,n609);
and (n597,n598,n606);
xor (n598,n599,n603);
nand (n599,n600,n602);
or (n600,n601,n382);
not (n601,n583);
nand (n602,n391,n384);
nand (n603,n604,n605);
or (n604,n17,n47);
nand (n605,n15,n424);
nand (n606,n607,n608);
or (n607,n112,n506);
nand (n608,n133,n151);
and (n609,n599,n603);
or (n610,n611,n625);
and (n611,n612,n621);
xor (n612,n613,n617);
nand (n613,n614,n616);
or (n614,n615,n489);
not (n615,n491);
nand (n616,n288,n273);
nand (n617,n618,n620);
or (n618,n306,n619);
not (n619,n501);
nand (n620,n321,n317);
nand (n621,n622,n624);
or (n622,n623,n351);
not (n623,n434);
nand (n624,n362,n341);
and (n625,n613,n617);
or (n626,n627,n634);
and (n627,n628,n633);
xor (n628,n629,n632);
or (n629,n630,n631);
and (n630,n573,n579);
and (n631,n574,n575);
xor (n632,n598,n606);
xor (n633,n612,n621);
and (n634,n629,n632);
not (n635,n636);
or (n636,n637,n697);
and (n637,n638,n696);
xor (n638,n639,n640);
xor (n639,n628,n633);
or (n640,n641,n695);
and (n641,n642,n645);
xor (n642,n643,n644);
xor (n643,n482,n504);
xor (n644,n416,n437);
or (n645,n646,n694);
and (n646,n647,n669);
xor (n647,n648,n649);
xor (n648,n438,n444);
or (n649,n650,n668);
and (n650,n651,n660);
xor (n651,n652,n653);
nor (n652,n206,n17);
nand (n653,n654,n659);
or (n654,n655,n489);
not (n655,n656);
nand (n656,n657,n658);
or (n657,n271,n323);
nand (n658,n323,n271);
nand (n659,n560,n273);
nand (n660,n661,n667);
or (n661,n662,n230);
not (n662,n663);
nand (n663,n664,n666);
or (n664,n218,n665);
not (n665,n136);
nand (n666,n665,n218);
nand (n667,n447,n232);
and (n668,n652,n653);
or (n669,n670,n693);
and (n670,n671,n686);
xor (n671,n672,n679);
nand (n672,n673,n678);
or (n673,n674,n112);
not (n674,n675);
nand (n675,n676,n677);
or (n676,n135,n188);
nand (n677,n135,n188);
nand (n678,n525,n151);
nand (n679,n680,n682);
or (n680,n681,n566);
not (n681,n317);
nand (n682,n683,n307);
nand (n683,n684,n685);
or (n684,n131,n50);
nand (n685,n50,n131);
nand (n686,n687,n692);
or (n687,n382,n688);
not (n688,n689);
nand (n689,n690,n691);
or (n690,n364,n290);
nand (n691,n290,n364);
nand (n692,n550,n384);
and (n693,n672,n679);
and (n694,n648,n649);
and (n695,n643,n644);
xor (n696,n413,n516);
and (n697,n639,n640);
nand (n698,n6,n636);
nand (n699,n700,n927);
nor (n700,n701,n921);
and (n701,n702,n808);
and (n702,n703,n770);
nand (n703,n704,n706);
not (n704,n705);
xor (n705,n638,n696);
not (n706,n707);
or (n707,n708,n769);
and (n708,n709,n712);
xor (n709,n710,n711);
xor (n710,n518,n572);
xor (n711,n642,n645);
or (n712,n713,n768);
and (n713,n714,n717);
xor (n714,n715,n716);
xor (n715,n521,n536);
xor (n716,n546,n564);
or (n717,n718,n767);
and (n718,n719,n742);
xor (n719,n720,n727);
nand (n720,n721,n726);
or (n721,n722,n351);
not (n722,n723);
nand (n723,n724,n725);
or (n724,n281,n223);
nand (n725,n223,n281);
nand (n726,n539,n362);
and (n727,n728,n736);
nand (n728,n729,n735);
or (n729,n730,n489);
not (n730,n731);
nand (n731,n732,n734);
or (n732,n234,n733);
not (n733,n145);
nand (n734,n733,n234);
nand (n735,n656,n273);
nor (n736,n737,n135);
and (n737,n738,n741);
nand (n738,n739,n131);
not (n739,n740);
and (n740,n207,n117);
nand (n741,n116,n206);
or (n742,n743,n766);
and (n743,n744,n759);
xor (n744,n745,n752);
nand (n745,n746,n747);
or (n746,n231,n662);
nand (n747,n748,n751);
nand (n748,n749,n750);
or (n749,n217,n104);
nand (n750,n104,n217);
not (n751,n230);
nand (n752,n753,n758);
or (n753,n754,n112);
not (n754,n755);
nand (n755,n756,n757);
or (n756,n135,n207);
nand (n757,n207,n135);
nand (n758,n675,n151);
nand (n759,n760,n762);
or (n760,n681,n761);
not (n761,n683);
nand (n762,n763,n307);
nand (n763,n764,n765);
or (n764,n131,n164);
nand (n765,n131,n164);
and (n766,n745,n752);
and (n767,n720,n727);
and (n768,n715,n716);
and (n769,n710,n711);
nand (n770,n771,n773);
not (n771,n772);
xor (n772,n709,n712);
not (n773,n774);
or (n774,n775,n807);
and (n775,n776,n806);
xor (n776,n777,n778);
xor (n777,n647,n669);
or (n778,n779,n805);
and (n779,n780,n783);
xor (n780,n781,n782);
xor (n781,n671,n686);
xor (n782,n651,n660);
or (n783,n784,n804);
and (n784,n785,n800);
xor (n785,n786,n793);
nand (n786,n787,n792);
or (n787,n788,n351);
not (n788,n789);
nand (n789,n790,n791);
or (n790,n350,n332);
nand (n791,n332,n350);
nand (n792,n723,n362);
nand (n793,n794,n799);
or (n794,n795,n382);
not (n795,n796);
nand (n796,n797,n798);
or (n797,n364,n258);
nand (n798,n258,n364);
nand (n799,n689,n384);
nand (n800,n801,n803);
or (n801,n736,n802);
not (n802,n728);
nand (n803,n802,n736);
and (n804,n786,n793);
and (n805,n781,n782);
xor (n806,n714,n717);
and (n807,n777,n778);
nand (n808,n809,n920);
or (n809,n810,n867);
nor (n810,n811,n812);
xor (n811,n776,n806);
or (n812,n813,n866);
and (n813,n814,n865);
xor (n814,n815,n816);
xor (n815,n719,n742);
or (n816,n817,n864);
and (n817,n818,n863);
xor (n818,n819,n844);
or (n819,n820,n843);
and (n820,n821,n836);
xor (n821,n822,n829);
nand (n822,n823,n828);
or (n823,n824,n306);
not (n824,n825);
nand (n825,n826,n827);
or (n826,n131,n188);
nand (n827,n131,n188);
nand (n828,n763,n317);
nand (n829,n830,n832);
or (n830,n231,n831);
not (n831,n748);
nand (n832,n833,n751);
nand (n833,n834,n835);
or (n834,n218,n514);
nand (n835,n514,n218);
nand (n836,n837,n842);
or (n837,n838,n351);
not (n838,n839);
nor (n839,n840,n841);
and (n840,n323,n281);
and (n841,n350,n453);
nand (n842,n789,n362);
and (n843,n822,n829);
or (n844,n845,n862);
and (n845,n846,n855);
xor (n846,n847,n848);
nor (n847,n206,n123);
nand (n848,n849,n854);
or (n849,n489,n850);
not (n850,n851);
nand (n851,n852,n853);
or (n852,n271,n136);
nand (n853,n136,n271);
nand (n854,n731,n273);
nand (n855,n856,n861);
or (n856,n857,n382);
not (n857,n858);
nand (n858,n859,n860);
or (n859,n364,n223);
nand (n860,n223,n364);
nand (n861,n796,n384);
and (n862,n847,n848);
xor (n863,n744,n759);
and (n864,n819,n844);
xor (n865,n780,n783);
and (n866,n815,n816);
nand (n867,n868,n869);
xor (n868,n814,n865);
or (n869,n870,n919);
and (n870,n871,n874);
xor (n871,n872,n873);
xor (n872,n785,n800);
xor (n873,n818,n863);
or (n874,n875,n918);
and (n875,n876,n917);
xor (n876,n877,n891);
and (n877,n878,n884);
nor (n878,n879,n131);
and (n879,n880,n883);
nand (n880,n881,n217);
not (n881,n882);
and (n882,n207,n310);
nand (n883,n206,n316);
nand (n884,n885,n890);
or (n885,n489,n886);
not (n886,n887);
nand (n887,n888,n889);
or (n888,n271,n104);
nand (n889,n104,n271);
nand (n890,n851,n273);
or (n891,n892,n916);
and (n892,n893,n909);
xor (n893,n894,n902);
nand (n894,n895,n901);
or (n895,n382,n896);
not (n896,n897);
nand (n897,n898,n900);
or (n898,n364,n899);
not (n899,n332);
nand (n900,n899,n364);
nand (n901,n858,n384);
nand (n902,n903,n908);
or (n903,n904,n351);
not (n904,n905);
nand (n905,n906,n907);
or (n906,n281,n733);
nand (n907,n733,n281);
nand (n908,n839,n362);
nand (n909,n910,n915);
or (n910,n911,n230);
not (n911,n912);
nand (n912,n913,n914);
or (n913,n217,n164);
nand (n914,n164,n217);
nand (n915,n833,n232);
and (n916,n894,n902);
xor (n917,n846,n855);
and (n918,n877,n891);
and (n919,n872,n873);
nand (n920,n811,n812);
nand (n921,n922,n926);
or (n922,n923,n925);
not (n923,n924);
nor (n924,n771,n773);
not (n925,n703);
nand (n926,n705,n707);
nand (n927,n703,n928,n1229,n770);
nand (n928,n929,n1217,n1223);
nand (n929,n930,n971,n1075);
nand (n930,n931,n933);
not (n931,n932);
xor (n932,n871,n874);
not (n933,n934);
or (n934,n935,n970);
and (n935,n936,n969);
xor (n936,n937,n938);
xor (n937,n821,n836);
or (n938,n939,n968);
and (n939,n940,n949);
xor (n940,n941,n948);
nand (n941,n942,n947);
or (n942,n306,n943);
not (n943,n944);
nor (n944,n945,n946);
and (n945,n131,n206);
and (n946,n207,n125);
nand (n947,n317,n825);
xor (n948,n878,n884);
or (n949,n950,n967);
and (n950,n951,n960);
xor (n951,n952,n953);
and (n952,n317,n207);
nand (n953,n954,n959);
or (n954,n955,n351);
not (n955,n956);
nand (n956,n957,n958);
or (n957,n281,n665);
nand (n958,n665,n281);
nand (n959,n905,n362);
nand (n960,n961,n966);
or (n961,n382,n962);
not (n962,n963);
nand (n963,n964,n965);
or (n964,n364,n453);
nand (n965,n453,n364);
nand (n966,n897,n384);
and (n967,n952,n953);
and (n968,n941,n948);
xor (n969,n876,n917);
and (n970,n937,n938);
nor (n971,n972,n1059,n1070);
nor (n972,n973,n1031);
xor (n973,n974,n1007);
xor (n974,n975,n1006);
or (n975,n976,n1005);
and (n976,n977,n995);
xor (n977,n978,n985);
nand (n978,n979,n984);
or (n979,n382,n980);
not (n980,n981);
nand (n981,n982,n983);
or (n982,n364,n733);
nand (n983,n733,n364);
nand (n984,n963,n384);
nand (n985,n986,n991);
or (n986,n987,n230);
not (n987,n988);
nand (n988,n989,n990);
or (n989,n218,n206);
or (n990,n207,n217);
nand (n991,n992,n232);
nand (n992,n993,n994);
or (n993,n217,n188);
nand (n994,n188,n217);
nand (n995,n996,n1001);
or (n996,n997,n489);
not (n997,n998);
nand (n998,n999,n1000);
or (n999,n271,n164);
nand (n1000,n164,n271);
nand (n1001,n1002,n273);
nand (n1002,n1003,n1004);
or (n1003,n271,n50);
nand (n1004,n50,n271);
and (n1005,n978,n985);
xor (n1006,n951,n960);
xor (n1007,n1008,n1017);
xor (n1008,n1009,n1013);
nand (n1009,n1010,n1012);
or (n1010,n1011,n230);
not (n1011,n992);
nand (n1012,n912,n232);
nand (n1013,n1014,n1016);
or (n1014,n1015,n489);
not (n1015,n1002);
nand (n1016,n887,n273);
and (n1017,n1018,n1025);
nand (n1018,n1019,n1024);
or (n1019,n1020,n351);
not (n1020,n1021);
nand (n1021,n1022,n1023);
or (n1022,n350,n104);
nand (n1023,n104,n350);
nand (n1024,n956,n362);
nor (n1025,n1026,n217);
and (n1026,n1027,n1030);
nand (n1027,n1028,n271);
not (n1028,n1029);
and (n1029,n207,n240);
nand (n1030,n206,n239);
or (n1031,n1032,n1058);
and (n1032,n1033,n1057);
xor (n1033,n1034,n1038);
nand (n1034,n1035,n1037);
or (n1035,n1025,n1036);
not (n1036,n1018);
nand (n1037,n1036,n1025);
or (n1038,n1039,n1056);
and (n1039,n1040,n1049);
xor (n1040,n1041,n1042);
and (n1041,n232,n207);
nand (n1042,n1043,n1048);
or (n1043,n1044,n351);
not (n1044,n1045);
nand (n1045,n1046,n1047);
or (n1046,n281,n514);
nand (n1047,n514,n281);
nand (n1048,n1021,n362);
nand (n1049,n1050,n1055);
or (n1050,n1051,n489);
not (n1051,n1052);
nand (n1052,n1053,n1054);
or (n1053,n271,n188);
nand (n1054,n188,n271);
nand (n1055,n998,n273);
and (n1056,n1041,n1042);
xor (n1057,n977,n995);
and (n1058,n1034,n1038);
nor (n1059,n1060,n1061);
xor (n1060,n936,n969);
or (n1061,n1062,n1069);
and (n1062,n1063,n1068);
xor (n1063,n1064,n1065);
xor (n1064,n893,n909);
or (n1065,n1066,n1067);
and (n1066,n1008,n1017);
and (n1067,n1009,n1013);
xor (n1068,n940,n949);
and (n1069,n1064,n1065);
nor (n1070,n1071,n1072);
xor (n1071,n1063,n1068);
or (n1072,n1073,n1074);
and (n1073,n974,n1007);
and (n1074,n975,n1006);
nand (n1075,n1076,n1216);
or (n1076,n1077,n1108);
not (n1077,n1078);
nand (n1078,n1079,n1081);
not (n1079,n1080);
xor (n1080,n1033,n1057);
not (n1081,n1082);
or (n1082,n1083,n1107);
and (n1083,n1084,n1106);
xor (n1084,n1085,n1092);
nand (n1085,n1086,n1091);
or (n1086,n382,n1087);
not (n1087,n1088);
nand (n1088,n1089,n1090);
or (n1089,n389,n136);
nand (n1090,n136,n389);
nand (n1091,n981,n384);
and (n1092,n1093,n1099);
nor (n1093,n1094,n271);
and (n1094,n1095,n1098);
nand (n1095,n1096,n350);
not (n1096,n1097);
and (n1097,n207,n276);
nand (n1098,n206,n275);
nand (n1099,n1100,n1105);
or (n1100,n1101,n351);
not (n1101,n1102);
nand (n1102,n1103,n1104);
or (n1103,n350,n164);
nand (n1104,n164,n350);
nand (n1105,n1045,n362);
xor (n1106,n1040,n1049);
and (n1107,n1085,n1092);
not (n1108,n1109);
nand (n1109,n1110,n1215);
or (n1110,n1111,n1210);
nor (n1111,n1112,n1209);
and (n1112,n1113,n1152);
nand (n1113,n1114,n1132);
not (n1114,n1115);
xor (n1115,n1116,n1131);
xor (n1116,n1117,n1124);
nand (n1117,n1118,n1123);
or (n1118,n1119,n489);
not (n1119,n1120);
nor (n1120,n1121,n1122);
and (n1121,n207,n234);
and (n1122,n271,n206);
nand (n1123,n273,n1052);
nand (n1124,n1125,n1126);
or (n1125,n410,n1087);
nand (n1126,n1127,n383);
nand (n1127,n1128,n1130);
or (n1128,n364,n1129);
not (n1129,n104);
nand (n1130,n364,n1129);
xor (n1131,n1093,n1099);
not (n1132,n1133);
or (n1133,n1134,n1151);
and (n1134,n1135,n1144);
xor (n1135,n1136,n1137);
and (n1136,n273,n207);
nand (n1137,n1138,n1140);
or (n1138,n410,n1139);
not (n1139,n1127);
nand (n1140,n1141,n383);
nand (n1141,n1142,n1143);
or (n1142,n364,n514);
nand (n1143,n514,n364);
nand (n1144,n1145,n1150);
or (n1145,n1146,n351);
not (n1146,n1147);
nand (n1147,n1148,n1149);
or (n1148,n350,n188);
nand (n1149,n188,n350);
nand (n1150,n1102,n362);
and (n1151,n1136,n1137);
nand (n1152,n1153,n1207);
or (n1153,n1154,n1172);
not (n1154,n1155);
nand (n1155,n1156,n1158);
not (n1156,n1157);
xor (n1157,n1135,n1144);
nand (n1158,n1159,n1166);
nand (n1159,n1160,n1162);
or (n1160,n410,n1161);
not (n1161,n1141);
nand (n1162,n1163,n383);
nand (n1163,n1164,n1165);
or (n1164,n389,n164);
nand (n1165,n164,n389);
nor (n1166,n1167,n350);
and (n1167,n1168,n1171);
nand (n1168,n1169,n389);
not (n1169,n1170);
and (n1170,n207,n355);
nand (n1171,n206,n361);
not (n1172,n1173);
or (n1173,n1174,n1206);
and (n1174,n1175,n1187);
xor (n1175,n1176,n1183);
nand (n1176,n1177,n1182);
or (n1177,n1178,n351);
not (n1178,n1179);
nor (n1179,n1180,n1181);
and (n1180,n207,n281);
and (n1181,n350,n206);
nand (n1182,n362,n1147);
nand (n1183,n1184,n1186);
or (n1184,n1185,n1159);
not (n1185,n1166);
nand (n1186,n1159,n1185);
or (n1187,n1188,n1205);
and (n1188,n1189,n1198);
xor (n1189,n1190,n1191);
and (n1190,n207,n362);
nand (n1191,n1192,n1194);
or (n1192,n410,n1193);
not (n1193,n1163);
nand (n1194,n1195,n383);
nand (n1195,n1196,n1197);
or (n1196,n389,n188);
nand (n1197,n188,n389);
nor (n1198,n1199,n1202);
nor (n1199,n1200,n1201);
and (n1200,n383,n206);
and (n1201,n1195,n384);
nand (n1202,n1203,n364);
not (n1203,n1204);
and (n1204,n207,n384);
and (n1205,n1190,n1191);
and (n1206,n1176,n1183);
nand (n1207,n1157,n1208);
not (n1208,n1158);
and (n1209,n1115,n1133);
nor (n1210,n1211,n1212);
xor (n1211,n1084,n1106);
or (n1212,n1213,n1214);
and (n1213,n1116,n1131);
and (n1214,n1117,n1124);
nand (n1215,n1211,n1212);
nand (n1216,n1080,n1082);
nand (n1217,n1218,n930);
or (n1218,n1219,n1221);
not (n1219,n1220);
nand (n1220,n1060,n1061);
not (n1221,n1222);
nand (n1222,n932,n934);
nand (n1223,n930,n1224,n1225);
not (n1224,n1059);
nand (n1225,n1226,n1228);
or (n1226,n1070,n1227);
nand (n1227,n973,n1031);
nand (n1228,n1071,n1072);
nor (n1229,n810,n1230);
nor (n1230,n868,n869);
nand (n1231,n699,n3);
xor (n1232,n1233,n1310);
xor (n1233,n1234,n1237);
xor (n1234,n1235,n1236);
and (n1235,n365,n207);
and (n1236,n385,n188);
not (n1237,n1238);
xor (n1238,n1239,n1301);
and (n1239,n1240,n1251);
wire s0n1240,s1n1240,notn1240;
or (n1240,s0n1240,s1n1240);
not(notn1240,n1243);
and (s0n1240,notn1240,n1241);
and (s1n1240,n1243,n1242);
and (n1243,n1244,n1249);
and (n1244,n1245,n1247);
not (n1245,n1246);
not (n1247,n1248);
not (n1249,n1250);
wire s0n1251,s1n1251,notn1251;
or (n1251,s0n1251,s1n1251);
not(notn1251,n1264);
and (s0n1251,notn1251,n1252);
and (s1n1251,n1264,n1263);
wire s0n1252,s1n1252,notn1252;
or (n1252,s0n1252,s1n1252);
not(notn1252,n1255);
and (s0n1252,notn1252,n1253);
and (s1n1252,n1255,n1254);
and (n1255,n1256,n1261);
and (n1256,n1257,n1259);
not (n1257,n1258);
not (n1259,n1260);
not (n1261,n1262);
and (n1264,n1265,n1267);
not (n1265,n1266);
or (n1267,n1268,n1269);
and (n1269,n1270,n1271);
or (n1271,n1272,n1273,n1274,n1275,n1276,n1277,n1278,n1279,n1280,n1281,n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,n1300);
and (n1301,n1302,n1305);
wire s0n1302,s1n1302,notn1302;
or (n1302,s0n1302,s1n1302);
not(notn1302,n1243);
and (s0n1302,notn1302,n1303);
and (s1n1302,n1243,n1304);
wire s0n1305,s1n1305,notn1305;
or (n1305,s0n1305,s1n1305);
not(notn1305,n1264);
and (s0n1305,notn1305,n1306);
and (s1n1305,n1264,n1309);
wire s0n1306,s1n1306,notn1306;
or (n1306,s0n1306,s1n1306);
not(notn1306,n1255);
and (s0n1306,notn1306,n1307);
and (s1n1306,n1255,n1308);
or (n1310,n1311,n1312);
and (n1311,n385,n207);
not (n1312,n1313);
and (n1313,n1302,n1251);
and (n1314,n1232,n1315);
xor (n1315,n1316,n2021);
xor (n1316,n1317,n2019);
xor (n1317,n1318,n2018);
xor (n1318,n1319,n2010);
xor (n1319,n1320,n2009);
xor (n1320,n1321,n1994);
xor (n1321,n1322,n1993);
xor (n1322,n1323,n1973);
xor (n1323,n1324,n1972);
xor (n1324,n1325,n1946);
xor (n1325,n1326,n1945);
xor (n1326,n1327,n1913);
xor (n1327,n1328,n1912);
xor (n1328,n1329,n1874);
xor (n1329,n1330,n1873);
xor (n1330,n1331,n1829);
xor (n1331,n1332,n1828);
xor (n1332,n1333,n1777);
xor (n1333,n1334,n229);
xor (n1334,n1335,n1721);
xor (n1335,n1336,n1720);
xor (n1336,n1337,n1658);
xor (n1337,n1338,n296);
xor (n1338,n1339,n1590);
xor (n1339,n1340,n1589);
xor (n1340,n1341,n1517);
xor (n1341,n1342,n1516);
xor (n1342,n1343,n1436);
xor (n1343,n1344,n1435);
xor (n1344,n1345,n1348);
xor (n1345,n1346,n1347);
and (n1346,n403,n384);
and (n1347,n394,n364);
or (n1348,n1349,n1352);
and (n1349,n1350,n1351);
and (n1350,n394,n384);
and (n1351,n373,n364);
and (n1352,n1353,n1354);
xor (n1353,n1350,n1351);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
and (n1356,n373,n384);
and (n1357,n344,n364);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
and (n1362,n344,n384);
and (n1363,n265,n364);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
and (n1368,n265,n384);
and (n1369,n291,n364);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
and (n1374,n291,n384);
and (n1375,n252,n364);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
and (n1380,n252,n384);
and (n1381,n224,n364);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
and (n1386,n224,n384);
and (n1387,n332,n364);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
and (n1392,n332,n384);
and (n1393,n323,n364);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
and (n1398,n323,n384);
and (n1399,n145,n364);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
and (n1404,n145,n384);
and (n1405,n136,n364);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
and (n1410,n136,n384);
and (n1411,n104,n364);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
and (n1416,n104,n384);
and (n1417,n50,n364);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
and (n1422,n50,n384);
and (n1423,n164,n364);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
and (n1428,n164,n384);
and (n1429,n188,n364);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
and (n1432,n1433,n1434);
and (n1433,n188,n384);
and (n1434,n207,n364);
and (n1435,n373,n355);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1353,n1354);
and (n1439,n344,n355);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1359,n1360);
and (n1445,n265,n355);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1365,n1366);
and (n1451,n291,n355);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1371,n1372);
and (n1457,n252,n355);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1377,n1378);
and (n1463,n224,n355);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
or (n1466,n1467,n1470);
and (n1467,n1468,n1469);
xor (n1468,n1383,n1384);
and (n1469,n332,n355);
and (n1470,n1471,n1472);
xor (n1471,n1468,n1469);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1389,n1390);
and (n1475,n323,n355);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1395,n1396);
and (n1481,n145,n355);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1401,n1402);
and (n1487,n136,n355);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1407,n1408);
and (n1493,n104,n355);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1413,n1414);
and (n1499,n50,n355);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1419,n1420);
and (n1505,n164,n355);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1425,n1426);
and (n1511,n188,n355);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
and (n1514,n1515,n1170);
xor (n1515,n1431,n1432);
and (n1516,n344,n281);
or (n1517,n1518,n1520);
and (n1518,n1519,n436);
xor (n1519,n1441,n1442);
and (n1520,n1521,n1522);
xor (n1521,n1519,n436);
or (n1522,n1523,n1526);
and (n1523,n1524,n1525);
xor (n1524,n1447,n1448);
and (n1525,n291,n281);
and (n1526,n1527,n1528);
xor (n1527,n1524,n1525);
or (n1528,n1529,n1532);
and (n1529,n1530,n1531);
xor (n1530,n1453,n1454);
and (n1531,n252,n281);
and (n1532,n1533,n1534);
xor (n1533,n1530,n1531);
or (n1534,n1535,n1538);
and (n1535,n1536,n1537);
xor (n1536,n1459,n1460);
and (n1537,n224,n281);
and (n1538,n1539,n1540);
xor (n1539,n1536,n1537);
or (n1540,n1541,n1544);
and (n1541,n1542,n1543);
xor (n1542,n1465,n1466);
and (n1543,n332,n281);
and (n1544,n1545,n1546);
xor (n1545,n1542,n1543);
or (n1546,n1547,n1549);
and (n1547,n1548,n840);
xor (n1548,n1471,n1472);
and (n1549,n1550,n1551);
xor (n1550,n1548,n840);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1477,n1478);
and (n1554,n145,n281);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1483,n1484);
and (n1560,n136,n281);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1489,n1490);
and (n1566,n104,n281);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
or (n1569,n1570,n1573);
and (n1570,n1571,n1572);
xor (n1571,n1495,n1496);
and (n1572,n50,n281);
and (n1573,n1574,n1575);
xor (n1574,n1571,n1572);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1501,n1502);
and (n1578,n164,n281);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1507,n1508);
and (n1584,n188,n281);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
and (n1587,n1588,n1180);
xor (n1588,n1513,n1514);
and (n1589,n265,n276);
or (n1590,n1591,n1594);
and (n1591,n1592,n1593);
xor (n1592,n1521,n1522);
and (n1593,n291,n276);
and (n1594,n1595,n1596);
xor (n1595,n1592,n1593);
or (n1596,n1597,n1600);
and (n1597,n1598,n1599);
xor (n1598,n1527,n1528);
and (n1599,n252,n276);
and (n1600,n1601,n1602);
xor (n1601,n1598,n1599);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1533,n1534);
and (n1605,n224,n276);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1539,n1540);
and (n1611,n332,n276);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1545,n1546);
and (n1617,n323,n276);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
or (n1620,n1621,n1624);
and (n1621,n1622,n1623);
xor (n1622,n1550,n1551);
and (n1623,n145,n276);
and (n1624,n1625,n1626);
xor (n1625,n1622,n1623);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1556,n1557);
and (n1629,n136,n276);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1562,n1563);
and (n1635,n104,n276);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1568,n1569);
and (n1641,n50,n276);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
xor (n1646,n1574,n1575);
and (n1647,n164,n276);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
or (n1650,n1651,n1654);
and (n1651,n1652,n1653);
xor (n1652,n1580,n1581);
and (n1653,n188,n276);
and (n1654,n1655,n1656);
xor (n1655,n1652,n1653);
and (n1656,n1657,n1097);
xor (n1657,n1586,n1587);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1595,n1596);
and (n1661,n252,n234);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1601,n1602);
and (n1667,n224,n234);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
or (n1670,n1671,n1674);
and (n1671,n1672,n1673);
xor (n1672,n1607,n1608);
and (n1673,n332,n234);
and (n1674,n1675,n1676);
xor (n1675,n1672,n1673);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1613,n1614);
and (n1679,n323,n234);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1619,n1620);
and (n1685,n145,n234);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1625,n1626);
and (n1691,n136,n234);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1631,n1632);
and (n1697,n104,n234);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1637,n1638);
and (n1703,n50,n234);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1643,n1644);
and (n1709,n164,n234);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1716);
and (n1713,n1714,n1715);
xor (n1714,n1649,n1650);
and (n1715,n188,n234);
and (n1716,n1717,n1718);
xor (n1717,n1714,n1715);
and (n1718,n1719,n1121);
xor (n1719,n1655,n1656);
and (n1720,n252,n240);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1663,n1664);
and (n1724,n224,n240);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1669,n1670);
and (n1730,n332,n240);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1675,n1676);
and (n1736,n323,n240);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1681,n1682);
and (n1742,n145,n240);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
or (n1745,n1746,n1749);
and (n1746,n1747,n1748);
xor (n1747,n1687,n1688);
and (n1748,n136,n240);
and (n1749,n1750,n1751);
xor (n1750,n1747,n1748);
or (n1751,n1752,n1755);
and (n1752,n1753,n1754);
xor (n1753,n1693,n1694);
and (n1754,n104,n240);
and (n1755,n1756,n1757);
xor (n1756,n1753,n1754);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
xor (n1759,n1699,n1700);
and (n1760,n50,n240);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1705,n1706);
and (n1766,n164,n240);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1711,n1712);
and (n1772,n188,n240);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
and (n1775,n1776,n1029);
xor (n1776,n1717,n1718);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1726,n1727);
and (n1780,n332,n218);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1732,n1733);
and (n1786,n323,n218);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1738,n1739);
and (n1792,n145,n218);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1744,n1745);
and (n1798,n136,n218);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1750,n1751);
and (n1804,n104,n218);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1756,n1757);
and (n1810,n50,n218);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1762,n1763);
and (n1816,n164,n218);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1768,n1769);
and (n1822,n188,n218);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
and (n1825,n1826,n1827);
xor (n1826,n1774,n1775);
and (n1827,n207,n218);
and (n1828,n332,n310);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1782,n1783);
and (n1832,n323,n310);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1788,n1789);
and (n1838,n145,n310);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
or (n1841,n1842,n1845);
and (n1842,n1843,n1844);
xor (n1843,n1794,n1795);
and (n1844,n136,n310);
and (n1845,n1846,n1847);
xor (n1846,n1843,n1844);
or (n1847,n1848,n1851);
and (n1848,n1849,n1850);
xor (n1849,n1800,n1801);
and (n1850,n104,n310);
and (n1851,n1852,n1853);
xor (n1852,n1849,n1850);
or (n1853,n1854,n1857);
and (n1854,n1855,n1856);
xor (n1855,n1806,n1807);
and (n1856,n50,n310);
and (n1857,n1858,n1859);
xor (n1858,n1855,n1856);
or (n1859,n1860,n1863);
and (n1860,n1861,n1862);
xor (n1861,n1812,n1813);
and (n1862,n164,n310);
and (n1863,n1864,n1865);
xor (n1864,n1861,n1862);
or (n1865,n1866,n1869);
and (n1866,n1867,n1868);
xor (n1867,n1818,n1819);
and (n1868,n188,n310);
and (n1869,n1870,n1871);
xor (n1870,n1867,n1868);
and (n1871,n1872,n882);
xor (n1872,n1824,n1825);
and (n1873,n323,n125);
or (n1874,n1875,n1878);
and (n1875,n1876,n1877);
xor (n1876,n1834,n1835);
and (n1877,n145,n125);
and (n1878,n1879,n1880);
xor (n1879,n1876,n1877);
or (n1880,n1881,n1884);
and (n1881,n1882,n1883);
xor (n1882,n1840,n1841);
and (n1883,n136,n125);
and (n1884,n1885,n1886);
xor (n1885,n1882,n1883);
or (n1886,n1887,n1890);
and (n1887,n1888,n1889);
xor (n1888,n1846,n1847);
and (n1889,n104,n125);
and (n1890,n1891,n1892);
xor (n1891,n1888,n1889);
or (n1892,n1893,n1896);
and (n1893,n1894,n1895);
xor (n1894,n1852,n1853);
and (n1895,n50,n125);
and (n1896,n1897,n1898);
xor (n1897,n1894,n1895);
or (n1898,n1899,n1902);
and (n1899,n1900,n1901);
xor (n1900,n1858,n1859);
and (n1901,n164,n125);
and (n1902,n1903,n1904);
xor (n1903,n1900,n1901);
or (n1904,n1905,n1908);
and (n1905,n1906,n1907);
xor (n1906,n1864,n1865);
and (n1907,n188,n125);
and (n1908,n1909,n1910);
xor (n1909,n1906,n1907);
and (n1910,n1911,n946);
xor (n1911,n1870,n1871);
and (n1912,n145,n117);
or (n1913,n1914,n1917);
and (n1914,n1915,n1916);
xor (n1915,n1879,n1880);
and (n1916,n136,n117);
and (n1917,n1918,n1919);
xor (n1918,n1915,n1916);
or (n1919,n1920,n1923);
and (n1920,n1921,n1922);
xor (n1921,n1885,n1886);
and (n1922,n104,n117);
and (n1923,n1924,n1925);
xor (n1924,n1921,n1922);
or (n1925,n1926,n1929);
and (n1926,n1927,n1928);
xor (n1927,n1891,n1892);
and (n1928,n50,n117);
and (n1929,n1930,n1931);
xor (n1930,n1927,n1928);
or (n1931,n1932,n1935);
and (n1932,n1933,n1934);
xor (n1933,n1897,n1898);
and (n1934,n164,n117);
and (n1935,n1936,n1937);
xor (n1936,n1933,n1934);
or (n1937,n1938,n1941);
and (n1938,n1939,n1940);
xor (n1939,n1903,n1904);
and (n1940,n188,n117);
and (n1941,n1942,n1943);
xor (n1942,n1939,n1940);
and (n1943,n1944,n740);
xor (n1944,n1909,n1910);
and (n1945,n136,n18);
or (n1946,n1947,n1950);
and (n1947,n1948,n1949);
xor (n1948,n1918,n1919);
and (n1949,n104,n18);
and (n1950,n1951,n1952);
xor (n1951,n1948,n1949);
or (n1952,n1953,n1955);
and (n1953,n1954,n512);
xor (n1954,n1924,n1925);
and (n1955,n1956,n1957);
xor (n1956,n1954,n512);
or (n1957,n1958,n1961);
and (n1958,n1959,n1960);
xor (n1959,n1930,n1931);
and (n1960,n164,n18);
and (n1961,n1962,n1963);
xor (n1962,n1959,n1960);
or (n1963,n1964,n1967);
and (n1964,n1965,n1966);
xor (n1965,n1936,n1937);
and (n1966,n188,n18);
and (n1967,n1968,n1969);
xor (n1968,n1965,n1966);
and (n1969,n1970,n1971);
xor (n1970,n1942,n1943);
and (n1971,n207,n18);
and (n1972,n104,n32);
or (n1973,n1974,n1977);
and (n1974,n1975,n1976);
xor (n1975,n1951,n1952);
and (n1976,n50,n32);
and (n1977,n1978,n1979);
xor (n1978,n1975,n1976);
or (n1979,n1980,n1983);
and (n1980,n1981,n1982);
xor (n1981,n1956,n1957);
and (n1982,n164,n32);
and (n1983,n1984,n1985);
xor (n1984,n1981,n1982);
or (n1985,n1986,n1989);
and (n1986,n1987,n1988);
xor (n1987,n1962,n1963);
and (n1988,n188,n32);
and (n1989,n1990,n1991);
xor (n1990,n1987,n1988);
and (n1991,n1992,n442);
xor (n1992,n1968,n1969);
and (n1993,n50,n40);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1978,n1979);
and (n1997,n164,n40);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
or (n2000,n2001,n2004);
and (n2001,n2002,n2003);
xor (n2002,n1984,n1985);
and (n2003,n188,n40);
and (n2004,n2005,n2006);
xor (n2005,n2002,n2003);
and (n2006,n2007,n2008);
xor (n2007,n1990,n1991);
and (n2008,n207,n40);
and (n2009,n164,n174);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1999,n2000);
and (n2013,n188,n174);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
and (n2016,n2017,n471);
xor (n2017,n2005,n2006);
and (n2018,n188,n158);
and (n2019,n2020,n463);
xor (n2020,n2015,n2016);
and (n2021,n207,n199);
endmodule
