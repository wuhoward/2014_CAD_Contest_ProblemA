module top (out,n7,n28,n30,n37,n44,n50,n58,n60,n68
        ,n69,n79,n86,n91,n92,n104,n119,n121,n125,n133
        ,n141,n168,n176,n180,n216,n237,n392,n414,n422,n428
        ,n465,n471,n525,n558,n597,n638,n643,n652,n695,n853
        ,n860,n867,n874,n881,n887,n889,n902,n932,n950,n977
        ,n1005,n1073);
output out;
input n7;
input n28;
input n30;
input n37;
input n44;
input n50;
input n58;
input n60;
input n68;
input n69;
input n79;
input n86;
input n91;
input n92;
input n104;
input n119;
input n121;
input n125;
input n133;
input n141;
input n168;
input n176;
input n180;
input n216;
input n237;
input n392;
input n414;
input n422;
input n428;
input n465;
input n471;
input n525;
input n558;
input n597;
input n638;
input n643;
input n652;
input n695;
input n853;
input n860;
input n867;
input n874;
input n881;
input n887;
input n889;
input n902;
input n932;
input n950;
input n977;
input n1005;
input n1073;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n639;
wire n640;
wire n641;
wire n642;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n888;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
xor (out,n0,n1077);
nand (n0,n1,n1076);
or (n1,n2,n909);
not (n2,n3);
nand (n3,n4,n903);
or (n4,n5,n689);
nor (n5,n6,n8);
not (n6,n7);
nand (n8,n9,n688);
or (n9,n10,n576);
nand (n10,n11,n575);
or (n11,n12,n445);
not (n12,n13);
nand (n13,n14,n444);
or (n14,n15,n359);
nor (n15,n16,n358);
and (n16,n17,n270);
nand (n17,n18,n239);
not (n18,n19);
xor (n19,n20,n150);
xor (n20,n21,n106);
xor (n21,n22,n81);
xor (n22,n23,n53);
nand (n23,n24,n46);
or (n24,n25,n33);
not (n25,n26);
nand (n26,n27,n31);
or (n27,n28,n29);
not (n29,n30);
or (n31,n32,n30);
not (n32,n28);
nand (n33,n34,n41);
or (n34,n35,n38);
not (n35,n36);
nand (n36,n29,n37);
not (n38,n39);
nand (n39,n40,n30);
not (n40,n37);
nor (n41,n42,n45);
and (n42,n43,n37);
not (n43,n44);
and (n45,n44,n40);
nand (n46,n47,n52);
nor (n47,n48,n51);
and (n48,n49,n29);
not (n49,n50);
and (n51,n50,n30);
not (n52,n41);
nand (n53,n54,n75);
or (n54,n55,n63);
not (n55,n56);
nor (n56,n57,n61);
and (n57,n58,n59);
not (n59,n60);
and (n61,n62,n60);
not (n62,n58);
nand (n63,n64,n71);
not (n64,n65);
nand (n65,n66,n70);
or (n66,n67,n69);
not (n67,n68);
nand (n70,n67,n69);
nand (n71,n72,n74);
or (n72,n73,n60);
not (n73,n69);
nand (n74,n60,n73);
or (n75,n64,n76);
nor (n76,n77,n80);
and (n77,n59,n78);
not (n78,n79);
and (n80,n60,n79);
nand (n81,n82,n95);
or (n82,n83,n88);
nor (n83,n84,n87);
and (n84,n85,n60);
not (n85,n86);
and (n87,n86,n59);
not (n88,n89);
nand (n89,n90,n93);
or (n90,n91,n92);
not (n93,n94);
and (n94,n92,n91);
or (n95,n96,n101);
nand (n96,n83,n97);
nand (n97,n98,n100);
or (n98,n86,n99);
not (n99,n91);
nand (n100,n99,n86);
nor (n101,n102,n105);
and (n102,n103,n99);
not (n103,n104);
and (n105,n104,n91);
or (n106,n107,n149);
and (n107,n108,n135);
xor (n108,n109,n116);
nand (n109,n110,n115);
or (n110,n111,n63);
nor (n111,n112,n113);
and (n112,n92,n60);
and (n113,n114,n59);
not (n114,n92);
nand (n115,n56,n65);
nand (n116,n117,n129);
or (n117,n118,n122);
nand (n118,n119,n120);
not (n120,n121);
not (n122,n123);
nor (n123,n124,n126);
and (n124,n125,n119);
and (n126,n127,n128);
not (n127,n125);
not (n128,n119);
or (n129,n130,n120);
not (n130,n131);
nand (n131,n132,n134);
or (n132,n133,n128);
nand (n134,n128,n133);
and (n135,n136,n144);
nor (n136,n137,n43);
and (n137,n138,n142);
nand (n138,n139,n128);
not (n139,n140);
and (n140,n28,n141);
nand (n142,n143,n32);
not (n143,n141);
nor (n144,n145,n60);
and (n145,n146,n148);
nand (n146,n147,n68);
or (n147,n103,n69);
nand (n148,n103,n69);
and (n149,n109,n116);
xor (n150,n151,n221);
xor (n151,n152,n198);
or (n152,n153,n197);
and (n153,n154,n190);
xor (n154,n155,n173);
nand (n155,n156,n165);
or (n156,n157,n161);
not (n157,n158);
nand (n158,n159,n160);
or (n159,n50,n43);
nand (n160,n43,n50);
not (n161,n162);
nand (n162,n163,n164);
nand (n163,n119,n141,n43);
nand (n164,n143,n128,n44);
nand (n165,n166,n170);
nand (n166,n167,n169);
or (n167,n168,n43);
nand (n169,n43,n168);
nand (n170,n171,n172);
or (n171,n143,n119);
nand (n172,n143,n119);
nand (n173,n174,n183);
or (n174,n175,n177);
not (n175,n176);
not (n177,n178);
nor (n178,n179,n181);
and (n179,n180,n67);
and (n181,n182,n68);
not (n182,n180);
nand (n183,n184,n188);
nand (n184,n185,n187);
not (n185,n186);
and (n186,n79,n68);
nand (n187,n67,n78);
not (n188,n189);
nand (n189,n175,n68);
nand (n190,n191,n196);
or (n191,n192,n194);
not (n192,n193);
nand (n193,n52,n28);
nand (n194,n195,n104);
not (n195,n83);
nand (n196,n192,n194);
and (n197,n155,n173);
xor (n198,n199,n211);
xor (n199,n200,n206);
nor (n200,n201,n29);
and (n201,n202,n205);
nand (n202,n203,n43);
not (n203,n204);
and (n204,n28,n37);
nand (n205,n32,n40);
and (n206,n207,n99);
nand (n207,n208,n209);
or (n208,n85,n104);
nand (n209,n210,n60);
or (n210,n86,n103);
nand (n211,n212,n219);
or (n212,n120,n213);
not (n213,n214);
nor (n214,n215,n217);
and (n215,n216,n119);
and (n217,n218,n128);
not (n218,n216);
nand (n219,n131,n220);
not (n220,n118);
xor (n221,n222,n231);
xor (n222,n223,n230);
nand (n223,n224,n226);
or (n224,n225,n161);
not (n225,n166);
nand (n226,n227,n170);
nand (n227,n228,n229);
or (n228,n127,n44);
nand (n229,n44,n127);
nor (n230,n194,n193);
nand (n231,n232,n233);
or (n232,n189,n177);
or (n233,n234,n175);
nor (n234,n235,n238);
and (n235,n67,n236);
not (n236,n237);
and (n238,n68,n237);
not (n239,n240);
or (n240,n241,n269);
and (n241,n242,n268);
xor (n242,n243,n267);
or (n243,n244,n266);
and (n244,n245,n260);
xor (n245,n246,n253);
nand (n246,n247,n252);
or (n247,n248,n161);
not (n248,n249);
nor (n249,n250,n251);
and (n250,n32,n43);
and (n251,n28,n44);
nand (n252,n158,n170);
nand (n253,n254,n259);
or (n254,n189,n255);
not (n255,n256);
nor (n256,n257,n258);
and (n257,n58,n67);
and (n258,n62,n68);
nand (n259,n184,n176);
nand (n260,n261,n265);
or (n261,n63,n262);
nor (n262,n263,n264);
and (n263,n59,n103);
and (n264,n104,n60);
or (n265,n64,n111);
and (n266,n246,n253);
xor (n267,n154,n190);
xor (n268,n108,n135);
and (n269,n243,n267);
nand (n270,n271,n357);
or (n271,n272,n316);
not (n272,n273);
nand (n273,n274,n276);
not (n274,n275);
xor (n275,n242,n268);
not (n276,n277);
or (n277,n278,n315);
and (n278,n279,n293);
xor (n279,n280,n288);
nand (n280,n281,n282);
or (n281,n120,n122);
or (n282,n118,n283);
not (n283,n284);
nor (n284,n285,n286);
and (n285,n168,n119);
and (n286,n287,n128);
not (n287,n168);
xor (n288,n289,n290);
xor (n289,n136,n144);
nor (n290,n291,n292);
nand (n291,n65,n104);
nand (n292,n170,n28);
or (n293,n294,n314);
and (n294,n295,n307);
xor (n295,n296,n303);
nand (n296,n297,n302);
or (n297,n118,n298);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n49,n128);
and (n301,n50,n119);
nand (n302,n284,n121);
nand (n303,n304,n306);
or (n304,n292,n305);
not (n305,n291);
nand (n306,n305,n292);
nand (n307,n308,n313);
or (n308,n189,n309);
not (n309,n310);
nor (n310,n311,n312);
and (n311,n92,n67);
and (n312,n114,n68);
nand (n313,n256,n176);
and (n314,n296,n303);
and (n315,n280,n288);
not (n316,n317);
nand (n317,n318,n356);
or (n318,n319,n322);
nor (n319,n320,n321);
xor (n320,n279,n293);
xor (n321,n245,n260);
nor (n322,n323,n354);
and (n323,n324,n341);
nand (n324,n325,n327);
not (n325,n326);
xor (n326,n295,n307);
not (n327,n328);
or (n328,n329,n340);
and (n329,n330,n334);
xor (n330,n331,n333);
nor (n331,n332,n128);
and (n332,n28,n121);
and (n333,n67,n103,n176);
nand (n334,n335,n336);
or (n335,n175,n309);
or (n336,n337,n189);
nor (n337,n338,n339);
and (n338,n67,n103);
and (n339,n104,n68);
and (n340,n331,n333);
or (n341,n342,n353);
and (n342,n343,n352);
xor (n343,n344,n346);
and (n344,n332,n345);
and (n345,n104,n176);
nand (n346,n347,n348);
or (n347,n120,n298);
nand (n348,n349,n220);
nand (n349,n350,n351);
or (n350,n128,n28);
or (n351,n32,n119);
xor (n352,n330,n334);
and (n353,n344,n346);
not (n354,n355);
nand (n355,n326,n328);
nand (n356,n320,n321);
nand (n357,n275,n277);
and (n358,n19,n240);
nor (n359,n360,n441);
xor (n360,n361,n379);
xor (n361,n362,n376);
xor (n362,n363,n373);
xor (n363,n364,n370);
nand (n364,n365,n366);
or (n365,n88,n96);
nand (n366,n195,n367);
nor (n367,n368,n369);
and (n368,n62,n91);
and (n369,n58,n99);
or (n370,n371,n372);
and (n371,n222,n231);
and (n372,n223,n230);
or (n373,n374,n375);
and (n374,n199,n211);
and (n375,n200,n206);
or (n376,n377,n378);
and (n377,n151,n221);
and (n378,n152,n198);
xor (n379,n380,n407);
xor (n380,n381,n384);
or (n381,n382,n383);
and (n382,n22,n81);
and (n383,n23,n53);
xor (n384,n385,n401);
xor (n385,n386,n394);
nand (n386,n387,n388);
or (n387,n234,n189);
or (n388,n389,n175);
nor (n389,n390,n393);
and (n390,n67,n391);
not (n391,n392);
and (n393,n68,n392);
nand (n394,n395,n397);
or (n395,n396,n33);
not (n396,n47);
nand (n397,n398,n52);
nand (n398,n399,n400);
or (n399,n168,n29);
or (n400,n30,n287);
nand (n401,n402,n403);
or (n402,n63,n76);
nand (n403,n65,n404);
nor (n404,n405,n406);
and (n405,n182,n60);
and (n406,n180,n59);
xor (n407,n408,n431);
xor (n408,n409,n416);
nand (n409,n410,n411);
or (n410,n213,n118);
nand (n411,n412,n121);
nand (n412,n413,n415);
or (n413,n414,n128);
nand (n415,n128,n414);
nand (n416,n417,n430);
or (n417,n418,n424);
not (n418,n419);
nand (n419,n420,n28);
nand (n420,n421,n423);
or (n421,n29,n422);
nand (n423,n29,n422);
nand (n424,n425,n104);
nand (n425,n426,n429);
or (n426,n427,n91);
not (n427,n428);
nand (n429,n427,n91);
nand (n430,n418,n424);
nand (n431,n432,n434);
or (n432,n161,n433);
not (n433,n227);
or (n434,n435,n436);
not (n435,n170);
not (n436,n437);
nand (n437,n438,n440);
or (n438,n439,n44);
not (n439,n133);
nand (n440,n44,n439);
or (n441,n442,n443);
and (n442,n20,n150);
and (n443,n21,n106);
nand (n444,n360,n441);
not (n445,n446);
nand (n446,n447,n571);
not (n447,n448);
xor (n448,n449,n528);
xor (n449,n450,n453);
or (n450,n451,n452);
and (n451,n380,n407);
and (n452,n381,n384);
xor (n453,n454,n490);
xor (n454,n455,n487);
xor (n455,n456,n472);
xor (n456,n457,n466);
nor (n457,n458,n464);
and (n458,n459,n462);
nand (n459,n460,n29);
not (n460,n461);
and (n461,n28,n422);
nand (n462,n463,n32);
not (n463,n422);
not (n464,n465);
nor (n466,n467,n471);
nor (n467,n468,n470);
and (n468,n469,n91);
nand (n469,n104,n427);
and (n470,n103,n428);
nand (n472,n473,n483);
or (n473,n474,n478);
not (n474,n475);
nor (n475,n476,n477);
and (n476,n464,n32);
and (n477,n28,n465);
nand (n478,n479,n482);
nand (n479,n480,n481);
or (n480,n422,n464);
nand (n481,n464,n422);
not (n482,n420);
nand (n483,n484,n420);
nand (n484,n485,n486);
or (n485,n50,n464);
nand (n486,n464,n50);
or (n487,n488,n489);
and (n488,n385,n401);
and (n489,n386,n394);
xor (n490,n491,n518);
xor (n491,n492,n499);
nand (n492,n493,n495);
or (n493,n494,n96);
not (n494,n367);
nand (n495,n195,n496);
nor (n496,n497,n498);
and (n497,n78,n91);
and (n498,n79,n99);
nand (n499,n500,n507);
or (n500,n501,n502);
not (n501,n425);
not (n502,n503);
nand (n503,n504,n505);
or (n504,n471,n92);
not (n505,n506);
and (n506,n92,n471);
nand (n507,n508,n513);
not (n508,n509);
nor (n509,n510,n512);
and (n510,n103,n511);
not (n511,n471);
and (n512,n104,n471);
not (n513,n514);
nand (n514,n501,n515);
nand (n515,n516,n517);
or (n516,n428,n511);
nand (n517,n511,n428);
nand (n518,n519,n521);
or (n519,n118,n520);
not (n520,n412);
or (n521,n522,n120);
not (n522,n523);
nor (n523,n524,n526);
and (n524,n525,n119);
and (n526,n527,n128);
not (n527,n525);
xor (n528,n529,n549);
xor (n529,n530,n546);
xor (n530,n531,n539);
xor (n531,n532,n538);
nand (n532,n533,n534);
or (n533,n436,n161);
nand (n534,n535,n170);
nor (n535,n536,n537);
and (n536,n218,n43);
and (n537,n216,n44);
nor (n538,n419,n424);
nand (n539,n540,n542);
or (n540,n541,n33);
not (n541,n398);
nand (n542,n52,n543);
nand (n543,n544,n545);
or (n544,n125,n29);
nand (n545,n29,n125);
or (n546,n547,n548);
and (n547,n363,n373);
and (n548,n364,n370);
xor (n549,n550,n568);
xor (n550,n551,n561);
nand (n551,n552,n553);
or (n552,n389,n189);
or (n553,n554,n175);
not (n554,n555);
nand (n555,n556,n559);
not (n556,n557);
and (n557,n558,n68);
nand (n559,n67,n560);
not (n560,n558);
nand (n561,n562,n564);
or (n562,n563,n63);
not (n563,n404);
nand (n564,n65,n565);
nor (n565,n566,n567);
and (n566,n236,n60);
and (n567,n237,n59);
or (n568,n569,n570);
and (n569,n408,n431);
and (n570,n409,n416);
not (n571,n572);
or (n572,n573,n574);
and (n573,n361,n379);
and (n574,n362,n376);
nand (n575,n448,n572);
nand (n576,n577,n687);
or (n577,n578,n684);
xor (n578,n579,n665);
xor (n579,n580,n662);
xor (n580,n581,n630);
xor (n581,n582,n607);
xor (n582,n583,n600);
xor (n583,n584,n591);
nand (n584,n585,n587);
nand (n585,n586,n543);
not (n586,n33);
nand (n587,n588,n52);
nor (n588,n589,n590);
and (n589,n439,n29);
and (n590,n133,n30);
nand (n591,n592,n599);
or (n592,n175,n593);
not (n593,n594);
nor (n594,n595,n598);
and (n595,n596,n68);
not (n596,n597);
and (n598,n597,n67);
nand (n599,n555,n188);
nand (n600,n601,n603);
or (n601,n602,n63);
not (n602,n565);
nand (n603,n65,n604);
nor (n604,n605,n606);
and (n605,n391,n60);
and (n606,n392,n59);
xor (n607,n608,n623);
xor (n608,n609,n616);
nand (n609,n610,n612);
or (n610,n611,n478);
not (n611,n484);
nand (n612,n613,n420);
nand (n613,n614,n615);
or (n614,n168,n464);
nand (n615,n464,n168);
nand (n616,n617,n619);
or (n617,n618,n96);
not (n618,n496);
nand (n619,n195,n620);
nor (n620,n621,n622);
and (n621,n182,n91);
and (n622,n180,n99);
nand (n623,n624,n625);
or (n624,n502,n514);
nand (n625,n425,n626);
nand (n626,n627,n628);
or (n627,n471,n58);
not (n628,n629);
and (n629,n58,n471);
xor (n630,n631,n654);
xor (n631,n632,n646);
nand (n632,n633,n645);
or (n633,n634,n640);
not (n634,n635);
nand (n635,n636,n28);
nand (n636,n637,n639);
or (n637,n464,n638);
nand (n639,n464,n638);
nand (n640,n641,n104);
nand (n641,n642,n644);
or (n642,n511,n643);
nand (n644,n511,n643);
nand (n645,n634,n640);
nand (n646,n647,n648);
or (n647,n118,n522);
nand (n648,n649,n121);
nand (n649,n650,n653);
or (n650,n651,n119);
not (n651,n652);
nand (n653,n119,n651);
nand (n654,n655,n657);
or (n655,n161,n656);
not (n656,n535);
or (n657,n435,n658);
nor (n658,n659,n660);
and (n659,n414,n43);
and (n660,n661,n44);
not (n661,n414);
or (n662,n663,n664);
and (n663,n529,n549);
and (n664,n530,n546);
xor (n665,n666,n673);
xor (n666,n667,n670);
or (n667,n668,n669);
and (n668,n550,n568);
and (n669,n551,n561);
or (n670,n671,n672);
and (n671,n454,n490);
and (n672,n455,n487);
xor (n673,n674,n681);
xor (n674,n675,n678);
or (n675,n676,n677);
and (n676,n531,n539);
and (n677,n532,n538);
or (n678,n679,n680);
and (n679,n456,n472);
and (n680,n457,n466);
or (n681,n682,n683);
and (n682,n491,n518);
and (n683,n492,n499);
or (n684,n685,n686);
and (n685,n449,n528);
and (n686,n450,n453);
nand (n687,n578,n684);
nand (n688,n576,n10);
not (n689,n690);
and (n690,n691,n898);
or (n691,n692,n897);
and (n692,n693,n702);
xor (n693,n694,n696);
not (n694,n695);
nand (n696,n697,n701);
or (n697,n698,n699);
not (n698,n15);
nand (n699,n700,n444);
not (n700,n359);
nand (n701,n699,n698);
or (n702,n703,n854,n896);
and (n703,n704,n852);
xor (n704,n705,n822);
xor (n705,n706,n763);
xor (n706,n707,n762);
xor (n707,n708,n760);
xor (n708,n709,n759);
xor (n709,n710,n751);
xor (n710,n711,n750);
xor (n711,n712,n736);
xor (n712,n713,n735);
xor (n713,n714,n717);
xor (n714,n715,n716);
and (n715,n216,n121);
and (n716,n133,n119);
or (n717,n718,n720);
and (n718,n719,n124);
and (n719,n133,n121);
and (n720,n721,n722);
xor (n721,n719,n124);
or (n722,n723,n725);
and (n723,n724,n285);
and (n724,n125,n121);
and (n725,n726,n727);
xor (n726,n724,n285);
or (n727,n728,n730);
and (n728,n729,n301);
and (n729,n168,n121);
and (n730,n731,n732);
xor (n731,n729,n301);
and (n732,n733,n734);
and (n733,n50,n121);
and (n734,n28,n119);
and (n735,n125,n141);
or (n736,n737,n740);
and (n737,n738,n739);
xor (n738,n721,n722);
and (n739,n168,n141);
and (n740,n741,n742);
xor (n741,n738,n739);
or (n742,n743,n746);
and (n743,n744,n745);
xor (n744,n726,n727);
and (n745,n50,n141);
and (n746,n747,n748);
xor (n747,n744,n745);
and (n748,n749,n140);
xor (n749,n731,n732);
and (n750,n168,n44);
or (n751,n752,n755);
and (n752,n753,n754);
xor (n753,n741,n742);
and (n754,n50,n44);
and (n755,n756,n757);
xor (n756,n753,n754);
and (n757,n758,n251);
xor (n758,n747,n748);
and (n759,n50,n37);
and (n760,n761,n204);
xor (n761,n756,n757);
and (n762,n28,n30);
not (n763,n764);
xor (n764,n765,n105);
xor (n765,n766,n819);
xor (n766,n767,n818);
xor (n767,n768,n811);
xor (n768,n769,n810);
xor (n769,n770,n795);
xor (n770,n771,n794);
xor (n771,n772,n775);
xor (n772,n773,n774);
and (n773,n237,n176);
and (n774,n180,n68);
or (n775,n776,n778);
and (n776,n777,n186);
and (n777,n180,n176);
and (n778,n779,n780);
xor (n779,n777,n186);
or (n780,n781,n784);
and (n781,n782,n783);
and (n782,n79,n176);
and (n783,n58,n68);
and (n784,n785,n786);
xor (n785,n782,n783);
or (n786,n787,n790);
and (n787,n788,n789);
and (n788,n58,n176);
and (n789,n92,n68);
and (n790,n791,n792);
xor (n791,n788,n789);
and (n792,n793,n339);
and (n793,n92,n176);
and (n794,n79,n69);
or (n795,n796,n799);
and (n796,n797,n798);
xor (n797,n779,n780);
and (n798,n58,n69);
and (n799,n800,n801);
xor (n800,n797,n798);
or (n801,n802,n805);
and (n802,n803,n804);
xor (n803,n785,n786);
and (n804,n92,n69);
and (n805,n806,n807);
xor (n806,n803,n804);
and (n807,n808,n809);
xor (n808,n791,n792);
and (n809,n104,n69);
and (n810,n58,n60);
or (n811,n812,n814);
and (n812,n813,n112);
xor (n813,n800,n801);
and (n814,n815,n816);
xor (n815,n813,n112);
and (n816,n817,n264);
xor (n817,n806,n807);
and (n818,n92,n86);
and (n819,n820,n821);
xor (n820,n815,n816);
and (n821,n104,n86);
or (n822,n823,n827,n851);
and (n823,n824,n825);
xor (n824,n761,n204);
not (n825,n826);
xor (n826,n820,n821);
and (n827,n825,n828);
or (n828,n829,n833,n850);
and (n829,n830,n831);
xor (n830,n758,n251);
not (n831,n832);
xor (n832,n817,n264);
and (n833,n831,n834);
or (n834,n835,n839,n849);
and (n835,n836,n837);
xor (n836,n749,n140);
not (n837,n838);
xor (n838,n808,n809);
and (n839,n837,n840);
or (n840,n841,n845,n848);
and (n841,n842,n843);
xor (n842,n733,n734);
not (n843,n844);
xor (n844,n793,n339);
and (n845,n843,n846);
or (n846,n332,n847);
not (n847,n345);
and (n848,n842,n846);
and (n849,n836,n840);
and (n850,n830,n834);
and (n851,n824,n828);
not (n852,n853);
and (n854,n852,n855);
or (n855,n856,n861,n895);
and (n856,n857,n859);
xor (n857,n858,n828);
xor (n858,n824,n825);
not (n859,n860);
and (n861,n859,n862);
or (n862,n863,n868,n894);
and (n863,n864,n866);
xor (n864,n865,n834);
xor (n865,n830,n831);
not (n866,n867);
and (n868,n866,n869);
or (n869,n870,n875,n893);
and (n870,n871,n873);
xor (n871,n872,n840);
xor (n872,n836,n837);
not (n873,n874);
and (n875,n873,n876);
or (n876,n877,n882,n892);
and (n877,n878,n880);
xor (n878,n879,n846);
xor (n879,n842,n843);
not (n880,n881);
and (n882,n883,n880);
or (n883,n884,n891);
and (n884,n885,n890);
xor (n885,n886,n888);
not (n886,n887);
not (n888,n889);
xor (n890,n332,n345);
and (n891,n888,n886);
and (n892,n878,n883);
and (n893,n871,n876);
and (n894,n864,n869);
and (n895,n857,n862);
and (n896,n704,n855);
and (n897,n694,n696);
nand (n898,n899,n902);
not (n899,n900);
xnor (n900,n13,n901);
nand (n901,n446,n575);
nor (n903,n904,n907);
nor (n904,n5,n905);
nand (n905,n906,n900);
not (n906,n902);
nor (n907,n908,n7);
not (n908,n8);
not (n909,n910);
nand (n910,n911,n1074);
nand (n911,n912,n1073);
not (n912,n913);
nand (n913,n914,n1072);
or (n914,n915,n1069);
not (n915,n916);
nand (n916,n917,n1068);
nand (n917,n918,n1064);
not (n918,n919);
xor (n919,n920,n995);
xor (n920,n921,n992);
xor (n921,n922,n989);
xor (n922,n923,n942);
xor (n923,n924,n941);
xor (n924,n925,n934);
nand (n925,n926,n928);
or (n926,n118,n927);
not (n927,n649);
or (n928,n929,n120);
nor (n929,n930,n933);
and (n930,n119,n931);
not (n931,n932);
nor (n933,n931,n119);
nand (n934,n935,n940);
or (n935,n936,n41);
not (n936,n937);
nor (n937,n938,n939);
and (n938,n29,n218);
and (n939,n30,n216);
nand (n940,n588,n586);
nor (n941,n635,n640);
xor (n942,n943,n970);
xor (n943,n944,n962);
nand (n944,n945,n952);
or (n945,n946,n947);
not (n946,n636);
not (n947,n948);
nand (n948,n949,n951);
or (n949,n950,n49);
nand (n951,n950,n49);
nand (n952,n946,n953,n956);
nand (n953,n954,n955);
or (n954,n950,n32);
nand (n955,n32,n950);
not (n956,n957);
nor (n957,n958,n960);
and (n958,n638,n959);
not (n959,n950);
and (n960,n950,n961);
not (n961,n638);
nand (n962,n963,n965);
or (n963,n964,n514);
not (n964,n626);
nand (n965,n425,n966);
nand (n966,n967,n969);
not (n967,n968);
and (n968,n79,n471);
nand (n969,n78,n511);
nand (n970,n971,n985);
or (n971,n972,n982);
nand (n972,n973,n981);
or (n973,n974,n978);
not (n974,n975);
nand (n975,n976,n643);
not (n976,n977);
not (n978,n979);
nand (n979,n980,n977);
not (n980,n643);
not (n981,n641);
nor (n982,n983,n984);
and (n983,n103,n976);
and (n984,n104,n977);
or (n985,n981,n986);
nor (n986,n987,n988);
and (n987,n976,n114);
and (n988,n977,n92);
or (n989,n990,n991);
and (n990,n674,n681);
and (n991,n675,n678);
or (n992,n993,n994);
and (n993,n666,n673);
and (n994,n667,n670);
xor (n995,n996,n1016);
xor (n996,n997,n1013);
xor (n997,n998,n1010);
xor (n998,n999,n1007);
nand (n999,n1000,n1001);
or (n1000,n189,n593);
or (n1001,n1002,n175);
nor (n1002,n1003,n1006);
and (n1003,n67,n1004);
not (n1004,n1005);
and (n1006,n68,n1005);
or (n1007,n1008,n1009);
and (n1008,n631,n654);
and (n1009,n632,n646);
or (n1010,n1011,n1012);
and (n1011,n583,n600);
and (n1012,n584,n591);
or (n1013,n1014,n1015);
and (n1014,n581,n630);
and (n1015,n582,n607);
xor (n1016,n1017,n1040);
xor (n1017,n1018,n1037);
xor (n1018,n1019,n1031);
xor (n1019,n1020,n1026);
nor (n1020,n1021,n959);
and (n1021,n1022,n1025);
nand (n1022,n1023,n464);
not (n1023,n1024);
and (n1024,n28,n638);
nand (n1025,n32,n961);
nor (n1026,n1027,n977);
nor (n1027,n1028,n1030);
and (n1028,n1029,n471);
nand (n1029,n104,n980);
and (n1030,n103,n643);
nand (n1031,n1032,n1033);
or (n1032,n658,n161);
nand (n1033,n1034,n170);
nor (n1034,n1035,n1036);
and (n1035,n527,n43);
and (n1036,n525,n44);
or (n1037,n1038,n1039);
and (n1038,n608,n623);
and (n1039,n609,n616);
xor (n1040,n1041,n1057);
xor (n1041,n1042,n1049);
nand (n1042,n1043,n1045);
or (n1043,n1044,n478);
not (n1044,n613);
nand (n1045,n420,n1046);
nor (n1046,n1047,n1048);
and (n1047,n127,n464);
and (n1048,n125,n465);
nand (n1049,n1050,n1052);
or (n1050,n63,n1051);
not (n1051,n604);
nand (n1052,n65,n1053);
nand (n1053,n1054,n1055);
or (n1054,n558,n60);
not (n1055,n1056);
and (n1056,n558,n60);
nand (n1057,n1058,n1060);
or (n1058,n1059,n96);
not (n1059,n620);
nand (n1060,n195,n1061);
nor (n1061,n1062,n1063);
and (n1062,n236,n91);
and (n1063,n237,n99);
not (n1064,n1065);
or (n1065,n1066,n1067);
and (n1066,n579,n665);
and (n1067,n580,n662);
nand (n1068,n919,n1065);
nor (n1069,n1070,n1071);
and (n1070,n10,n577);
not (n1071,n687);
nand (n1072,n915,n1069);
nand (n1074,n1075,n913);
not (n1075,n1073);
or (n1076,n910,n3);
xor (n1077,n1078,n1404);
xor (n1078,n1079,n1075);
xor (n1079,n1080,n1379);
xor (n1080,n1081,n1230);
xor (n1081,n1082,n1229);
xor (n1082,n1083,n1227);
xor (n1083,n1084,n1226);
xor (n1084,n1085,n1218);
xor (n1085,n1086,n1217);
xor (n1086,n1087,n1203);
xor (n1087,n1088,n1202);
xor (n1088,n1089,n1184);
xor (n1089,n1090,n590);
xor (n1090,n1091,n1163);
xor (n1091,n1092,n1162);
xor (n1092,n1093,n1142);
xor (n1093,n1094,n1141);
xor (n1094,n1095,n1120);
xor (n1095,n1096,n1119);
xor (n1096,n1097,n1100);
xor (n1097,n1098,n1099);
and (n1098,n932,n121);
and (n1099,n652,n119);
or (n1100,n1101,n1103);
and (n1101,n1102,n524);
and (n1102,n652,n121);
and (n1103,n1104,n1105);
xor (n1104,n1102,n524);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
and (n1107,n525,n121);
and (n1108,n414,n119);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1114);
and (n1112,n1113,n215);
and (n1113,n414,n121);
and (n1114,n1115,n1116);
xor (n1115,n1113,n215);
or (n1116,n1117,n1118);
and (n1117,n715,n716);
and (n1118,n714,n717);
and (n1119,n525,n141);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1104,n1105);
and (n1123,n414,n141);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1110,n1111);
and (n1129,n216,n141);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
xor (n1134,n1115,n1116);
and (n1135,n133,n141);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1140);
and (n1139,n713,n735);
and (n1140,n712,n736);
and (n1141,n414,n44);
or (n1142,n1143,n1145);
and (n1143,n1144,n537);
xor (n1144,n1125,n1126);
and (n1145,n1146,n1147);
xor (n1146,n1144,n537);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
xor (n1149,n1131,n1132);
and (n1150,n133,n44);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
xor (n1155,n1137,n1138);
and (n1156,n125,n44);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1161);
and (n1160,n711,n750);
and (n1161,n710,n751);
and (n1162,n216,n37);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
xor (n1165,n1146,n1147);
and (n1166,n133,n37);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1152,n1153);
and (n1172,n125,n37);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1158,n1159);
and (n1178,n168,n37);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1183);
and (n1182,n709,n759);
and (n1183,n708,n760);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1168,n1169);
and (n1187,n125,n30);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1174,n1175);
and (n1193,n168,n30);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
or (n1196,n1197,n1199);
and (n1197,n1198,n51);
xor (n1198,n1180,n1181);
and (n1199,n1200,n1201);
xor (n1200,n1198,n51);
and (n1201,n707,n762);
and (n1202,n125,n422);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1189,n1190);
and (n1206,n168,n422);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1195,n1196);
and (n1212,n50,n422);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
and (n1215,n1216,n461);
xor (n1216,n1200,n1201);
and (n1217,n168,n465);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1208,n1209);
and (n1221,n50,n465);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
and (n1224,n1225,n477);
xor (n1225,n1214,n1215);
and (n1226,n50,n638);
and (n1227,n1228,n1024);
xor (n1228,n1223,n1224);
and (n1229,n28,n950);
not (n1230,n1231);
xor (n1231,n1232,n984);
xor (n1232,n1233,n1376);
xor (n1233,n1234,n1375);
xor (n1234,n1235,n1368);
xor (n1235,n1236,n629);
xor (n1236,n1237,n1353);
xor (n1237,n1238,n1352);
xor (n1238,n1239,n1334);
xor (n1239,n1240,n1333);
xor (n1240,n1241,n1312);
xor (n1241,n1242,n1311);
xor (n1242,n1243,n1291);
xor (n1243,n1244,n1290);
xor (n1244,n1245,n1269);
xor (n1245,n1246,n1268);
xor (n1246,n1247,n1250);
xor (n1247,n1248,n1249);
and (n1248,n1005,n176);
and (n1249,n597,n68);
or (n1250,n1251,n1253);
and (n1251,n1252,n557);
and (n1252,n597,n176);
and (n1253,n1254,n1255);
xor (n1254,n1252,n557);
or (n1255,n1256,n1258);
and (n1256,n1257,n393);
and (n1257,n558,n176);
and (n1258,n1259,n1260);
xor (n1259,n1257,n393);
or (n1260,n1261,n1263);
and (n1261,n1262,n238);
and (n1262,n392,n176);
and (n1263,n1264,n1265);
xor (n1264,n1262,n238);
or (n1265,n1266,n1267);
and (n1266,n773,n774);
and (n1267,n772,n775);
and (n1268,n558,n69);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1254,n1255);
and (n1272,n392,n69);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1259,n1260);
and (n1278,n237,n69);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1264,n1265);
and (n1284,n180,n69);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1289);
and (n1288,n771,n794);
and (n1289,n770,n795);
and (n1290,n392,n60);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1274,n1275);
and (n1294,n237,n60);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
or (n1297,n1298,n1301);
and (n1298,n1299,n1300);
xor (n1299,n1280,n1281);
and (n1300,n180,n60);
and (n1301,n1302,n1303);
xor (n1302,n1299,n1300);
or (n1303,n1304,n1306);
and (n1304,n1305,n80);
xor (n1305,n1286,n1287);
and (n1306,n1307,n1308);
xor (n1307,n1305,n80);
or (n1308,n1309,n1310);
and (n1309,n769,n810);
and (n1310,n768,n811);
and (n1311,n237,n86);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1296,n1297);
and (n1315,n180,n86);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1322);
and (n1319,n1320,n1321);
xor (n1320,n1302,n1303);
and (n1321,n79,n86);
and (n1322,n1323,n1324);
xor (n1323,n1320,n1321);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1307,n1308);
and (n1327,n58,n86);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1332);
and (n1331,n767,n818);
and (n1332,n766,n819);
and (n1333,n180,n91);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1317,n1318);
and (n1337,n79,n91);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1323,n1324);
and (n1343,n58,n91);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
or (n1346,n1347,n1349);
and (n1347,n1348,n94);
xor (n1348,n1329,n1330);
and (n1349,n1350,n1351);
xor (n1350,n1348,n94);
and (n1351,n765,n105);
and (n1352,n79,n428);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1339,n1340);
and (n1356,n58,n428);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
or (n1359,n1360,n1363);
and (n1360,n1361,n1362);
xor (n1361,n1345,n1346);
and (n1362,n92,n428);
and (n1363,n1364,n1365);
xor (n1364,n1361,n1362);
and (n1365,n1366,n1367);
xor (n1366,n1350,n1351);
and (n1367,n104,n428);
or (n1368,n1369,n1371);
and (n1369,n1370,n506);
xor (n1370,n1358,n1359);
and (n1371,n1372,n1373);
xor (n1372,n1370,n506);
and (n1373,n1374,n512);
xor (n1374,n1364,n1365);
and (n1375,n92,n643);
and (n1376,n1377,n1378);
xor (n1377,n1372,n1373);
and (n1378,n104,n643);
or (n1379,n1380,n1384,n1403);
and (n1380,n1381,n1382);
xor (n1381,n1228,n1024);
not (n1382,n1383);
xor (n1383,n1377,n1378);
and (n1384,n1382,n1385);
or (n1385,n1386,n1390,n1402);
and (n1386,n1387,n1388);
xor (n1387,n1225,n477);
not (n1388,n1389);
xor (n1389,n1374,n512);
and (n1390,n1388,n1391);
or (n1391,n1392,n1396,n1401);
and (n1392,n1393,n1394);
xor (n1393,n1216,n461);
not (n1394,n1395);
xor (n1395,n1366,n1367);
and (n1396,n1394,n1397);
or (n1397,n1398,n1399,n1400);
and (n1398,n706,n763);
and (n1399,n763,n822);
and (n1400,n706,n822);
and (n1401,n1393,n1397);
and (n1402,n1387,n1391);
and (n1403,n1381,n1385);
or (n1404,n1405,n1408,n1421);
and (n1405,n1406,n6);
xor (n1406,n1407,n1385);
xor (n1407,n1381,n1382);
and (n1408,n6,n1409);
or (n1409,n1410,n1413,n1420);
and (n1410,n1411,n906);
xor (n1411,n1412,n1391);
xor (n1412,n1387,n1388);
and (n1413,n906,n1414);
or (n1414,n1415,n1418,n1419);
and (n1415,n1416,n694);
xor (n1416,n1417,n1397);
xor (n1417,n1393,n1394);
and (n1418,n694,n702);
and (n1419,n1416,n702);
and (n1420,n1411,n1414);
and (n1421,n1406,n1409);
endmodule
