module top (out,n3,n20,n21,n24,n25,n32,n33,n35,n36
        ,n53,n71,n72,n74,n75,n94,n134,n140,n149,n158
        ,n159,n165,n166,n171,n178,n184,n197,n198,n202,n207
        ,n225,n268,n349,n399,n598,n1026);
output out;
input n3;
input n20;
input n21;
input n24;
input n25;
input n32;
input n33;
input n35;
input n36;
input n53;
input n71;
input n72;
input n74;
input n75;
input n94;
input n134;
input n140;
input n149;
input n158;
input n159;
input n165;
input n166;
input n171;
input n178;
input n184;
input n197;
input n198;
input n202;
input n207;
input n225;
input n268;
input n349;
input n399;
input n598;
input n1026;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n167;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
xnor (out,n0,n1027);
nand (n0,n1,n1026);
nand (n1,n2,n1017);
or (n2,n3,n4);
not (n4,n5);
nand (n5,n6,n1016);
or (n6,n7,n111);
not (n7,n8);
nor (n8,n9,n110);
and (n9,n10,n98);
not (n10,n11);
or (n11,n12,n97);
and (n12,n13,n59);
xor (n13,n14,n48);
nand (n14,n15,n39);
or (n15,n16,n28);
not (n16,n17);
nand (n17,n18,n26);
or (n18,n19,n22);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n3);
and (s0n19,notn19,n20);
and (s1n19,n3,n21);
not (n22,n23);
and (n23,n24,n25);
or (n26,n27,n23);
not (n27,n19);
nor (n28,n29,n37);
and (n29,n30,n34);
not (n30,n31);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n3);
and (s0n31,notn31,n32);
and (s1n31,n3,n33);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n3);
and (s0n34,notn34,n35);
and (s1n34,n3,n36);
and (n37,n31,n38);
not (n38,n34);
or (n39,n40,n44);
nand (n40,n28,n41);
nand (n41,n42,n43);
or (n42,n30,n19);
nand (n43,n19,n30);
nor (n44,n45,n46);
and (n45,n27,n25);
and (n46,n19,n47);
not (n47,n25);
nand (n48,n49,n54,n56);
or (n49,n50,n53);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n3);
and (s0n50,notn50,1'b0);
and (s1n50,n3,n52);
and (n52,n24,n21);
not (n54,n55);
and (n55,n53,n50);
not (n56,n57);
nand (n57,n19,n58);
not (n58,n50);
or (n59,n60,n96);
and (n60,n61,n90);
xor (n61,n62,n83);
nand (n62,n63,n80);
or (n63,n64,n67);
not (n64,n65);
nand (n65,n66,n77);
not (n66,n67);
nand (n67,n68,n76);
or (n68,n69,n73);
not (n69,n70);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n3);
and (s0n70,notn70,n71);
and (s1n70,n3,n72);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n3);
and (s0n73,notn73,n74);
and (s1n73,n3,n75);
nand (n76,n73,n69);
nand (n77,n78,n79);
or (n78,n69,n34);
nand (n79,n34,n69);
nand (n80,n81,n82);
or (n81,n34,n22);
or (n82,n38,n23);
nand (n83,n84,n89);
or (n84,n40,n85);
nor (n85,n86,n87);
and (n86,n27,n53);
and (n87,n19,n88);
not (n88,n53);
or (n89,n28,n44);
nor (n90,n57,n91);
nor (n91,n92,n95);
and (n92,n50,n93);
not (n93,n94);
and (n95,n58,n94);
and (n96,n62,n83);
and (n97,n14,n48);
not (n98,n99);
xor (n99,n100,n109);
xor (n100,n101,n105);
nand (n101,n102,n17);
or (n102,n103,n104);
not (n103,n40);
not (n104,n28);
nor (n105,n57,n106);
nor (n106,n107,n108);
and (n107,n50,n47);
and (n108,n58,n25);
not (n109,n48);
and (n110,n11,n99);
nand (n111,n112,n992,n1015);
nand (n112,n113,n769);
nand (n113,n114,n758,n768);
nand (n114,n115,n561);
nand (n115,n116,n417,n560);
nand (n116,n117,n368);
nand (n117,n118,n367);
or (n118,n119,n320);
nor (n119,n120,n319);
and (n120,n121,n291);
not (n121,n122);
nor (n122,n123,n249);
or (n123,n124,n248);
and (n124,n125,n217);
xor (n125,n126,n188);
or (n126,n127,n187);
and (n127,n128,n174);
xor (n128,n129,n143);
nand (n129,n130,n137);
or (n130,n131,n40);
not (n131,n132);
nand (n132,n133,n135);
or (n133,n27,n134);
or (n135,n19,n136);
not (n136,n134);
or (n137,n28,n138);
nor (n138,n139,n141);
and (n139,n140,n27);
and (n141,n142,n19);
not (n142,n140);
nand (n143,n144,n168);
or (n144,n145,n152);
not (n145,n146);
nand (n146,n147,n150);
or (n147,n73,n148);
not (n148,n149);
or (n150,n151,n149);
not (n151,n73);
not (n152,n153);
and (n153,n154,n161);
nand (n154,n155,n160);
or (n155,n156,n73);
not (n156,n157);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n3);
and (s0n157,notn157,n158);
and (s1n157,n3,n159);
nand (n160,n73,n156);
not (n161,n162);
nand (n162,n163,n167);
or (n163,n156,n164);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n3);
and (s0n164,notn164,n165);
and (s1n164,n3,n166);
nand (n167,n164,n156);
nand (n168,n162,n169);
nor (n169,n170,n172);
and (n170,n171,n73);
and (n172,n173,n151);
not (n173,n171);
nand (n174,n175,n181);
or (n175,n65,n176);
nor (n176,n177,n179);
and (n177,n38,n178);
and (n179,n34,n180);
not (n180,n178);
or (n181,n66,n182);
nor (n182,n183,n185);
and (n183,n38,n184);
and (n185,n34,n186);
not (n186,n184);
and (n187,n129,n143);
xor (n188,n189,n211);
xor (n189,n190,n191);
and (n190,n56,n134);
nand (n191,n192,n204);
or (n192,n193,n199);
not (n193,n194);
nor (n194,n195,n196);
not (n195,n164);
wire s0n196,s1n196,notn196;
or (n196,s0n196,s1n196);
not(notn196,n3);
and (s0n196,notn196,n197);
and (s1n196,n3,n198);
nor (n199,n200,n203);
and (n200,n201,n164);
not (n201,n202);
and (n203,n202,n195);
or (n204,n205,n210);
nor (n205,n206,n208);
and (n206,n195,n207);
and (n208,n164,n209);
not (n209,n207);
not (n210,n196);
nand (n211,n212,n213);
or (n212,n40,n138);
or (n213,n28,n214);
nor (n214,n215,n216);
and (n215,n178,n27);
and (n216,n180,n19);
xor (n217,n218,n234);
xor (n218,n219,n228);
nand (n219,n220,n222);
or (n220,n152,n221);
not (n221,n169);
or (n222,n161,n223);
nor (n223,n224,n226);
and (n224,n151,n225);
and (n226,n73,n227);
not (n227,n225);
nand (n228,n229,n230);
or (n229,n65,n182);
or (n230,n66,n231);
nor (n231,n232,n233);
and (n232,n38,n149);
and (n233,n34,n148);
and (n234,n235,n240);
nor (n235,n236,n27);
nor (n236,n237,n239);
and (n237,n38,n238);
nand (n238,n31,n134);
and (n239,n30,n136);
nand (n240,n241,n246);
or (n241,n242,n193);
not (n242,n243);
nor (n243,n244,n245);
and (n244,n225,n164);
and (n245,n227,n195);
nand (n246,n247,n196);
not (n247,n199);
and (n248,n126,n188);
xor (n249,n250,n274);
xor (n250,n251,n271);
xor (n251,n252,n263);
xor (n252,n253,n259);
nand (n253,n254,n255);
or (n254,n214,n40);
nand (n255,n256,n104);
nor (n256,n257,n258);
and (n257,n184,n19);
and (n258,n186,n27);
nor (n259,n57,n260);
nor (n260,n261,n262);
and (n261,n50,n142);
and (n262,n58,n140);
nand (n263,n264,n265);
or (n264,n193,n205);
or (n265,n266,n210);
nor (n266,n267,n269);
and (n267,n195,n268);
and (n269,n164,n270);
not (n270,n268);
or (n271,n272,n273);
and (n272,n218,n234);
and (n273,n219,n228);
xor (n274,n275,n288);
xor (n275,n276,n282);
nand (n276,n277,n278);
or (n277,n65,n231);
or (n278,n66,n279);
nor (n279,n280,n281);
and (n280,n38,n171);
and (n281,n34,n173);
nand (n282,n283,n284);
or (n283,n152,n223);
or (n284,n285,n161);
nor (n285,n286,n287);
and (n286,n151,n202);
and (n287,n73,n201);
or (n288,n289,n290);
and (n289,n189,n211);
and (n290,n190,n191);
not (n291,n292);
nand (n292,n293,n294);
xor (n293,n125,n217);
or (n294,n295,n318);
and (n295,n296,n317);
xor (n296,n297,n298);
xor (n297,n235,n240);
or (n298,n299,n316);
and (n299,n300,n309);
xor (n300,n301,n302);
and (n301,n104,n134);
nand (n302,n303,n304);
or (n303,n210,n242);
nand (n304,n305,n194);
not (n305,n306);
nor (n306,n307,n308);
and (n307,n171,n195);
and (n308,n173,n164);
nand (n309,n310,n315);
or (n310,n311,n152);
not (n311,n312);
nor (n312,n313,n314);
and (n313,n184,n73);
and (n314,n151,n186);
nand (n315,n162,n146);
and (n316,n301,n302);
xor (n317,n128,n174);
and (n318,n297,n298);
and (n319,n123,n249);
nor (n320,n321,n364);
xor (n321,n322,n361);
xor (n322,n323,n342);
xor (n323,n324,n336);
xor (n324,n325,n332);
nand (n325,n326,n328);
or (n326,n327,n40);
not (n327,n256);
nand (n328,n104,n329);
nor (n329,n330,n331);
and (n330,n149,n19);
and (n331,n148,n27);
nor (n332,n57,n333);
nor (n333,n334,n335);
and (n334,n50,n180);
and (n335,n58,n178);
nand (n336,n337,n338);
or (n337,n65,n279);
or (n338,n66,n339);
nor (n339,n340,n341);
and (n340,n38,n225);
and (n341,n34,n227);
xor (n342,n343,n358);
xor (n343,n344,n352);
nand (n344,n345,n346);
or (n345,n193,n266);
or (n346,n347,n210);
nor (n347,n348,n350);
and (n348,n195,n349);
and (n350,n164,n351);
not (n351,n349);
nand (n352,n353,n354);
or (n353,n152,n285);
or (n354,n355,n161);
nor (n355,n356,n357);
and (n356,n151,n207);
and (n357,n73,n209);
or (n358,n359,n360);
and (n359,n252,n263);
and (n360,n253,n259);
or (n361,n362,n363);
and (n362,n275,n288);
and (n363,n276,n282);
or (n364,n365,n366);
and (n365,n250,n274);
and (n366,n251,n271);
nand (n367,n321,n364);
nand (n368,n369,n413);
not (n369,n370);
xor (n370,n371,n412);
xor (n371,n372,n391);
xor (n372,n373,n385);
xor (n373,n374,n381);
nand (n374,n375,n377);
or (n375,n376,n40);
not (n376,n329);
nand (n377,n104,n378);
nor (n378,n379,n380);
and (n379,n171,n19);
and (n380,n173,n27);
nor (n381,n57,n382);
nor (n382,n383,n384);
and (n383,n50,n186);
and (n384,n58,n184);
nand (n385,n386,n387);
or (n386,n65,n339);
or (n387,n66,n388);
nor (n388,n389,n390);
and (n389,n38,n202);
and (n390,n34,n201);
xor (n391,n392,n409);
xor (n392,n393,n408);
xor (n393,n394,n402);
nand (n394,n395,n396);
or (n395,n193,n347);
or (n396,n397,n210);
nor (n397,n398,n400);
and (n398,n195,n399);
and (n400,n164,n401);
not (n401,n399);
nand (n402,n403,n404);
or (n403,n152,n355);
or (n404,n161,n405);
nor (n405,n406,n407);
and (n406,n151,n268);
and (n407,n73,n270);
and (n408,n344,n352);
or (n409,n410,n411);
and (n410,n324,n336);
and (n411,n325,n332);
and (n412,n343,n358);
not (n413,n414);
or (n414,n415,n416);
and (n415,n322,n361);
and (n416,n323,n342);
nand (n417,n368,n418,n559);
nor (n418,n419,n556);
nor (n419,n420,n554);
and (n420,n421,n549);
or (n421,n422,n548);
and (n422,n423,n464);
xor (n423,n424,n457);
or (n424,n425,n456);
and (n425,n426,n444);
xor (n426,n427,n434);
nand (n427,n428,n433);
or (n428,n429,n152);
not (n429,n430);
nor (n430,n431,n432);
and (n431,n180,n151);
and (n432,n178,n73);
nand (n433,n162,n312);
nand (n434,n435,n440);
or (n435,n436,n66);
not (n436,n437);
nor (n437,n438,n439);
and (n438,n140,n34);
and (n439,n142,n38);
nand (n440,n64,n441);
nand (n441,n442,n443);
or (n442,n38,n134);
or (n443,n34,n136);
xor (n444,n445,n450);
and (n445,n446,n34);
nand (n446,n447,n449);
or (n447,n73,n448);
and (n448,n134,n70);
or (n449,n70,n134);
nand (n450,n451,n455);
or (n451,n193,n452);
nor (n452,n453,n454);
and (n453,n195,n149);
and (n454,n164,n148);
or (n455,n306,n210);
and (n456,n427,n434);
xor (n457,n458,n463);
xor (n458,n459,n462);
nand (n459,n460,n461);
or (n460,n436,n65);
or (n461,n66,n176);
and (n462,n445,n450);
xor (n463,n300,n309);
or (n464,n465,n547);
and (n465,n466,n487);
xor (n466,n467,n486);
or (n467,n468,n485);
and (n468,n469,n478);
xor (n469,n470,n471);
and (n470,n67,n134);
nand (n471,n472,n477);
or (n472,n473,n152);
not (n473,n474);
nor (n474,n475,n476);
and (n475,n140,n73);
and (n476,n142,n151);
nand (n477,n430,n162);
nand (n478,n479,n484);
or (n479,n193,n480);
not (n480,n481);
nor (n481,n482,n483);
and (n482,n186,n195);
and (n483,n184,n164);
or (n484,n452,n210);
and (n485,n470,n471);
xor (n486,n426,n444);
or (n487,n488,n546);
and (n488,n489,n545);
xor (n489,n490,n504);
nor (n490,n491,n499);
not (n491,n492);
nand (n492,n493,n498);
or (n493,n494,n193);
not (n494,n495);
nand (n495,n496,n497);
or (n496,n180,n164);
nand (n497,n164,n180);
nand (n498,n481,n196);
nand (n499,n500,n73);
nand (n500,n501,n503);
or (n501,n164,n502);
and (n502,n134,n157);
or (n503,n157,n134);
nand (n504,n505,n543);
or (n505,n506,n529);
not (n506,n507);
nand (n507,n508,n528);
or (n508,n509,n518);
nor (n509,n510,n517);
nand (n510,n511,n516);
or (n511,n512,n193);
not (n512,n513);
nand (n513,n514,n515);
or (n514,n142,n164);
nand (n515,n164,n142);
nand (n516,n495,n196);
nor (n517,n161,n136);
nand (n518,n519,n526);
nand (n519,n520,n525);
or (n520,n521,n193);
not (n521,n522);
nand (n522,n523,n524);
or (n523,n195,n134);
or (n524,n164,n136);
nand (n525,n513,n196);
nor (n526,n527,n195);
and (n527,n134,n196);
nand (n528,n510,n517);
not (n529,n530);
nand (n530,n531,n539);
not (n531,n532);
nand (n532,n533,n538);
or (n533,n534,n152);
not (n534,n535);
nand (n535,n536,n537);
or (n536,n151,n134);
or (n537,n73,n136);
nand (n538,n162,n474);
nor (n539,n540,n542);
and (n540,n491,n541);
not (n541,n499);
and (n542,n492,n499);
nand (n543,n544,n532);
not (n544,n539);
xor (n545,n469,n478);
and (n546,n490,n504);
and (n547,n467,n486);
and (n548,n424,n457);
or (n549,n550,n551);
xor (n550,n296,n317);
or (n551,n552,n553);
and (n552,n458,n463);
and (n553,n459,n462);
not (n554,n555);
nand (n555,n550,n551);
nand (n556,n557,n121);
not (n557,n558);
nor (n558,n293,n294);
not (n559,n320);
nand (n560,n370,n414);
nor (n561,n562,n662);
nand (n562,n563,n655);
not (n563,n564);
nor (n564,n565,n646);
xor (n565,n566,n637);
xor (n566,n567,n591);
xor (n567,n568,n582);
xor (n568,n569,n578);
nand (n569,n570,n574);
or (n570,n40,n571);
nor (n571,n572,n573);
and (n572,n27,n225);
and (n573,n19,n227);
or (n574,n28,n575);
nor (n575,n576,n577);
and (n576,n202,n27);
and (n577,n201,n19);
nor (n578,n57,n579);
nor (n579,n580,n581);
and (n580,n50,n173);
and (n581,n58,n171);
nand (n582,n583,n587);
or (n583,n584,n66);
nor (n584,n585,n586);
and (n585,n38,n268);
and (n586,n34,n270);
or (n587,n65,n588);
nor (n588,n589,n590);
and (n589,n38,n207);
and (n590,n34,n209);
xor (n591,n592,n621);
xor (n592,n593,n614);
xor (n593,n594,n605);
nand (n594,n595,n601);
or (n595,n193,n596);
nor (n596,n597,n599);
and (n597,n195,n598);
and (n599,n164,n600);
not (n600,n598);
or (n601,n602,n210);
nor (n602,n603,n604);
and (n603,n195,n94);
and (n604,n164,n93);
nand (n605,n606,n610);
or (n606,n152,n607);
nor (n607,n608,n609);
and (n608,n151,n349);
and (n609,n73,n351);
or (n610,n611,n161);
nor (n611,n612,n613);
and (n612,n151,n399);
and (n613,n73,n401);
and (n614,n615,n618);
nand (n615,n616,n617);
or (n616,n193,n397);
or (n617,n596,n210);
nand (n618,n619,n620);
or (n619,n152,n405);
or (n620,n607,n161);
or (n621,n622,n636);
and (n622,n623,n633);
xor (n623,n624,n629);
nand (n624,n625,n627);
or (n625,n626,n40);
not (n626,n378);
nand (n627,n628,n104);
not (n628,n571);
nor (n629,n57,n630);
nor (n630,n631,n632);
and (n631,n50,n148);
and (n632,n58,n149);
nand (n633,n634,n635);
or (n634,n65,n388);
or (n635,n66,n588);
and (n636,n624,n629);
or (n637,n638,n645);
and (n638,n639,n642);
xor (n639,n640,n641);
xor (n640,n615,n618);
and (n641,n394,n402);
or (n642,n643,n644);
and (n643,n373,n385);
and (n644,n374,n381);
and (n645,n640,n641);
or (n646,n647,n654);
and (n647,n648,n651);
xor (n648,n649,n650);
xor (n649,n623,n633);
xor (n650,n639,n642);
or (n651,n652,n653);
and (n652,n392,n409);
and (n653,n393,n408);
and (n654,n649,n650);
nand (n655,n656,n658);
not (n656,n657);
xor (n657,n648,n651);
not (n658,n659);
or (n659,n660,n661);
and (n660,n371,n412);
and (n661,n372,n391);
nand (n662,n663,n711);
nand (n663,n664,n707);
not (n664,n665);
xor (n665,n666,n704);
xor (n666,n667,n685);
xor (n667,n668,n679);
xor (n668,n669,n675);
nand (n669,n670,n671);
or (n670,n575,n40);
nand (n671,n104,n672);
nor (n672,n673,n674);
and (n673,n207,n19);
and (n674,n209,n27);
nor (n675,n57,n676);
nor (n676,n677,n678);
and (n677,n50,n227);
and (n678,n58,n225);
nand (n679,n680,n681);
or (n680,n65,n584);
or (n681,n66,n682);
nor (n682,n683,n684);
and (n683,n38,n349);
and (n684,n34,n351);
xor (n685,n686,n701);
xor (n686,n687,n700);
xor (n687,n688,n694);
nand (n688,n689,n690);
or (n689,n193,n602);
or (n690,n691,n210);
nor (n691,n692,n693);
and (n692,n195,n53);
and (n693,n164,n88);
nand (n694,n695,n696);
or (n695,n152,n611);
or (n696,n161,n697);
nor (n697,n698,n699);
and (n698,n151,n598);
and (n699,n73,n600);
and (n700,n594,n605);
or (n701,n702,n703);
and (n702,n568,n582);
and (n703,n569,n578);
or (n704,n705,n706);
and (n705,n592,n621);
and (n706,n593,n614);
not (n707,n708);
or (n708,n709,n710);
and (n709,n566,n637);
and (n710,n567,n591);
nand (n711,n712,n754);
not (n712,n713);
xor (n713,n714,n751);
xor (n714,n715,n734);
xor (n715,n716,n728);
xor (n716,n717,n724);
nand (n717,n718,n720);
or (n718,n719,n40);
not (n719,n672);
nand (n720,n104,n721);
nor (n721,n722,n723);
and (n722,n268,n19);
and (n723,n270,n27);
nor (n724,n57,n725);
nor (n725,n726,n727);
and (n726,n50,n201);
and (n727,n58,n202);
nand (n728,n729,n730);
or (n729,n65,n682);
or (n730,n66,n731);
nor (n731,n732,n733);
and (n732,n38,n399);
and (n733,n34,n401);
xor (n734,n735,n748);
xor (n735,n736,n747);
xor (n736,n737,n743);
nand (n737,n738,n739);
or (n738,n193,n691);
or (n739,n740,n210);
nor (n740,n741,n742);
and (n741,n195,n25);
and (n742,n164,n47);
nand (n743,n744,n745);
or (n744,n152,n697);
or (n745,n746,n161);
xor (n746,n94,n151);
and (n747,n688,n694);
or (n748,n749,n750);
and (n749,n668,n679);
and (n750,n669,n675);
or (n751,n752,n753);
and (n752,n686,n701);
and (n753,n687,n700);
not (n754,n755);
or (n755,n756,n757);
and (n756,n666,n704);
and (n757,n667,n685);
nand (n758,n759,n711);
nand (n759,n760,n767);
or (n760,n761,n762);
not (n761,n663);
not (n762,n763);
nand (n763,n764,n766);
or (n764,n564,n765);
nand (n765,n657,n659);
nand (n766,n565,n646);
nand (n767,n665,n708);
nand (n768,n755,n713);
and (n769,n770,n948,n987);
and (n770,n771,n870,n942);
nor (n771,n772,n819);
nor (n772,n773,n776);
or (n773,n774,n775);
and (n774,n714,n751);
and (n775,n715,n734);
xor (n776,n777,n816);
xor (n777,n778,n797);
xor (n778,n779,n791);
xor (n779,n780,n787);
nand (n780,n781,n783);
or (n781,n782,n40);
not (n782,n721);
or (n783,n28,n784);
nor (n784,n785,n786);
and (n785,n27,n349);
and (n786,n19,n351);
nor (n787,n57,n788);
nor (n788,n789,n790);
and (n789,n50,n209);
and (n790,n58,n207);
nand (n791,n792,n793);
or (n792,n65,n731);
or (n793,n66,n794);
nor (n794,n795,n796);
and (n795,n38,n598);
and (n796,n34,n600);
xor (n797,n798,n813);
xor (n798,n799,n812);
xor (n799,n800,n806);
nand (n800,n801,n802);
or (n801,n193,n740);
or (n802,n803,n210);
nor (n803,n804,n805);
and (n804,n195,n23);
and (n805,n164,n22);
nand (n806,n807,n808);
or (n807,n746,n152);
nand (n808,n162,n809);
nand (n809,n810,n811);
or (n810,n73,n88);
or (n811,n151,n53);
and (n812,n737,n743);
or (n813,n814,n815);
and (n814,n716,n728);
and (n815,n717,n724);
or (n816,n817,n818);
and (n817,n735,n748);
and (n818,n736,n747);
not (n819,n820);
nand (n820,n821,n866);
not (n821,n822);
xor (n822,n823,n842);
xor (n823,n824,n839);
xor (n824,n825,n833);
xor (n825,n826,n830);
nor (n826,n57,n827);
nor (n827,n828,n829);
and (n828,n50,n270);
and (n829,n58,n268);
nand (n830,n831,n832);
or (n831,n196,n194);
not (n832,n803);
nand (n833,n834,n838);
or (n834,n835,n66);
nor (n835,n836,n837);
and (n836,n94,n38);
and (n837,n93,n34);
or (n838,n65,n794);
or (n839,n840,n841);
and (n840,n798,n813);
and (n841,n799,n812);
xor (n842,n843,n848);
xor (n843,n844,n845);
and (n844,n800,n806);
or (n845,n846,n847);
and (n846,n779,n791);
and (n847,n780,n787);
nand (n848,n849,n865);
or (n849,n850,n858);
not (n850,n851);
nand (n851,n852,n854);
or (n852,n152,n853);
not (n853,n809);
or (n854,n161,n855);
nor (n855,n856,n857);
and (n856,n151,n25);
and (n857,n73,n47);
not (n858,n859);
nand (n859,n860,n861);
or (n860,n40,n784);
or (n861,n28,n862);
nor (n862,n863,n864);
and (n863,n27,n399);
and (n864,n19,n401);
or (n865,n859,n851);
not (n866,n867);
or (n867,n868,n869);
and (n868,n777,n816);
and (n869,n778,n797);
nand (n870,n871,n932);
not (n871,n872);
xor (n872,n873,n924);
xor (n873,n874,n894);
xor (n874,n875,n890);
xor (n875,n876,n881);
nand (n876,n877,n878);
or (n877,n153,n162);
nand (n878,n879,n880);
or (n879,n73,n22);
or (n880,n151,n23);
nand (n881,n882,n886);
or (n882,n65,n883);
nor (n883,n884,n885);
and (n884,n38,n53);
and (n885,n34,n88);
or (n886,n66,n887);
nor (n887,n888,n889);
and (n888,n38,n25);
and (n889,n34,n47);
nor (n890,n57,n891);
nor (n891,n892,n893);
and (n892,n50,n401);
and (n893,n58,n399);
xor (n894,n895,n910);
xor (n895,n896,n905);
nand (n896,n897,n901);
or (n897,n40,n898);
nor (n898,n899,n900);
and (n899,n27,n598);
and (n900,n19,n600);
or (n901,n28,n902);
nor (n902,n903,n904);
and (n903,n27,n94);
and (n904,n19,n93);
nand (n905,n906,n908);
or (n906,n907,n161);
not (n907,n878);
nand (n908,n909,n153);
not (n909,n855);
or (n910,n911,n923);
and (n911,n912,n920);
xor (n912,n913,n917);
nor (n913,n57,n914);
nor (n914,n915,n916);
and (n915,n50,n351);
and (n916,n58,n349);
nand (n917,n918,n919);
or (n918,n65,n835);
or (n919,n66,n883);
nand (n920,n921,n922);
or (n921,n40,n862);
or (n922,n28,n898);
and (n923,n913,n917);
or (n924,n925,n931);
and (n925,n926,n928);
xor (n926,n927,n865);
not (n927,n905);
or (n928,n929,n930);
and (n929,n825,n833);
and (n930,n826,n830);
and (n931,n927,n865);
not (n932,n933);
or (n933,n934,n941);
and (n934,n935,n938);
xor (n935,n936,n937);
xor (n936,n912,n920);
xor (n937,n926,n928);
or (n938,n939,n940);
and (n939,n843,n848);
and (n940,n844,n845);
and (n941,n936,n937);
not (n942,n943);
nor (n943,n944,n945);
xor (n944,n935,n938);
or (n945,n946,n947);
and (n946,n823,n842);
and (n947,n824,n839);
nor (n948,n949,n974);
nor (n949,n950,n953);
or (n950,n951,n952);
and (n951,n873,n924);
and (n952,n874,n894);
xor (n953,n954,n971);
xor (n954,n955,n958);
or (n955,n956,n957);
and (n956,n875,n890);
and (n957,n876,n881);
xor (n958,n959,n967);
xor (n959,n960,n963);
nand (n960,n961,n962);
or (n961,n40,n902);
or (n962,n28,n85);
nor (n963,n57,n964);
nor (n964,n965,n966);
and (n965,n50,n600);
and (n966,n58,n598);
nor (n967,n968,n970);
and (n968,n64,n969);
not (n969,n887);
and (n970,n67,n80);
or (n971,n972,n973);
and (n972,n895,n910);
and (n973,n896,n905);
and (n974,n975,n979);
not (n975,n976);
or (n976,n977,n978);
and (n977,n954,n971);
and (n978,n955,n958);
not (n979,n980);
xor (n980,n981,n984);
xor (n981,n982,n983);
not (n982,n967);
xor (n983,n61,n90);
or (n984,n985,n986);
and (n985,n959,n967);
and (n986,n960,n963);
or (n987,n988,n991);
or (n988,n989,n990);
and (n989,n981,n984);
and (n990,n982,n983);
xor (n991,n13,n59);
nand (n992,n993,n987);
nand (n993,n994,n1009);
or (n994,n995,n996);
not (n995,n948);
not (n996,n997);
nand (n997,n998,n1008);
or (n998,n999,n1000);
not (n999,n870);
not (n1000,n1001);
nand (n1001,n1002,n1007);
or (n1002,n1003,n943);
nor (n1003,n1004,n1006);
and (n1004,n1005,n820);
and (n1005,n773,n776);
nor (n1006,n821,n866);
nand (n1007,n944,n945);
or (n1008,n871,n932);
nor (n1009,n1010,n1014);
and (n1010,n1011,n1013);
not (n1011,n1012);
nand (n1012,n950,n953);
not (n1013,n974);
nor (n1014,n975,n979);
nand (n1015,n988,n991);
nand (n1016,n7,n111);
nand (n1017,n1018,n3);
xor (n1018,n1019,n1020);
nand (n1019,n711,n768);
nor (n1020,n1021,n1025);
and (n1021,n1022,n663);
nand (n1022,n1023,n762);
or (n1023,n562,n1024);
not (n1024,n115);
not (n1025,n767);
and (n1027,n1026,n1028);
wire s0n1028,s1n1028,notn1028;
or (n1028,s0n1028,s1n1028);
not(notn1028,n3);
and (s0n1028,notn1028,n1029);
and (s1n1028,n3,n2328);
xor (n1029,n1030,n1844);
xor (n1030,n1031,n2326);
xor (n1031,n1032,n1839);
xor (n1032,n1033,n2319);
xor (n1033,n1034,n1833);
xor (n1034,n1035,n2307);
xor (n1035,n1036,n1827);
xor (n1036,n1037,n2290);
xor (n1037,n1038,n1821);
xor (n1038,n1039,n2268);
xor (n1039,n1040,n1815);
xor (n1040,n1041,n2241);
xor (n1041,n1042,n1809);
xor (n1042,n1043,n2209);
xor (n1043,n1044,n1803);
xor (n1044,n1045,n2172);
xor (n1045,n1046,n1797);
xor (n1046,n1047,n2130);
xor (n1047,n1048,n1791);
xor (n1048,n1049,n2083);
xor (n1049,n1050,n1785);
xor (n1050,n1051,n2031);
xor (n1051,n1052,n1779);
xor (n1052,n1053,n1974);
xor (n1053,n1054,n1773);
xor (n1054,n1055,n1912);
xor (n1055,n1056,n1767);
xor (n1056,n1057,n1845);
xor (n1057,n1058,n55);
xor (n1058,n1059,n1759);
xor (n1059,n1060,n1758);
xor (n1060,n1061,n1670);
xor (n1061,n1062,n1669);
xor (n1062,n1063,n1571);
xor (n1063,n1064,n1570);
xor (n1064,n1065,n1468);
xor (n1065,n1066,n1467);
xor (n1066,n1067,n1360);
xor (n1067,n1068,n1359);
xor (n1068,n1069,n1080);
xor (n1069,n1070,n1079);
xor (n1070,n1071,n1078);
xor (n1071,n1072,n1077);
xor (n1072,n1073,n1076);
xor (n1073,n1074,n1075);
and (n1074,n23,n196);
and (n1075,n23,n164);
and (n1076,n1074,n1075);
and (n1077,n23,n157);
and (n1078,n1072,n1077);
and (n1079,n23,n73);
or (n1080,n1081,n1082);
and (n1081,n1070,n1079);
and (n1082,n1069,n1083);
or (n1083,n1081,n1084);
and (n1084,n1069,n1085);
or (n1085,n1081,n1086);
and (n1086,n1069,n1087);
or (n1087,n1081,n1088);
and (n1088,n1069,n1089);
or (n1089,n1090,n1274);
and (n1090,n1091,n1273);
xor (n1091,n1071,n1092);
or (n1092,n1093,n1185);
and (n1093,n1094,n1184);
xor (n1094,n1073,n1095);
or (n1095,n1076,n1096);
and (n1096,n1097,n1099);
xor (n1097,n1074,n1098);
and (n1098,n25,n164);
or (n1099,n1100,n1103);
and (n1100,n1101,n1102);
and (n1101,n25,n196);
and (n1102,n53,n164);
and (n1103,n1104,n1105);
xor (n1104,n1101,n1102);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
and (n1107,n53,n196);
and (n1108,n94,n164);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
and (n1113,n94,n196);
and (n1114,n598,n164);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
and (n1119,n598,n196);
and (n1120,n399,n164);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
and (n1125,n399,n196);
and (n1126,n349,n164);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
and (n1131,n349,n196);
and (n1132,n268,n164);
and (n1133,n1134,n1135);
xor (n1134,n1131,n1132);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
and (n1137,n268,n196);
and (n1138,n207,n164);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
and (n1143,n207,n196);
and (n1144,n202,n164);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1150);
and (n1148,n1149,n244);
and (n1149,n202,n196);
and (n1150,n1151,n1152);
xor (n1151,n1149,n244);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
and (n1154,n225,n196);
and (n1155,n171,n164);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
and (n1160,n171,n196);
and (n1161,n149,n164);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1167);
and (n1165,n1166,n483);
and (n1166,n149,n196);
and (n1167,n1168,n1169);
xor (n1168,n1166,n483);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
and (n1171,n184,n196);
and (n1172,n178,n164);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
and (n1177,n178,n196);
and (n1178,n140,n164);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
and (n1181,n1182,n1183);
and (n1182,n140,n196);
and (n1183,n134,n164);
and (n1184,n25,n157);
and (n1185,n1186,n1187);
xor (n1186,n1094,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1097,n1099);
and (n1190,n53,n157);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1104,n1105);
and (n1196,n94,n157);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1203);
and (n1200,n1201,n1202);
xor (n1201,n1110,n1111);
and (n1202,n598,n157);
and (n1203,n1204,n1205);
xor (n1204,n1201,n1202);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1116,n1117);
and (n1208,n399,n157);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1122,n1123);
and (n1214,n349,n157);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1128,n1129);
and (n1220,n268,n157);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
or (n1223,n1224,n1227);
and (n1224,n1225,n1226);
xor (n1225,n1134,n1135);
and (n1226,n207,n157);
and (n1227,n1228,n1229);
xor (n1228,n1225,n1226);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1140,n1141);
and (n1232,n202,n157);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1146,n1147);
and (n1238,n225,n157);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1151,n1152);
and (n1244,n171,n157);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1157,n1158);
and (n1250,n149,n157);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1163,n1164);
and (n1256,n184,n157);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1168,n1169);
and (n1262,n178,n157);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1174,n1175);
and (n1268,n140,n157);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
and (n1271,n1272,n502);
xor (n1272,n1180,n1181);
and (n1273,n25,n73);
and (n1274,n1275,n1276);
xor (n1275,n1091,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
xor (n1278,n1186,n1187);
and (n1279,n53,n73);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1192,n1193);
and (n1285,n94,n73);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1198,n1199);
and (n1291,n598,n73);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1204,n1205);
and (n1297,n399,n73);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1210,n1211);
and (n1303,n349,n73);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1216,n1217);
and (n1309,n268,n73);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1222,n1223);
and (n1315,n207,n73);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1322);
and (n1319,n1320,n1321);
xor (n1320,n1228,n1229);
and (n1321,n202,n73);
and (n1322,n1323,n1324);
xor (n1323,n1320,n1321);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1234,n1235);
and (n1327,n225,n73);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1333);
and (n1331,n1332,n170);
xor (n1332,n1240,n1241);
and (n1333,n1334,n1335);
xor (n1334,n1332,n170);
or (n1335,n1336,n1339);
and (n1336,n1337,n1338);
xor (n1337,n1246,n1247);
and (n1338,n149,n73);
and (n1339,n1340,n1341);
xor (n1340,n1337,n1338);
or (n1341,n1342,n1344);
and (n1342,n1343,n313);
xor (n1343,n1252,n1253);
and (n1344,n1345,n1346);
xor (n1345,n1343,n313);
or (n1346,n1347,n1349);
and (n1347,n1348,n432);
xor (n1348,n1258,n1259);
and (n1349,n1350,n1351);
xor (n1350,n1348,n432);
or (n1351,n1352,n1354);
and (n1352,n1353,n475);
xor (n1353,n1264,n1265);
and (n1354,n1355,n1356);
xor (n1355,n1353,n475);
and (n1356,n1357,n1358);
xor (n1357,n1270,n1271);
and (n1358,n134,n73);
and (n1359,n23,n70);
or (n1360,n1361,n1363);
and (n1361,n1362,n1359);
xor (n1362,n1069,n1083);
and (n1363,n1364,n1365);
xor (n1364,n1362,n1359);
or (n1365,n1366,n1368);
and (n1366,n1367,n1359);
xor (n1367,n1069,n1085);
and (n1368,n1369,n1370);
xor (n1369,n1367,n1359);
or (n1370,n1371,n1373);
and (n1371,n1372,n1359);
xor (n1372,n1069,n1087);
and (n1373,n1374,n1375);
xor (n1374,n1372,n1359);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1069,n1089);
and (n1378,n25,n70);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1275,n1276);
and (n1384,n53,n70);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1281,n1282);
and (n1390,n94,n70);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1287,n1288);
and (n1396,n598,n70);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1293,n1294);
and (n1402,n399,n70);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1299,n1300);
and (n1408,n349,n70);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1305,n1306);
and (n1414,n268,n70);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1311,n1312);
and (n1420,n207,n70);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1317,n1318);
and (n1426,n202,n70);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1323,n1324);
and (n1432,n225,n70);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1329,n1330);
and (n1438,n171,n70);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1334,n1335);
and (n1444,n149,n70);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1340,n1341);
and (n1450,n184,n70);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1345,n1346);
and (n1456,n178,n70);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
or (n1459,n1460,n1463);
and (n1460,n1461,n1462);
xor (n1461,n1350,n1351);
and (n1462,n140,n70);
and (n1463,n1464,n1465);
xor (n1464,n1461,n1462);
and (n1465,n1466,n448);
xor (n1466,n1355,n1356);
and (n1467,n23,n34);
or (n1468,n1469,n1471);
and (n1469,n1470,n1467);
xor (n1470,n1364,n1365);
and (n1471,n1472,n1473);
xor (n1472,n1470,n1467);
or (n1473,n1474,n1476);
and (n1474,n1475,n1467);
xor (n1475,n1369,n1370);
and (n1476,n1477,n1478);
xor (n1477,n1475,n1467);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1374,n1375);
and (n1481,n25,n34);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1380,n1381);
and (n1487,n53,n34);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1386,n1387);
and (n1493,n94,n34);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1392,n1393);
and (n1499,n598,n34);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1398,n1399);
and (n1505,n399,n34);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1404,n1405);
and (n1511,n349,n34);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1410,n1411);
and (n1517,n268,n34);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
or (n1520,n1521,n1524);
and (n1521,n1522,n1523);
xor (n1522,n1416,n1417);
and (n1523,n207,n34);
and (n1524,n1525,n1526);
xor (n1525,n1522,n1523);
or (n1526,n1527,n1530);
and (n1527,n1528,n1529);
xor (n1528,n1422,n1423);
and (n1529,n202,n34);
and (n1530,n1531,n1532);
xor (n1531,n1528,n1529);
or (n1532,n1533,n1536);
and (n1533,n1534,n1535);
xor (n1534,n1428,n1429);
and (n1535,n225,n34);
and (n1536,n1537,n1538);
xor (n1537,n1534,n1535);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1434,n1435);
and (n1541,n171,n34);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
or (n1544,n1545,n1548);
and (n1545,n1546,n1547);
xor (n1546,n1440,n1441);
and (n1547,n149,n34);
and (n1548,n1549,n1550);
xor (n1549,n1546,n1547);
or (n1550,n1551,n1554);
and (n1551,n1552,n1553);
xor (n1552,n1446,n1447);
and (n1553,n184,n34);
and (n1554,n1555,n1556);
xor (n1555,n1552,n1553);
or (n1556,n1557,n1560);
and (n1557,n1558,n1559);
xor (n1558,n1452,n1453);
and (n1559,n178,n34);
and (n1560,n1561,n1562);
xor (n1561,n1558,n1559);
or (n1562,n1563,n1565);
and (n1563,n1564,n438);
xor (n1564,n1458,n1459);
and (n1565,n1566,n1567);
xor (n1566,n1564,n438);
and (n1567,n1568,n1569);
xor (n1568,n1464,n1465);
and (n1569,n134,n34);
and (n1570,n23,n31);
or (n1571,n1572,n1574);
and (n1572,n1573,n1570);
xor (n1573,n1472,n1473);
and (n1574,n1575,n1576);
xor (n1575,n1573,n1570);
or (n1576,n1577,n1580);
and (n1577,n1578,n1579);
xor (n1578,n1477,n1478);
and (n1579,n25,n31);
and (n1580,n1581,n1582);
xor (n1581,n1578,n1579);
or (n1582,n1583,n1586);
and (n1583,n1584,n1585);
xor (n1584,n1483,n1484);
and (n1585,n53,n31);
and (n1586,n1587,n1588);
xor (n1587,n1584,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n1489,n1490);
and (n1591,n94,n31);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1495,n1496);
and (n1597,n598,n31);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1501,n1502);
and (n1603,n399,n31);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1507,n1508);
and (n1609,n349,n31);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1513,n1514);
and (n1615,n268,n31);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1519,n1520);
and (n1621,n207,n31);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1525,n1526);
and (n1627,n202,n31);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1531,n1532);
and (n1633,n225,n31);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1537,n1538);
and (n1639,n171,n31);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1543,n1544);
and (n1645,n149,n31);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1549,n1550);
and (n1651,n184,n31);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1555,n1556);
and (n1657,n178,n31);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1561,n1562);
and (n1663,n140,n31);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
and (n1666,n1667,n1668);
xor (n1667,n1566,n1567);
not (n1668,n238);
and (n1669,n23,n19);
or (n1670,n1671,n1674);
and (n1671,n1672,n1673);
xor (n1672,n1575,n1576);
and (n1673,n25,n19);
and (n1674,n1675,n1676);
xor (n1675,n1672,n1673);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1581,n1582);
and (n1679,n53,n19);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1587,n1588);
and (n1685,n94,n19);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1593,n1594);
and (n1691,n598,n19);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1599,n1600);
and (n1697,n399,n19);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1605,n1606);
and (n1703,n349,n19);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1709);
and (n1707,n1708,n722);
xor (n1708,n1611,n1612);
and (n1709,n1710,n1711);
xor (n1710,n1708,n722);
or (n1711,n1712,n1714);
and (n1712,n1713,n673);
xor (n1713,n1617,n1618);
and (n1714,n1715,n1716);
xor (n1715,n1713,n673);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
xor (n1718,n1623,n1624);
and (n1719,n202,n19);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
xor (n1724,n1629,n1630);
and (n1725,n225,n19);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
or (n1728,n1729,n1731);
and (n1729,n1730,n379);
xor (n1730,n1635,n1636);
and (n1731,n1732,n1733);
xor (n1732,n1730,n379);
or (n1733,n1734,n1736);
and (n1734,n1735,n330);
xor (n1735,n1641,n1642);
and (n1736,n1737,n1738);
xor (n1737,n1735,n330);
or (n1738,n1739,n1741);
and (n1739,n1740,n257);
xor (n1740,n1647,n1648);
and (n1741,n1742,n1743);
xor (n1742,n1740,n257);
or (n1743,n1744,n1747);
and (n1744,n1745,n1746);
xor (n1745,n1653,n1654);
and (n1746,n178,n19);
and (n1747,n1748,n1749);
xor (n1748,n1745,n1746);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
xor (n1751,n1659,n1660);
and (n1752,n140,n19);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
and (n1755,n1756,n1757);
xor (n1756,n1665,n1666);
and (n1757,n134,n19);
and (n1758,n25,n50);
or (n1759,n1760,n1762);
and (n1760,n1761,n55);
xor (n1761,n1675,n1676);
and (n1762,n1763,n1764);
xor (n1763,n1761,n55);
or (n1764,n1765,n1768);
and (n1765,n1766,n1767);
xor (n1766,n1681,n1682);
and (n1767,n94,n50);
and (n1768,n1769,n1770);
xor (n1769,n1766,n1767);
or (n1770,n1771,n1774);
and (n1771,n1772,n1773);
xor (n1772,n1687,n1688);
and (n1773,n598,n50);
and (n1774,n1775,n1776);
xor (n1775,n1772,n1773);
or (n1776,n1777,n1780);
and (n1777,n1778,n1779);
xor (n1778,n1693,n1694);
and (n1779,n399,n50);
and (n1780,n1781,n1782);
xor (n1781,n1778,n1779);
or (n1782,n1783,n1786);
and (n1783,n1784,n1785);
xor (n1784,n1699,n1700);
and (n1785,n349,n50);
and (n1786,n1787,n1788);
xor (n1787,n1784,n1785);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1705,n1706);
and (n1791,n268,n50);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1710,n1711);
and (n1797,n207,n50);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
xor (n1802,n1715,n1716);
and (n1803,n202,n50);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
xor (n1808,n1721,n1722);
and (n1809,n225,n50);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
xor (n1814,n1727,n1728);
and (n1815,n171,n50);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
xor (n1820,n1732,n1733);
and (n1821,n149,n50);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
xor (n1826,n1737,n1738);
and (n1827,n184,n50);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1742,n1743);
and (n1833,n178,n50);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1748,n1749);
and (n1839,n140,n50);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
and (n1842,n1843,n1844);
xor (n1843,n1754,n1755);
and (n1844,n134,n50);
or (n1845,n1846,n1848);
and (n1846,n1847,n1767);
xor (n1847,n1763,n1764);
and (n1848,n1849,n1850);
xor (n1849,n1847,n1767);
or (n1850,n1851,n1853);
and (n1851,n1852,n1773);
xor (n1852,n1769,n1770);
and (n1853,n1854,n1855);
xor (n1854,n1852,n1773);
or (n1855,n1856,n1858);
and (n1856,n1857,n1779);
xor (n1857,n1775,n1776);
and (n1858,n1859,n1860);
xor (n1859,n1857,n1779);
or (n1860,n1861,n1863);
and (n1861,n1862,n1785);
xor (n1862,n1781,n1782);
and (n1863,n1864,n1865);
xor (n1864,n1862,n1785);
or (n1865,n1866,n1868);
and (n1866,n1867,n1791);
xor (n1867,n1787,n1788);
and (n1868,n1869,n1870);
xor (n1869,n1867,n1791);
or (n1870,n1871,n1873);
and (n1871,n1872,n1797);
xor (n1872,n1793,n1794);
and (n1873,n1874,n1875);
xor (n1874,n1872,n1797);
or (n1875,n1876,n1878);
and (n1876,n1877,n1803);
xor (n1877,n1799,n1800);
and (n1878,n1879,n1880);
xor (n1879,n1877,n1803);
or (n1880,n1881,n1883);
and (n1881,n1882,n1809);
xor (n1882,n1805,n1806);
and (n1883,n1884,n1885);
xor (n1884,n1882,n1809);
or (n1885,n1886,n1888);
and (n1886,n1887,n1815);
xor (n1887,n1811,n1812);
and (n1888,n1889,n1890);
xor (n1889,n1887,n1815);
or (n1890,n1891,n1893);
and (n1891,n1892,n1821);
xor (n1892,n1817,n1818);
and (n1893,n1894,n1895);
xor (n1894,n1892,n1821);
or (n1895,n1896,n1898);
and (n1896,n1897,n1827);
xor (n1897,n1823,n1824);
and (n1898,n1899,n1900);
xor (n1899,n1897,n1827);
or (n1900,n1901,n1903);
and (n1901,n1902,n1833);
xor (n1902,n1829,n1830);
and (n1903,n1904,n1905);
xor (n1904,n1902,n1833);
or (n1905,n1906,n1908);
and (n1906,n1907,n1839);
xor (n1907,n1835,n1836);
and (n1908,n1909,n1910);
xor (n1909,n1907,n1839);
and (n1910,n1911,n1844);
xor (n1911,n1841,n1842);
or (n1912,n1913,n1915);
and (n1913,n1914,n1773);
xor (n1914,n1849,n1850);
and (n1915,n1916,n1917);
xor (n1916,n1914,n1773);
or (n1917,n1918,n1920);
and (n1918,n1919,n1779);
xor (n1919,n1854,n1855);
and (n1920,n1921,n1922);
xor (n1921,n1919,n1779);
or (n1922,n1923,n1925);
and (n1923,n1924,n1785);
xor (n1924,n1859,n1860);
and (n1925,n1926,n1927);
xor (n1926,n1924,n1785);
or (n1927,n1928,n1930);
and (n1928,n1929,n1791);
xor (n1929,n1864,n1865);
and (n1930,n1931,n1932);
xor (n1931,n1929,n1791);
or (n1932,n1933,n1935);
and (n1933,n1934,n1797);
xor (n1934,n1869,n1870);
and (n1935,n1936,n1937);
xor (n1936,n1934,n1797);
or (n1937,n1938,n1940);
and (n1938,n1939,n1803);
xor (n1939,n1874,n1875);
and (n1940,n1941,n1942);
xor (n1941,n1939,n1803);
or (n1942,n1943,n1945);
and (n1943,n1944,n1809);
xor (n1944,n1879,n1880);
and (n1945,n1946,n1947);
xor (n1946,n1944,n1809);
or (n1947,n1948,n1950);
and (n1948,n1949,n1815);
xor (n1949,n1884,n1885);
and (n1950,n1951,n1952);
xor (n1951,n1949,n1815);
or (n1952,n1953,n1955);
and (n1953,n1954,n1821);
xor (n1954,n1889,n1890);
and (n1955,n1956,n1957);
xor (n1956,n1954,n1821);
or (n1957,n1958,n1960);
and (n1958,n1959,n1827);
xor (n1959,n1894,n1895);
and (n1960,n1961,n1962);
xor (n1961,n1959,n1827);
or (n1962,n1963,n1965);
and (n1963,n1964,n1833);
xor (n1964,n1899,n1900);
and (n1965,n1966,n1967);
xor (n1966,n1964,n1833);
or (n1967,n1968,n1970);
and (n1968,n1969,n1839);
xor (n1969,n1904,n1905);
and (n1970,n1971,n1972);
xor (n1971,n1969,n1839);
and (n1972,n1973,n1844);
xor (n1973,n1909,n1910);
or (n1974,n1975,n1977);
and (n1975,n1976,n1779);
xor (n1976,n1916,n1917);
and (n1977,n1978,n1979);
xor (n1978,n1976,n1779);
or (n1979,n1980,n1982);
and (n1980,n1981,n1785);
xor (n1981,n1921,n1922);
and (n1982,n1983,n1984);
xor (n1983,n1981,n1785);
or (n1984,n1985,n1987);
and (n1985,n1986,n1791);
xor (n1986,n1926,n1927);
and (n1987,n1988,n1989);
xor (n1988,n1986,n1791);
or (n1989,n1990,n1992);
and (n1990,n1991,n1797);
xor (n1991,n1931,n1932);
and (n1992,n1993,n1994);
xor (n1993,n1991,n1797);
or (n1994,n1995,n1997);
and (n1995,n1996,n1803);
xor (n1996,n1936,n1937);
and (n1997,n1998,n1999);
xor (n1998,n1996,n1803);
or (n1999,n2000,n2002);
and (n2000,n2001,n1809);
xor (n2001,n1941,n1942);
and (n2002,n2003,n2004);
xor (n2003,n2001,n1809);
or (n2004,n2005,n2007);
and (n2005,n2006,n1815);
xor (n2006,n1946,n1947);
and (n2007,n2008,n2009);
xor (n2008,n2006,n1815);
or (n2009,n2010,n2012);
and (n2010,n2011,n1821);
xor (n2011,n1951,n1952);
and (n2012,n2013,n2014);
xor (n2013,n2011,n1821);
or (n2014,n2015,n2017);
and (n2015,n2016,n1827);
xor (n2016,n1956,n1957);
and (n2017,n2018,n2019);
xor (n2018,n2016,n1827);
or (n2019,n2020,n2022);
and (n2020,n2021,n1833);
xor (n2021,n1961,n1962);
and (n2022,n2023,n2024);
xor (n2023,n2021,n1833);
or (n2024,n2025,n2027);
and (n2025,n2026,n1839);
xor (n2026,n1966,n1967);
and (n2027,n2028,n2029);
xor (n2028,n2026,n1839);
and (n2029,n2030,n1844);
xor (n2030,n1971,n1972);
or (n2031,n2032,n2034);
and (n2032,n2033,n1785);
xor (n2033,n1978,n1979);
and (n2034,n2035,n2036);
xor (n2035,n2033,n1785);
or (n2036,n2037,n2039);
and (n2037,n2038,n1791);
xor (n2038,n1983,n1984);
and (n2039,n2040,n2041);
xor (n2040,n2038,n1791);
or (n2041,n2042,n2044);
and (n2042,n2043,n1797);
xor (n2043,n1988,n1989);
and (n2044,n2045,n2046);
xor (n2045,n2043,n1797);
or (n2046,n2047,n2049);
and (n2047,n2048,n1803);
xor (n2048,n1993,n1994);
and (n2049,n2050,n2051);
xor (n2050,n2048,n1803);
or (n2051,n2052,n2054);
and (n2052,n2053,n1809);
xor (n2053,n1998,n1999);
and (n2054,n2055,n2056);
xor (n2055,n2053,n1809);
or (n2056,n2057,n2059);
and (n2057,n2058,n1815);
xor (n2058,n2003,n2004);
and (n2059,n2060,n2061);
xor (n2060,n2058,n1815);
or (n2061,n2062,n2064);
and (n2062,n2063,n1821);
xor (n2063,n2008,n2009);
and (n2064,n2065,n2066);
xor (n2065,n2063,n1821);
or (n2066,n2067,n2069);
and (n2067,n2068,n1827);
xor (n2068,n2013,n2014);
and (n2069,n2070,n2071);
xor (n2070,n2068,n1827);
or (n2071,n2072,n2074);
and (n2072,n2073,n1833);
xor (n2073,n2018,n2019);
and (n2074,n2075,n2076);
xor (n2075,n2073,n1833);
or (n2076,n2077,n2079);
and (n2077,n2078,n1839);
xor (n2078,n2023,n2024);
and (n2079,n2080,n2081);
xor (n2080,n2078,n1839);
and (n2081,n2082,n1844);
xor (n2082,n2028,n2029);
or (n2083,n2084,n2086);
and (n2084,n2085,n1791);
xor (n2085,n2035,n2036);
and (n2086,n2087,n2088);
xor (n2087,n2085,n1791);
or (n2088,n2089,n2091);
and (n2089,n2090,n1797);
xor (n2090,n2040,n2041);
and (n2091,n2092,n2093);
xor (n2092,n2090,n1797);
or (n2093,n2094,n2096);
and (n2094,n2095,n1803);
xor (n2095,n2045,n2046);
and (n2096,n2097,n2098);
xor (n2097,n2095,n1803);
or (n2098,n2099,n2101);
and (n2099,n2100,n1809);
xor (n2100,n2050,n2051);
and (n2101,n2102,n2103);
xor (n2102,n2100,n1809);
or (n2103,n2104,n2106);
and (n2104,n2105,n1815);
xor (n2105,n2055,n2056);
and (n2106,n2107,n2108);
xor (n2107,n2105,n1815);
or (n2108,n2109,n2111);
and (n2109,n2110,n1821);
xor (n2110,n2060,n2061);
and (n2111,n2112,n2113);
xor (n2112,n2110,n1821);
or (n2113,n2114,n2116);
and (n2114,n2115,n1827);
xor (n2115,n2065,n2066);
and (n2116,n2117,n2118);
xor (n2117,n2115,n1827);
or (n2118,n2119,n2121);
and (n2119,n2120,n1833);
xor (n2120,n2070,n2071);
and (n2121,n2122,n2123);
xor (n2122,n2120,n1833);
or (n2123,n2124,n2126);
and (n2124,n2125,n1839);
xor (n2125,n2075,n2076);
and (n2126,n2127,n2128);
xor (n2127,n2125,n1839);
and (n2128,n2129,n1844);
xor (n2129,n2080,n2081);
or (n2130,n2131,n2133);
and (n2131,n2132,n1797);
xor (n2132,n2087,n2088);
and (n2133,n2134,n2135);
xor (n2134,n2132,n1797);
or (n2135,n2136,n2138);
and (n2136,n2137,n1803);
xor (n2137,n2092,n2093);
and (n2138,n2139,n2140);
xor (n2139,n2137,n1803);
or (n2140,n2141,n2143);
and (n2141,n2142,n1809);
xor (n2142,n2097,n2098);
and (n2143,n2144,n2145);
xor (n2144,n2142,n1809);
or (n2145,n2146,n2148);
and (n2146,n2147,n1815);
xor (n2147,n2102,n2103);
and (n2148,n2149,n2150);
xor (n2149,n2147,n1815);
or (n2150,n2151,n2153);
and (n2151,n2152,n1821);
xor (n2152,n2107,n2108);
and (n2153,n2154,n2155);
xor (n2154,n2152,n1821);
or (n2155,n2156,n2158);
and (n2156,n2157,n1827);
xor (n2157,n2112,n2113);
and (n2158,n2159,n2160);
xor (n2159,n2157,n1827);
or (n2160,n2161,n2163);
and (n2161,n2162,n1833);
xor (n2162,n2117,n2118);
and (n2163,n2164,n2165);
xor (n2164,n2162,n1833);
or (n2165,n2166,n2168);
and (n2166,n2167,n1839);
xor (n2167,n2122,n2123);
and (n2168,n2169,n2170);
xor (n2169,n2167,n1839);
and (n2170,n2171,n1844);
xor (n2171,n2127,n2128);
or (n2172,n2173,n2175);
and (n2173,n2174,n1803);
xor (n2174,n2134,n2135);
and (n2175,n2176,n2177);
xor (n2176,n2174,n1803);
or (n2177,n2178,n2180);
and (n2178,n2179,n1809);
xor (n2179,n2139,n2140);
and (n2180,n2181,n2182);
xor (n2181,n2179,n1809);
or (n2182,n2183,n2185);
and (n2183,n2184,n1815);
xor (n2184,n2144,n2145);
and (n2185,n2186,n2187);
xor (n2186,n2184,n1815);
or (n2187,n2188,n2190);
and (n2188,n2189,n1821);
xor (n2189,n2149,n2150);
and (n2190,n2191,n2192);
xor (n2191,n2189,n1821);
or (n2192,n2193,n2195);
and (n2193,n2194,n1827);
xor (n2194,n2154,n2155);
and (n2195,n2196,n2197);
xor (n2196,n2194,n1827);
or (n2197,n2198,n2200);
and (n2198,n2199,n1833);
xor (n2199,n2159,n2160);
and (n2200,n2201,n2202);
xor (n2201,n2199,n1833);
or (n2202,n2203,n2205);
and (n2203,n2204,n1839);
xor (n2204,n2164,n2165);
and (n2205,n2206,n2207);
xor (n2206,n2204,n1839);
and (n2207,n2208,n1844);
xor (n2208,n2169,n2170);
or (n2209,n2210,n2212);
and (n2210,n2211,n1809);
xor (n2211,n2176,n2177);
and (n2212,n2213,n2214);
xor (n2213,n2211,n1809);
or (n2214,n2215,n2217);
and (n2215,n2216,n1815);
xor (n2216,n2181,n2182);
and (n2217,n2218,n2219);
xor (n2218,n2216,n1815);
or (n2219,n2220,n2222);
and (n2220,n2221,n1821);
xor (n2221,n2186,n2187);
and (n2222,n2223,n2224);
xor (n2223,n2221,n1821);
or (n2224,n2225,n2227);
and (n2225,n2226,n1827);
xor (n2226,n2191,n2192);
and (n2227,n2228,n2229);
xor (n2228,n2226,n1827);
or (n2229,n2230,n2232);
and (n2230,n2231,n1833);
xor (n2231,n2196,n2197);
and (n2232,n2233,n2234);
xor (n2233,n2231,n1833);
or (n2234,n2235,n2237);
and (n2235,n2236,n1839);
xor (n2236,n2201,n2202);
and (n2237,n2238,n2239);
xor (n2238,n2236,n1839);
and (n2239,n2240,n1844);
xor (n2240,n2206,n2207);
or (n2241,n2242,n2244);
and (n2242,n2243,n1815);
xor (n2243,n2213,n2214);
and (n2244,n2245,n2246);
xor (n2245,n2243,n1815);
or (n2246,n2247,n2249);
and (n2247,n2248,n1821);
xor (n2248,n2218,n2219);
and (n2249,n2250,n2251);
xor (n2250,n2248,n1821);
or (n2251,n2252,n2254);
and (n2252,n2253,n1827);
xor (n2253,n2223,n2224);
and (n2254,n2255,n2256);
xor (n2255,n2253,n1827);
or (n2256,n2257,n2259);
and (n2257,n2258,n1833);
xor (n2258,n2228,n2229);
and (n2259,n2260,n2261);
xor (n2260,n2258,n1833);
or (n2261,n2262,n2264);
and (n2262,n2263,n1839);
xor (n2263,n2233,n2234);
and (n2264,n2265,n2266);
xor (n2265,n2263,n1839);
and (n2266,n2267,n1844);
xor (n2267,n2238,n2239);
or (n2268,n2269,n2271);
and (n2269,n2270,n1821);
xor (n2270,n2245,n2246);
and (n2271,n2272,n2273);
xor (n2272,n2270,n1821);
or (n2273,n2274,n2276);
and (n2274,n2275,n1827);
xor (n2275,n2250,n2251);
and (n2276,n2277,n2278);
xor (n2277,n2275,n1827);
or (n2278,n2279,n2281);
and (n2279,n2280,n1833);
xor (n2280,n2255,n2256);
and (n2281,n2282,n2283);
xor (n2282,n2280,n1833);
or (n2283,n2284,n2286);
and (n2284,n2285,n1839);
xor (n2285,n2260,n2261);
and (n2286,n2287,n2288);
xor (n2287,n2285,n1839);
and (n2288,n2289,n1844);
xor (n2289,n2265,n2266);
or (n2290,n2291,n2293);
and (n2291,n2292,n1827);
xor (n2292,n2272,n2273);
and (n2293,n2294,n2295);
xor (n2294,n2292,n1827);
or (n2295,n2296,n2298);
and (n2296,n2297,n1833);
xor (n2297,n2277,n2278);
and (n2298,n2299,n2300);
xor (n2299,n2297,n1833);
or (n2300,n2301,n2303);
and (n2301,n2302,n1839);
xor (n2302,n2282,n2283);
and (n2303,n2304,n2305);
xor (n2304,n2302,n1839);
and (n2305,n2306,n1844);
xor (n2306,n2287,n2288);
or (n2307,n2308,n2310);
and (n2308,n2309,n1833);
xor (n2309,n2294,n2295);
and (n2310,n2311,n2312);
xor (n2311,n2309,n1833);
or (n2312,n2313,n2315);
and (n2313,n2314,n1839);
xor (n2314,n2299,n2300);
and (n2315,n2316,n2317);
xor (n2316,n2314,n1839);
and (n2317,n2318,n1844);
xor (n2318,n2304,n2305);
or (n2319,n2320,n2322);
and (n2320,n2321,n1839);
xor (n2321,n2311,n2312);
and (n2322,n2323,n2324);
xor (n2323,n2321,n1839);
and (n2324,n2325,n1844);
xor (n2325,n2316,n2317);
and (n2326,n2327,n1844);
xor (n2327,n2323,n2324);
xor (n2328,n2208,n1844);
endmodule
