module top (out,n8,n9,n11,n12,n19,n21,n27,n36,n46
        ,n47,n49,n56,n85,n87,n100,n109,n119,n127);
output out;
input n8;
input n9;
input n11;
input n12;
input n19;
input n21;
input n27;
input n36;
input n46;
input n47;
input n49;
input n56;
input n85;
input n87;
input n100;
input n109;
input n119;
input n127;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n10;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n20;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
xor (out,n0,n181);
xor (n0,n1,n150);
xor (n1,n2,n79);
xor (n2,n3,n76);
xor (n3,n4,n57);
xor (n4,n5,n38);
xor (n5,n6,n13);
and (n6,n7,n10);
and (n7,n8,n9);
and (n10,n11,n12);
or (n13,n14,n30,n37);
and (n14,n15,n29);
or (n15,n16,n23,n28);
and (n16,n17,n22);
and (n17,n18,n20);
and (n18,n8,n19);
and (n20,n11,n21);
and (n22,n8,n12);
and (n23,n22,n24);
xor (n24,n25,n26);
and (n25,n11,n19);
and (n26,n27,n21);
and (n28,n17,n24);
xor (n29,n7,n10);
and (n30,n29,n31);
xor (n31,n32,n35);
xor (n32,n33,n34);
and (n33,n25,n26);
and (n34,n27,n19);
and (n35,n36,n21);
and (n37,n15,n31);
xor (n38,n39,n51);
xor (n39,n40,n43);
or (n40,n33,n41,n42);
and (n41,n34,n35);
and (n42,n33,n35);
xor (n43,n44,n50);
xor (n44,n45,n48);
and (n45,n46,n47);
and (n48,n8,n49);
and (n50,n11,n9);
xor (n51,n52,n53);
and (n52,n27,n12);
xor (n53,n54,n55);
and (n54,n36,n19);
and (n55,n56,n21);
and (n57,n58,n74);
or (n58,n59,n70,n73);
and (n59,n60,n69);
or (n60,n61,n66,n68);
and (n61,n62,n65);
and (n62,n63,n64);
and (n63,n46,n19);
and (n64,n8,n21);
and (n65,n46,n12);
and (n66,n65,n67);
xor (n67,n18,n20);
and (n68,n62,n67);
and (n69,n46,n9);
and (n70,n69,n71);
xor (n71,n72,n24);
xor (n72,n17,n22);
and (n73,n60,n71);
xor (n74,n75,n31);
xor (n75,n15,n29);
and (n76,n77,n78);
and (n77,n46,n49);
xor (n78,n58,n74);
xor (n79,n80,n147);
xor (n80,n81,n128);
xor (n81,n82,n111);
xor (n82,n83,n88);
and (n83,n84,n86);
and (n84,n85,n9);
and (n86,n87,n12);
or (n88,n89,n103,n110);
and (n89,n90,n102);
or (n90,n91,n96,n101);
and (n91,n92,n95);
and (n92,n93,n94);
and (n93,n85,n19);
and (n94,n87,n21);
and (n95,n85,n12);
and (n96,n95,n97);
xor (n97,n98,n99);
and (n98,n87,n19);
and (n99,n100,n21);
and (n101,n92,n97);
xor (n102,n84,n86);
and (n103,n102,n104);
xor (n104,n105,n108);
xor (n105,n106,n107);
and (n106,n98,n99);
and (n107,n100,n19);
and (n108,n109,n21);
and (n110,n90,n104);
xor (n111,n112,n122);
xor (n112,n113,n116);
or (n113,n106,n114,n115);
and (n114,n107,n108);
and (n115,n106,n108);
xor (n116,n117,n121);
xor (n117,n118,n120);
and (n118,n119,n47);
and (n120,n85,n49);
and (n121,n87,n9);
xor (n122,n123,n124);
and (n123,n100,n12);
xor (n124,n125,n126);
and (n125,n109,n19);
and (n126,n127,n21);
and (n128,n129,n145);
or (n129,n130,n141,n144);
and (n130,n131,n140);
or (n131,n132,n137,n139);
and (n132,n133,n136);
and (n133,n134,n135);
and (n134,n119,n19);
and (n135,n85,n21);
and (n136,n119,n12);
and (n137,n136,n138);
xor (n138,n93,n94);
and (n139,n133,n138);
and (n140,n119,n9);
and (n141,n140,n142);
xor (n142,n143,n97);
xor (n143,n92,n95);
and (n144,n131,n142);
xor (n145,n146,n104);
xor (n146,n90,n102);
and (n147,n148,n149);
and (n148,n119,n49);
xor (n149,n129,n145);
or (n150,n151,n154,n180);
and (n151,n152,n153);
xor (n152,n77,n78);
xor (n153,n148,n149);
and (n154,n153,n155);
or (n155,n156,n161,n179);
and (n156,n157,n159);
xor (n157,n158,n71);
xor (n158,n60,n69);
xor (n159,n160,n142);
xor (n160,n131,n140);
and (n161,n159,n162);
or (n162,n163,n168,n178);
and (n163,n164,n166);
xor (n164,n165,n67);
xor (n165,n62,n65);
xor (n166,n167,n138);
xor (n167,n133,n136);
and (n168,n166,n169);
or (n169,n170,n173,n177);
and (n170,n171,n172);
xor (n171,n63,n64);
xor (n172,n134,n135);
and (n173,n172,n174);
and (n174,n175,n176);
and (n175,n46,n21);
and (n176,n119,n21);
and (n177,n171,n174);
and (n178,n164,n169);
and (n179,n157,n162);
and (n180,n152,n155);
xor (n181,n182,n271);
xor (n182,n183,n252);
xor (n183,n184,n230);
xor (n184,n185,n197);
and (n185,n186,n190);
and (n186,n187,n9);
xor (n187,n188,n189);
xor (n188,n8,n85);
and (n189,n46,n119);
and (n190,n191,n12);
xor (n191,n192,n193);
xor (n192,n11,n87);
or (n193,n194,n195,n196);
and (n194,n8,n85);
and (n195,n85,n189);
and (n196,n8,n189);
or (n197,n198,n217,n229);
and (n198,n199,n216);
or (n199,n200,n205,n215);
and (n200,n201,n204);
and (n201,n202,n203);
and (n202,n187,n19);
and (n203,n191,n21);
and (n204,n187,n12);
and (n205,n204,n206);
xor (n206,n207,n208);
and (n207,n191,n19);
and (n208,n209,n21);
xor (n209,n210,n211);
xor (n210,n27,n100);
or (n211,n212,n213,n214);
and (n212,n11,n87);
and (n213,n87,n193);
and (n214,n11,n193);
and (n215,n201,n206);
xor (n216,n186,n190);
and (n217,n216,n218);
xor (n218,n219,n222);
xor (n219,n220,n221);
and (n220,n207,n208);
and (n221,n209,n19);
and (n222,n223,n21);
xor (n223,n224,n225);
xor (n224,n36,n109);
or (n225,n226,n227,n228);
and (n226,n27,n100);
and (n227,n100,n211);
and (n228,n27,n211);
and (n229,n199,n218);
xor (n230,n231,n241);
xor (n231,n232,n235);
or (n232,n220,n233,n234);
and (n233,n221,n222);
and (n234,n220,n222);
xor (n235,n236,n240);
xor (n236,n237,n239);
and (n237,n238,n47);
xor (n238,n46,n119);
and (n239,n187,n49);
and (n240,n191,n9);
xor (n241,n242,n243);
and (n242,n209,n12);
xor (n243,n244,n245);
and (n244,n223,n19);
and (n245,n246,n21);
xor (n246,n247,n248);
xor (n247,n56,n127);
or (n248,n249,n250,n251);
and (n249,n36,n109);
and (n250,n109,n225);
and (n251,n36,n225);
and (n252,n253,n269);
or (n253,n254,n265,n268);
and (n254,n255,n264);
or (n255,n256,n261,n263);
and (n256,n257,n260);
and (n257,n258,n259);
and (n258,n238,n19);
and (n259,n187,n21);
and (n260,n238,n12);
and (n261,n260,n262);
xor (n262,n202,n203);
and (n263,n257,n262);
and (n264,n238,n9);
and (n265,n264,n266);
xor (n266,n267,n206);
xor (n267,n201,n204);
and (n268,n255,n266);
xor (n269,n270,n218);
xor (n270,n199,n216);
and (n271,n272,n273);
and (n272,n238,n49);
xor (n273,n253,n269);
endmodule
