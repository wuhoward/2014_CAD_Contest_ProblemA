module top (out,n18,n20,n26,n30,n36,n45,n47,n52,n57
        ,n65,n74,n79,n83,n89,n102,n110,n117,n127,n128
        ,n137,n143,n152,n153,n159,n170,n179,n185,n188,n194
        ,n202);
output out;
input n18;
input n20;
input n26;
input n30;
input n36;
input n45;
input n47;
input n52;
input n57;
input n65;
input n74;
input n79;
input n83;
input n89;
input n102;
input n110;
input n117;
input n127;
input n128;
input n137;
input n143;
input n152;
input n153;
input n159;
input n170;
input n179;
input n185;
input n188;
input n194;
input n202;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
xor (out,n0,n803);
nand (n0,n1,n802);
or (n1,n2,n389);
not (n2,n3);
nor (n3,n4,n385);
not (n4,n5);
nand (n5,n6,n353);
xor (n6,n7,n301);
xor (n7,n8,n205);
xor (n8,n9,n173);
xor (n9,n10,n93);
or (n10,n11,n92);
and (n11,n12,n68);
xor (n12,n13,n39);
nand (n13,n14,n33);
or (n14,n15,n28);
nand (n15,n16,n23);
nor (n16,n17,n21);
and (n17,n18,n19);
not (n19,n20);
and (n21,n22,n20);
not (n22,n18);
nand (n23,n24,n27);
or (n24,n20,n25);
not (n25,n26);
nand (n27,n25,n20);
nor (n28,n29,n31);
and (n29,n25,n30);
and (n31,n26,n32);
not (n32,n30);
or (n33,n16,n34);
nor (n34,n35,n37);
and (n35,n25,n36);
and (n37,n26,n38);
not (n38,n36);
nand (n39,n40,n60);
or (n40,n41,n55);
not (n41,n42);
nor (n42,n43,n49);
nand (n43,n44,n48);
or (n44,n45,n46);
not (n46,n47);
nand (n48,n45,n46);
nor (n49,n50,n53);
and (n50,n51,n45);
not (n51,n52);
and (n53,n52,n54);
not (n54,n45);
nor (n55,n56,n58);
and (n56,n51,n57);
and (n58,n52,n59);
not (n59,n57);
or (n60,n61,n62);
not (n61,n43);
not (n62,n63);
nor (n63,n64,n66);
and (n64,n65,n52);
and (n66,n67,n51);
not (n67,n65);
nand (n68,n69,n86);
or (n69,n70,n81);
nand (n70,n71,n76);
and (n71,n72,n75);
nand (n72,n52,n73);
not (n73,n74);
nand (n75,n74,n51);
nand (n76,n77,n80);
or (n77,n74,n78);
not (n78,n79);
nand (n80,n78,n74);
nor (n81,n82,n84);
and (n82,n78,n83);
and (n84,n79,n85);
not (n85,n83);
or (n86,n71,n87);
nor (n87,n88,n90);
and (n88,n78,n89);
and (n90,n79,n91);
not (n91,n89);
and (n92,n13,n39);
or (n93,n94,n172);
and (n94,n95,n146);
xor (n95,n96,n120);
nand (n96,n97,n113);
or (n97,n98,n108);
not (n98,n99);
nor (n99,n100,n105);
nand (n100,n101,n103);
or (n101,n102,n25);
or (n103,n26,n104);
not (n104,n102);
nor (n105,n106,n107);
and (n106,n46,n102);
and (n107,n47,n104);
nor (n108,n109,n111);
and (n109,n46,n110);
and (n111,n47,n112);
not (n112,n110);
or (n113,n114,n115);
not (n114,n100);
nor (n115,n116,n118);
and (n116,n46,n117);
and (n118,n47,n119);
not (n119,n117);
nand (n120,n121,n140);
or (n121,n122,n135);
not (n122,n123);
nor (n123,n124,n131);
nor (n124,n125,n129);
and (n125,n126,n128);
not (n126,n127);
and (n129,n127,n130);
not (n130,n128);
not (n131,n132);
nor (n132,n133,n134);
and (n133,n78,n128);
and (n134,n79,n130);
nor (n135,n136,n138);
and (n136,n126,n137);
and (n138,n127,n139);
not (n139,n137);
or (n140,n132,n141);
nor (n141,n142,n144);
and (n142,n126,n143);
and (n144,n127,n145);
not (n145,n143);
nand (n146,n147,n161);
or (n147,n148,n156);
not (n148,n149);
nand (n149,n150,n154);
or (n150,n151,n153);
not (n151,n152);
or (n154,n155,n152);
not (n155,n153);
not (n156,n157);
nand (n157,n158,n160);
or (n158,n159,n126);
nand (n160,n126,n159);
or (n161,n162,n167);
nand (n162,n156,n163);
nand (n163,n164,n166);
or (n164,n153,n165);
not (n165,n159);
nand (n166,n153,n165);
nor (n167,n168,n171);
and (n168,n169,n153);
not (n169,n170);
and (n171,n170,n155);
and (n172,n96,n120);
xor (n173,n174,n197);
xor (n174,n175,n181);
nor (n175,n176,n169);
not (n176,n177);
nand (n177,n178,n180);
or (n178,n155,n179);
nand (n180,n179,n155);
nand (n181,n182,n191);
or (n182,n183,n186);
nand (n183,n184,n18);
not (n184,n185);
nor (n186,n187,n189);
and (n187,n22,n188);
and (n189,n18,n190);
not (n190,n188);
or (n191,n192,n184);
nor (n192,n193,n195);
and (n193,n22,n194);
and (n195,n18,n196);
not (n196,n194);
nand (n197,n198,n199);
or (n198,n15,n34);
or (n199,n16,n200);
nor (n200,n201,n203);
and (n201,n25,n202);
and (n203,n26,n204);
not (n204,n202);
xor (n205,n206,n255);
xor (n206,n207,n228);
xor (n207,n208,n222);
xor (n208,n209,n216);
nand (n209,n210,n211);
or (n210,n62,n41);
nand (n211,n212,n43);
not (n212,n213);
nor (n213,n214,n215);
and (n214,n51,n110);
and (n215,n52,n112);
nand (n216,n217,n218);
or (n217,n70,n87);
or (n218,n71,n219);
nor (n219,n220,n221);
and (n220,n59,n79);
and (n221,n57,n78);
nand (n222,n223,n224);
or (n223,n98,n115);
or (n224,n114,n225);
nor (n225,n226,n227);
and (n226,n46,n30);
and (n227,n47,n32);
xor (n228,n229,n242);
xor (n229,n230,n236);
nand (n230,n231,n232);
or (n231,n122,n141);
or (n232,n132,n233);
nor (n233,n234,n235);
and (n234,n126,n83);
and (n235,n127,n85);
nand (n236,n237,n238);
or (n237,n148,n162);
or (n238,n156,n239);
nor (n239,n240,n241);
and (n240,n155,n137);
and (n241,n153,n139);
and (n242,n243,n249);
nor (n243,n244,n155);
nor (n244,n245,n248);
and (n245,n246,n126);
not (n246,n247);
and (n247,n170,n159);
and (n248,n169,n165);
nand (n249,n250,n254);
or (n250,n251,n183);
nor (n251,n252,n253);
and (n252,n22,n202);
and (n253,n18,n204);
or (n254,n186,n184);
or (n255,n256,n300);
and (n256,n257,n277);
xor (n257,n258,n259);
xor (n258,n243,n249);
or (n259,n260,n276);
and (n260,n261,n270);
xor (n261,n262,n263);
nor (n262,n156,n169);
nand (n263,n264,n269);
or (n264,n265,n15);
not (n265,n266);
nand (n266,n267,n268);
or (n267,n26,n119);
or (n268,n25,n117);
or (n269,n16,n28);
nand (n270,n271,n275);
or (n271,n41,n272);
nor (n272,n273,n274);
and (n273,n51,n89);
and (n274,n52,n91);
or (n275,n61,n55);
and (n276,n262,n263);
or (n277,n278,n299);
and (n278,n279,n293);
xor (n279,n280,n286);
nand (n280,n281,n285);
or (n281,n70,n282);
nor (n282,n283,n284);
and (n283,n78,n143);
and (n284,n79,n145);
or (n285,n71,n81);
nand (n286,n287,n292);
or (n287,n183,n288);
not (n288,n289);
nor (n289,n290,n291);
and (n290,n36,n18);
and (n291,n38,n22);
or (n292,n251,n184);
nand (n293,n294,n298);
or (n294,n122,n295);
nor (n295,n296,n297);
and (n296,n126,n152);
and (n297,n127,n151);
or (n298,n132,n135);
and (n299,n280,n286);
and (n300,n258,n259);
or (n301,n302,n352);
and (n302,n303,n306);
xor (n303,n304,n305);
xor (n304,n95,n146);
xor (n305,n12,n68);
or (n306,n307,n351);
and (n307,n308,n329);
xor (n308,n309,n315);
nand (n309,n310,n314);
or (n310,n98,n311);
nor (n311,n312,n313);
and (n312,n46,n65);
and (n313,n47,n67);
or (n314,n114,n108);
and (n315,n316,n322);
nand (n316,n317,n321);
or (n317,n15,n318);
nor (n318,n319,n320);
and (n319,n25,n110);
and (n320,n26,n112);
or (n321,n16,n265);
not (n322,n323);
nand (n323,n324,n127);
nand (n324,n325,n326);
or (n325,n170,n128);
nand (n326,n327,n78);
not (n327,n328);
and (n328,n170,n128);
or (n329,n330,n350);
and (n330,n331,n344);
xor (n331,n332,n338);
nand (n332,n333,n337);
or (n333,n41,n334);
nor (n334,n335,n336);
and (n335,n51,n83);
and (n336,n52,n85);
or (n337,n61,n272);
nand (n338,n339,n343);
or (n339,n70,n340);
nor (n340,n341,n342);
and (n341,n78,n137);
and (n342,n79,n139);
or (n343,n71,n282);
nand (n344,n345,n346);
or (n345,n184,n288);
or (n346,n347,n183);
nor (n347,n348,n349);
and (n348,n22,n30);
and (n349,n18,n32);
and (n350,n332,n338);
and (n351,n309,n315);
and (n352,n304,n305);
or (n353,n354,n384);
and (n354,n355,n383);
xor (n355,n356,n357);
xor (n356,n257,n277);
or (n357,n358,n382);
and (n358,n359,n362);
xor (n359,n360,n361);
xor (n360,n279,n293);
xor (n361,n261,n270);
or (n362,n363,n381);
and (n363,n364,n377);
xor (n364,n365,n371);
nand (n365,n366,n370);
or (n366,n122,n367);
nor (n367,n368,n369);
and (n368,n169,n127);
and (n369,n126,n170);
or (n370,n132,n295);
nand (n371,n372,n376);
or (n372,n98,n373);
nor (n373,n374,n375);
and (n374,n46,n57);
and (n375,n47,n59);
or (n376,n114,n311);
nand (n377,n378,n380);
or (n378,n322,n379);
not (n379,n316);
or (n380,n316,n323);
and (n381,n365,n371);
and (n382,n360,n361);
xor (n383,n303,n306);
and (n384,n356,n357);
not (n385,n386);
nand (n386,n387,n388);
not (n387,n6);
not (n388,n353);
not (n389,n390);
nor (n390,n391,n798);
and (n391,n392,n779);
or (n392,n393,n778);
and (n393,n394,n519);
xor (n394,n395,n504);
or (n395,n396,n503);
and (n396,n397,n470);
xor (n397,n398,n418);
xor (n398,n399,n412);
xor (n399,n400,n406);
nand (n400,n401,n405);
or (n401,n70,n402);
nor (n402,n403,n404);
and (n403,n78,n152);
and (n404,n79,n151);
or (n405,n71,n340);
nand (n406,n407,n411);
or (n407,n408,n183);
nor (n408,n409,n410);
and (n409,n22,n117);
and (n410,n18,n119);
or (n411,n347,n184);
nand (n412,n413,n417);
or (n413,n98,n414);
nor (n414,n415,n416);
and (n415,n46,n89);
and (n416,n47,n91);
or (n417,n114,n373);
or (n418,n419,n469);
and (n419,n420,n443);
xor (n420,n421,n427);
nand (n421,n422,n426);
or (n422,n98,n423);
nor (n423,n424,n425);
and (n424,n46,n83);
and (n425,n47,n85);
or (n426,n114,n414);
xor (n427,n428,n434);
and (n428,n429,n79);
nand (n429,n430,n431);
or (n430,n170,n74);
nand (n431,n432,n51);
not (n432,n433);
and (n433,n170,n74);
nand (n434,n435,n439);
or (n435,n15,n436);
nor (n436,n437,n438);
and (n437,n25,n57);
and (n438,n26,n59);
or (n439,n16,n440);
nor (n440,n441,n442);
and (n441,n25,n65);
and (n442,n26,n67);
or (n443,n444,n468);
and (n444,n445,n457);
xor (n445,n446,n448);
and (n446,n447,n170);
not (n447,n71);
nand (n448,n449,n453);
or (n449,n183,n450);
nor (n450,n451,n452);
and (n451,n22,n65);
and (n452,n18,n67);
or (n453,n454,n184);
nor (n454,n455,n456);
and (n455,n22,n110);
and (n456,n18,n112);
nand (n457,n458,n463);
or (n458,n459,n41);
not (n459,n460);
nor (n460,n461,n462);
and (n461,n152,n52);
and (n462,n151,n51);
nand (n463,n464,n43);
not (n464,n465);
nor (n465,n466,n467);
and (n466,n51,n137);
and (n467,n52,n139);
and (n468,n446,n448);
and (n469,n421,n427);
xor (n470,n471,n494);
xor (n471,n472,n473);
and (n472,n428,n434);
or (n473,n474,n493);
and (n474,n475,n490);
xor (n475,n476,n482);
nand (n476,n477,n478);
or (n477,n41,n465);
or (n478,n61,n479);
nor (n479,n480,n481);
and (n480,n51,n143);
and (n481,n52,n145);
nand (n482,n483,n488);
or (n483,n484,n70);
not (n484,n485);
nand (n485,n486,n487);
or (n486,n78,n170);
or (n487,n169,n79);
nand (n488,n489,n447);
not (n489,n402);
nand (n490,n491,n492);
or (n491,n183,n454);
or (n492,n408,n184);
and (n493,n476,n482);
xor (n494,n495,n500);
xor (n495,n496,n497);
nor (n496,n132,n169);
nand (n497,n498,n499);
or (n498,n15,n440);
or (n499,n16,n318);
nand (n500,n501,n502);
or (n501,n41,n479);
or (n502,n61,n334);
and (n503,n398,n418);
xor (n504,n505,n516);
xor (n505,n506,n507);
xor (n506,n364,n377);
xor (n507,n508,n515);
xor (n508,n509,n512);
or (n509,n510,n511);
and (n510,n495,n500);
and (n511,n496,n497);
or (n512,n513,n514);
and (n513,n399,n412);
and (n514,n400,n406);
xor (n515,n331,n344);
or (n516,n517,n518);
and (n517,n471,n494);
and (n518,n472,n473);
or (n519,n520,n777);
and (n520,n521,n561);
xor (n521,n522,n560);
or (n522,n523,n559);
and (n523,n524,n558);
xor (n524,n525,n526);
xor (n525,n475,n490);
or (n526,n527,n557);
and (n527,n528,n543);
xor (n528,n529,n535);
nand (n529,n530,n534);
or (n530,n15,n531);
nor (n531,n532,n533);
and (n532,n91,n26);
and (n533,n89,n25);
or (n534,n16,n436);
nand (n535,n536,n541);
or (n536,n537,n98);
not (n537,n538);
nand (n538,n539,n540);
or (n539,n47,n145);
or (n540,n46,n143);
nand (n541,n542,n100);
not (n542,n423);
and (n543,n544,n550);
nor (n544,n545,n51);
nor (n545,n546,n549);
and (n546,n547,n46);
not (n547,n548);
and (n548,n170,n45);
and (n549,n169,n54);
nand (n550,n551,n556);
or (n551,n183,n552);
not (n552,n553);
nor (n553,n554,n555);
and (n554,n59,n22);
and (n555,n57,n18);
or (n556,n450,n184);
and (n557,n529,n535);
xor (n558,n420,n443);
and (n559,n525,n526);
xor (n560,n397,n470);
or (n561,n562,n776);
and (n562,n563,n598);
xor (n563,n564,n597);
or (n564,n565,n596);
and (n565,n566,n595);
xor (n566,n567,n594);
or (n567,n568,n593);
and (n568,n569,n586);
xor (n569,n570,n577);
nand (n570,n571,n576);
or (n571,n572,n41);
not (n572,n573);
nand (n573,n574,n575);
or (n574,n51,n170);
or (n575,n169,n52);
nand (n576,n43,n460);
nand (n577,n578,n583);
or (n578,n579,n15);
not (n579,n580);
nor (n580,n581,n582);
and (n581,n85,n25);
and (n582,n83,n26);
nand (n583,n584,n585);
not (n584,n531);
not (n585,n16);
nand (n586,n587,n592);
or (n587,n588,n98);
not (n588,n589);
nor (n589,n590,n591);
and (n590,n137,n47);
and (n591,n139,n46);
nand (n592,n100,n538);
and (n593,n570,n577);
xor (n594,n445,n457);
xor (n595,n528,n543);
and (n596,n567,n594);
xor (n597,n524,n558);
nand (n598,n599,n775);
or (n599,n600,n630);
not (n600,n601);
nand (n601,n602,n604);
not (n602,n603);
xor (n603,n566,n595);
not (n604,n605);
or (n605,n606,n629);
and (n606,n607,n628);
xor (n607,n608,n609);
xor (n608,n544,n550);
or (n609,n610,n627);
and (n610,n611,n620);
xor (n611,n612,n613);
and (n612,n43,n170);
nand (n613,n614,n619);
or (n614,n183,n615);
not (n615,n616);
nor (n616,n617,n618);
and (n617,n89,n18);
and (n618,n91,n22);
nand (n619,n553,n185);
nand (n620,n621,n626);
or (n621,n622,n15);
not (n622,n623);
nor (n623,n624,n625);
and (n624,n145,n25);
and (n625,n143,n26);
nand (n626,n585,n580);
and (n627,n612,n613);
xor (n628,n569,n586);
and (n629,n608,n609);
not (n630,n631);
nand (n631,n632,n774);
or (n632,n633,n664);
not (n633,n634);
nand (n634,n635,n637);
not (n635,n636);
xor (n636,n607,n628);
not (n637,n638);
or (n638,n639,n663);
and (n639,n640,n662);
xor (n640,n641,n648);
nand (n641,n642,n647);
or (n642,n643,n98);
not (n643,n644);
nor (n644,n645,n646);
and (n645,n152,n47);
and (n646,n151,n46);
nand (n647,n100,n589);
and (n648,n649,n654);
and (n649,n650,n47);
nand (n650,n651,n653);
or (n651,n652,n26);
and (n652,n170,n102);
or (n653,n170,n102);
nand (n654,n655,n656);
or (n655,n184,n615);
nand (n656,n657,n661);
not (n657,n658);
nor (n658,n659,n660);
and (n659,n83,n22);
and (n660,n85,n18);
not (n661,n183);
xor (n662,n611,n620);
and (n663,n641,n648);
not (n664,n665);
nand (n665,n666,n773);
or (n666,n667,n691);
not (n667,n668);
nand (n668,n669,n671);
not (n669,n670);
xor (n670,n640,n662);
not (n671,n672);
or (n672,n673,n690);
and (n673,n674,n689);
xor (n674,n675,n682);
nand (n675,n676,n681);
or (n676,n677,n15);
not (n677,n678);
nor (n678,n679,n680);
and (n679,n139,n25);
and (n680,n137,n26);
nand (n681,n585,n623);
nand (n682,n683,n688);
or (n683,n684,n98);
not (n684,n685);
nand (n685,n686,n687);
or (n686,n46,n170);
or (n687,n47,n169);
nand (n688,n100,n644);
xor (n689,n649,n654);
and (n690,n675,n682);
not (n691,n692);
nand (n692,n693,n772);
or (n693,n694,n718);
not (n694,n695);
nand (n695,n696,n698);
not (n696,n697);
xor (n697,n674,n689);
not (n698,n699);
or (n699,n700,n717);
and (n700,n701,n710);
xor (n701,n702,n703);
and (n702,n100,n170);
nand (n703,n704,n709);
or (n704,n705,n15);
not (n705,n706);
nor (n706,n707,n708);
and (n707,n152,n26);
and (n708,n151,n25);
nand (n709,n585,n678);
nand (n710,n711,n716);
or (n711,n183,n712);
not (n712,n713);
nor (n713,n714,n715);
and (n714,n145,n22);
and (n715,n143,n18);
or (n716,n658,n184);
and (n717,n702,n703);
not (n718,n719);
nand (n719,n720,n771);
or (n720,n721,n737);
nor (n721,n722,n723);
xor (n722,n701,n710);
and (n723,n724,n730);
nor (n724,n725,n25);
nor (n725,n726,n727);
and (n726,n19,n169);
and (n727,n728,n22);
not (n728,n729);
and (n729,n170,n20);
nand (n730,n731,n732);
or (n731,n184,n712);
nand (n732,n733,n661);
not (n733,n734);
nor (n734,n735,n736);
and (n735,n22,n137);
and (n736,n18,n139);
not (n737,n738);
or (n738,n739,n770);
and (n739,n740,n749);
xor (n740,n741,n748);
nand (n741,n742,n747);
or (n742,n743,n15);
not (n743,n744);
nand (n744,n745,n746);
or (n745,n25,n170);
or (n746,n26,n169);
nand (n747,n585,n706);
xor (n748,n724,n730);
or (n749,n750,n769);
and (n750,n751,n759);
xor (n751,n752,n753);
nor (n752,n16,n169);
nand (n753,n754,n758);
or (n754,n755,n183);
nor (n755,n756,n757);
and (n756,n22,n152);
and (n757,n18,n151);
or (n758,n734,n184);
nor (n759,n760,n767);
nor (n760,n761,n763);
and (n761,n762,n185);
not (n762,n755);
nor (n763,n764,n183);
nor (n764,n765,n766);
and (n765,n170,n22);
and (n766,n169,n18);
or (n767,n768,n22);
and (n768,n170,n185);
and (n769,n752,n753);
and (n770,n741,n748);
nand (n771,n722,n723);
nand (n772,n697,n699);
nand (n773,n670,n672);
nand (n774,n636,n638);
nand (n775,n603,n605);
and (n776,n564,n597);
and (n777,n522,n560);
and (n778,n395,n504);
not (n779,n780);
nand (n780,n781,n793);
not (n781,n782);
nor (n782,n783,n784);
xor (n783,n355,n383);
or (n784,n785,n792);
and (n785,n786,n791);
xor (n786,n787,n788);
xor (n787,n308,n329);
or (n788,n789,n790);
and (n789,n508,n515);
and (n790,n509,n512);
xor (n791,n359,n362);
and (n792,n787,n788);
or (n793,n794,n797);
or (n794,n795,n796);
and (n795,n505,n516);
and (n796,n506,n507);
xor (n797,n786,n791);
nand (n798,n799,n801);
or (n799,n782,n800);
nand (n800,n794,n797);
nand (n801,n783,n784);
or (n802,n390,n3);
xor (n803,n804,n1333);
xor (n804,n805,n1330);
xor (n805,n806,n1329);
xor (n806,n807,n1321);
xor (n807,n808,n1320);
xor (n808,n809,n1305);
xor (n809,n810,n1304);
xor (n810,n811,n1284);
xor (n811,n812,n1283);
xor (n812,n813,n1256);
xor (n813,n814,n1255);
xor (n814,n815,n1223);
xor (n815,n816,n1222);
xor (n816,n817,n1184);
xor (n817,n818,n64);
xor (n818,n819,n1140);
xor (n819,n820,n1139);
xor (n820,n821,n1090);
xor (n821,n822,n1089);
xor (n822,n823,n1033);
xor (n823,n824,n1032);
xor (n824,n825,n973);
xor (n825,n826,n972);
xor (n826,n827,n904);
xor (n827,n828,n903);
xor (n828,n829,n832);
xor (n829,n830,n831);
and (n830,n194,n185);
and (n831,n188,n18);
or (n832,n833,n836);
and (n833,n834,n835);
and (n834,n188,n185);
and (n835,n202,n18);
and (n836,n837,n838);
xor (n837,n834,n835);
or (n838,n839,n841);
and (n839,n840,n290);
and (n840,n202,n185);
and (n841,n842,n843);
xor (n842,n840,n290);
or (n843,n844,n847);
and (n844,n845,n846);
and (n845,n36,n185);
and (n846,n30,n18);
and (n847,n848,n849);
xor (n848,n845,n846);
or (n849,n850,n853);
and (n850,n851,n852);
and (n851,n30,n185);
and (n852,n117,n18);
and (n853,n854,n855);
xor (n854,n851,n852);
or (n855,n856,n859);
and (n856,n857,n858);
and (n857,n117,n185);
and (n858,n110,n18);
and (n859,n860,n861);
xor (n860,n857,n858);
or (n861,n862,n865);
and (n862,n863,n864);
and (n863,n110,n185);
and (n864,n65,n18);
and (n865,n866,n867);
xor (n866,n863,n864);
or (n867,n868,n870);
and (n868,n869,n555);
and (n869,n65,n185);
and (n870,n871,n872);
xor (n871,n869,n555);
or (n872,n873,n875);
and (n873,n874,n617);
and (n874,n57,n185);
and (n875,n876,n877);
xor (n876,n874,n617);
or (n877,n878,n881);
and (n878,n879,n880);
and (n879,n89,n185);
and (n880,n83,n18);
and (n881,n882,n883);
xor (n882,n879,n880);
or (n883,n884,n886);
and (n884,n885,n715);
and (n885,n83,n185);
and (n886,n887,n888);
xor (n887,n885,n715);
or (n888,n889,n892);
and (n889,n890,n891);
and (n890,n143,n185);
and (n891,n137,n18);
and (n892,n893,n894);
xor (n893,n890,n891);
or (n894,n895,n898);
and (n895,n896,n897);
and (n896,n137,n185);
and (n897,n152,n18);
and (n898,n899,n900);
xor (n899,n896,n897);
and (n900,n901,n902);
and (n901,n152,n185);
and (n902,n170,n18);
and (n903,n202,n20);
or (n904,n905,n908);
and (n905,n906,n907);
xor (n906,n837,n838);
and (n907,n36,n20);
and (n908,n909,n910);
xor (n909,n906,n907);
or (n910,n911,n914);
and (n911,n912,n913);
xor (n912,n842,n843);
and (n913,n30,n20);
and (n914,n915,n916);
xor (n915,n912,n913);
or (n916,n917,n920);
and (n917,n918,n919);
xor (n918,n848,n849);
and (n919,n117,n20);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
xor (n924,n854,n855);
and (n925,n110,n20);
and (n926,n927,n928);
xor (n927,n924,n925);
or (n928,n929,n932);
and (n929,n930,n931);
xor (n930,n860,n861);
and (n931,n65,n20);
and (n932,n933,n934);
xor (n933,n930,n931);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n866,n867);
and (n937,n57,n20);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n871,n872);
and (n943,n89,n20);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
xor (n948,n876,n877);
and (n949,n83,n20);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n956);
and (n953,n954,n955);
xor (n954,n882,n883);
and (n955,n143,n20);
and (n956,n957,n958);
xor (n957,n954,n955);
or (n958,n959,n962);
and (n959,n960,n961);
xor (n960,n887,n888);
and (n961,n137,n20);
and (n962,n963,n964);
xor (n963,n960,n961);
or (n964,n965,n968);
and (n965,n966,n967);
xor (n966,n893,n894);
and (n967,n152,n20);
and (n968,n969,n970);
xor (n969,n966,n967);
and (n970,n971,n729);
xor (n971,n899,n900);
and (n972,n36,n26);
or (n973,n974,n977);
and (n974,n975,n976);
xor (n975,n909,n910);
and (n976,n30,n26);
and (n977,n978,n979);
xor (n978,n975,n976);
or (n979,n980,n983);
and (n980,n981,n982);
xor (n981,n915,n916);
and (n982,n117,n26);
and (n983,n984,n985);
xor (n984,n981,n982);
or (n985,n986,n989);
and (n986,n987,n988);
xor (n987,n921,n922);
and (n988,n110,n26);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
xor (n993,n927,n928);
and (n994,n65,n26);
and (n995,n996,n997);
xor (n996,n993,n994);
or (n997,n998,n1001);
and (n998,n999,n1000);
xor (n999,n933,n934);
and (n1000,n57,n26);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n939,n940);
and (n1006,n89,n26);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1012);
and (n1010,n1011,n582);
xor (n1011,n945,n946);
and (n1012,n1013,n1014);
xor (n1013,n1011,n582);
or (n1014,n1015,n1017);
and (n1015,n1016,n625);
xor (n1016,n951,n952);
and (n1017,n1018,n1019);
xor (n1018,n1016,n625);
or (n1019,n1020,n1022);
and (n1020,n1021,n680);
xor (n1021,n957,n958);
and (n1022,n1023,n1024);
xor (n1023,n1021,n680);
or (n1024,n1025,n1027);
and (n1025,n1026,n707);
xor (n1026,n963,n964);
and (n1027,n1028,n1029);
xor (n1028,n1026,n707);
and (n1029,n1030,n1031);
xor (n1030,n969,n970);
and (n1031,n170,n26);
and (n1032,n30,n102);
or (n1033,n1034,n1037);
and (n1034,n1035,n1036);
xor (n1035,n978,n979);
and (n1036,n117,n102);
and (n1037,n1038,n1039);
xor (n1038,n1035,n1036);
or (n1039,n1040,n1043);
and (n1040,n1041,n1042);
xor (n1041,n984,n985);
and (n1042,n110,n102);
and (n1043,n1044,n1045);
xor (n1044,n1041,n1042);
or (n1045,n1046,n1049);
and (n1046,n1047,n1048);
xor (n1047,n990,n991);
and (n1048,n65,n102);
and (n1049,n1050,n1051);
xor (n1050,n1047,n1048);
or (n1051,n1052,n1055);
and (n1052,n1053,n1054);
xor (n1053,n996,n997);
and (n1054,n57,n102);
and (n1055,n1056,n1057);
xor (n1056,n1053,n1054);
or (n1057,n1058,n1061);
and (n1058,n1059,n1060);
xor (n1059,n1002,n1003);
and (n1060,n89,n102);
and (n1061,n1062,n1063);
xor (n1062,n1059,n1060);
or (n1063,n1064,n1067);
and (n1064,n1065,n1066);
xor (n1065,n1008,n1009);
and (n1066,n83,n102);
and (n1067,n1068,n1069);
xor (n1068,n1065,n1066);
or (n1069,n1070,n1073);
and (n1070,n1071,n1072);
xor (n1071,n1013,n1014);
and (n1072,n143,n102);
and (n1073,n1074,n1075);
xor (n1074,n1071,n1072);
or (n1075,n1076,n1079);
and (n1076,n1077,n1078);
xor (n1077,n1018,n1019);
and (n1078,n137,n102);
and (n1079,n1080,n1081);
xor (n1080,n1077,n1078);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
xor (n1083,n1023,n1024);
and (n1084,n152,n102);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
and (n1087,n1088,n652);
xor (n1088,n1028,n1029);
and (n1089,n117,n47);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
xor (n1092,n1038,n1039);
and (n1093,n110,n47);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
or (n1096,n1097,n1100);
and (n1097,n1098,n1099);
xor (n1098,n1044,n1045);
and (n1099,n65,n47);
and (n1100,n1101,n1102);
xor (n1101,n1098,n1099);
or (n1102,n1103,n1106);
and (n1103,n1104,n1105);
xor (n1104,n1050,n1051);
and (n1105,n57,n47);
and (n1106,n1107,n1108);
xor (n1107,n1104,n1105);
or (n1108,n1109,n1112);
and (n1109,n1110,n1111);
xor (n1110,n1056,n1057);
and (n1111,n89,n47);
and (n1112,n1113,n1114);
xor (n1113,n1110,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
xor (n1116,n1062,n1063);
and (n1117,n83,n47);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1068,n1069);
and (n1123,n143,n47);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1129);
and (n1127,n1128,n590);
xor (n1128,n1074,n1075);
and (n1129,n1130,n1131);
xor (n1130,n1128,n590);
or (n1131,n1132,n1134);
and (n1132,n1133,n645);
xor (n1133,n1080,n1081);
and (n1134,n1135,n1136);
xor (n1135,n1133,n645);
and (n1136,n1137,n1138);
xor (n1137,n1086,n1087);
and (n1138,n170,n47);
and (n1139,n110,n45);
or (n1140,n1141,n1144);
and (n1141,n1142,n1143);
xor (n1142,n1095,n1096);
and (n1143,n65,n45);
and (n1144,n1145,n1146);
xor (n1145,n1142,n1143);
or (n1146,n1147,n1150);
and (n1147,n1148,n1149);
xor (n1148,n1101,n1102);
and (n1149,n57,n45);
and (n1150,n1151,n1152);
xor (n1151,n1148,n1149);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
xor (n1154,n1107,n1108);
and (n1155,n89,n45);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
xor (n1160,n1113,n1114);
and (n1161,n83,n45);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
xor (n1166,n1119,n1120);
and (n1167,n143,n45);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1125,n1126);
and (n1173,n137,n45);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1130,n1131);
and (n1179,n152,n45);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
and (n1182,n1183,n548);
xor (n1183,n1135,n1136);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1145,n1146);
and (n1187,n57,n52);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1151,n1152);
and (n1193,n89,n52);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
or (n1196,n1197,n1200);
and (n1197,n1198,n1199);
xor (n1198,n1157,n1158);
and (n1199,n83,n52);
and (n1200,n1201,n1202);
xor (n1201,n1198,n1199);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
xor (n1204,n1163,n1164);
and (n1205,n143,n52);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
or (n1208,n1209,n1212);
and (n1209,n1210,n1211);
xor (n1210,n1169,n1170);
and (n1211,n137,n52);
and (n1212,n1213,n1214);
xor (n1213,n1210,n1211);
or (n1214,n1215,n1217);
and (n1215,n1216,n461);
xor (n1216,n1175,n1176);
and (n1217,n1218,n1219);
xor (n1218,n1216,n461);
and (n1219,n1220,n1221);
xor (n1220,n1181,n1182);
and (n1221,n170,n52);
and (n1222,n57,n74);
or (n1223,n1224,n1227);
and (n1224,n1225,n1226);
xor (n1225,n1189,n1190);
and (n1226,n89,n74);
and (n1227,n1228,n1229);
xor (n1228,n1225,n1226);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1195,n1196);
and (n1232,n83,n74);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1201,n1202);
and (n1238,n143,n74);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1207,n1208);
and (n1244,n137,n74);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1213,n1214);
and (n1250,n152,n74);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
and (n1253,n1254,n433);
xor (n1254,n1218,n1219);
and (n1255,n89,n79);
or (n1256,n1257,n1260);
and (n1257,n1258,n1259);
xor (n1258,n1228,n1229);
and (n1259,n83,n79);
and (n1260,n1261,n1262);
xor (n1261,n1258,n1259);
or (n1262,n1263,n1266);
and (n1263,n1264,n1265);
xor (n1264,n1234,n1235);
and (n1265,n143,n79);
and (n1266,n1267,n1268);
xor (n1267,n1264,n1265);
or (n1268,n1269,n1272);
and (n1269,n1270,n1271);
xor (n1270,n1240,n1241);
and (n1271,n137,n79);
and (n1272,n1273,n1274);
xor (n1273,n1270,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1246,n1247);
and (n1277,n152,n79);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
and (n1280,n1281,n1282);
xor (n1281,n1252,n1253);
and (n1282,n170,n79);
and (n1283,n83,n128);
or (n1284,n1285,n1288);
and (n1285,n1286,n1287);
xor (n1286,n1261,n1262);
and (n1287,n143,n128);
and (n1288,n1289,n1290);
xor (n1289,n1286,n1287);
or (n1290,n1291,n1294);
and (n1291,n1292,n1293);
xor (n1292,n1267,n1268);
and (n1293,n137,n128);
and (n1294,n1295,n1296);
xor (n1295,n1292,n1293);
or (n1296,n1297,n1300);
and (n1297,n1298,n1299);
xor (n1298,n1273,n1274);
and (n1299,n152,n128);
and (n1300,n1301,n1302);
xor (n1301,n1298,n1299);
and (n1302,n1303,n328);
xor (n1303,n1279,n1280);
and (n1304,n143,n127);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1289,n1290);
and (n1308,n137,n127);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1295,n1296);
and (n1314,n152,n127);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
and (n1317,n1318,n1319);
xor (n1318,n1301,n1302);
and (n1319,n170,n127);
and (n1320,n137,n159);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1310,n1311);
and (n1324,n152,n159);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
and (n1327,n1328,n247);
xor (n1328,n1316,n1317);
and (n1329,n152,n153);
and (n1330,n1331,n1332);
xor (n1331,n1326,n1327);
and (n1332,n170,n153);
and (n1333,n170,n179);
endmodule
