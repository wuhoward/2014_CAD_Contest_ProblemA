module top (out,n17,n19,n20,n24,n29,n31,n34,n39,n41
        ,n43,n46,n53,n55,n57,n60,n65,n67,n69,n72
        ,n88,n90,n93,n148,n180,n365,n379,n380,n452,n461
        ,n462,n498,n570,n600,n601,n791,n795,n797,n823,n824
        ,n931,n948,n949,n1135,n1139,n1141,n1152,n1164,n1178);
output out;
input n17;
input n19;
input n20;
input n24;
input n29;
input n31;
input n34;
input n39;
input n41;
input n43;
input n46;
input n53;
input n55;
input n57;
input n60;
input n65;
input n67;
input n69;
input n72;
input n88;
input n90;
input n93;
input n148;
input n180;
input n365;
input n379;
input n380;
input n452;
input n461;
input n462;
input n498;
input n570;
input n600;
input n601;
input n791;
input n795;
input n797;
input n823;
input n824;
input n931;
input n948;
input n949;
input n1135;
input n1139;
input n1141;
input n1152;
input n1164;
input n1178;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n42;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n56;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n68;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n792;
wire n793;
wire n794;
wire n796;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1136;
wire n1137;
wire n1138;
wire n1140;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
xor (out,n0,n3104);
xnor (n0,n1,n3078);
nand (n1,n2,n340);
nor (n2,n3,n334);
nor (n3,n4,n270);
nor (n4,n5,n268);
nor (n5,n6,n231);
nand (n6,n7,n191);
nand (n7,n8,n137,n190);
nand (n8,n9,n95);
nand (n9,n10,n74,n94);
nand (n10,n11,n48);
nand (n11,n12,n35,n47);
nand (n12,n13,n25);
not (n13,n14);
xor (n14,n15,n24);
or (n15,n16,n21);
and (n16,n17,n18);
xor (n18,n19,n20);
and (n21,n17,n22);
nor (n22,n18,n23);
xnor (n23,n24,n19);
xor (n25,n26,n34);
or (n26,n27,n30);
and (n27,n17,n28);
xor (n28,n29,n24);
and (n30,n31,n32);
nor (n32,n28,n33);
xnor (n33,n34,n29);
nand (n35,n36,n25);
xor (n36,n37,n46);
or (n37,n38,n42);
and (n38,n39,n40);
xor (n40,n41,n34);
and (n42,n43,n44);
nor (n44,n40,n45);
xnor (n45,n46,n41);
nand (n47,n13,n36);
nand (n48,n49,n61,n73);
nand (n49,n50,n14);
xor (n50,n51,n60);
or (n51,n52,n56);
and (n52,n53,n54);
xor (n54,n55,n46);
and (n56,n57,n58);
nor (n58,n54,n59);
xnor (n59,n60,n55);
nand (n61,n62,n14);
xor (n62,n63,n72);
or (n63,n64,n68);
and (n64,n65,n66);
xor (n66,n67,n60);
and (n68,n69,n70);
nor (n70,n66,n71);
xnor (n71,n72,n67);
nand (n73,n50,n62);
nand (n74,n75,n48);
xor (n75,n76,n84);
xor (n76,n77,n80);
xor (n77,n78,n34);
or (n78,n27,n79);
and (n79,n17,n32);
xor (n80,n81,n72);
or (n81,n82,n83);
and (n82,n57,n66);
and (n83,n65,n70);
xor (n84,n85,n93);
or (n85,n86,n89);
and (n86,n69,n87);
xor (n87,n88,n72);
and (n89,n90,n91);
nor (n91,n87,n92);
xnor (n92,n93,n88);
nand (n94,n11,n75);
xor (n95,n96,n120);
xor (n96,n97,n110);
nand (n97,n98,n108,n109);
nand (n98,n99,n103);
xor (n99,n100,n60);
or (n100,n101,n102);
and (n101,n43,n54);
and (n102,n53,n58);
not (n103,n104);
xor (n104,n105,n46);
or (n105,n106,n107);
and (n106,n31,n40);
and (n107,n39,n44);
nand (n108,n93,n103);
nand (n109,n99,n93);
xor (n110,n111,n93);
xor (n111,n112,n116);
xor (n112,n113,n93);
or (n113,n114,n115);
and (n114,n65,n87);
and (n115,n69,n91);
xor (n116,n117,n60);
or (n117,n118,n119);
and (n118,n39,n54);
and (n119,n43,n58);
xor (n120,n121,n126);
xor (n121,n104,n122);
nand (n122,n123,n124,n125);
nand (n123,n77,n80);
nand (n124,n84,n80);
nand (n125,n77,n84);
xor (n126,n127,n133);
xor (n127,n128,n129);
not (n128,n77);
xor (n129,n130,n46);
or (n130,n131,n132);
and (n131,n17,n40);
and (n132,n31,n44);
xor (n133,n134,n72);
or (n134,n135,n136);
and (n135,n53,n66);
and (n136,n57,n70);
nand (n137,n138,n95);
nand (n138,n139,n167,n189);
nand (n139,n140,n142);
xor (n140,n141,n93);
xor (n141,n99,n103);
nand (n142,n143,n149,n166);
nand (n143,n144,n93);
xor (n144,n145,n93);
or (n145,n146,n147);
and (n146,n90,n87);
and (n147,n148,n91);
nand (n149,n150,n93);
nand (n150,n151,n160,n165);
nand (n151,n152,n156);
xor (n152,n153,n34);
or (n153,n154,n155);
and (n154,n31,n28);
and (n155,n39,n32);
xor (n156,n157,n46);
or (n157,n158,n159);
and (n158,n43,n40);
and (n159,n53,n44);
nand (n160,n161,n156);
xor (n161,n162,n60);
or (n162,n163,n164);
and (n163,n57,n54);
and (n164,n65,n58);
nand (n165,n152,n161);
nand (n166,n144,n150);
nand (n167,n168,n142);
nand (n168,n169,n185,n188);
nand (n169,n170,n183);
nand (n170,n171,n181,n182);
nand (n171,n172,n176);
xor (n172,n173,n72);
or (n173,n174,n175);
and (n174,n69,n66);
and (n175,n90,n70);
xor (n176,n177,n93);
or (n177,n178,n179);
and (n178,n148,n87);
and (n179,n180,n91);
nand (n181,n13,n176);
nand (n182,n172,n13);
xor (n183,n184,n36);
xor (n184,n13,n25);
nand (n185,n186,n183);
xor (n186,n187,n62);
xor (n187,n50,n14);
nand (n188,n170,n186);
nand (n189,n140,n168);
nand (n190,n9,n138);
xor (n191,n192,n227);
xor (n192,n193,n197);
nand (n193,n194,n195,n196);
nand (n194,n104,n122);
nand (n195,n126,n122);
nand (n196,n104,n126);
xor (n197,n198,n217);
xor (n198,n199,n213);
xor (n199,n200,n209);
xor (n200,n201,n205);
xor (n201,n202,n60);
or (n202,n203,n204);
and (n203,n31,n54);
and (n204,n39,n58);
xor (n205,n206,n93);
or (n206,n207,n208);
and (n207,n57,n87);
and (n208,n65,n91);
xor (n209,n210,n72);
or (n210,n211,n212);
and (n211,n43,n66);
and (n212,n53,n70);
nand (n213,n214,n215,n216);
nand (n214,n112,n116);
nand (n215,n93,n116);
nand (n216,n112,n93);
xor (n217,n218,n223);
xor (n218,n219,n93);
not (n219,n220);
xor (n220,n221,n46);
or (n221,n131,n222);
and (n222,n17,n44);
nand (n223,n224,n225,n226);
nand (n224,n128,n129);
nand (n225,n133,n129);
nand (n226,n128,n133);
nand (n227,n228,n229,n230);
nand (n228,n97,n110);
nand (n229,n120,n110);
nand (n230,n97,n120);
nor (n231,n232,n264);
xor (n232,n233,n260);
xor (n233,n234,n238);
nand (n234,n235,n236,n237);
nand (n235,n219,n93);
nand (n236,n223,n93);
nand (n237,n219,n223);
xor (n238,n239,n254);
xor (n239,n240,n244);
nand (n240,n241,n242,n243);
nand (n241,n201,n205);
nand (n242,n209,n205);
nand (n243,n201,n209);
xor (n244,n245,n250);
xor (n245,n219,n246);
xor (n246,n247,n60);
or (n247,n248,n249);
and (n248,n17,n54);
and (n249,n31,n58);
xor (n250,n251,n93);
or (n251,n252,n253);
and (n252,n53,n87);
and (n253,n57,n91);
xor (n254,n255,n220);
xor (n255,n256,n93);
xor (n256,n257,n72);
or (n257,n258,n259);
and (n258,n39,n66);
and (n259,n43,n70);
nand (n260,n261,n262,n263);
nand (n261,n199,n213);
nand (n262,n217,n213);
nand (n263,n199,n217);
nand (n264,n265,n266,n267);
nand (n265,n193,n197);
nand (n266,n227,n197);
nand (n267,n193,n227);
not (n268,n269);
nand (n269,n232,n264);
not (n270,n271);
nor (n271,n272,n307);
nor (n272,n273,n303);
xor (n273,n274,n299);
xor (n274,n275,n285);
xor (n275,n276,n93);
xor (n276,n277,n281);
xor (n277,n278,n72);
or (n278,n279,n280);
and (n279,n31,n66);
and (n280,n39,n70);
xor (n281,n282,n93);
or (n282,n283,n284);
and (n283,n43,n87);
and (n284,n53,n91);
xor (n285,n286,n295);
xor (n286,n287,n291);
not (n287,n288);
xor (n288,n289,n60);
or (n289,n248,n290);
and (n290,n17,n58);
nand (n291,n292,n293,n294);
nand (n292,n219,n246);
nand (n293,n250,n246);
nand (n294,n219,n250);
nand (n295,n296,n297,n298);
nand (n296,n256,n93);
nand (n297,n220,n93);
nand (n298,n256,n220);
nand (n299,n300,n301,n302);
nand (n300,n240,n244);
nand (n301,n254,n244);
nand (n302,n240,n254);
nand (n303,n304,n305,n306);
nand (n304,n234,n238);
nand (n305,n260,n238);
nand (n306,n234,n260);
nor (n307,n308,n312);
nand (n308,n309,n310,n311);
nand (n309,n275,n285);
nand (n310,n299,n285);
nand (n311,n275,n299);
xor (n312,n313,n330);
xor (n313,n314,n318);
nand (n314,n315,n316,n317);
nand (n315,n277,n281);
nand (n316,n93,n281);
nand (n317,n277,n93);
xor (n318,n319,n320);
xor (n319,n93,n288);
xor (n320,n321,n326);
xor (n321,n287,n322);
xor (n322,n323,n72);
or (n323,n324,n325);
and (n324,n17,n66);
and (n325,n31,n70);
xor (n326,n327,n93);
or (n327,n328,n329);
and (n328,n39,n87);
and (n329,n43,n91);
nand (n330,n331,n332,n333);
nand (n331,n287,n291);
nand (n332,n295,n291);
nand (n333,n287,n295);
not (n334,n335);
nor (n335,n336,n338);
nor (n336,n337,n307);
nand (n337,n273,n303);
not (n338,n339);
nand (n339,n308,n312);
nand (n340,n341,n3074);
nand (n341,n342,n1112);
nor (n342,n343,n1097);
nor (n343,n344,n690);
nand (n344,n345,n667);
nor (n345,n346,n643);
nor (n346,n347,n520);
xor (n347,n348,n477);
xor (n348,n349,n368);
xor (n349,n350,n355);
xor (n350,n351,n353);
xor (n351,n352,n161);
xor (n352,n152,n156);
xor (n353,n354,n13);
xor (n354,n172,n176);
nand (n355,n356,n366,n367);
nand (n356,n357,n361);
xor (n357,n358,n72);
or (n358,n359,n360);
and (n359,n90,n66);
and (n360,n148,n70);
xor (n361,n362,n93);
or (n362,n363,n364);
and (n363,n180,n87);
and (n364,n365,n91);
nand (n366,n93,n361);
nand (n367,n357,n93);
xor (n368,n369,n439);
xor (n369,n370,n405);
xor (n370,n371,n393);
xor (n371,n93,n372);
nand (n372,n373,n387,n392);
nand (n373,n374,n384);
not (n374,n375);
xor (n375,n376,n20);
or (n376,n377,n381);
and (n377,n17,n378);
xor (n378,n379,n380);
and (n381,n17,n382);
nor (n382,n378,n383);
xnor (n383,n20,n379);
xor (n384,n385,n24);
or (n385,n16,n386);
and (n386,n31,n22);
nand (n387,n388,n384);
xor (n388,n389,n46);
or (n389,n390,n391);
and (n390,n53,n40);
and (n391,n57,n44);
nand (n392,n374,n388);
nand (n393,n394,n399,n404);
nand (n394,n395,n375);
xor (n395,n396,n34);
or (n396,n397,n398);
and (n397,n39,n28);
and (n398,n43,n32);
nand (n399,n400,n375);
xor (n400,n401,n60);
or (n401,n402,n403);
and (n402,n65,n54);
and (n403,n69,n58);
nand (n404,n395,n400);
nand (n405,n406,n425,n438);
nand (n406,n407,n409);
xor (n407,n408,n388);
xor (n408,n374,n384);
nand (n409,n410,n419,n424);
nand (n410,n411,n415);
xor (n411,n412,n24);
or (n412,n413,n414);
and (n413,n31,n18);
and (n414,n39,n22);
xor (n415,n416,n46);
or (n416,n417,n418);
and (n417,n57,n40);
and (n418,n65,n44);
nand (n419,n420,n415);
xor (n420,n421,n34);
or (n421,n422,n423);
and (n422,n43,n28);
and (n423,n53,n32);
nand (n424,n411,n420);
nand (n425,n426,n409);
nand (n426,n427,n432,n437);
nand (n427,n374,n428);
xor (n428,n429,n60);
or (n429,n430,n431);
and (n430,n69,n54);
and (n431,n90,n58);
nand (n432,n433,n428);
xor (n433,n434,n72);
or (n434,n435,n436);
and (n435,n148,n66);
and (n436,n180,n70);
nand (n437,n374,n433);
nand (n438,n407,n426);
nand (n439,n440,n445,n476);
nand (n440,n441,n443);
xor (n441,n442,n93);
xor (n442,n357,n361);
xor (n443,n444,n400);
xor (n444,n395,n375);
nand (n445,n446,n443);
nand (n446,n447,n453,n475);
nand (n447,n448,n93);
xor (n448,n449,n93);
or (n449,n450,n451);
and (n450,n365,n87);
and (n451,n452,n91);
nand (n453,n454,n93);
nand (n454,n455,n469,n474);
nand (n455,n456,n466);
not (n456,n457);
xor (n457,n458,n380);
or (n458,n459,n463);
and (n459,n17,n460);
xor (n460,n461,n462);
and (n463,n17,n464);
nor (n464,n460,n465);
xnor (n465,n380,n461);
xor (n466,n467,n20);
or (n467,n377,n468);
and (n468,n31,n382);
nand (n469,n470,n466);
xor (n470,n471,n24);
or (n471,n472,n473);
and (n472,n39,n18);
and (n473,n43,n22);
nand (n474,n456,n470);
nand (n475,n448,n454);
nand (n476,n441,n446);
nand (n477,n478,n516,n519);
nand (n478,n479,n514);
nand (n479,n480,n500,n513);
nand (n480,n481,n483);
xor (n481,n482,n420);
xor (n482,n411,n415);
nand (n483,n484,n493,n499);
nand (n484,n485,n489);
xor (n485,n486,n34);
or (n486,n487,n488);
and (n487,n53,n28);
and (n488,n57,n32);
xor (n489,n490,n46);
or (n490,n491,n492);
and (n491,n65,n40);
and (n492,n69,n44);
nand (n493,n494,n489);
xor (n494,n495,n93);
or (n495,n496,n497);
and (n496,n452,n87);
and (n497,n498,n91);
nand (n499,n485,n494);
nand (n500,n501,n483);
nand (n501,n502,n507,n512);
nand (n502,n457,n503);
xor (n503,n504,n60);
or (n504,n505,n506);
and (n505,n90,n54);
and (n506,n148,n58);
nand (n507,n508,n503);
xor (n508,n509,n72);
or (n509,n510,n511);
and (n510,n180,n66);
and (n511,n365,n70);
nand (n512,n457,n508);
nand (n513,n481,n501);
xor (n514,n515,n426);
xor (n515,n407,n409);
nand (n516,n517,n514);
xor (n517,n518,n446);
xor (n518,n441,n443);
nand (n519,n479,n517);
nand (n520,n521,n553,n642);
nand (n521,n522,n551);
nand (n522,n523,n527,n550);
nand (n523,n524,n526);
xor (n524,n525,n433);
xor (n525,n374,n428);
xor (n526,n449,n454);
nand (n527,n528,n526);
nand (n528,n529,n532,n549);
nand (n529,n93,n530);
xor (n530,n531,n470);
xor (n531,n456,n466);
nand (n532,n533,n530);
nand (n533,n534,n543,n548);
nand (n534,n535,n539);
xor (n535,n536,n20);
or (n536,n537,n538);
and (n537,n31,n378);
and (n538,n39,n382);
xor (n539,n540,n24);
or (n540,n541,n542);
and (n541,n43,n18);
and (n542,n53,n22);
nand (n543,n544,n539);
xor (n544,n545,n34);
or (n545,n546,n547);
and (n546,n57,n28);
and (n547,n65,n32);
nand (n548,n535,n544);
nand (n549,n93,n533);
nand (n550,n524,n528);
xor (n551,n552,n517);
xor (n552,n479,n514);
nand (n553,n554,n551);
nand (n554,n555,n579,n641);
nand (n555,n556,n558);
xor (n556,n557,n501);
xor (n557,n481,n483);
nand (n558,n559,n575,n578);
nand (n559,n560,n573);
nand (n560,n561,n571,n572);
nand (n561,n562,n566);
xor (n562,n563,n46);
or (n563,n564,n565);
and (n564,n69,n40);
and (n565,n90,n44);
xor (n566,n567,n93);
or (n567,n568,n569);
and (n568,n498,n87);
and (n569,n570,n91);
nand (n571,n456,n566);
nand (n572,n562,n456);
xor (n573,n574,n494);
xor (n574,n485,n489);
nand (n575,n576,n573);
xor (n576,n577,n508);
xor (n577,n457,n503);
nand (n578,n560,n576);
nand (n579,n580,n558);
nand (n580,n581,n637,n640);
nand (n581,n582,n615);
nand (n582,n583,n592,n614);
nand (n583,n584,n588);
xor (n584,n585,n60);
or (n585,n586,n587);
and (n586,n148,n54);
and (n587,n180,n58);
xor (n588,n589,n72);
or (n589,n590,n591);
and (n590,n365,n66);
and (n591,n452,n70);
nand (n592,n593,n588);
nand (n593,n594,n608,n613);
nand (n594,n595,n605);
not (n595,n596);
xor (n596,n597,n462);
or (n597,n598,n602);
and (n598,n17,n599);
xor (n599,n600,n601);
and (n602,n17,n603);
nor (n603,n599,n604);
xnor (n604,n462,n600);
xor (n605,n606,n380);
or (n606,n459,n607);
and (n607,n31,n464);
nand (n608,n609,n605);
xor (n609,n610,n24);
or (n610,n611,n612);
and (n611,n53,n18);
and (n612,n57,n22);
nand (n613,n595,n609);
nand (n614,n584,n593);
nand (n615,n616,n619,n636);
nand (n616,n93,n617);
xor (n617,n618,n544);
xor (n618,n535,n539);
nand (n619,n620,n617);
nand (n620,n621,n630,n635);
nand (n621,n622,n626);
xor (n622,n623,n20);
or (n623,n624,n625);
and (n624,n39,n378);
and (n625,n43,n382);
xor (n626,n627,n34);
or (n627,n628,n629);
and (n628,n65,n28);
and (n629,n69,n32);
nand (n630,n631,n626);
xor (n631,n632,n46);
or (n632,n633,n634);
and (n633,n90,n40);
and (n634,n148,n44);
nand (n635,n622,n631);
nand (n636,n93,n620);
nand (n637,n638,n615);
xor (n638,n639,n533);
xor (n639,n93,n530);
nand (n640,n582,n638);
nand (n641,n556,n580);
nand (n642,n522,n554);
nor (n643,n644,n648);
nand (n644,n645,n646,n647);
nand (n645,n349,n368);
nand (n646,n477,n368);
nand (n647,n349,n477);
xor (n648,n649,n663);
xor (n649,n650,n654);
nand (n650,n651,n652,n653);
nand (n651,n351,n353);
nand (n652,n355,n353);
nand (n653,n351,n355);
xor (n654,n655,n661);
xor (n655,n656,n660);
nand (n656,n657,n658,n659);
nand (n657,n93,n372);
nand (n658,n393,n372);
nand (n659,n93,n393);
xor (n660,n145,n150);
xor (n661,n662,n186);
xor (n662,n170,n183);
nand (n663,n664,n665,n666);
nand (n664,n370,n405);
nand (n665,n439,n405);
nand (n666,n370,n439);
nor (n667,n668,n683);
nor (n668,n669,n673);
nand (n669,n670,n671,n672);
nand (n670,n650,n654);
nand (n671,n663,n654);
nand (n672,n650,n663);
xor (n673,n674,n679);
xor (n674,n675,n677);
xor (n675,n676,n75);
xor (n676,n11,n48);
xor (n677,n678,n168);
xor (n678,n140,n142);
nand (n679,n680,n681,n682);
nand (n680,n656,n660);
nand (n681,n661,n660);
nand (n682,n656,n661);
nor (n683,n684,n688);
nand (n684,n685,n686,n687);
nand (n685,n675,n677);
nand (n686,n679,n677);
nand (n687,n675,n679);
xor (n688,n689,n138);
xor (n689,n9,n95);
nor (n690,n691,n1091);
nor (n691,n692,n1067);
nor (n692,n693,n1065);
nor (n693,n694,n1040);
nand (n694,n695,n1002);
nand (n695,n696,n918,n1001);
nand (n696,n697,n781);
xor (n697,n698,n771);
xor (n698,n699,n721);
xor (n699,n700,n705);
xor (n700,n701,n93);
xor (n701,n702,n60);
or (n702,n703,n704);
and (n703,n180,n54);
and (n704,n365,n58);
nand (n705,n706,n715,n720);
nand (n706,n707,n711);
xor (n707,n708,n24);
or (n708,n709,n710);
and (n709,n57,n18);
and (n710,n65,n22);
xor (n711,n712,n380);
or (n712,n713,n714);
and (n713,n31,n460);
and (n714,n39,n464);
nand (n715,n716,n711);
xor (n716,n717,n20);
or (n717,n718,n719);
and (n718,n43,n378);
and (n719,n53,n382);
nand (n720,n707,n716);
nand (n721,n722,n753,n770);
nand (n722,n723,n739);
nand (n723,n724,n733,n738);
nand (n724,n725,n729);
xor (n725,n726,n24);
or (n726,n727,n728);
and (n727,n65,n18);
and (n728,n69,n22);
xor (n729,n730,n380);
or (n730,n731,n732);
and (n731,n39,n460);
and (n732,n43,n464);
nand (n733,n734,n729);
xor (n734,n735,n34);
or (n735,n736,n737);
and (n736,n90,n28);
and (n737,n148,n32);
nand (n738,n725,n734);
xor (n739,n740,n749);
xor (n740,n741,n745);
xor (n741,n742,n34);
or (n742,n743,n744);
and (n743,n69,n28);
and (n744,n90,n32);
xor (n745,n746,n46);
or (n746,n747,n748);
and (n747,n148,n40);
and (n748,n180,n44);
xor (n749,n750,n72);
or (n750,n751,n752);
and (n751,n498,n66);
and (n752,n570,n70);
nand (n753,n754,n739);
nand (n754,n755,n764,n769);
nand (n755,n756,n760);
xor (n756,n757,n462);
or (n757,n758,n759);
and (n758,n31,n599);
and (n759,n39,n603);
xor (n760,n761,n46);
or (n761,n762,n763);
and (n762,n180,n40);
and (n763,n365,n44);
nand (n764,n765,n760);
xor (n765,n766,n60);
or (n766,n767,n768);
and (n767,n452,n54);
and (n768,n498,n58);
nand (n769,n756,n765);
nand (n770,n723,n754);
xor (n771,n772,n777);
xor (n772,n773,n775);
xor (n773,n774,n609);
xor (n774,n595,n605);
xor (n775,n776,n631);
xor (n776,n622,n626);
nand (n777,n778,n779,n780);
nand (n778,n741,n745);
nand (n779,n749,n745);
nand (n780,n741,n749);
xor (n781,n782,n857);
xor (n782,n783,n837);
nand (n783,n784,n810,n836);
nand (n784,n785,n800);
nand (n785,n786,n798,n799);
nand (n786,n787,n792);
xor (n787,n788,n72);
or (n788,n789,n790);
and (n789,n570,n66);
and (n790,n791,n70);
xor (n792,n793,n93);
or (n793,n794,n796);
and (n794,n795,n87);
and (n796,n797,n91);
nand (n798,n93,n792);
nand (n799,n787,n93);
xor (n800,n801,n806);
xor (n801,n802,n595);
xor (n802,n803,n93);
or (n803,n804,n805);
and (n804,n791,n87);
and (n805,n795,n91);
xor (n806,n807,n60);
or (n807,n808,n809);
and (n808,n365,n54);
and (n809,n452,n58);
nand (n810,n811,n800);
xor (n811,n812,n834);
xor (n812,n93,n813);
nand (n813,n814,n828,n833);
nand (n814,n815,n818);
xor (n815,n816,n462);
or (n816,n598,n817);
and (n817,n31,n603);
not (n818,n819);
xor (n819,n820,n601);
or (n820,n821,n825);
and (n821,n17,n822);
xor (n822,n823,n824);
and (n825,n17,n826);
nor (n826,n822,n827);
xnor (n827,n601,n823);
nand (n828,n829,n818);
xor (n829,n830,n20);
or (n830,n831,n832);
and (n831,n53,n378);
and (n832,n57,n382);
nand (n833,n815,n829);
xor (n834,n835,n716);
xor (n835,n707,n711);
nand (n836,n785,n811);
xor (n837,n838,n853);
xor (n838,n839,n843);
nand (n839,n840,n841,n842);
nand (n840,n802,n595);
nand (n841,n806,n595);
nand (n842,n802,n806);
xor (n843,n844,n596);
xor (n844,n845,n849);
xor (n845,n846,n72);
or (n846,n847,n848);
and (n847,n452,n66);
and (n848,n498,n70);
xor (n849,n850,n93);
or (n850,n851,n852);
and (n851,n570,n87);
and (n852,n791,n91);
nand (n853,n854,n855,n856);
nand (n854,n93,n813);
nand (n855,n834,n813);
nand (n856,n93,n834);
nand (n857,n858,n914,n917);
nand (n858,n859,n879);
nand (n859,n860,n875,n878);
nand (n860,n861,n873);
nand (n861,n862,n867,n872);
nand (n862,n819,n863);
xor (n863,n864,n20);
or (n864,n865,n866);
and (n865,n57,n378);
and (n866,n65,n382);
nand (n867,n868,n863);
xor (n868,n869,n24);
or (n869,n870,n871);
and (n870,n69,n18);
and (n871,n90,n22);
nand (n872,n819,n868);
xor (n873,n874,n734);
xor (n874,n725,n729);
nand (n875,n876,n873);
xor (n876,n877,n829);
xor (n877,n815,n818);
nand (n878,n861,n876);
nand (n879,n880,n910,n913);
nand (n880,n881,n894);
nand (n881,n882,n888,n893);
nand (n882,n883,n887);
xor (n883,n884,n380);
or (n884,n885,n886);
and (n885,n43,n460);
and (n886,n53,n464);
not (n887,n756);
nand (n888,n889,n887);
xor (n889,n890,n34);
or (n890,n891,n892);
and (n891,n148,n28);
and (n892,n180,n32);
nand (n893,n883,n889);
nand (n894,n895,n904,n909);
nand (n895,n896,n900);
xor (n896,n897,n46);
or (n897,n898,n899);
and (n898,n365,n40);
and (n899,n452,n44);
xor (n900,n901,n60);
or (n901,n902,n903);
and (n902,n498,n54);
and (n903,n570,n58);
nand (n904,n905,n900);
xor (n905,n906,n72);
or (n906,n907,n908);
and (n907,n791,n66);
and (n908,n795,n70);
nand (n909,n896,n905);
nand (n910,n911,n894);
xor (n911,n912,n765);
xor (n912,n756,n760);
nand (n913,n881,n911);
nand (n914,n915,n879);
xor (n915,n916,n754);
xor (n916,n723,n739);
nand (n917,n859,n915);
nand (n918,n919,n781);
nand (n919,n920,n997,n1000);
nand (n920,n921,n923);
xor (n921,n922,n811);
xor (n922,n785,n800);
nand (n923,n924,n957,n996);
nand (n924,n925,n955);
nand (n925,n926,n932,n954);
nand (n926,n927,n93);
xor (n927,n928,n93);
or (n928,n929,n930);
and (n929,n797,n87);
and (n930,n931,n91);
nand (n932,n933,n93);
nand (n933,n934,n942,n953);
nand (n934,n935,n938);
xor (n935,n936,n601);
or (n936,n821,n937);
and (n937,n31,n826);
xor (n938,n939,n462);
or (n939,n940,n941);
and (n940,n39,n599);
and (n941,n43,n603);
nand (n942,n943,n938);
not (n943,n944);
xor (n944,n945,n824);
or (n945,n946,n950);
and (n946,n17,n947);
xor (n947,n948,n949);
and (n950,n17,n951);
nor (n951,n947,n952);
xnor (n952,n824,n948);
nand (n953,n935,n943);
nand (n954,n927,n933);
xor (n955,n956,n93);
xor (n956,n787,n792);
nand (n957,n958,n955);
nand (n958,n959,n978,n995);
nand (n959,n960,n976);
nand (n960,n961,n970,n975);
nand (n961,n962,n966);
xor (n962,n963,n380);
or (n963,n964,n965);
and (n964,n53,n460);
and (n965,n57,n464);
xor (n966,n967,n20);
or (n967,n968,n969);
and (n968,n65,n378);
and (n969,n69,n382);
nand (n970,n971,n966);
xor (n971,n972,n24);
or (n972,n973,n974);
and (n973,n90,n18);
and (n974,n148,n22);
nand (n975,n962,n971);
xor (n976,n977,n868);
xor (n977,n819,n863);
nand (n978,n979,n976);
nand (n979,n980,n989,n994);
nand (n980,n981,n985);
xor (n981,n982,n46);
or (n982,n983,n984);
and (n983,n452,n40);
and (n984,n498,n44);
xor (n985,n986,n601);
or (n986,n987,n988);
and (n987,n31,n822);
and (n988,n39,n826);
nand (n989,n990,n985);
xor (n990,n991,n34);
or (n991,n992,n993);
and (n992,n180,n28);
and (n993,n365,n32);
nand (n994,n981,n990);
nand (n995,n960,n979);
nand (n996,n925,n958);
nand (n997,n998,n923);
xor (n998,n999,n915);
xor (n999,n859,n879);
nand (n1000,n921,n998);
nand (n1001,n697,n919);
xor (n1002,n1003,n1036);
xor (n1003,n1004,n1008);
nand (n1004,n1005,n1006,n1007);
nand (n1005,n699,n721);
nand (n1006,n771,n721);
nand (n1007,n699,n771);
xor (n1008,n1009,n1024);
xor (n1009,n1010,n1014);
nand (n1010,n1011,n1012,n1013);
nand (n1011,n839,n843);
nand (n1012,n853,n843);
nand (n1013,n839,n853);
xor (n1014,n1015,n1022);
xor (n1015,n1016,n1020);
nand (n1016,n1017,n1018,n1019);
nand (n1017,n845,n849);
nand (n1018,n596,n849);
nand (n1019,n845,n596);
xor (n1020,n1021,n593);
xor (n1021,n584,n588);
xor (n1022,n1023,n456);
xor (n1023,n562,n566);
xor (n1024,n1025,n1032);
xor (n1025,n1026,n1030);
nand (n1026,n1027,n1028,n1029);
nand (n1027,n701,n93);
nand (n1028,n705,n93);
nand (n1029,n701,n705);
xor (n1030,n1031,n620);
xor (n1031,n93,n617);
nand (n1032,n1033,n1034,n1035);
nand (n1033,n773,n775);
nand (n1034,n777,n775);
nand (n1035,n773,n777);
nand (n1036,n1037,n1038,n1039);
nand (n1037,n783,n837);
nand (n1038,n857,n837);
nand (n1039,n783,n857);
nor (n1040,n1041,n1045);
nand (n1041,n1042,n1043,n1044);
nand (n1042,n1004,n1008);
nand (n1043,n1036,n1008);
nand (n1044,n1004,n1036);
xor (n1045,n1046,n1061);
xor (n1046,n1047,n1049);
xor (n1047,n1048,n638);
xor (n1048,n582,n615);
xor (n1049,n1050,n1057);
xor (n1050,n1051,n1053);
xor (n1051,n1052,n576);
xor (n1052,n560,n573);
nand (n1053,n1054,n1055,n1056);
nand (n1054,n1016,n1020);
nand (n1055,n1022,n1020);
nand (n1056,n1016,n1022);
nand (n1057,n1058,n1059,n1060);
nand (n1058,n1026,n1030);
nand (n1059,n1032,n1030);
nand (n1060,n1026,n1032);
nand (n1061,n1062,n1063,n1064);
nand (n1062,n1010,n1014);
nand (n1063,n1024,n1014);
nand (n1064,n1010,n1024);
not (n1065,n1066);
nand (n1066,n1041,n1045);
not (n1067,n1068);
nor (n1068,n1069,n1084);
nor (n1069,n1070,n1074);
nand (n1070,n1071,n1072,n1073);
nand (n1071,n1047,n1049);
nand (n1072,n1061,n1049);
nand (n1073,n1047,n1061);
xor (n1074,n1075,n1080);
xor (n1075,n1076,n1078);
xor (n1076,n1077,n528);
xor (n1077,n524,n526);
xor (n1078,n1079,n580);
xor (n1079,n556,n558);
nand (n1080,n1081,n1082,n1083);
nand (n1081,n1051,n1053);
nand (n1082,n1057,n1053);
nand (n1083,n1051,n1057);
nor (n1084,n1085,n1089);
nand (n1085,n1086,n1087,n1088);
nand (n1086,n1076,n1078);
nand (n1087,n1080,n1078);
nand (n1088,n1076,n1080);
xor (n1089,n1090,n554);
xor (n1090,n522,n551);
not (n1091,n1092);
nor (n1092,n1093,n1095);
nor (n1093,n1094,n1084);
nand (n1094,n1070,n1074);
not (n1095,n1096);
nand (n1096,n1085,n1089);
not (n1097,n1098);
nor (n1098,n1099,n1106);
nor (n1099,n1100,n1105);
nor (n1100,n1101,n1103);
nor (n1101,n1102,n643);
nand (n1102,n347,n520);
not (n1103,n1104);
nand (n1104,n644,n648);
not (n1105,n667);
not (n1106,n1107);
nor (n1107,n1108,n1110);
nor (n1108,n1109,n683);
nand (n1109,n669,n673);
not (n1110,n1111);
nand (n1111,n684,n688);
nand (n1112,n1113,n1117);
nor (n1113,n1114,n344);
nand (n1114,n1115,n1068);
nor (n1115,n1116,n1040);
nor (n1116,n695,n1002);
nand (n1117,n1118,n2648);
nor (n1118,n1119,n2616);
nor (n1119,n1120,n2089);
nor (n1120,n1121,n2074);
nor (n1121,n1122,n1795);
nand (n1122,n1123,n1578);
nor (n1123,n1124,n1477);
nor (n1124,n1125,n1387);
nand (n1125,n1126,n1302,n1386);
nand (n1126,n1127,n1204);
xor (n1127,n1128,n1180);
xor (n1128,n1129,n1154);
xor (n1129,n1130,n1142);
xor (n1130,n1131,n1136);
xor (n1131,n1132,n34);
or (n1132,n1133,n1134);
and (n1133,n931,n28);
and (n1134,n1135,n32);
xor (n1136,n1137,n46);
or (n1137,n1138,n1140);
and (n1138,n1139,n40);
and (n1140,n1141,n44);
xor (n1142,n1143,n1147);
xor (n1143,n1144,n824);
or (n1144,n1145,n1146);
and (n1145,n65,n947);
and (n1146,n69,n951);
xnor (n1147,n1148,n949);
nor (n1148,n1149,n1153);
and (n1149,n57,n1150);
and (n1150,n1151,n949);
not (n1151,n1152);
and (n1153,n53,n1152);
nand (n1154,n1155,n1165,n1179);
nand (n1155,n1156,n1160);
xor (n1156,n1157,n34);
or (n1157,n1158,n1159);
and (n1158,n1135,n28);
and (n1159,n1139,n32);
xor (n1160,n1161,n46);
or (n1161,n1162,n1163);
and (n1162,n1141,n40);
and (n1163,n1164,n44);
nand (n1165,n1166,n1160);
xor (n1166,n1167,n1176);
xor (n1167,n1168,n1172);
xor (n1168,n1169,n824);
or (n1169,n1170,n1171);
and (n1170,n69,n947);
and (n1171,n90,n951);
xor (n1172,n1173,n462);
or (n1173,n1174,n1175);
and (n1174,n365,n599);
and (n1175,n452,n603);
xnor (n1176,n1177,n60);
nand (n1177,n1178,n54);
nand (n1179,n1156,n1166);
xor (n1180,n1181,n1190);
xor (n1181,n1182,n1186);
xor (n1182,n1183,n60);
or (n1183,n1184,n1185);
and (n1184,n1164,n54);
and (n1185,n1178,n58);
nand (n1186,n1187,n1188,n1189);
nand (n1187,n1168,n1172);
nand (n1188,n1176,n1172);
nand (n1189,n1168,n1176);
xor (n1190,n1191,n1200);
xor (n1191,n1192,n1196);
xor (n1192,n1193,n462);
or (n1193,n1194,n1195);
and (n1194,n180,n599);
and (n1195,n365,n603);
xor (n1196,n1197,n601);
or (n1197,n1198,n1199);
and (n1198,n90,n822);
and (n1199,n148,n826);
xor (n1200,n1201,n380);
or (n1201,n1202,n1203);
and (n1202,n452,n460);
and (n1203,n498,n464);
nand (n1204,n1205,n1259,n1301);
nand (n1205,n1206,n1208);
xor (n1206,n1207,n1166);
xor (n1207,n1156,n1160);
xor (n1208,n1209,n1248);
xor (n1209,n1210,n1226);
nand (n1210,n1211,n1220,n1225);
nand (n1211,n1212,n1216);
xor (n1212,n1213,n462);
or (n1213,n1214,n1215);
and (n1214,n452,n599);
and (n1215,n498,n603);
xor (n1216,n1217,n601);
or (n1217,n1218,n1219);
and (n1218,n180,n822);
and (n1219,n365,n826);
nand (n1220,n1221,n1216);
xor (n1221,n1222,n380);
or (n1222,n1223,n1224);
and (n1223,n570,n460);
and (n1224,n791,n464);
nand (n1225,n1212,n1221);
nand (n1226,n1227,n1242,n1247);
nand (n1227,n1228,n1237);
xor (n1228,n1229,n1233);
xnor (n1229,n1230,n949);
nor (n1230,n1231,n1232);
and (n1231,n69,n1150);
and (n1232,n65,n1152);
xor (n1233,n1234,n824);
or (n1234,n1235,n1236);
and (n1235,n90,n947);
and (n1236,n148,n951);
and (n1237,n1238,n46);
xnor (n1238,n1239,n949);
nor (n1239,n1240,n1241);
and (n1240,n90,n1150);
and (n1241,n69,n1152);
nand (n1242,n1243,n1237);
xor (n1243,n1244,n20);
or (n1244,n1245,n1246);
and (n1245,n795,n378);
and (n1246,n797,n382);
nand (n1247,n1228,n1243);
xor (n1248,n1249,n1255);
xor (n1249,n1250,n1254);
xor (n1250,n1251,n20);
or (n1251,n1252,n1253);
and (n1252,n791,n378);
and (n1253,n795,n382);
and (n1254,n1229,n1233);
xor (n1255,n1256,n24);
or (n1256,n1257,n1258);
and (n1257,n797,n18);
and (n1258,n931,n22);
nand (n1259,n1260,n1208);
nand (n1260,n1261,n1285,n1300);
nand (n1261,n1262,n1283);
nand (n1262,n1263,n1277,n1282);
nand (n1263,n1264,n1273);
and (n1264,n1265,n1269);
xnor (n1265,n1266,n949);
nor (n1266,n1267,n1268);
and (n1267,n148,n1150);
and (n1268,n90,n1152);
xor (n1269,n1270,n824);
or (n1270,n1271,n1272);
and (n1271,n180,n947);
and (n1272,n365,n951);
xor (n1273,n1274,n20);
or (n1274,n1275,n1276);
and (n1275,n797,n378);
and (n1276,n931,n382);
nand (n1277,n1278,n1273);
xor (n1278,n1279,n24);
or (n1279,n1280,n1281);
and (n1280,n1135,n18);
and (n1281,n1139,n22);
nand (n1282,n1264,n1278);
xor (n1283,n1284,n1243);
xor (n1284,n1228,n1237);
nand (n1285,n1286,n1283);
xor (n1286,n1287,n1296);
xor (n1287,n1288,n1292);
xor (n1288,n1289,n24);
or (n1289,n1290,n1291);
and (n1290,n931,n18);
and (n1291,n1135,n22);
xor (n1292,n1293,n34);
or (n1293,n1294,n1295);
and (n1294,n1139,n28);
and (n1295,n1141,n32);
xor (n1296,n1297,n46);
or (n1297,n1298,n1299);
and (n1298,n1164,n40);
and (n1299,n1178,n44);
nand (n1300,n1262,n1286);
nand (n1301,n1206,n1260);
nand (n1302,n1303,n1204);
xor (n1303,n1304,n1343);
xor (n1304,n1305,n1309);
nand (n1305,n1306,n1307,n1308);
nand (n1306,n1210,n1226);
nand (n1307,n1248,n1226);
nand (n1308,n1210,n1248);
xor (n1309,n1310,n1332);
xor (n1310,n1311,n1328);
nand (n1311,n1312,n1322,n1327);
nand (n1312,n1313,n1317);
xor (n1313,n1314,n601);
or (n1314,n1315,n1316);
and (n1315,n148,n822);
and (n1316,n180,n826);
xor (n1317,n1318,n60);
xnor (n1318,n1319,n949);
nor (n1319,n1320,n1321);
and (n1320,n65,n1150);
and (n1321,n57,n1152);
nand (n1322,n1323,n1317);
xor (n1323,n1324,n380);
or (n1324,n1325,n1326);
and (n1325,n498,n460);
and (n1326,n570,n464);
nand (n1327,n1313,n1323);
nand (n1328,n1329,n1330,n1331);
nand (n1329,n1250,n1254);
nand (n1330,n1255,n1254);
nand (n1331,n1250,n1255);
xor (n1332,n1333,n1339);
xor (n1333,n1334,n1335);
and (n1334,n1318,n60);
xor (n1335,n1336,n20);
or (n1336,n1337,n1338);
and (n1337,n570,n378);
and (n1338,n791,n382);
xor (n1339,n1340,n24);
or (n1340,n1341,n1342);
and (n1341,n795,n18);
and (n1342,n797,n22);
nand (n1343,n1344,n1351,n1385);
nand (n1344,n1345,n1349);
nand (n1345,n1346,n1347,n1348);
nand (n1346,n1288,n1292);
nand (n1347,n1296,n1292);
nand (n1348,n1288,n1296);
xor (n1349,n1350,n1323);
xor (n1350,n1313,n1317);
nand (n1351,n1352,n1349);
nand (n1352,n1353,n1370,n1384);
nand (n1353,n1354,n1368);
nand (n1354,n1355,n1364,n1367);
nand (n1355,n1356,n1360);
xor (n1356,n1357,n824);
or (n1357,n1358,n1359);
and (n1358,n148,n947);
and (n1359,n180,n951);
xor (n1360,n1361,n462);
or (n1361,n1362,n1363);
and (n1362,n498,n599);
and (n1363,n570,n603);
nand (n1364,n1365,n1360);
xnor (n1365,n1366,n46);
nand (n1366,n1178,n40);
nand (n1367,n1356,n1365);
xor (n1368,n1369,n1221);
xor (n1369,n1212,n1216);
nand (n1370,n1371,n1368);
nand (n1371,n1372,n1378,n1383);
nand (n1372,n1373,n1377);
xor (n1373,n1374,n601);
or (n1374,n1375,n1376);
and (n1375,n365,n822);
and (n1376,n452,n826);
xor (n1377,n1238,n46);
nand (n1378,n1379,n1377);
xor (n1379,n1380,n380);
or (n1380,n1381,n1382);
and (n1381,n791,n460);
and (n1382,n795,n464);
nand (n1383,n1373,n1379);
nand (n1384,n1354,n1371);
nand (n1385,n1345,n1352);
nand (n1386,n1127,n1303);
xor (n1387,n1388,n1473);
xor (n1388,n1389,n1410);
xor (n1389,n1390,n1406);
xor (n1390,n1391,n1402);
xor (n1391,n1392,n1398);
xor (n1392,n1393,n1397);
xor (n1393,n1394,n46);
or (n1394,n1395,n1396);
and (n1395,n1135,n40);
and (n1396,n1139,n44);
and (n1397,n1143,n1147);
xor (n1398,n1399,n60);
or (n1399,n1400,n1401);
and (n1400,n1141,n54);
and (n1401,n1164,n58);
nand (n1402,n1403,n1404,n1405);
nand (n1403,n1182,n1186);
nand (n1404,n1190,n1186);
nand (n1405,n1182,n1190);
nand (n1406,n1407,n1408,n1409);
nand (n1407,n1311,n1328);
nand (n1408,n1332,n1328);
nand (n1409,n1311,n1332);
xor (n1410,n1411,n1469);
xor (n1411,n1412,n1436);
xor (n1412,n1413,n1432);
xor (n1413,n1414,n1418);
nand (n1414,n1415,n1416,n1417);
nand (n1415,n1334,n1335);
nand (n1416,n1339,n1335);
nand (n1417,n1334,n1339);
xor (n1418,n1419,n1428);
xor (n1419,n1420,n1424);
xnor (n1420,n1421,n949);
nor (n1421,n1422,n1423);
and (n1422,n53,n1150);
and (n1423,n43,n1152);
xor (n1424,n1425,n462);
or (n1425,n1426,n1427);
and (n1426,n148,n599);
and (n1427,n180,n603);
xor (n1428,n1429,n601);
or (n1429,n1430,n1431);
and (n1430,n69,n822);
and (n1431,n90,n826);
nand (n1432,n1433,n1434,n1435);
nand (n1433,n1192,n1196);
nand (n1434,n1200,n1196);
nand (n1435,n1192,n1200);
xor (n1436,n1437,n1455);
xor (n1437,n1438,n1442);
nand (n1438,n1439,n1440,n1441);
nand (n1439,n1131,n1136);
nand (n1440,n1142,n1136);
nand (n1441,n1131,n1142);
xor (n1442,n1443,n1453);
xor (n1443,n1444,n1448);
xor (n1444,n1445,n380);
or (n1445,n1446,n1447);
and (n1446,n365,n460);
and (n1447,n452,n464);
xor (n1448,n72,n1449);
xor (n1449,n1450,n824);
or (n1450,n1451,n1452);
and (n1451,n57,n947);
and (n1452,n65,n951);
xnor (n1453,n1454,n72);
nand (n1454,n1178,n66);
xor (n1455,n1456,n1465);
xor (n1456,n1457,n1461);
xor (n1457,n1458,n20);
or (n1458,n1459,n1460);
and (n1459,n498,n378);
and (n1460,n570,n382);
xor (n1461,n1462,n24);
or (n1462,n1463,n1464);
and (n1463,n791,n18);
and (n1464,n795,n22);
xor (n1465,n1466,n34);
or (n1466,n1467,n1468);
and (n1467,n797,n28);
and (n1468,n931,n32);
nand (n1469,n1470,n1471,n1472);
nand (n1470,n1129,n1154);
nand (n1471,n1180,n1154);
nand (n1472,n1129,n1180);
nand (n1473,n1474,n1475,n1476);
nand (n1474,n1305,n1309);
nand (n1475,n1343,n1309);
nand (n1476,n1305,n1343);
nor (n1477,n1478,n1482);
nand (n1478,n1479,n1480,n1481);
nand (n1479,n1389,n1410);
nand (n1480,n1473,n1410);
nand (n1481,n1389,n1473);
xor (n1482,n1483,n1492);
xor (n1483,n1484,n1488);
nand (n1484,n1485,n1486,n1487);
nand (n1485,n1391,n1402);
nand (n1486,n1406,n1402);
nand (n1487,n1391,n1406);
nand (n1488,n1489,n1490,n1491);
nand (n1489,n1412,n1436);
nand (n1490,n1469,n1436);
nand (n1491,n1412,n1469);
xor (n1492,n1493,n1554);
xor (n1493,n1494,n1525);
xor (n1494,n1495,n1514);
xor (n1495,n1496,n1510);
xor (n1496,n1497,n1506);
xor (n1497,n1498,n1502);
xor (n1498,n1499,n462);
or (n1499,n1500,n1501);
and (n1500,n90,n599);
and (n1501,n148,n603);
xor (n1502,n1503,n601);
or (n1503,n1504,n1505);
and (n1504,n65,n822);
and (n1505,n69,n826);
xor (n1506,n1507,n380);
or (n1507,n1508,n1509);
and (n1508,n180,n460);
and (n1509,n365,n464);
nand (n1510,n1511,n1512,n1513);
nand (n1511,n1444,n1448);
nand (n1512,n1453,n1448);
nand (n1513,n1444,n1453);
xor (n1514,n1515,n1521);
xor (n1515,n1516,n1520);
xor (n1516,n1517,n20);
or (n1517,n1518,n1519);
and (n1518,n452,n378);
and (n1519,n498,n382);
and (n1520,n72,n1449);
xor (n1521,n1522,n24);
or (n1522,n1523,n1524);
and (n1523,n570,n18);
and (n1524,n791,n22);
xor (n1525,n1526,n1550);
xor (n1526,n1527,n1531);
nand (n1527,n1528,n1529,n1530);
nand (n1528,n1457,n1461);
nand (n1529,n1465,n1461);
nand (n1530,n1457,n1465);
xor (n1531,n1532,n1541);
xor (n1532,n1533,n1537);
xor (n1533,n1534,n34);
or (n1534,n1535,n1536);
and (n1535,n795,n28);
and (n1536,n797,n32);
xor (n1537,n1538,n46);
or (n1538,n1539,n1540);
and (n1539,n931,n40);
and (n1540,n1135,n44);
xor (n1541,n1542,n1546);
xnor (n1542,n1543,n949);
nor (n1543,n1544,n1545);
and (n1544,n43,n1150);
and (n1545,n39,n1152);
xor (n1546,n1547,n824);
or (n1547,n1548,n1549);
and (n1548,n53,n947);
and (n1549,n57,n951);
nand (n1550,n1551,n1552,n1553);
nand (n1551,n1393,n1397);
nand (n1552,n1398,n1397);
nand (n1553,n1393,n1398);
xor (n1554,n1555,n1574);
xor (n1555,n1556,n1570);
xor (n1556,n1557,n1566);
xor (n1557,n1558,n1562);
xor (n1558,n1559,n60);
or (n1559,n1560,n1561);
and (n1560,n1139,n54);
and (n1561,n1141,n58);
xor (n1562,n1563,n72);
or (n1563,n1564,n1565);
and (n1564,n1164,n66);
and (n1565,n1178,n70);
nand (n1566,n1567,n1568,n1569);
nand (n1567,n1420,n1424);
nand (n1568,n1428,n1424);
nand (n1569,n1420,n1428);
nand (n1570,n1571,n1572,n1573);
nand (n1571,n1414,n1418);
nand (n1572,n1432,n1418);
nand (n1573,n1414,n1432);
nand (n1574,n1575,n1576,n1577);
nand (n1575,n1438,n1442);
nand (n1576,n1455,n1442);
nand (n1577,n1438,n1455);
nor (n1578,n1579,n1684);
nor (n1579,n1580,n1584);
nand (n1580,n1581,n1582,n1583);
nand (n1581,n1484,n1488);
nand (n1582,n1492,n1488);
nand (n1583,n1484,n1492);
xor (n1584,n1585,n1680);
xor (n1585,n1586,n1620);
xor (n1586,n1587,n1616);
xor (n1587,n1588,n1592);
nand (n1588,n1589,n1590,n1591);
nand (n1589,n1496,n1510);
nand (n1590,n1514,n1510);
nand (n1591,n1496,n1514);
xor (n1592,n1593,n1602);
xor (n1593,n1594,n1598);
xor (n1594,n1595,n72);
or (n1595,n1596,n1597);
and (n1596,n1141,n66);
and (n1597,n1164,n70);
nand (n1598,n1599,n1600,n1601);
nand (n1599,n1516,n1520);
nand (n1600,n1521,n1520);
nand (n1601,n1516,n1521);
xor (n1602,n1603,n1612);
xor (n1603,n1604,n1608);
xor (n1604,n1605,n462);
or (n1605,n1606,n1607);
and (n1606,n69,n599);
and (n1607,n90,n603);
xnor (n1608,n1609,n949);
nor (n1609,n1610,n1611);
and (n1610,n39,n1150);
and (n1611,n31,n1152);
xor (n1612,n1613,n601);
or (n1613,n1614,n1615);
and (n1614,n57,n822);
and (n1615,n65,n826);
nand (n1616,n1617,n1618,n1619);
nand (n1617,n1527,n1531);
nand (n1618,n1550,n1531);
nand (n1619,n1527,n1550);
xor (n1620,n1621,n1676);
xor (n1621,n1622,n1644);
xor (n1622,n1623,n1632);
xor (n1623,n1624,n1628);
nand (n1624,n1625,n1626,n1627);
nand (n1625,n1498,n1502);
nand (n1626,n1506,n1502);
nand (n1627,n1498,n1506);
nand (n1628,n1629,n1630,n1631);
nand (n1629,n1533,n1537);
nand (n1630,n1541,n1537);
nand (n1631,n1533,n1541);
xor (n1632,n1633,n1640);
xor (n1633,n1634,n1638);
xor (n1634,n1635,n380);
or (n1635,n1636,n1637);
and (n1636,n148,n460);
and (n1637,n180,n464);
xnor (n1638,n1639,n93);
nand (n1639,n1178,n87);
xor (n1640,n1641,n20);
or (n1641,n1642,n1643);
and (n1642,n365,n378);
and (n1643,n452,n382);
xor (n1644,n1645,n1664);
xor (n1645,n1646,n1650);
nand (n1646,n1647,n1648,n1649);
nand (n1647,n1558,n1562);
nand (n1648,n1566,n1562);
nand (n1649,n1558,n1566);
xor (n1650,n1651,n1660);
xor (n1651,n1652,n1656);
xor (n1652,n1653,n24);
or (n1653,n1654,n1655);
and (n1654,n498,n18);
and (n1655,n570,n22);
xor (n1656,n1657,n34);
or (n1657,n1658,n1659);
and (n1658,n791,n28);
and (n1659,n795,n32);
xor (n1660,n1661,n46);
or (n1661,n1662,n1663);
and (n1662,n797,n40);
and (n1663,n931,n44);
xor (n1664,n1665,n1672);
xor (n1665,n1666,n1671);
xor (n1666,n93,n1667);
xor (n1667,n1668,n824);
or (n1668,n1669,n1670);
and (n1669,n43,n947);
and (n1670,n53,n951);
and (n1671,n1542,n1546);
xor (n1672,n1673,n60);
or (n1673,n1674,n1675);
and (n1674,n1135,n54);
and (n1675,n1139,n58);
nand (n1676,n1677,n1678,n1679);
nand (n1677,n1556,n1570);
nand (n1678,n1574,n1570);
nand (n1679,n1556,n1574);
nand (n1680,n1681,n1682,n1683);
nand (n1681,n1494,n1525);
nand (n1682,n1554,n1525);
nand (n1683,n1494,n1554);
nor (n1684,n1685,n1689);
nand (n1685,n1686,n1687,n1688);
nand (n1686,n1586,n1620);
nand (n1687,n1680,n1620);
nand (n1688,n1586,n1680);
xor (n1689,n1690,n1699);
xor (n1690,n1691,n1695);
nand (n1691,n1692,n1693,n1694);
nand (n1692,n1588,n1592);
nand (n1693,n1616,n1592);
nand (n1694,n1588,n1616);
nand (n1695,n1696,n1697,n1698);
nand (n1696,n1622,n1644);
nand (n1697,n1676,n1644);
nand (n1698,n1622,n1676);
xor (n1699,n1700,n1761);
xor (n1700,n1701,n1725);
xor (n1701,n1702,n1721);
xor (n1702,n1703,n1707);
nand (n1703,n1704,n1705,n1706);
nand (n1704,n1652,n1656);
nand (n1705,n1660,n1656);
nand (n1706,n1652,n1660);
xor (n1707,n1708,n1717);
xor (n1708,n1709,n1713);
xor (n1709,n1710,n20);
or (n1710,n1711,n1712);
and (n1711,n180,n378);
and (n1712,n365,n382);
xor (n1713,n1714,n24);
or (n1714,n1715,n1716);
and (n1715,n452,n18);
and (n1716,n498,n22);
xor (n1717,n1718,n34);
or (n1718,n1719,n1720);
and (n1719,n570,n28);
and (n1720,n791,n32);
nand (n1721,n1722,n1723,n1724);
nand (n1722,n1666,n1671);
nand (n1723,n1672,n1671);
nand (n1724,n1666,n1672);
xor (n1725,n1726,n1747);
xor (n1726,n1727,n1743);
xor (n1727,n1728,n1742);
xor (n1728,n1729,n1733);
xor (n1729,n1730,n46);
or (n1730,n1731,n1732);
and (n1731,n795,n40);
and (n1732,n797,n44);
xor (n1733,n1734,n1738);
xnor (n1734,n1735,n949);
nor (n1735,n1736,n1737);
and (n1736,n31,n1150);
and (n1737,n17,n1152);
xor (n1738,n1739,n824);
or (n1739,n1740,n1741);
and (n1740,n39,n947);
and (n1741,n43,n951);
and (n1742,n93,n1667);
nand (n1743,n1744,n1745,n1746);
nand (n1744,n1594,n1598);
nand (n1745,n1602,n1598);
nand (n1746,n1594,n1602);
xor (n1747,n1748,n1757);
xor (n1748,n1749,n1753);
xor (n1749,n1750,n60);
or (n1750,n1751,n1752);
and (n1751,n931,n54);
and (n1752,n1135,n58);
xor (n1753,n1754,n93);
or (n1754,n1755,n1756);
and (n1755,n1164,n87);
and (n1756,n1178,n91);
xor (n1757,n1758,n72);
or (n1758,n1759,n1760);
and (n1759,n1139,n66);
and (n1760,n1141,n70);
xor (n1761,n1762,n1791);
xor (n1762,n1763,n1787);
xor (n1763,n1764,n1783);
xor (n1764,n1765,n1769);
nand (n1765,n1766,n1767,n1768);
nand (n1766,n1604,n1608);
nand (n1767,n1612,n1608);
nand (n1768,n1604,n1612);
xor (n1769,n1770,n1779);
xor (n1770,n1771,n1775);
xor (n1771,n1772,n462);
or (n1772,n1773,n1774);
and (n1773,n65,n599);
and (n1774,n69,n603);
xor (n1775,n1776,n601);
or (n1776,n1777,n1778);
and (n1777,n53,n822);
and (n1778,n57,n826);
xor (n1779,n1780,n380);
or (n1780,n1781,n1782);
and (n1781,n90,n460);
and (n1782,n148,n464);
nand (n1783,n1784,n1785,n1786);
nand (n1784,n1634,n1638);
nand (n1785,n1640,n1638);
nand (n1786,n1634,n1640);
nand (n1787,n1788,n1789,n1790);
nand (n1788,n1624,n1628);
nand (n1789,n1632,n1628);
nand (n1790,n1624,n1632);
nand (n1791,n1792,n1793,n1794);
nand (n1792,n1646,n1650);
nand (n1793,n1664,n1650);
nand (n1794,n1646,n1664);
nor (n1795,n1796,n2068);
nor (n1796,n1797,n2044);
nor (n1797,n1798,n2042);
nor (n1798,n1799,n2017);
nand (n1799,n1800,n1979);
nand (n1800,n1801,n1926,n1978);
nand (n1801,n1802,n1853);
xor (n1802,n1803,n1840);
xor (n1803,n1804,n1825);
nand (n1804,n1805,n1819,n1824);
nand (n1805,n1806,n1815);
and (n1806,n1807,n1811);
xnor (n1807,n1808,n949);
nor (n1808,n1809,n1810);
and (n1809,n365,n1150);
and (n1810,n180,n1152);
xor (n1811,n1812,n824);
or (n1812,n1813,n1814);
and (n1813,n452,n947);
and (n1814,n498,n951);
xor (n1815,n1816,n20);
or (n1816,n1817,n1818);
and (n1817,n1135,n378);
and (n1818,n1139,n382);
nand (n1819,n1820,n1815);
xor (n1820,n1821,n24);
or (n1821,n1822,n1823);
and (n1822,n1141,n18);
and (n1823,n1164,n22);
nand (n1824,n1806,n1820);
xor (n1825,n1826,n1835);
xor (n1826,n1827,n1831);
xor (n1827,n1828,n462);
or (n1828,n1829,n1830);
and (n1829,n570,n599);
and (n1830,n791,n603);
xor (n1831,n1832,n601);
or (n1832,n1833,n1834);
and (n1833,n452,n822);
and (n1834,n498,n826);
and (n1835,n1836,n34);
xnor (n1836,n1837,n949);
nor (n1837,n1838,n1839);
and (n1838,n180,n1150);
and (n1839,n148,n1152);
nand (n1840,n1841,n1847,n1852);
nand (n1841,n1842,n1846);
xor (n1842,n1843,n601);
or (n1843,n1844,n1845);
and (n1844,n498,n822);
and (n1845,n570,n826);
xor (n1846,n1836,n34);
nand (n1847,n1848,n1846);
xor (n1848,n1849,n380);
or (n1849,n1850,n1851);
and (n1850,n797,n460);
and (n1851,n931,n464);
nand (n1852,n1842,n1848);
xor (n1853,n1854,n1890);
xor (n1854,n1855,n1866);
xor (n1855,n1856,n1862);
xor (n1856,n1857,n1861);
xor (n1857,n1858,n380);
or (n1858,n1859,n1860);
and (n1859,n795,n460);
and (n1860,n797,n464);
xor (n1861,n1265,n1269);
xor (n1862,n1863,n20);
or (n1863,n1864,n1865);
and (n1864,n931,n378);
and (n1865,n1135,n382);
xor (n1866,n1867,n1876);
xor (n1867,n1868,n1872);
xor (n1868,n1869,n24);
or (n1869,n1870,n1871);
and (n1870,n1139,n18);
and (n1871,n1141,n22);
xor (n1872,n1873,n34);
or (n1873,n1874,n1875);
and (n1874,n1164,n28);
and (n1875,n1178,n32);
nand (n1876,n1877,n1884,n1889);
nand (n1877,n1878,n1882);
xor (n1878,n1879,n824);
or (n1879,n1880,n1881);
and (n1880,n365,n947);
and (n1881,n452,n951);
xnor (n1882,n1883,n34);
nand (n1883,n1178,n28);
nand (n1884,n1885,n1882);
xor (n1885,n1886,n462);
or (n1886,n1887,n1888);
and (n1887,n791,n599);
and (n1888,n795,n603);
nand (n1889,n1878,n1885);
nand (n1890,n1891,n1911,n1925);
nand (n1891,n1892,n1894);
xor (n1892,n1893,n1885);
xor (n1893,n1878,n1882);
nand (n1894,n1895,n1904,n1910);
nand (n1895,n1896,n1900);
xor (n1896,n1897,n462);
or (n1897,n1898,n1899);
and (n1898,n795,n599);
and (n1899,n797,n603);
xor (n1900,n1901,n601);
or (n1901,n1902,n1903);
and (n1902,n570,n822);
and (n1903,n791,n826);
nand (n1904,n1905,n1900);
and (n1905,n1906,n24);
xnor (n1906,n1907,n949);
nor (n1907,n1908,n1909);
and (n1908,n452,n1150);
and (n1909,n365,n1152);
nand (n1910,n1896,n1905);
nand (n1911,n1912,n1894);
nand (n1912,n1913,n1919,n1924);
nand (n1913,n1914,n1918);
xor (n1914,n1915,n380);
or (n1915,n1916,n1917);
and (n1916,n931,n460);
and (n1917,n1135,n464);
xor (n1918,n1807,n1811);
nand (n1919,n1920,n1918);
xor (n1920,n1921,n20);
or (n1921,n1922,n1923);
and (n1922,n1139,n378);
and (n1923,n1141,n382);
nand (n1924,n1914,n1920);
nand (n1925,n1892,n1912);
nand (n1926,n1927,n1853);
nand (n1927,n1928,n1933,n1977);
nand (n1928,n1929,n1931);
xor (n1929,n1930,n1820);
xor (n1930,n1806,n1815);
xor (n1931,n1932,n1848);
xor (n1932,n1842,n1846);
nand (n1933,n1934,n1931);
nand (n1934,n1935,n1954,n1976);
nand (n1935,n1936,n1940);
xor (n1936,n1937,n24);
or (n1937,n1938,n1939);
and (n1938,n1164,n18);
and (n1939,n1178,n22);
nand (n1940,n1941,n1948,n1953);
nand (n1941,n1942,n1946);
xor (n1942,n1943,n824);
or (n1943,n1944,n1945);
and (n1944,n498,n947);
and (n1945,n570,n951);
xnor (n1946,n1947,n24);
nand (n1947,n1178,n18);
nand (n1948,n1949,n1946);
xor (n1949,n1950,n462);
or (n1950,n1951,n1952);
and (n1951,n797,n599);
and (n1952,n931,n603);
nand (n1953,n1942,n1949);
nand (n1954,n1955,n1940);
nand (n1955,n1956,n1970,n1975);
nand (n1956,n1957,n1961);
xor (n1957,n1958,n601);
or (n1958,n1959,n1960);
and (n1959,n791,n822);
and (n1960,n795,n826);
and (n1961,n1962,n1966);
xnor (n1962,n1963,n949);
nor (n1963,n1964,n1965);
and (n1964,n498,n1150);
and (n1965,n452,n1152);
xor (n1966,n1967,n824);
or (n1967,n1968,n1969);
and (n1968,n570,n947);
and (n1969,n791,n951);
nand (n1970,n1971,n1961);
xor (n1971,n1972,n380);
or (n1972,n1973,n1974);
and (n1973,n1135,n460);
and (n1974,n1139,n464);
nand (n1975,n1957,n1971);
nand (n1976,n1936,n1955);
nand (n1977,n1929,n1934);
nand (n1978,n1802,n1927);
xor (n1979,n1980,n1995);
xor (n1980,n1981,n1991);
xor (n1981,n1982,n1989);
xor (n1982,n1983,n1987);
nand (n1983,n1984,n1985,n1986);
nand (n1984,n1827,n1831);
nand (n1985,n1835,n1831);
nand (n1986,n1827,n1835);
xor (n1987,n1988,n1278);
xor (n1988,n1264,n1273);
xor (n1989,n1990,n1379);
xor (n1990,n1373,n1377);
nand (n1991,n1992,n1993,n1994);
nand (n1992,n1855,n1866);
nand (n1993,n1890,n1866);
nand (n1994,n1855,n1890);
xor (n1995,n1996,n2005);
xor (n1996,n1997,n2001);
nand (n1997,n1998,n1999,n2000);
nand (n1998,n1868,n1872);
nand (n1999,n1876,n1872);
nand (n2000,n1868,n1876);
nand (n2001,n2002,n2003,n2004);
nand (n2002,n1804,n1825);
nand (n2003,n1840,n1825);
nand (n2004,n1804,n1840);
xor (n2005,n2006,n2015);
xor (n2006,n2007,n2011);
xor (n2007,n2008,n34);
or (n2008,n2009,n2010);
and (n2009,n1141,n28);
and (n2010,n1164,n32);
nand (n2011,n2012,n2013,n2014);
nand (n2012,n1857,n1861);
nand (n2013,n1862,n1861);
nand (n2014,n1857,n1862);
xor (n2015,n2016,n1365);
xor (n2016,n1356,n1360);
nor (n2017,n2018,n2022);
nand (n2018,n2019,n2020,n2021);
nand (n2019,n1981,n1991);
nand (n2020,n1995,n1991);
nand (n2021,n1981,n1995);
xor (n2022,n2023,n2030);
xor (n2023,n2024,n2026);
xor (n2024,n2025,n1286);
xor (n2025,n1262,n1283);
nand (n2026,n2027,n2028,n2029);
nand (n2027,n1997,n2001);
nand (n2028,n2005,n2001);
nand (n2029,n1997,n2005);
xor (n2030,n2031,n2040);
xor (n2031,n2032,n2036);
nand (n2032,n2033,n2034,n2035);
nand (n2033,n2007,n2011);
nand (n2034,n2015,n2011);
nand (n2035,n2007,n2015);
nand (n2036,n2037,n2038,n2039);
nand (n2037,n1983,n1987);
nand (n2038,n1989,n1987);
nand (n2039,n1983,n1989);
xor (n2040,n2041,n1371);
xor (n2041,n1354,n1368);
not (n2042,n2043);
nand (n2043,n2018,n2022);
not (n2044,n2045);
nor (n2045,n2046,n2061);
nor (n2046,n2047,n2051);
nand (n2047,n2048,n2049,n2050);
nand (n2048,n2024,n2026);
nand (n2049,n2030,n2026);
nand (n2050,n2024,n2030);
xor (n2051,n2052,n2059);
xor (n2052,n2053,n2055);
xor (n2053,n2054,n1352);
xor (n2054,n1345,n1349);
nand (n2055,n2056,n2057,n2058);
nand (n2056,n2032,n2036);
nand (n2057,n2040,n2036);
nand (n2058,n2032,n2040);
xor (n2059,n2060,n1260);
xor (n2060,n1206,n1208);
nor (n2061,n2062,n2066);
nand (n2062,n2063,n2064,n2065);
nand (n2063,n2053,n2055);
nand (n2064,n2059,n2055);
nand (n2065,n2053,n2059);
xor (n2066,n2067,n1303);
xor (n2067,n1127,n1204);
not (n2068,n2069);
nor (n2069,n2070,n2072);
nor (n2070,n2071,n2061);
nand (n2071,n2047,n2051);
not (n2072,n2073);
nand (n2073,n2062,n2066);
not (n2074,n2075);
nor (n2075,n2076,n2083);
nor (n2076,n2077,n2082);
nor (n2077,n2078,n2080);
nor (n2078,n2079,n1477);
nand (n2079,n1125,n1387);
not (n2080,n2081);
nand (n2081,n1478,n1482);
not (n2082,n1578);
not (n2083,n2084);
nor (n2084,n2085,n2087);
nor (n2085,n2086,n1684);
nand (n2086,n1580,n1584);
not (n2087,n2088);
nand (n2088,n1685,n1689);
not (n2089,n2090);
nor (n2090,n2091,n2506);
nand (n2091,n2092,n2319);
nor (n2092,n2093,n2205);
nor (n2093,n2094,n2098);
nand (n2094,n2095,n2096,n2097);
nand (n2095,n1691,n1695);
nand (n2096,n1699,n1695);
nand (n2097,n1691,n1699);
xor (n2098,n2099,n2201);
xor (n2099,n2100,n2133);
xor (n2100,n2101,n2129);
xor (n2101,n2102,n2125);
xor (n2102,n2103,n2121);
xor (n2103,n2104,n2117);
xor (n2104,n2105,n2114);
xor (n2105,n2106,n2110);
xor (n2106,n2107,n824);
or (n2107,n2108,n2109);
and (n2108,n31,n947);
and (n2109,n39,n951);
xor (n2110,n2111,n601);
or (n2111,n2112,n2113);
and (n2112,n43,n822);
and (n2113,n53,n826);
xnor (n2114,n2115,n949);
nor (n2115,n2116,n1737);
and (n2116,n17,n1150);
nand (n2117,n2118,n2119,n2120);
nand (n2118,n1709,n1713);
nand (n2119,n1717,n1713);
nand (n2120,n1709,n1717);
nand (n2121,n2122,n2123,n2124);
nand (n2122,n1729,n1733);
nand (n2123,n1742,n1733);
nand (n2124,n1729,n1742);
nand (n2125,n2126,n2127,n2128);
nand (n2126,n1703,n1707);
nand (n2127,n1721,n1707);
nand (n2128,n1703,n1721);
nand (n2129,n2130,n2131,n2132);
nand (n2130,n1727,n1743);
nand (n2131,n1747,n1743);
nand (n2132,n1727,n1747);
xor (n2133,n2134,n2197);
xor (n2134,n2135,n2173);
xor (n2135,n2136,n2158);
xor (n2136,n2137,n2151);
xor (n2137,n2138,n2147);
xor (n2138,n2139,n2143);
xor (n2139,n2140,n380);
or (n2140,n2141,n2142);
and (n2141,n69,n460);
and (n2142,n90,n464);
xor (n2143,n2144,n20);
or (n2144,n2145,n2146);
and (n2145,n148,n378);
and (n2146,n180,n382);
xor (n2147,n2148,n24);
or (n2148,n2149,n2150);
and (n2149,n365,n18);
and (n2150,n452,n22);
xor (n2151,n2152,n2154);
xor (n2152,n93,n2153);
and (n2153,n1734,n1738);
xor (n2154,n2155,n60);
or (n2155,n2156,n2157);
and (n2156,n797,n54);
and (n2157,n931,n58);
xor (n2158,n2159,n2168);
xor (n2159,n2160,n2164);
xor (n2160,n2161,n34);
or (n2161,n2162,n2163);
and (n2162,n498,n28);
and (n2163,n570,n32);
xor (n2164,n2165,n46);
or (n2165,n2166,n2167);
and (n2166,n791,n40);
and (n2167,n795,n44);
xor (n2168,n93,n2169);
xor (n2169,n2170,n462);
or (n2170,n2171,n2172);
and (n2171,n57,n599);
and (n2172,n65,n603);
xor (n2173,n2174,n2183);
xor (n2174,n2175,n2179);
nand (n2175,n2176,n2177,n2178);
nand (n2176,n1749,n1753);
nand (n2177,n1757,n1753);
nand (n2178,n1749,n1757);
nand (n2179,n2180,n2181,n2182);
nand (n2180,n1765,n1769);
nand (n2181,n1783,n1769);
nand (n2182,n1765,n1783);
xor (n2183,n2184,n2193);
xor (n2184,n2185,n2189);
xor (n2185,n2186,n72);
or (n2186,n2187,n2188);
and (n2187,n1135,n66);
and (n2188,n1139,n70);
xor (n2189,n2190,n93);
or (n2190,n2191,n2192);
and (n2191,n1141,n87);
and (n2192,n1164,n91);
nand (n2193,n2194,n2195,n2196);
nand (n2194,n1771,n1775);
nand (n2195,n1779,n1775);
nand (n2196,n1771,n1779);
nand (n2197,n2198,n2199,n2200);
nand (n2198,n1763,n1787);
nand (n2199,n1791,n1787);
nand (n2200,n1763,n1791);
nand (n2201,n2202,n2203,n2204);
nand (n2202,n1701,n1725);
nand (n2203,n1761,n1725);
nand (n2204,n1701,n1761);
nor (n2205,n2206,n2210);
nand (n2206,n2207,n2208,n2209);
nand (n2207,n2100,n2133);
nand (n2208,n2201,n2133);
nand (n2209,n2100,n2201);
xor (n2210,n2211,n2220);
xor (n2211,n2212,n2216);
nand (n2212,n2213,n2214,n2215);
nand (n2213,n2102,n2125);
nand (n2214,n2129,n2125);
nand (n2215,n2102,n2129);
nand (n2216,n2217,n2218,n2219);
nand (n2217,n2135,n2173);
nand (n2218,n2197,n2173);
nand (n2219,n2135,n2197);
xor (n2220,n2221,n2278);
xor (n2221,n2222,n2253);
xor (n2222,n2223,n2239);
xor (n2223,n2224,n2228);
nand (n2224,n2225,n2226,n2227);
nand (n2225,n93,n2153);
nand (n2226,n2154,n2153);
nand (n2227,n93,n2154);
xor (n2228,n2229,n2235);
xor (n2229,n2230,n2234);
xor (n2230,n2231,n46);
or (n2231,n2232,n2233);
and (n2232,n570,n40);
and (n2233,n791,n44);
and (n2234,n93,n2169);
xor (n2235,n2236,n60);
or (n2236,n2237,n2238);
and (n2237,n795,n54);
and (n2238,n797,n58);
xor (n2239,n2240,n2249);
xor (n2240,n2241,n2245);
xor (n2241,n2242,n72);
or (n2242,n2243,n2244);
and (n2243,n931,n66);
and (n2244,n1135,n70);
xor (n2245,n2246,n93);
or (n2246,n2247,n2248);
and (n2247,n1139,n87);
and (n2248,n1141,n91);
nand (n2249,n2250,n2251,n2252);
nand (n2250,n2106,n2110);
nand (n2251,n2114,n2110);
nand (n2252,n2106,n2114);
xor (n2253,n2254,n2263);
xor (n2254,n2255,n2259);
nand (n2255,n2256,n2257,n2258);
nand (n2256,n2185,n2189);
nand (n2257,n2193,n2189);
nand (n2258,n2185,n2193);
nand (n2259,n2260,n2261,n2262);
nand (n2260,n2104,n2117);
nand (n2261,n2121,n2117);
nand (n2262,n2104,n2121);
xor (n2263,n2264,n93);
xor (n2264,n2265,n2269);
nand (n2265,n2266,n2267,n2268);
nand (n2266,n2139,n2143);
nand (n2267,n2147,n2143);
nand (n2268,n2139,n2147);
xor (n2269,n2270,n2275);
not (n2270,n2271);
xor (n2271,n2272,n462);
or (n2272,n2273,n2274);
and (n2273,n53,n599);
and (n2274,n57,n603);
xor (n2275,n2276,n824);
or (n2276,n946,n2277);
and (n2277,n31,n951);
xor (n2278,n2279,n2315);
xor (n2279,n2280,n2284);
nand (n2280,n2281,n2282,n2283);
nand (n2281,n2137,n2151);
nand (n2282,n2158,n2151);
nand (n2283,n2137,n2158);
xor (n2284,n2285,n2304);
xor (n2285,n2286,n2290);
nand (n2286,n2287,n2288,n2289);
nand (n2287,n2160,n2164);
nand (n2288,n2168,n2164);
nand (n2289,n2160,n2168);
xor (n2290,n2291,n2300);
xor (n2291,n2292,n2296);
xor (n2292,n2293,n20);
or (n2293,n2294,n2295);
and (n2294,n90,n378);
and (n2295,n148,n382);
xor (n2296,n2297,n24);
or (n2297,n2298,n2299);
and (n2298,n180,n18);
and (n2299,n365,n22);
xor (n2300,n2301,n34);
or (n2301,n2302,n2303);
and (n2302,n452,n28);
and (n2303,n498,n32);
xor (n2304,n2305,n2311);
xor (n2305,n2306,n2310);
xor (n2306,n2307,n601);
or (n2307,n2308,n2309);
and (n2308,n39,n822);
and (n2309,n43,n826);
not (n2310,n2114);
xor (n2311,n2312,n380);
or (n2312,n2313,n2314);
and (n2313,n65,n460);
and (n2314,n69,n464);
nand (n2315,n2316,n2317,n2318);
nand (n2316,n2175,n2179);
nand (n2317,n2183,n2179);
nand (n2318,n2175,n2183);
nor (n2319,n2320,n2427);
nor (n2320,n2321,n2325);
nand (n2321,n2322,n2323,n2324);
nand (n2322,n2212,n2216);
nand (n2323,n2220,n2216);
nand (n2324,n2212,n2220);
xor (n2325,n2326,n2423);
xor (n2326,n2327,n2367);
xor (n2327,n2328,n2363);
xor (n2328,n2329,n2359);
xor (n2329,n2330,n2355);
xor (n2330,n2331,n2345);
xor (n2331,n2332,n2341);
xor (n2332,n2333,n2337);
xor (n2333,n2334,n20);
or (n2334,n2335,n2336);
and (n2335,n69,n378);
and (n2336,n90,n382);
xor (n2337,n2338,n24);
or (n2338,n2339,n2340);
and (n2339,n148,n18);
and (n2340,n180,n22);
xor (n2341,n2342,n46);
or (n2342,n2343,n2344);
and (n2343,n498,n40);
and (n2344,n570,n44);
xor (n2345,n2346,n2351);
xor (n2346,n2347,n944);
xor (n2347,n2348,n462);
or (n2348,n2349,n2350);
and (n2349,n43,n599);
and (n2350,n53,n603);
xor (n2351,n2352,n380);
or (n2352,n2353,n2354);
and (n2353,n57,n460);
and (n2354,n65,n464);
nand (n2355,n2356,n2357,n2358);
nand (n2356,n2230,n2234);
nand (n2357,n2235,n2234);
nand (n2358,n2230,n2235);
nand (n2359,n2360,n2361,n2362);
nand (n2360,n2224,n2228);
nand (n2361,n2239,n2228);
nand (n2362,n2224,n2239);
nand (n2363,n2364,n2365,n2366);
nand (n2364,n2255,n2259);
nand (n2365,n2263,n2259);
nand (n2366,n2255,n2263);
xor (n2367,n2368,n2419);
xor (n2368,n2369,n2390);
xor (n2369,n2370,n2386);
xor (n2370,n2371,n2382);
xor (n2371,n2372,n2378);
xor (n2372,n2373,n2374);
not (n2373,n985);
xor (n2374,n2375,n34);
or (n2375,n2376,n2377);
and (n2376,n365,n28);
and (n2377,n452,n32);
xor (n2378,n2379,n60);
or (n2379,n2380,n2381);
and (n2380,n791,n54);
and (n2381,n795,n58);
nand (n2382,n2383,n2384,n2385);
nand (n2383,n2241,n2245);
nand (n2384,n2249,n2245);
nand (n2385,n2241,n2249);
nand (n2386,n2387,n2388,n2389);
nand (n2387,n2265,n2269);
nand (n2388,n93,n2269);
nand (n2389,n2265,n93);
xor (n2390,n2391,n2415);
xor (n2391,n2392,n2405);
xor (n2392,n2393,n2402);
xor (n2393,n2394,n2398);
xor (n2394,n2395,n72);
or (n2395,n2396,n2397);
and (n2396,n797,n66);
and (n2397,n931,n70);
xor (n2398,n2399,n93);
or (n2399,n2400,n2401);
and (n2400,n1135,n87);
and (n2401,n1139,n91);
nand (n2402,n2270,n2403,n2404);
nand (n2403,n2275,n2271);
not (n2404,n2275);
xor (n2405,n2406,n2411);
xor (n2406,n93,n2407);
nand (n2407,n2408,n2409,n2410);
nand (n2408,n2306,n2310);
nand (n2409,n2311,n2310);
nand (n2410,n2306,n2311);
nand (n2411,n2412,n2413,n2414);
nand (n2412,n2292,n2296);
nand (n2413,n2300,n2296);
nand (n2414,n2292,n2300);
nand (n2415,n2416,n2417,n2418);
nand (n2416,n2286,n2290);
nand (n2417,n2304,n2290);
nand (n2418,n2286,n2304);
nand (n2419,n2420,n2421,n2422);
nand (n2420,n2280,n2284);
nand (n2421,n2315,n2284);
nand (n2422,n2280,n2315);
nand (n2423,n2424,n2425,n2426);
nand (n2424,n2222,n2253);
nand (n2425,n2278,n2253);
nand (n2426,n2222,n2278);
nor (n2427,n2428,n2432);
nand (n2428,n2429,n2430,n2431);
nand (n2429,n2327,n2367);
nand (n2430,n2423,n2367);
nand (n2431,n2327,n2423);
xor (n2432,n2433,n2442);
xor (n2433,n2434,n2438);
nand (n2434,n2435,n2436,n2437);
nand (n2435,n2329,n2359);
nand (n2436,n2363,n2359);
nand (n2437,n2329,n2363);
nand (n2438,n2439,n2440,n2441);
nand (n2439,n2369,n2390);
nand (n2440,n2419,n2390);
nand (n2441,n2369,n2419);
xor (n2442,n2443,n2474);
xor (n2443,n2444,n2448);
nand (n2444,n2445,n2446,n2447);
nand (n2445,n2392,n2405);
nand (n2446,n2415,n2405);
nand (n2447,n2392,n2415);
xor (n2448,n2449,n2462);
xor (n2449,n2450,n2454);
nand (n2450,n2451,n2452,n2453);
nand (n2451,n93,n2407);
nand (n2452,n2411,n2407);
nand (n2453,n93,n2411);
xor (n2454,n2455,n2458);
xor (n2455,n2456,n93);
xor (n2456,n2457,n943);
xor (n2457,n935,n938);
nand (n2458,n2459,n2460,n2461);
nand (n2459,n2347,n944);
nand (n2460,n2351,n944);
nand (n2461,n2347,n2351);
xor (n2462,n2463,n2470);
xor (n2463,n2464,n2466);
xor (n2464,n2465,n971);
xor (n2465,n962,n966);
nand (n2466,n2467,n2468,n2469);
nand (n2467,n2333,n2337);
nand (n2468,n2341,n2337);
nand (n2469,n2333,n2341);
nand (n2470,n2471,n2472,n2473);
nand (n2471,n2394,n2398);
nand (n2472,n2402,n2398);
nand (n2473,n2394,n2402);
xor (n2474,n2475,n2484);
xor (n2475,n2476,n2480);
nand (n2476,n2477,n2478,n2479);
nand (n2477,n2331,n2345);
nand (n2478,n2355,n2345);
nand (n2479,n2331,n2355);
nand (n2480,n2481,n2482,n2483);
nand (n2481,n2371,n2382);
nand (n2482,n2386,n2382);
nand (n2483,n2371,n2386);
xor (n2484,n2485,n2492);
xor (n2485,n2486,n2490);
nand (n2486,n2487,n2488,n2489);
nand (n2487,n2373,n2374);
nand (n2488,n2378,n2374);
nand (n2489,n2373,n2378);
xor (n2490,n2491,n990);
xor (n2491,n981,n985);
xor (n2492,n2493,n2502);
xor (n2493,n2494,n2498);
xor (n2494,n2495,n60);
or (n2495,n2496,n2497);
and (n2496,n570,n54);
and (n2497,n791,n58);
xor (n2498,n2499,n72);
or (n2499,n2500,n2501);
and (n2500,n795,n66);
and (n2501,n797,n70);
xor (n2502,n2503,n93);
or (n2503,n2504,n2505);
and (n2504,n931,n87);
and (n2505,n1135,n91);
nand (n2506,n2507,n2591);
nor (n2507,n2508,n2558);
nor (n2508,n2509,n2513);
nand (n2509,n2510,n2511,n2512);
nand (n2510,n2434,n2438);
nand (n2511,n2442,n2438);
nand (n2512,n2434,n2442);
xor (n2513,n2514,n2554);
xor (n2514,n2515,n2535);
xor (n2515,n2516,n2523);
xor (n2516,n2517,n2519);
xor (n2517,n2518,n979);
xor (n2518,n960,n976);
nand (n2519,n2520,n2521,n2522);
nand (n2520,n2486,n2490);
nand (n2521,n2492,n2490);
nand (n2522,n2486,n2492);
xor (n2523,n2524,n2531);
xor (n2524,n2525,n2529);
nand (n2525,n2526,n2527,n2528);
nand (n2526,n2494,n2498);
nand (n2527,n2502,n2498);
nand (n2528,n2494,n2502);
xor (n2529,n2530,n889);
xor (n2530,n883,n887);
nand (n2531,n2532,n2533,n2534);
nand (n2532,n2456,n93);
nand (n2533,n2458,n93);
nand (n2534,n2456,n2458);
xor (n2535,n2536,n2550);
xor (n2536,n2537,n2541);
nand (n2537,n2538,n2539,n2540);
nand (n2538,n2450,n2454);
nand (n2539,n2462,n2454);
nand (n2540,n2450,n2462);
xor (n2541,n2542,n2546);
xor (n2542,n2543,n2545);
xor (n2543,n2544,n905);
xor (n2544,n896,n900);
xor (n2545,n928,n933);
nand (n2546,n2547,n2548,n2549);
nand (n2547,n2464,n2466);
nand (n2548,n2470,n2466);
nand (n2549,n2464,n2470);
nand (n2550,n2551,n2552,n2553);
nand (n2551,n2476,n2480);
nand (n2552,n2484,n2480);
nand (n2553,n2476,n2484);
nand (n2554,n2555,n2556,n2557);
nand (n2555,n2444,n2448);
nand (n2556,n2474,n2448);
nand (n2557,n2444,n2474);
nor (n2558,n2559,n2563);
nand (n2559,n2560,n2561,n2562);
nand (n2560,n2515,n2535);
nand (n2561,n2554,n2535);
nand (n2562,n2515,n2554);
xor (n2563,n2564,n2587);
xor (n2564,n2565,n2575);
xor (n2565,n2566,n2573);
xor (n2566,n2567,n2569);
xor (n2567,n2568,n876);
xor (n2568,n861,n873);
nand (n2569,n2570,n2571,n2572);
nand (n2570,n2525,n2529);
nand (n2571,n2531,n2529);
nand (n2572,n2525,n2531);
xor (n2573,n2574,n911);
xor (n2574,n881,n894);
xor (n2575,n2576,n2583);
xor (n2576,n2577,n2579);
xor (n2577,n2578,n958);
xor (n2578,n925,n955);
nand (n2579,n2580,n2581,n2582);
nand (n2580,n2543,n2545);
nand (n2581,n2546,n2545);
nand (n2582,n2543,n2546);
nand (n2583,n2584,n2585,n2586);
nand (n2584,n2517,n2519);
nand (n2585,n2523,n2519);
nand (n2586,n2517,n2523);
nand (n2587,n2588,n2589,n2590);
nand (n2588,n2537,n2541);
nand (n2589,n2550,n2541);
nand (n2590,n2537,n2550);
nor (n2591,n2592,n2609);
nor (n2592,n2593,n2597);
nand (n2593,n2594,n2595,n2596);
nand (n2594,n2565,n2575);
nand (n2595,n2587,n2575);
nand (n2596,n2565,n2587);
xor (n2597,n2598,n2605);
xor (n2598,n2599,n2603);
nand (n2599,n2600,n2601,n2602);
nand (n2600,n2567,n2569);
nand (n2601,n2573,n2569);
nand (n2602,n2567,n2573);
xor (n2603,n2604,n998);
xor (n2604,n921,n923);
nand (n2605,n2606,n2607,n2608);
nand (n2606,n2577,n2579);
nand (n2607,n2583,n2579);
nand (n2608,n2577,n2583);
nor (n2609,n2610,n2614);
nand (n2610,n2611,n2612,n2613);
nand (n2611,n2599,n2603);
nand (n2612,n2605,n2603);
nand (n2613,n2599,n2605);
xor (n2614,n2615,n919);
xor (n2615,n697,n781);
not (n2616,n2617);
nor (n2617,n2618,n2633);
nor (n2618,n2506,n2619);
nor (n2619,n2620,n2627);
nor (n2620,n2621,n2626);
nor (n2621,n2622,n2624);
nor (n2622,n2623,n2205);
nand (n2623,n2094,n2098);
not (n2624,n2625);
nand (n2625,n2206,n2210);
not (n2626,n2319);
not (n2627,n2628);
nor (n2628,n2629,n2631);
nor (n2629,n2630,n2427);
nand (n2630,n2321,n2325);
not (n2631,n2632);
nand (n2632,n2428,n2432);
not (n2633,n2634);
nor (n2634,n2635,n2642);
nor (n2635,n2636,n2641);
nor (n2636,n2637,n2639);
nor (n2637,n2638,n2558);
nand (n2638,n2509,n2513);
not (n2639,n2640);
nand (n2640,n2559,n2563);
not (n2641,n2591);
not (n2642,n2643);
nor (n2643,n2644,n2646);
nor (n2644,n2645,n2609);
nand (n2645,n2593,n2597);
not (n2646,n2647);
nand (n2647,n2610,n2614);
nand (n2648,n2649,n3068);
nand (n2649,n2650,n2961);
nor (n2650,n2651,n2946);
nor (n2651,n2652,n2817);
nand (n2652,n2653,n2794);
nor (n2653,n2654,n2771);
nor (n2654,n2655,n2744);
nand (n2655,n2656,n2701,n2743);
nand (n2656,n2657,n2669);
xor (n2657,n2658,n2664);
xor (n2658,n2659,n2660);
xor (n2659,n1962,n1966);
xor (n2660,n2661,n20);
or (n2661,n2662,n2663);
and (n2662,n1164,n378);
and (n2663,n1178,n382);
and (n2664,n20,n2665);
xor (n2665,n2666,n824);
or (n2666,n2667,n2668);
and (n2667,n791,n947);
and (n2668,n795,n951);
nand (n2669,n2670,n2687,n2700);
nand (n2670,n2671,n2672);
xor (n2671,n20,n2665);
nand (n2672,n2673,n2682,n2686);
nand (n2673,n2674,n2678);
xor (n2674,n2675,n462);
or (n2675,n2676,n2677);
and (n2676,n1139,n599);
and (n2677,n1141,n603);
xor (n2678,n2679,n601);
or (n2679,n2680,n2681);
and (n2680,n931,n822);
and (n2681,n1135,n826);
nand (n2682,n2683,n2678);
and (n2683,n380,n2684);
xnor (n2684,n2685,n380);
nand (n2685,n1178,n460);
nand (n2686,n2674,n2683);
nand (n2687,n2688,n2672);
xor (n2688,n2689,n2696);
xor (n2689,n2690,n2694);
xnor (n2690,n2691,n949);
nor (n2691,n2692,n2693);
and (n2692,n570,n1150);
and (n2693,n498,n1152);
xnor (n2694,n2695,n20);
nand (n2695,n1178,n378);
xor (n2696,n2697,n462);
or (n2697,n2698,n2699);
and (n2698,n1135,n599);
and (n2699,n1139,n603);
nand (n2700,n2671,n2688);
nand (n2701,n2702,n2669);
xor (n2702,n2703,n2722);
xor (n2703,n2704,n2708);
nand (n2704,n2705,n2706,n2707);
nand (n2705,n2690,n2694);
nand (n2706,n2696,n2694);
nand (n2707,n2690,n2696);
xor (n2708,n2709,n2718);
xor (n2709,n2710,n2714);
xor (n2710,n2711,n462);
or (n2711,n2712,n2713);
and (n2712,n931,n599);
and (n2713,n1135,n603);
xor (n2714,n2715,n601);
or (n2715,n2716,n2717);
and (n2716,n795,n822);
and (n2717,n797,n826);
xor (n2718,n2719,n380);
or (n2719,n2720,n2721);
and (n2720,n1139,n460);
and (n2721,n1141,n464);
nand (n2722,n2723,n2737,n2742);
nand (n2723,n2724,n2728);
xor (n2724,n2725,n601);
or (n2725,n2726,n2727);
and (n2726,n797,n822);
and (n2727,n931,n826);
and (n2728,n2729,n2733);
xnor (n2729,n2730,n949);
nor (n2730,n2731,n2732);
and (n2731,n791,n1150);
and (n2732,n570,n1152);
xor (n2733,n2734,n824);
or (n2734,n2735,n2736);
and (n2735,n795,n947);
and (n2736,n797,n951);
nand (n2737,n2738,n2728);
xor (n2738,n2739,n380);
or (n2739,n2740,n2741);
and (n2740,n1141,n460);
and (n2741,n1164,n464);
nand (n2742,n2724,n2738);
nand (n2743,n2657,n2702);
xor (n2744,n2745,n2759);
xor (n2745,n2746,n2755);
xor (n2746,n2747,n2753);
xor (n2747,n2748,n2752);
xor (n2748,n2749,n20);
or (n2749,n2750,n2751);
and (n2750,n1141,n378);
and (n2751,n1164,n382);
xor (n2752,n1906,n24);
xor (n2753,n2754,n1949);
xor (n2754,n1942,n1946);
nand (n2755,n2756,n2757,n2758);
nand (n2756,n2704,n2708);
nand (n2757,n2722,n2708);
nand (n2758,n2704,n2722);
xor (n2759,n2760,n2769);
xor (n2760,n2761,n2765);
nand (n2761,n2762,n2763,n2764);
nand (n2762,n2659,n2660);
nand (n2763,n2664,n2660);
nand (n2764,n2659,n2664);
nand (n2765,n2766,n2767,n2768);
nand (n2766,n2710,n2714);
nand (n2767,n2718,n2714);
nand (n2768,n2710,n2718);
xor (n2769,n2770,n1971);
xor (n2770,n1957,n1961);
nor (n2771,n2772,n2776);
nand (n2772,n2773,n2774,n2775);
nand (n2773,n2746,n2755);
nand (n2774,n2759,n2755);
nand (n2775,n2746,n2759);
xor (n2776,n2777,n2784);
xor (n2777,n2778,n2780);
xor (n2778,n2779,n1955);
xor (n2779,n1936,n1940);
nand (n2780,n2781,n2782,n2783);
nand (n2781,n2761,n2765);
nand (n2782,n2769,n2765);
nand (n2783,n2761,n2769);
xor (n2784,n2785,n2790);
xor (n2785,n2786,n2788);
xor (n2786,n2787,n1905);
xor (n2787,n1896,n1900);
xor (n2788,n2789,n1920);
xor (n2789,n1914,n1918);
nand (n2790,n2791,n2792,n2793);
nand (n2791,n2748,n2752);
nand (n2792,n2753,n2752);
nand (n2793,n2748,n2753);
nor (n2794,n2795,n2810);
nor (n2795,n2796,n2800);
nand (n2796,n2797,n2798,n2799);
nand (n2797,n2778,n2780);
nand (n2798,n2784,n2780);
nand (n2799,n2778,n2784);
xor (n2800,n2801,n2808);
xor (n2801,n2802,n2804);
xor (n2802,n2803,n1912);
xor (n2803,n1892,n1894);
nand (n2804,n2805,n2806,n2807);
nand (n2805,n2786,n2788);
nand (n2806,n2790,n2788);
nand (n2807,n2786,n2790);
xor (n2808,n2809,n1934);
xor (n2809,n1929,n1931);
nor (n2810,n2811,n2815);
nand (n2811,n2812,n2813,n2814);
nand (n2812,n2802,n2804);
nand (n2813,n2808,n2804);
nand (n2814,n2802,n2808);
xor (n2815,n2816,n1927);
xor (n2816,n1802,n1853);
nor (n2817,n2818,n2940);
nor (n2818,n2819,n2916);
nor (n2819,n2820,n2913);
nor (n2820,n2821,n2889);
nand (n2821,n2822,n2861);
or (n2822,n2823,n2847,n2860);
and (n2823,n2824,n2833);
xor (n2824,n2825,n2829);
xnor (n2825,n2826,n949);
nor (n2826,n2827,n2828);
and (n2827,n797,n1150);
and (n2828,n795,n1152);
xnor (n2829,n2830,n824);
nor (n2830,n2831,n2832);
and (n2831,n1135,n951);
and (n2832,n931,n947);
or (n2833,n2834,n2841,n2846);
and (n2834,n2835,n2837);
not (n2835,n2836);
nand (n2836,n1178,n599);
xnor (n2837,n2838,n949);
nor (n2838,n2839,n2840);
and (n2839,n931,n1150);
and (n2840,n797,n1152);
and (n2841,n2837,n2842);
xnor (n2842,n2843,n824);
nor (n2843,n2844,n2845);
and (n2844,n1139,n951);
and (n2845,n1135,n947);
and (n2846,n2835,n2842);
and (n2847,n2833,n2848);
xor (n2848,n2849,n2856);
xor (n2849,n2850,n2852);
and (n2850,n462,n2851);
xnor (n2851,n2836,n462);
xnor (n2852,n2853,n601);
nor (n2853,n2854,n2855);
and (n2854,n1141,n826);
and (n2855,n1139,n822);
xnor (n2856,n2857,n462);
nor (n2857,n2858,n2859);
and (n2858,n1178,n603);
and (n2859,n1164,n599);
and (n2860,n2824,n2848);
xor (n2861,n2862,n2878);
xor (n2862,n2863,n2867);
or (n2863,n2864,n2865,n2866);
and (n2864,n2850,n2852);
and (n2865,n2852,n2856);
and (n2866,n2850,n2856);
xor (n2867,n2868,n2874);
xor (n2868,n2869,n2870);
and (n2869,n2825,n2829);
xnor (n2870,n2871,n601);
nor (n2871,n2872,n2873);
and (n2872,n1139,n826);
and (n2873,n1135,n822);
xnor (n2874,n2875,n462);
nor (n2875,n2876,n2877);
and (n2876,n1164,n603);
and (n2877,n1141,n599);
xor (n2878,n2879,n2885);
xor (n2879,n2880,n2881);
not (n2880,n2685);
xnor (n2881,n2882,n949);
nor (n2882,n2883,n2884);
and (n2883,n795,n1150);
and (n2884,n791,n1152);
xnor (n2885,n2886,n824);
nor (n2886,n2887,n2888);
and (n2887,n931,n951);
and (n2888,n797,n947);
nor (n2889,n2890,n2894);
or (n2890,n2891,n2892,n2893);
and (n2891,n2863,n2867);
and (n2892,n2867,n2878);
and (n2893,n2863,n2878);
xor (n2894,n2895,n2902);
xor (n2895,n2896,n2900);
or (n2896,n2897,n2898,n2899);
and (n2897,n2869,n2870);
and (n2898,n2870,n2874);
and (n2899,n2869,n2874);
xor (n2900,n2901,n2683);
xor (n2901,n2674,n2678);
xor (n2902,n2903,n2909);
xor (n2903,n2904,n2908);
xor (n2904,n2905,n380);
or (n2905,n2906,n2907);
and (n2906,n1164,n460);
and (n2907,n1178,n464);
xor (n2908,n2729,n2733);
or (n2909,n2910,n2911,n2912);
and (n2910,n2880,n2881);
and (n2911,n2881,n2885);
and (n2912,n2880,n2885);
not (n2913,n2914);
not (n2914,n2915);
and (n2915,n2890,n2894);
not (n2916,n2917);
nor (n2917,n2918,n2933);
nor (n2918,n2919,n2923);
nand (n2919,n2920,n2921,n2922);
nand (n2920,n2896,n2900);
nand (n2921,n2902,n2900);
nand (n2922,n2896,n2902);
xor (n2923,n2924,n2931);
xor (n2924,n2925,n2927);
xor (n2925,n2926,n2738);
xor (n2926,n2724,n2728);
nand (n2927,n2928,n2929,n2930);
nand (n2928,n2904,n2908);
nand (n2929,n2909,n2908);
nand (n2930,n2904,n2909);
xor (n2931,n2932,n2688);
xor (n2932,n2671,n2672);
nor (n2933,n2934,n2938);
nand (n2934,n2935,n2936,n2937);
nand (n2935,n2925,n2927);
nand (n2936,n2931,n2927);
nand (n2937,n2925,n2931);
xor (n2938,n2939,n2702);
xor (n2939,n2657,n2669);
not (n2940,n2941);
nor (n2941,n2942,n2944);
nor (n2942,n2943,n2933);
nand (n2943,n2919,n2923);
not (n2944,n2945);
nand (n2945,n2934,n2938);
not (n2946,n2947);
nor (n2947,n2948,n2955);
nor (n2948,n2949,n2954);
nor (n2949,n2950,n2952);
nor (n2950,n2951,n2771);
nand (n2951,n2655,n2744);
not (n2952,n2953);
nand (n2953,n2772,n2776);
not (n2954,n2794);
not (n2955,n2956);
nor (n2956,n2957,n2959);
nor (n2957,n2958,n2810);
nand (n2958,n2796,n2800);
not (n2959,n2960);
nand (n2960,n2811,n2815);
nand (n2961,n2962,n2966);
nor (n2962,n2963,n2652);
nand (n2963,n2964,n2917);
nor (n2964,n2965,n2889);
nor (n2965,n2822,n2861);
or (n2966,n2967,n2989);
and (n2967,n2968,n2970);
xor (n2968,n2969,n2848);
xor (n2969,n2824,n2833);
or (n2970,n2971,n2985,n2988);
and (n2971,n2972,n2981);
and (n2972,n2973,n2977);
xnor (n2973,n2974,n949);
nor (n2974,n2975,n2976);
and (n2975,n1135,n1150);
and (n2976,n931,n1152);
xnor (n2977,n2978,n824);
nor (n2978,n2979,n2980);
and (n2979,n1141,n951);
and (n2980,n1139,n947);
xnor (n2981,n2982,n601);
nor (n2982,n2983,n2984);
and (n2983,n1164,n826);
and (n2984,n1141,n822);
and (n2985,n2981,n2986);
xor (n2986,n2987,n2842);
xor (n2987,n2835,n2837);
and (n2988,n2972,n2986);
and (n2989,n2990,n2991);
xor (n2990,n2968,n2970);
or (n2991,n2992,n3007);
and (n2992,n2993,n3005);
or (n2993,n2994,n2999,n3004);
and (n2994,n2995,n2996);
xor (n2995,n2973,n2977);
and (n2996,n601,n2997);
xnor (n2997,n2998,n601);
nand (n2998,n1178,n822);
and (n2999,n2996,n3000);
xnor (n3000,n3001,n601);
nor (n3001,n3002,n3003);
and (n3002,n1178,n826);
and (n3003,n1164,n822);
and (n3004,n2995,n3000);
xor (n3005,n3006,n2986);
xor (n3006,n2972,n2981);
and (n3007,n3008,n3009);
xor (n3008,n2993,n3005);
or (n3009,n3010,n3026);
and (n3010,n3011,n3013);
xor (n3011,n3012,n3000);
xor (n3012,n2995,n2996);
or (n3013,n3014,n3020,n3025);
and (n3014,n3015,n3016);
not (n3015,n2998);
xnor (n3016,n3017,n949);
nor (n3017,n3018,n3019);
and (n3018,n1139,n1150);
and (n3019,n1135,n1152);
and (n3020,n3016,n3021);
xnor (n3021,n3022,n824);
nor (n3022,n3023,n3024);
and (n3023,n1164,n951);
and (n3024,n1141,n947);
and (n3025,n3015,n3021);
and (n3026,n3027,n3028);
xor (n3027,n3011,n3013);
or (n3028,n3029,n3040);
and (n3029,n3030,n3032);
xor (n3030,n3031,n3021);
xor (n3031,n3015,n3016);
and (n3032,n3033,n3036);
and (n3033,n824,n3034);
xnor (n3034,n3035,n824);
nand (n3035,n1178,n947);
xnor (n3036,n3037,n949);
nor (n3037,n3038,n3039);
and (n3038,n1141,n1150);
and (n3039,n1139,n1152);
and (n3040,n3041,n3042);
xor (n3041,n3030,n3032);
or (n3042,n3043,n3049);
and (n3043,n3044,n3048);
xnor (n3044,n3045,n824);
nor (n3045,n3046,n3047);
and (n3046,n1178,n951);
and (n3047,n1164,n947);
xor (n3048,n3033,n3036);
and (n3049,n3050,n3051);
xor (n3050,n3044,n3048);
or (n3051,n3052,n3058);
and (n3052,n3053,n3057);
xnor (n3053,n3054,n949);
nor (n3054,n3055,n3056);
and (n3055,n1164,n1150);
and (n3056,n1141,n1152);
not (n3057,n3035);
and (n3058,n3059,n3060);
xor (n3059,n3053,n3057);
and (n3060,n3061,n3065);
xnor (n3061,n3062,n949);
nor (n3062,n3063,n3064);
and (n3063,n1178,n1150);
and (n3064,n1164,n1152);
and (n3065,n3066,n949);
xnor (n3066,n3067,n949);
nand (n3067,n1178,n1152);
not (n3068,n3069);
nand (n3069,n3070,n2090);
nor (n3070,n3071,n1122);
nand (n3071,n3072,n2045);
nor (n3072,n3073,n2017);
nor (n3073,n1800,n1979);
not (n3074,n3075);
nand (n3075,n3076,n271);
nor (n3076,n3077,n231);
nor (n3077,n7,n191);
nand (n3078,n3079,n3103);
not (n3079,n3080);
nor (n3080,n3081,n3085);
nand (n3081,n3082,n3083,n3084);
nand (n3082,n314,n318);
nand (n3083,n330,n318);
nand (n3084,n314,n330);
xor (n3085,n3086,n3099);
xor (n3086,n3087,n3091);
nand (n3087,n3088,n3089,n3090);
nand (n3088,n287,n322);
nand (n3089,n326,n322);
nand (n3090,n287,n326);
xor (n3091,n3092,n3095);
or (n3092,n3093,n3094);
and (n3093,n31,n87);
and (n3094,n39,n91);
not (n3095,n3096);
xor (n3096,n3097,n72);
or (n3097,n324,n3098);
and (n3098,n17,n70);
nand (n3099,n3100,n3101,n3102);
nand (n3100,n93,n288);
nand (n3101,n320,n288);
nand (n3102,n93,n320);
nand (n3103,n3081,n3085);
xor (n3104,n3105,n3407);
not (n3105,n3106);
xor (n3106,n3107,n3124);
xor (n3107,n3108,n3111);
xor (n3108,n3109,n3087);
xor (n3109,n3096,n3110);
xor (n3110,n3092,n93);
or (n3111,n3112,n3114,n3123);
and (n3112,n3113,n320);
not (n3113,n315);
and (n3114,n320,n3115);
or (n3115,n3116,n3117,n3122);
and (n3116,n288,n276);
and (n3117,n276,n3118);
or (n3118,n3119,n3120,n3121);
not (n3119,n292);
and (n3120,n246,n256);
and (n3121,n219,n256);
and (n3122,n288,n3118);
and (n3123,n3113,n3115);
or (n3124,n3125,n3165,n3406);
and (n3125,n3126,n3128);
xor (n3126,n3127,n3115);
xor (n3127,n3113,n320);
or (n3128,n3129,n3137,n3164);
and (n3129,n3130,n3135);
or (n3130,n3131,n3132,n3134);
and (n3131,n250,n240);
and (n3132,n240,n3133);
xor (n3133,n245,n256);
and (n3134,n250,n3133);
xor (n3135,n3136,n3118);
xor (n3136,n288,n276);
and (n3137,n3135,n3138);
or (n3138,n3139,n3147,n3163);
and (n3139,n3140,n3145);
or (n3140,n3141,n3142,n3144);
and (n3141,n220,n199);
and (n3142,n199,n3143);
not (n3143,n214);
and (n3144,n220,n3143);
xor (n3145,n3146,n3133);
xor (n3146,n250,n240);
and (n3147,n3145,n3148);
or (n3148,n3149,n3159,n3162);
and (n3149,n3150,n3154);
or (n3150,n3151,n3152,n3153);
and (n3151,n77,n129);
not (n3152,n225);
and (n3153,n77,n133);
or (n3154,n3155,n3156,n3158);
and (n3155,n128,n111);
and (n3156,n111,n3157);
not (n3157,n98);
and (n3158,n128,n3157);
and (n3159,n3154,n3160);
xor (n3160,n3161,n3143);
xor (n3161,n220,n199);
and (n3162,n3150,n3160);
and (n3163,n3140,n3148);
and (n3164,n3130,n3138);
and (n3165,n3128,n3166);
or (n3166,n3167,n3169);
xor (n3167,n3168,n3138);
xor (n3168,n3130,n3135);
or (n3169,n3170,n3201,n3405);
and (n3170,n3171,n3173);
xor (n3171,n3172,n3148);
xor (n3172,n3140,n3145);
or (n3173,n3174,n3186,n3200);
and (n3174,n3175,n3184);
or (n3175,n3176,n3181,n3183);
and (n3176,n3177,n104);
or (n3177,n3178,n3179,n3180);
and (n3178,n128,n80);
not (n3179,n124);
and (n3180,n128,n84);
and (n3181,n104,n3182);
not (n3182,n126);
and (n3183,n3177,n3182);
xor (n3184,n3185,n3160);
xor (n3185,n3150,n3154);
and (n3186,n3184,n3187);
or (n3187,n3188,n3196,n3199);
and (n3188,n3189,n3194);
or (n3189,n3190,n3192,n3193);
and (n3190,n3191,n141);
not (n3191,n75);
and (n3192,n141,n11);
and (n3193,n3191,n11);
xor (n3194,n3195,n3157);
xor (n3195,n128,n111);
and (n3196,n3194,n3197);
xor (n3197,n3198,n3182);
xor (n3198,n3177,n104);
and (n3199,n3189,n3197);
and (n3200,n3175,n3187);
and (n3201,n3173,n3202);
or (n3202,n3203,n3291,n3404);
and (n3203,n3204,n3206);
xor (n3204,n3205,n3187);
xor (n3205,n3175,n3184);
or (n3206,n3207,n3228,n3290);
and (n3207,n3208,n3226);
or (n3208,n3209,n3222,n3225);
and (n3209,n3210,n3214);
or (n3210,n3211,n3212,n3213);
not (n3211,n73);
and (n3212,n62,n144);
and (n3213,n50,n144);
or (n3214,n3215,n3220,n3221);
and (n3215,n150,n3216);
or (n3216,n3217,n3218,n3219);
and (n3217,n14,n172);
not (n3218,n171);
and (n3219,n14,n176);
and (n3220,n3216,n183);
and (n3221,n150,n183);
and (n3222,n3214,n3223);
xor (n3223,n3224,n11);
xor (n3224,n3191,n141);
and (n3225,n3210,n3223);
xor (n3226,n3227,n3197);
xor (n3227,n3189,n3194);
and (n3228,n3226,n3229);
or (n3229,n3230,n3243,n3289);
and (n3230,n3231,n3241);
or (n3231,n3232,n3237,n3240);
and (n3232,n3233,n3235);
xor (n3233,n3234,n144);
xor (n3234,n50,n62);
and (n3235,n351,n3236);
not (n3236,n353);
and (n3237,n3235,n3238);
xor (n3238,n3239,n183);
xor (n3239,n150,n3216);
and (n3240,n3233,n3238);
xor (n3241,n3242,n3223);
xor (n3242,n3210,n3214);
and (n3243,n3241,n3244);
or (n3244,n3245,n3258,n3288);
and (n3245,n3246,n3256);
or (n3246,n3247,n3253,n3255);
and (n3247,n3248,n3249);
not (n3248,n356);
or (n3249,n3250,n3251,n3252);
not (n3250,n373);
and (n3251,n384,n395);
and (n3252,n374,n395);
and (n3253,n3249,n3254);
not (n3254,n350);
and (n3255,n3248,n3254);
xor (n3256,n3257,n3238);
xor (n3257,n3233,n3235);
and (n3258,n3256,n3259);
or (n3259,n3260,n3274,n3287);
and (n3260,n3261,n3265);
or (n3261,n3262,n3263,n3264);
and (n3262,n388,n400);
and (n3263,n400,n442);
and (n3264,n388,n442);
or (n3265,n3266,n3271,n3273);
and (n3266,n409,n3267);
or (n3267,n3268,n3269,n3270);
and (n3268,n375,n428);
not (n3269,n432);
and (n3270,n375,n433);
and (n3271,n3267,n3272);
xor (n3272,n408,n395);
and (n3273,n409,n3272);
and (n3274,n3265,n3275);
or (n3275,n3276,n3283,n3286);
and (n3276,n3277,n3278);
not (n3277,n480);
or (n3278,n3279,n3281,n3282);
and (n3279,n448,n3280);
not (n3280,n524);
and (n3281,n3280,n454);
not (n3282,n475);
and (n3283,n3278,n3284);
xor (n3284,n3285,n442);
xor (n3285,n388,n400);
and (n3286,n3277,n3284);
and (n3287,n3261,n3275);
and (n3288,n3246,n3259);
and (n3289,n3231,n3244);
and (n3290,n3208,n3229);
and (n3291,n3206,n3292);
or (n3292,n3293,n3295);
xor (n3293,n3294,n3229);
xor (n3294,n3208,n3226);
or (n3295,n3296,n3298);
xor (n3296,n3297,n3244);
xor (n3297,n3231,n3241);
or (n3298,n3299,n3331,n3403);
and (n3299,n3300,n3329);
or (n3300,n3301,n3325,n3328);
and (n3301,n3302,n3304);
xor (n3302,n3303,n3254);
xor (n3303,n3248,n3249);
or (n3304,n3305,n3321,n3324);
and (n3305,n3306,n3308);
xor (n3306,n3307,n3272);
xor (n3307,n409,n3267);
or (n3308,n3309,n3315,n3320);
and (n3309,n557,n3310);
and (n3310,n3311,n573);
or (n3311,n3312,n3313,n3314);
and (n3312,n457,n562);
not (n3313,n561);
and (n3314,n457,n566);
and (n3315,n3310,n3316);
or (n3316,n3317,n3318,n3319);
not (n3317,n507);
and (n3318,n508,n533);
and (n3319,n503,n533);
and (n3320,n557,n3316);
and (n3321,n3308,n3322);
xor (n3322,n3323,n3284);
xor (n3323,n3277,n3278);
and (n3324,n3306,n3322);
and (n3325,n3304,n3326);
xor (n3326,n3327,n3275);
xor (n3327,n3261,n3265);
and (n3328,n3302,n3326);
xor (n3329,n3330,n3259);
xor (n3330,n3246,n3256);
and (n3331,n3329,n3332);
or (n3332,n3333,n3335);
xor (n3333,n3334,n3326);
xor (n3334,n3302,n3304);
or (n3335,n3336,n3367,n3402);
and (n3336,n3337,n3365);
or (n3337,n3338,n3347,n3364);
and (n3338,n3339,n3341);
xor (n3339,n3340,n454);
xor (n3340,n448,n3280);
or (n3341,n3342,n3344,n3346);
and (n3342,n3343,n530);
not (n3343,n583);
and (n3344,n530,n3345);
xor (n3345,n3311,n573);
and (n3346,n3343,n3345);
and (n3347,n3341,n3348);
or (n3348,n3349,n3360,n3363);
and (n3349,n3350,n3355);
or (n3350,n3351,n3353,n3354);
and (n3351,n617,n3352);
not (n3352,n1022);
and (n3353,n3352,n1021);
and (n3354,n617,n1021);
or (n3355,n3356,n3358,n3359);
and (n3356,n620,n3357);
not (n3357,n1017);
and (n3358,n3357,n593);
and (n3359,n620,n593);
and (n3360,n3355,n3361);
xor (n3361,n3362,n533);
xor (n3362,n503,n508);
and (n3363,n3350,n3361);
and (n3364,n3339,n3348);
xor (n3365,n3366,n3322);
xor (n3366,n3306,n3308);
and (n3367,n3365,n3368);
or (n3368,n3369,n3398,n3401);
and (n3369,n3370,n3372);
xor (n3370,n3371,n3316);
xor (n3371,n557,n3310);
or (n3372,n3373,n3394,n3397);
and (n3373,n3374,n3392);
or (n3374,n3375,n3388,n3391);
and (n3375,n3376,n3380);
or (n3376,n3377,n3378,n3379);
and (n3377,n701,n775);
and (n3378,n775,n844);
and (n3379,n701,n844);
or (n3380,n3381,n3382,n3387);
and (n3381,n705,n777);
and (n3382,n777,n3383);
or (n3383,n3384,n3385,n3386);
and (n3384,n596,n806);
not (n3385,n842);
and (n3386,n596,n802);
and (n3387,n705,n3383);
and (n3388,n3380,n3389);
xor (n3389,n3390,n1021);
xor (n3390,n617,n3352);
and (n3391,n3376,n3389);
xor (n3392,n3393,n3345);
xor (n3393,n3343,n530);
and (n3394,n3392,n3395);
xor (n3395,n3396,n3361);
xor (n3396,n3350,n3355);
and (n3397,n3374,n3395);
and (n3398,n3372,n3399);
xor (n3399,n3400,n3348);
xor (n3400,n3339,n3341);
and (n3401,n3370,n3399);
and (n3402,n3337,n3368);
and (n3403,n3300,n3332);
and (n3404,n3204,n3292);
and (n3405,n3171,n3202);
and (n3406,n3126,n3166);
and (n3407,n3408,n3410);
xor (n3408,n3409,n3166);
xor (n3409,n3126,n3128);
and (n3410,n3411,n3412);
xnor (n3411,n3167,n3169);
and (n3412,n3413,n3415);
xor (n3413,n3414,n3202);
xor (n3414,n3171,n3173);
and (n3415,n3416,n3418);
xor (n3416,n3417,n3292);
xor (n3417,n3204,n3206);
and (n3418,n3419,n3420);
xnor (n3419,n3293,n3295);
and (n3420,n3421,n3422);
xnor (n3421,n3296,n3298);
and (n3422,n3423,n3425);
xor (n3423,n3424,n3332);
xor (n3424,n3300,n3329);
and (n3425,n3426,n3427);
xnor (n3426,n3333,n3335);
or (n3427,n3428,n3508);
and (n3428,n3429,n3431);
xor (n3429,n3430,n3368);
xor (n3430,n3337,n3365);
or (n3431,n3432,n3434);
xor (n3432,n3433,n3399);
xor (n3433,n3370,n3372);
or (n3434,n3435,n3458,n3507);
and (n3435,n3436,n3456);
or (n3436,n3437,n3452,n3455);
and (n3437,n3438,n3440);
xor (n3438,n3439,n593);
xor (n3439,n620,n3357);
or (n3440,n3441,n3448,n3451);
and (n3441,n773,n3442);
or (n3442,n3443,n3445,n3447);
and (n3443,n834,n3444);
not (n3444,n800);
and (n3445,n3444,n3446);
not (n3446,n786);
and (n3447,n834,n3446);
and (n3448,n3442,n3449);
xor (n3449,n3450,n844);
xor (n3450,n701,n775);
and (n3451,n773,n3449);
and (n3452,n3440,n3453);
xor (n3453,n3454,n3389);
xor (n3454,n3376,n3380);
and (n3455,n3438,n3453);
xor (n3456,n3457,n3395);
xor (n3457,n3374,n3392);
and (n3458,n3456,n3459);
or (n3459,n3460,n3471,n3506);
and (n3460,n3461,n3469);
or (n3461,n3462,n3465,n3468);
and (n3462,n3463,n721);
xor (n3463,n3464,n3383);
xor (n3464,n705,n777);
and (n3465,n721,n3466);
xor (n3466,n3467,n3449);
xor (n3467,n773,n3442);
and (n3468,n3463,n3466);
xor (n3469,n3470,n3453);
xor (n3470,n3438,n3440);
and (n3471,n3469,n3472);
or (n3472,n3473,n3502,n3505);
and (n3473,n3474,n3487);
or (n3474,n3475,n3485,n3486);
and (n3475,n3476,n879);
or (n3476,n3477,n3482,n3484);
and (n3477,n3478,n873);
or (n3478,n3479,n3480,n3481);
and (n3479,n818,n863);
not (n3480,n867);
and (n3481,n818,n868);
and (n3482,n873,n3483);
not (n3483,n876);
and (n3484,n3478,n3483);
not (n3485,n914);
and (n3486,n3476,n915);
or (n3487,n3488,n3495,n3501);
and (n3488,n3489,n3493);
or (n3489,n3490,n3491,n3492);
and (n3490,n819,n815);
not (n3491,n833);
and (n3492,n819,n829);
xor (n3493,n3494,n3446);
xor (n3494,n834,n3444);
and (n3495,n3493,n3496);
or (n3496,n3497,n3498,n3500);
and (n3497,n818,n956);
and (n3498,n956,n3499);
not (n3499,n2570);
and (n3500,n818,n3499);
and (n3501,n3489,n3496);
and (n3502,n3487,n3503);
xor (n3503,n3504,n3466);
xor (n3504,n3463,n721);
and (n3505,n3474,n3503);
and (n3506,n3461,n3472);
and (n3507,n3436,n3459);
and (n3508,n3509,n3510);
xor (n3509,n3429,n3431);
and (n3510,n3511,n3512);
xnor (n3511,n3432,n3434);
or (n3512,n3513,n3598);
and (n3513,n3514,n3516);
xor (n3514,n3515,n3459);
xor (n3515,n3436,n3456);
or (n3516,n3517,n3519);
xor (n3517,n3518,n3472);
xor (n3518,n3461,n3469);
or (n3519,n3520,n3542,n3597);
and (n3520,n3521,n3540);
or (n3521,n3522,n3536,n3539);
and (n3522,n3523,n3525);
xor (n3523,n3524,n915);
xor (n3524,n3476,n879);
or (n3525,n3526,n3529,n3535);
and (n3526,n3527,n2573);
xor (n3527,n3528,n3483);
xor (n3528,n3478,n873);
and (n3529,n2573,n3530);
or (n3530,n3531,n3532,n3534);
not (n3531,n995);
and (n3532,n979,n3533);
not (n3533,n976);
and (n3534,n960,n3533);
and (n3535,n3527,n3530);
and (n3536,n3525,n3537);
xor (n3537,n3538,n3496);
xor (n3538,n3489,n3493);
and (n3539,n3523,n3537);
xor (n3540,n3541,n3503);
xor (n3541,n3474,n3487);
and (n3542,n3540,n3543);
or (n3543,n3544,n3559,n3596);
and (n3544,n3545,n3557);
or (n3545,n3546,n3553,n3556);
and (n3546,n3547,n3551);
or (n3547,n3548,n3549,n3550);
and (n3548,n927,n2543);
and (n3549,n2543,n2524);
and (n3550,n927,n2524);
xor (n3551,n3552,n3499);
xor (n3552,n818,n956);
and (n3553,n3551,n3554);
and (n3554,n2519,n3555);
not (n3555,n2517);
and (n3556,n3547,n3554);
xor (n3557,n3558,n3537);
xor (n3558,n3523,n3525);
and (n3559,n3557,n3560);
or (n3560,n3561,n3581,n3595);
and (n3561,n3562,n3579);
or (n3562,n3563,n3568,n3578);
and (n3563,n3564,n2546);
or (n3564,n3565,n3566,n3567);
and (n3565,n944,n935);
not (n3566,n934);
and (n3567,n944,n938);
and (n3568,n2546,n3569);
or (n3569,n3570,n3575,n3577);
and (n3570,n943,n3571);
or (n3571,n3572,n3573,n3574);
and (n3572,n943,n2347);
not (n3573,n2461);
and (n3574,n943,n2351);
and (n3575,n3571,n3576);
not (n3576,n2456);
and (n3577,n943,n3576);
and (n3578,n3564,n3569);
xor (n3579,n3580,n3530);
xor (n3580,n3527,n2573);
and (n3581,n3579,n3582);
or (n3582,n3583,n3587,n3594);
and (n3583,n3584,n3586);
xor (n3584,n3585,n2524);
xor (n3585,n927,n2543);
not (n3586,n2516);
and (n3587,n3586,n3588);
or (n3588,n3589,n3592,n3593);
and (n3589,n3590,n2462);
and (n3590,n2331,n3591);
not (n3591,n2345);
and (n3592,n2462,n2484);
and (n3593,n3590,n2484);
and (n3594,n3584,n3588);
and (n3595,n3562,n3582);
and (n3596,n3545,n3560);
and (n3597,n3521,n3543);
and (n3598,n3599,n3600);
xor (n3599,n3514,n3516);
and (n3600,n3601,n3602);
xnor (n3601,n3517,n3519);
or (n3602,n3603,n3807);
and (n3603,n3604,n3606);
xor (n3604,n3605,n3543);
xor (n3605,n3521,n3540);
or (n3606,n3607,n3682,n3806);
and (n3607,n3608,n3680);
or (n3608,n3609,n3676,n3679);
and (n3609,n3610,n3612);
xor (n3610,n3611,n3554);
xor (n3611,n3547,n3551);
or (n3612,n3613,n3647,n3675);
and (n3613,n3614,n3645);
or (n3614,n3615,n3633,n3644);
and (n3615,n3616,n3625);
and (n3616,n3617,n2371);
or (n3617,n3618,n3623,n3624);
and (n3618,n3619,n2241);
or (n3619,n3620,n3621,n3622);
and (n3620,n2310,n2106);
not (n3621,n2250);
and (n3622,n2310,n2110);
not (n3623,n2383);
and (n3624,n3619,n2245);
or (n3625,n3626,n3631,n3632);
and (n3626,n2411,n3627);
or (n3627,n3628,n3629,n3630);
and (n3628,n2310,n2230);
not (n3629,n2358);
and (n3630,n2310,n2235);
and (n3631,n3627,n2392);
and (n3632,n2411,n2392);
and (n3633,n3625,n3634);
or (n3634,n3635,n3641,n3643);
and (n3635,n3636,n3637);
not (n3636,n2330);
or (n3637,n3638,n3639,n3640);
and (n3638,n2114,n2306);
not (n3639,n2410);
and (n3640,n2114,n2311);
and (n3641,n3637,n3642);
not (n3642,n2387);
and (n3643,n3636,n3642);
and (n3644,n3616,n3634);
xor (n3645,n3646,n3569);
xor (n3646,n3564,n2546);
and (n3647,n3645,n3648);
or (n3648,n3649,n3671,n3674);
and (n3649,n3650,n3652);
xor (n3650,n3651,n3576);
xor (n3651,n943,n3571);
or (n3652,n3653,n3662,n3670);
and (n3653,n3654,n3661);
or (n3654,n3655,n3657,n3660);
and (n3655,n2290,n3656);
not (n3656,n2287);
and (n3657,n3656,n3658);
xor (n3658,n3659,n2235);
xor (n3659,n2310,n2230);
and (n3660,n2290,n3658);
xor (n3661,n3617,n2371);
and (n3662,n3661,n3663);
or (n3663,n3664,n3668,n3669);
and (n3664,n3665,n3666);
not (n3665,n2304);
xor (n3666,n3667,n2245);
xor (n3667,n3619,n2241);
and (n3668,n3666,n2264);
and (n3669,n3665,n2264);
and (n3670,n3654,n3663);
and (n3671,n3652,n3672);
xor (n3672,n3673,n2484);
xor (n3673,n3590,n2462);
and (n3674,n3650,n3672);
and (n3675,n3614,n3648);
and (n3676,n3612,n3677);
xor (n3677,n3678,n3582);
xor (n3678,n3562,n3579);
and (n3679,n3610,n3677);
xor (n3680,n3681,n3560);
xor (n3681,n3545,n3557);
and (n3682,n3680,n3683);
or (n3683,n3684,n3717,n3805);
and (n3684,n3685,n3715);
or (n3685,n3686,n3711,n3714);
and (n3686,n3687,n3689);
xor (n3687,n3688,n3588);
xor (n3688,n3584,n3586);
or (n3689,n3690,n3707,n3710);
and (n3690,n3691,n3693);
xor (n3691,n3692,n3634);
xor (n3692,n3616,n3625);
or (n3693,n3694,n3699,n3706);
and (n3694,n3695,n3697);
xor (n3695,n3696,n2392);
xor (n3696,n2411,n3627);
xor (n3697,n3698,n3642);
xor (n3698,n3636,n3637);
and (n3699,n3697,n3700);
and (n3700,n2255,n3701);
or (n3701,n3702,n3703,n3705);
not (n3702,n2261);
and (n3703,n2121,n3704);
not (n3704,n2104);
and (n3705,n2117,n3704);
and (n3706,n3695,n3700);
and (n3707,n3693,n3708);
xor (n3708,n3709,n3672);
xor (n3709,n3650,n3652);
and (n3710,n3691,n3708);
and (n3711,n3689,n3712);
xor (n3712,n3713,n3648);
xor (n3713,n3614,n3645);
and (n3714,n3687,n3712);
xor (n3715,n3716,n3677);
xor (n3716,n3610,n3612);
and (n3717,n3715,n3718);
or (n3718,n3719,n3776,n3804);
and (n3719,n3720,n3722);
xor (n3720,n3721,n3712);
xor (n3721,n3687,n3689);
or (n3722,n3723,n3755,n3775);
and (n3723,n3724,n3753);
or (n3724,n3725,n3738,n3752);
and (n3725,n3726,n3736);
or (n3726,n3727,n3734,n3735);
and (n3727,n3728,n3732);
or (n3728,n3729,n3730,n3731);
and (n3729,n2169,n2154);
and (n3730,n2154,n2137);
and (n3731,n2169,n2137);
xor (n3732,n3733,n3658);
xor (n3733,n2290,n3656);
and (n3734,n3732,n2315);
and (n3735,n3728,n2315);
xor (n3736,n3737,n3663);
xor (n3737,n3654,n3661);
and (n3738,n3736,n3739);
or (n3739,n3740,n3749,n3751);
and (n3740,n3741,n3747);
or (n3741,n3742,n3743,n3746);
and (n3742,n2159,n2153);
and (n3743,n2153,n3744);
xor (n3744,n3745,n2137);
xor (n3745,n2169,n2154);
and (n3746,n2159,n3744);
xor (n3747,n3748,n2264);
xor (n3748,n3665,n3666);
and (n3749,n3747,n3750);
xor (n3750,n2255,n3701);
and (n3751,n3741,n3750);
and (n3752,n3726,n3739);
xor (n3753,n3754,n3708);
xor (n3754,n3691,n3693);
and (n3755,n3753,n3756);
or (n3756,n3757,n3771,n3774);
and (n3757,n3758,n3760);
xor (n3758,n3759,n3700);
xor (n3759,n3695,n3697);
or (n3760,n3761,n3769,n3770);
and (n3761,n3762,n3764);
xor (n3762,n3763,n2315);
xor (n3763,n3728,n3732);
or (n3764,n3765,n3766,n3768);
not (n3765,n2214);
and (n3766,n2129,n3767);
not (n3767,n2102);
and (n3768,n2125,n3767);
and (n3769,n3764,n2216);
and (n3770,n3762,n2216);
and (n3771,n3760,n3772);
xor (n3772,n3773,n3739);
xor (n3773,n3726,n3736);
and (n3774,n3758,n3772);
and (n3775,n3724,n3756);
and (n3776,n3722,n3777);
or (n3777,n3778,n3780);
xor (n3778,n3779,n3756);
xor (n3779,n3724,n3753);
or (n3780,n3781,n3797,n3803);
and (n3781,n3782,n3795);
or (n3782,n3783,n3791,n3794);
and (n3783,n3784,n3786);
xor (n3784,n3785,n3750);
xor (n3785,n3741,n3747);
or (n3786,n3787,n3789,n3790);
and (n3787,n3788,n2201);
not (n3788,n2100);
not (n3789,n2208);
and (n3790,n3788,n2133);
and (n3791,n3786,n3792);
xor (n3792,n3793,n2216);
xor (n3793,n3762,n3764);
and (n3794,n3784,n3792);
xor (n3795,n3796,n3772);
xor (n3796,n3758,n3760);
and (n3797,n3795,n3798);
or (n3798,n3799,n3801);
or (n3799,n2094,n3800);
not (n3800,n2098);
xor (n3801,n3802,n3792);
xor (n3802,n3784,n3786);
and (n3803,n3782,n3798);
and (n3804,n3720,n3777);
and (n3805,n3685,n3718);
and (n3806,n3608,n3683);
and (n3807,n3808,n3809);
xor (n3808,n3604,n3606);
and (n3809,n3810,n3812);
xor (n3810,n3811,n3683);
xor (n3811,n3608,n3680);
or (n3812,n3813,n3815);
xor (n3813,n3814,n3718);
xor (n3814,n3685,n3715);
and (n3815,n3816,n3817);
not (n3816,n3813);
and (n3817,n3818,n3820);
xor (n3818,n3819,n3777);
xor (n3819,n3720,n3722);
and (n3820,n3821,n3822);
xnor (n3821,n3778,n3780);
and (n3822,n3823,n3825);
xor (n3823,n3824,n3798);
xor (n3824,n3782,n3795);
and (n3825,n3826,n3827);
xnor (n3826,n3799,n3801);
and (n3827,n3828,n3831);
not (n3828,n3829);
nand (n3829,n3830,n2623);
not (n3830,n2093);
nand (n3831,n1120,n3832);
nand (n3832,n3070,n2649);
endmodule
