module top (out,n12,n16,n19,n20,n30,n33,n34,n38,n48
        ,n51,n52,n55,n57,n64,n67,n68,n72,n78,n86
        ,n89,n90,n94,n101,n104,n105,n109,n117,n120,n124
        ,n360,n431,n516);
output out;
input n12;
input n16;
input n19;
input n20;
input n30;
input n33;
input n34;
input n38;
input n48;
input n51;
input n52;
input n55;
input n57;
input n64;
input n67;
input n68;
input n72;
input n78;
input n86;
input n89;
input n90;
input n94;
input n101;
input n104;
input n105;
input n109;
input n117;
input n120;
input n124;
input n360;
input n431;
input n516;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n53;
wire n54;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n102;
wire n103;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
xor (out,n0,n1173);
xor (n0,n1,n382);
xor (n1,n2,n312);
xor (n2,n3,n258);
or (n3,n4,n209,n257);
and (n4,n5,n198);
or (n5,n6,n164,n197);
and (n6,n7,n130);
or (n7,n8,n80,n129);
and (n8,n9,n43);
or (n9,n10,n26,n42);
and (n10,n11,n13);
not (n11,n12);
xnor (n13,n14,n23);
not (n14,n15);
and (n15,n16,n17);
and (n17,n18,n21);
xor (n18,n19,n20);
not (n21,n22);
xor (n22,n20,n12);
and (n23,n19,n24);
not (n24,n25);
and (n25,n20,n12);
and (n26,n13,n27);
xnor (n27,n28,n39);
nor (n28,n29,n37);
and (n29,n30,n31);
and (n31,n32,n35);
xor (n32,n33,n34);
not (n35,n36);
xor (n36,n34,n19);
and (n37,n38,n36);
and (n39,n33,n40);
not (n40,n41);
and (n41,n34,n19);
and (n42,n11,n27);
or (n43,n44,n76,n79);
and (n44,n45,n61);
xnor (n45,n46,n58);
nor (n46,n47,n56);
and (n47,n48,n49);
and (n49,n50,n53);
xor (n50,n51,n52);
not (n53,n54);
xor (n54,n52,n55);
and (n56,n57,n54);
and (n58,n51,n59);
not (n59,n60);
and (n60,n52,n55);
xnor (n61,n62,n73);
nor (n62,n63,n71);
and (n63,n64,n65);
and (n65,n66,n69);
xor (n66,n67,n68);
not (n69,n70);
xor (n70,n68,n51);
and (n71,n72,n70);
and (n73,n67,n74);
not (n74,n75);
and (n75,n68,n51);
and (n76,n61,n77);
and (n77,n78,n67);
and (n79,n45,n77);
and (n80,n43,n81);
or (n81,n82,n113,n128);
and (n82,n83,n98);
xnor (n83,n84,n95);
nor (n84,n85,n93);
and (n85,n86,n87);
and (n87,n88,n91);
xor (n88,n89,n90);
not (n91,n92);
xor (n92,n90,n33);
and (n93,n94,n92);
and (n95,n89,n96);
not (n96,n97);
and (n97,n90,n33);
xnor (n98,n99,n110);
nor (n99,n100,n108);
and (n100,n101,n102);
and (n102,n103,n106);
xor (n103,n104,n105);
not (n106,n107);
xor (n107,n105,n89);
and (n108,n109,n107);
and (n110,n104,n111);
not (n111,n112);
and (n112,n105,n89);
and (n113,n98,n114);
xnor (n114,n115,n125);
nor (n115,n116,n123);
and (n116,n117,n118);
and (n118,n119,n121);
xor (n119,n55,n120);
not (n121,n122);
xor (n122,n120,n104);
and (n123,n124,n122);
and (n125,n55,n126);
not (n126,n127);
and (n127,n120,n104);
and (n128,n83,n114);
and (n129,n9,n81);
or (n130,n131,n156,n163);
and (n131,n132,n142);
xor (n132,n133,n138);
xor (n133,n23,n134);
xnor (n134,n135,n39);
nor (n135,n136,n137);
and (n136,n38,n31);
and (n137,n16,n36);
xnor (n138,n139,n95);
nor (n139,n140,n141);
and (n140,n94,n87);
and (n141,n30,n92);
xor (n142,n143,n152);
xor (n143,n144,n148);
xnor (n144,n145,n110);
nor (n145,n146,n147);
and (n146,n109,n102);
and (n147,n86,n107);
xnor (n148,n149,n125);
nor (n149,n150,n151);
and (n150,n124,n118);
and (n151,n101,n122);
xnor (n152,n153,n58);
nor (n153,n154,n155);
and (n154,n57,n49);
and (n155,n117,n54);
and (n156,n142,n157);
xnor (n157,n158,n162);
xnor (n158,n159,n73);
nor (n159,n160,n161);
and (n160,n72,n65);
and (n161,n48,n70);
and (n162,n64,n67);
and (n163,n132,n157);
and (n164,n130,n165);
xor (n165,n166,n191);
xor (n166,n167,n177);
xor (n167,n168,n173);
xor (n168,n169,n170);
not (n169,n23);
xnor (n170,n171,n39);
not (n171,n172);
and (n172,n16,n31);
xnor (n173,n174,n95);
nor (n174,n175,n176);
and (n175,n30,n87);
and (n176,n38,n92);
xor (n177,n178,n187);
xor (n178,n179,n183);
xnor (n179,n180,n110);
nor (n180,n181,n182);
and (n181,n86,n102);
and (n182,n94,n107);
xnor (n183,n184,n125);
nor (n184,n185,n186);
and (n185,n101,n118);
and (n186,n109,n122);
xnor (n187,n188,n58);
nor (n188,n189,n190);
and (n189,n117,n49);
and (n190,n124,n54);
xor (n191,n192,n196);
xnor (n192,n193,n73);
nor (n193,n194,n195);
and (n194,n48,n65);
and (n195,n57,n70);
and (n196,n72,n67);
and (n197,n7,n165);
xor (n198,n199,n208);
xor (n199,n200,n204);
or (n200,n201,n202,n203);
and (n201,n169,n170);
and (n202,n170,n173);
and (n203,n169,n173);
or (n204,n205,n206,n207);
and (n205,n179,n183);
and (n206,n183,n187);
and (n207,n179,n187);
and (n208,n192,n196);
and (n209,n198,n210);
xor (n210,n211,n229);
xor (n211,n212,n225);
or (n212,n213,n222,n224);
and (n213,n214,n218);
or (n214,n215,n216,n217);
and (n215,n23,n134);
and (n216,n134,n138);
and (n217,n23,n138);
or (n218,n219,n220,n221);
and (n219,n144,n148);
and (n220,n148,n152);
and (n221,n144,n152);
and (n222,n218,n223);
or (n223,n158,n162);
and (n224,n214,n223);
or (n225,n226,n227,n228);
and (n226,n167,n177);
and (n227,n177,n191);
and (n228,n167,n191);
xor (n229,n230,n243);
xor (n230,n231,n232);
and (n231,n48,n67);
not (n232,n233);
xor (n233,n234,n239);
xor (n234,n39,n235);
xnor (n235,n236,n95);
nor (n236,n237,n238);
and (n237,n38,n87);
and (n238,n16,n92);
xnor (n239,n240,n110);
nor (n240,n241,n242);
and (n241,n94,n102);
and (n242,n30,n107);
xor (n243,n244,n253);
xor (n244,n245,n249);
xnor (n245,n246,n125);
nor (n246,n247,n248);
and (n247,n109,n118);
and (n248,n86,n122);
xnor (n249,n250,n58);
nor (n250,n251,n252);
and (n251,n124,n49);
and (n252,n101,n54);
xnor (n253,n254,n73);
nor (n254,n255,n256);
and (n255,n57,n65);
and (n256,n117,n70);
and (n257,n5,n210);
xor (n258,n259,n274);
xor (n259,n260,n264);
or (n260,n261,n262,n263);
and (n261,n212,n225);
and (n262,n225,n229);
and (n263,n212,n229);
xor (n264,n265,n231);
xor (n265,n266,n270);
or (n266,n267,n268,n269);
and (n267,n39,n235);
and (n268,n235,n239);
and (n269,n39,n239);
or (n270,n271,n272,n273);
and (n271,n245,n249);
and (n272,n249,n253);
and (n273,n245,n253);
xor (n274,n275,n285);
xor (n275,n276,n280);
or (n276,n277,n278,n279);
and (n277,n200,n204);
and (n278,n204,n208);
and (n279,n200,n208);
or (n280,n281,n282,n284);
and (n281,n233,n243);
and (n282,n243,n283);
not (n283,n231);
and (n284,n233,n283);
xor (n285,n286,n302);
xor (n286,n287,n288);
and (n287,n57,n67);
xor (n288,n289,n298);
xor (n289,n290,n294);
xnor (n290,n291,n125);
nor (n291,n292,n293);
and (n292,n86,n118);
and (n293,n94,n122);
xnor (n294,n295,n58);
nor (n295,n296,n297);
and (n296,n101,n49);
and (n297,n109,n54);
xnor (n298,n299,n73);
nor (n299,n300,n301);
and (n300,n117,n65);
and (n301,n124,n70);
xor (n302,n303,n308);
xor (n303,n304,n305);
not (n304,n39);
xnor (n305,n306,n95);
not (n306,n307);
and (n307,n16,n87);
xnor (n308,n309,n110);
nor (n309,n310,n311);
and (n310,n30,n102);
and (n311,n38,n107);
and (n312,n313,n380);
or (n313,n314,n376,n379);
and (n314,n315,n374);
or (n315,n316,n368,n373);
and (n316,n317,n363);
or (n317,n318,n347,n362);
and (n318,n319,n335);
or (n319,n320,n329,n334);
and (n320,n321,n325);
xnor (n321,n322,n95);
nor (n322,n323,n324);
and (n323,n109,n87);
and (n324,n86,n92);
xnor (n325,n326,n110);
nor (n326,n327,n328);
and (n327,n124,n102);
and (n328,n101,n107);
and (n329,n325,n330);
xnor (n330,n331,n125);
nor (n331,n332,n333);
and (n332,n57,n118);
and (n333,n117,n122);
and (n334,n321,n330);
or (n335,n336,n341,n346);
and (n336,n12,n337);
xnor (n337,n338,n23);
nor (n338,n339,n340);
and (n339,n38,n17);
and (n340,n16,n22);
and (n341,n337,n342);
xnor (n342,n343,n39);
nor (n343,n344,n345);
and (n344,n94,n31);
and (n345,n30,n36);
and (n346,n12,n342);
and (n347,n335,n348);
or (n348,n349,n358,n361);
and (n349,n350,n354);
xnor (n350,n351,n58);
nor (n351,n352,n353);
and (n352,n72,n49);
and (n353,n48,n54);
xnor (n354,n355,n73);
nor (n355,n356,n357);
and (n356,n78,n65);
and (n357,n64,n70);
and (n358,n354,n359);
and (n359,n360,n67);
and (n361,n350,n359);
and (n362,n319,n348);
or (n363,n364,n366);
xor (n364,n365,n77);
xor (n365,n45,n61);
xor (n366,n367,n114);
xor (n367,n83,n98);
and (n368,n363,n369);
xor (n369,n370,n372);
xor (n370,n371,n142);
not (n371,n132);
not (n372,n157);
and (n373,n317,n369);
xor (n374,n375,n223);
xor (n375,n214,n218);
and (n376,n374,n377);
xor (n377,n378,n165);
xor (n378,n7,n130);
and (n379,n315,n377);
xor (n380,n381,n210);
xor (n381,n5,n198);
or (n382,n383,n462);
and (n383,n384,n385);
xor (n384,n313,n380);
and (n385,n386,n460);
or (n386,n387,n456,n459);
and (n387,n388,n452);
or (n388,n389,n448,n451);
and (n389,n390,n438);
or (n390,n391,n424,n437);
and (n391,n392,n408);
or (n392,n393,n402,n407);
and (n393,n394,n398);
xnor (n394,n395,n39);
nor (n395,n396,n397);
and (n396,n86,n31);
and (n397,n94,n36);
xnor (n398,n399,n95);
nor (n399,n400,n401);
and (n400,n101,n87);
and (n401,n109,n92);
and (n402,n398,n403);
xnor (n403,n404,n110);
nor (n404,n405,n406);
and (n405,n117,n102);
and (n406,n124,n107);
and (n407,n394,n403);
or (n408,n409,n418,n423);
and (n409,n410,n414);
xnor (n410,n411,n125);
nor (n411,n412,n413);
and (n412,n48,n118);
and (n413,n57,n122);
xnor (n414,n415,n58);
nor (n415,n416,n417);
and (n416,n64,n49);
and (n417,n72,n54);
and (n418,n414,n419);
xnor (n419,n420,n73);
nor (n420,n421,n422);
and (n421,n360,n65);
and (n422,n78,n70);
and (n423,n410,n419);
and (n424,n408,n425);
and (n425,n426,n433);
xnor (n426,n427,n12);
not (n427,n428);
and (n428,n16,n429);
and (n429,n430,n432);
xor (n430,n12,n431);
not (n432,n431);
xnor (n433,n434,n23);
nor (n434,n435,n436);
and (n435,n30,n17);
and (n436,n38,n22);
and (n437,n392,n425);
or (n438,n439,n444,n447);
and (n439,n440,n442);
xor (n440,n441,n330);
xor (n441,n321,n325);
xor (n442,n443,n342);
xor (n443,n12,n337);
and (n444,n442,n445);
xor (n445,n446,n359);
xor (n446,n350,n354);
and (n447,n440,n445);
and (n448,n438,n449);
xor (n449,n450,n27);
xor (n450,n11,n13);
and (n451,n390,n449);
and (n452,n453,n455);
xor (n453,n454,n348);
xor (n454,n319,n335);
xnor (n455,n364,n366);
and (n456,n452,n457);
xor (n457,n458,n81);
xor (n458,n9,n43);
and (n459,n388,n457);
xor (n460,n461,n377);
xor (n461,n315,n374);
and (n462,n463,n464);
xor (n463,n384,n385);
or (n464,n465,n544);
and (n465,n466,n467);
xor (n466,n386,n460);
or (n467,n468,n540,n543);
and (n468,n469,n538);
or (n469,n470,n535,n537);
and (n470,n471,n533);
or (n471,n472,n529,n532);
and (n472,n473,n519);
or (n473,n474,n507,n518);
and (n474,n475,n491);
or (n475,n476,n485,n490);
and (n476,n477,n481);
xnor (n477,n478,n12);
nor (n478,n479,n480);
and (n479,n38,n429);
and (n480,n16,n431);
xnor (n481,n482,n23);
nor (n482,n483,n484);
and (n483,n94,n17);
and (n484,n30,n22);
and (n485,n481,n486);
xnor (n486,n487,n39);
nor (n487,n488,n489);
and (n488,n109,n31);
and (n489,n86,n36);
and (n490,n477,n486);
or (n491,n492,n501,n506);
and (n492,n493,n497);
xnor (n493,n494,n95);
nor (n494,n495,n496);
and (n495,n124,n87);
and (n496,n101,n92);
xnor (n497,n498,n110);
nor (n498,n499,n500);
and (n499,n57,n102);
and (n500,n117,n107);
and (n501,n497,n502);
xnor (n502,n503,n125);
nor (n503,n504,n505);
and (n504,n72,n118);
and (n505,n48,n122);
and (n506,n493,n502);
and (n507,n491,n508);
and (n508,n509,n513);
xnor (n509,n510,n58);
nor (n510,n511,n512);
and (n511,n78,n49);
and (n512,n64,n54);
xnor (n513,n514,n73);
nor (n514,n515,n517);
and (n515,n516,n65);
and (n517,n360,n70);
and (n518,n475,n508);
or (n519,n520,n525,n528);
and (n520,n521,n523);
not (n521,n522);
nand (n522,n516,n67);
xor (n523,n524,n403);
xor (n524,n394,n398);
and (n525,n523,n526);
xor (n526,n527,n419);
xor (n527,n410,n414);
and (n528,n521,n526);
and (n529,n519,n530);
xor (n530,n531,n445);
xor (n531,n440,n442);
and (n532,n473,n530);
xor (n533,n534,n449);
xor (n534,n390,n438);
and (n535,n533,n536);
xor (n536,n453,n455);
and (n537,n471,n536);
xor (n538,n539,n457);
xor (n539,n388,n452);
and (n540,n538,n541);
xor (n541,n542,n369);
xor (n542,n317,n363);
and (n543,n469,n541);
and (n544,n545,n546);
xor (n545,n466,n467);
or (n546,n547,n624);
and (n547,n548,n550);
xor (n548,n549,n541);
xor (n549,n469,n538);
and (n550,n551,n622);
or (n551,n552,n618,n621);
and (n552,n553,n613);
or (n553,n554,n610,n612);
and (n554,n555,n601);
or (n555,n556,n583,n600);
and (n556,n557,n571);
or (n557,n558,n567,n570);
and (n558,n559,n563);
xnor (n559,n560,n125);
nor (n560,n561,n562);
and (n561,n64,n118);
and (n562,n72,n122);
xnor (n563,n564,n58);
nor (n564,n565,n566);
and (n565,n360,n49);
and (n566,n78,n54);
and (n567,n563,n568);
xnor (n568,n569,n73);
nand (n569,n516,n70);
and (n570,n559,n568);
or (n571,n572,n581,n582);
and (n572,n573,n577);
xnor (n573,n574,n12);
nor (n574,n575,n576);
and (n575,n30,n429);
and (n576,n38,n431);
xnor (n577,n578,n23);
nor (n578,n579,n580);
and (n579,n86,n17);
and (n580,n94,n22);
and (n581,n577,n73);
and (n582,n573,n73);
and (n583,n571,n584);
or (n584,n585,n594,n599);
and (n585,n586,n590);
xnor (n586,n587,n39);
nor (n587,n588,n589);
and (n588,n101,n31);
and (n589,n109,n36);
xnor (n590,n591,n95);
nor (n591,n592,n593);
and (n592,n117,n87);
and (n593,n124,n92);
and (n594,n590,n595);
xnor (n595,n596,n110);
nor (n596,n597,n598);
and (n597,n48,n102);
and (n598,n57,n107);
and (n599,n586,n595);
and (n600,n557,n584);
or (n601,n602,n607,n609);
and (n602,n603,n605);
xor (n603,n604,n486);
xor (n604,n477,n481);
xor (n605,n606,n502);
xor (n606,n493,n497);
and (n607,n605,n608);
xor (n608,n509,n513);
and (n609,n603,n608);
and (n610,n601,n611);
xor (n611,n426,n433);
and (n612,n555,n611);
and (n613,n614,n616);
xor (n614,n615,n508);
xor (n615,n475,n491);
xor (n616,n617,n526);
xor (n617,n521,n523);
and (n618,n613,n619);
xor (n619,n620,n425);
xor (n620,n392,n408);
and (n621,n553,n619);
xor (n622,n623,n536);
xor (n623,n471,n533);
and (n624,n625,n626);
xor (n625,n548,n550);
or (n626,n627,n634);
and (n627,n628,n629);
xor (n628,n551,n622);
and (n629,n630,n632);
xor (n630,n631,n619);
xor (n631,n553,n613);
xor (n632,n633,n530);
xor (n633,n473,n519);
and (n634,n635,n636);
xor (n635,n628,n629);
or (n636,n637,n700);
and (n637,n638,n644);
xor (n638,n639,n642);
xor (n639,n619,n640);
xor (n640,n633,n641);
not (n641,n442);
xor (n642,n631,n643);
xnor (n643,n440,n445);
or (n644,n645,n697,n699);
and (n645,n646,n695);
or (n646,n647,n691,n694);
and (n647,n648,n686);
or (n648,n649,n682,n685);
and (n649,n650,n666);
or (n650,n651,n660,n665);
and (n651,n652,n656);
xnor (n652,n653,n12);
nor (n653,n654,n655);
and (n654,n94,n429);
and (n655,n30,n431);
xnor (n656,n657,n23);
nor (n657,n658,n659);
and (n658,n109,n17);
and (n659,n86,n22);
and (n660,n656,n661);
xnor (n661,n662,n39);
nor (n662,n663,n664);
and (n663,n124,n31);
and (n664,n101,n36);
and (n665,n652,n661);
or (n666,n667,n676,n681);
and (n667,n668,n672);
xnor (n668,n669,n95);
nor (n669,n670,n671);
and (n670,n57,n87);
and (n671,n117,n92);
xnor (n672,n673,n110);
nor (n673,n674,n675);
and (n674,n72,n102);
and (n675,n48,n107);
and (n676,n672,n677);
xnor (n677,n678,n125);
nor (n678,n679,n680);
and (n679,n78,n118);
and (n680,n64,n122);
and (n681,n668,n677);
and (n682,n666,n683);
xor (n683,n684,n568);
xor (n684,n559,n563);
and (n685,n650,n683);
and (n686,n687,n689);
xor (n687,n688,n73);
xor (n688,n573,n577);
xor (n689,n690,n595);
xor (n690,n586,n590);
and (n691,n686,n692);
xor (n692,n693,n608);
xor (n693,n603,n605);
and (n694,n648,n692);
xor (n695,n696,n611);
xor (n696,n555,n601);
and (n697,n695,n698);
xor (n698,n614,n616);
and (n699,n646,n698);
and (n700,n701,n702);
xor (n701,n638,n644);
or (n702,n703,n757);
and (n703,n704,n706);
xor (n704,n705,n698);
xor (n705,n646,n695);
or (n706,n707,n753,n756);
and (n707,n708,n751);
or (n708,n709,n748,n750);
and (n709,n710,n746);
or (n710,n711,n740,n745);
and (n711,n712,n724);
or (n712,n713,n722,n723);
and (n713,n714,n718);
xnor (n714,n715,n12);
nor (n715,n716,n717);
and (n716,n86,n429);
and (n717,n94,n431);
xnor (n718,n719,n23);
nor (n719,n720,n721);
and (n720,n101,n17);
and (n721,n109,n22);
and (n722,n718,n58);
and (n723,n714,n58);
or (n724,n725,n734,n739);
and (n725,n726,n730);
xnor (n726,n727,n39);
nor (n727,n728,n729);
and (n728,n117,n31);
and (n729,n124,n36);
xnor (n730,n731,n95);
nor (n731,n732,n733);
and (n732,n48,n87);
and (n733,n57,n92);
and (n734,n730,n735);
xnor (n735,n736,n110);
nor (n736,n737,n738);
and (n737,n64,n102);
and (n738,n72,n107);
and (n739,n726,n735);
and (n740,n724,n741);
xnor (n741,n742,n58);
nor (n742,n743,n744);
and (n743,n516,n49);
and (n744,n360,n54);
and (n745,n712,n741);
xor (n746,n747,n683);
xor (n747,n650,n666);
and (n748,n746,n749);
xor (n749,n687,n689);
and (n750,n710,n749);
xor (n751,n752,n584);
xor (n752,n557,n571);
and (n753,n751,n754);
xor (n754,n755,n692);
xor (n755,n648,n686);
and (n756,n708,n754);
and (n757,n758,n759);
xor (n758,n704,n706);
or (n759,n760,n830);
and (n760,n761,n763);
xor (n761,n762,n754);
xor (n762,n708,n751);
or (n763,n764,n826,n829);
and (n764,n765,n821);
or (n765,n766,n817,n820);
and (n766,n767,n807);
or (n767,n768,n801,n806);
and (n768,n769,n785);
or (n769,n770,n779,n784);
and (n770,n771,n775);
xnor (n771,n772,n95);
nor (n772,n773,n774);
and (n773,n72,n87);
and (n774,n48,n92);
xnor (n775,n776,n110);
nor (n776,n777,n778);
and (n777,n78,n102);
and (n778,n64,n107);
and (n779,n775,n780);
xnor (n780,n781,n125);
nor (n781,n782,n783);
and (n782,n516,n118);
and (n783,n360,n122);
and (n784,n771,n780);
or (n785,n786,n795,n800);
and (n786,n787,n791);
xnor (n787,n788,n12);
nor (n788,n789,n790);
and (n789,n109,n429);
and (n790,n86,n431);
xnor (n791,n792,n23);
nor (n792,n793,n794);
and (n793,n124,n17);
and (n794,n101,n22);
and (n795,n791,n796);
xnor (n796,n797,n39);
nor (n797,n798,n799);
and (n798,n57,n31);
and (n799,n117,n36);
and (n800,n787,n796);
and (n801,n785,n802);
xnor (n802,n803,n125);
nor (n803,n804,n805);
and (n804,n360,n118);
and (n805,n78,n122);
and (n806,n769,n802);
or (n807,n808,n813,n816);
and (n808,n809,n811);
xnor (n809,n810,n58);
nand (n810,n516,n54);
xor (n811,n812,n58);
xor (n812,n714,n718);
and (n813,n811,n814);
xor (n814,n815,n735);
xor (n815,n726,n730);
and (n816,n809,n814);
and (n817,n807,n818);
xor (n818,n819,n677);
xor (n819,n668,n672);
and (n820,n767,n818);
and (n821,n822,n824);
xor (n822,n823,n661);
xor (n823,n652,n656);
xor (n824,n825,n741);
xor (n825,n712,n724);
and (n826,n821,n827);
xor (n827,n828,n749);
xor (n828,n710,n746);
and (n829,n765,n827);
and (n830,n831,n832);
xor (n831,n761,n763);
or (n832,n833,n885);
and (n833,n834,n836);
xor (n834,n835,n827);
xor (n835,n765,n821);
or (n836,n837,n882,n884);
and (n837,n838,n880);
or (n838,n839,n876,n879);
and (n839,n840,n874);
or (n840,n841,n870,n873);
and (n841,n842,n858);
or (n842,n843,n852,n857);
and (n843,n844,n848);
xnor (n844,n845,n39);
nor (n845,n846,n847);
and (n846,n48,n31);
and (n847,n57,n36);
xnor (n848,n849,n95);
nor (n849,n850,n851);
and (n850,n64,n87);
and (n851,n72,n92);
and (n852,n848,n853);
xnor (n853,n854,n110);
nor (n854,n855,n856);
and (n855,n360,n102);
and (n856,n78,n107);
and (n857,n844,n853);
or (n858,n859,n868,n869);
and (n859,n860,n864);
xnor (n860,n861,n12);
nor (n861,n862,n863);
and (n862,n101,n429);
and (n863,n109,n431);
xnor (n864,n865,n23);
nor (n865,n866,n867);
and (n866,n117,n17);
and (n867,n124,n22);
and (n868,n864,n125);
and (n869,n860,n125);
and (n870,n858,n871);
xor (n871,n872,n780);
xor (n872,n771,n775);
and (n873,n842,n871);
xor (n874,n875,n802);
xor (n875,n769,n785);
and (n876,n874,n877);
xor (n877,n878,n814);
xor (n878,n809,n811);
and (n879,n840,n877);
xor (n880,n881,n818);
xor (n881,n767,n807);
and (n882,n880,n883);
xor (n883,n822,n824);
and (n884,n838,n883);
and (n885,n886,n887);
xor (n886,n834,n836);
or (n887,n888,n926);
and (n888,n889,n891);
xor (n889,n890,n883);
xor (n890,n838,n880);
and (n891,n892,n924);
or (n892,n893,n920,n923);
and (n893,n894,n918);
or (n894,n895,n914,n917);
and (n895,n896,n912);
or (n896,n897,n906,n911);
and (n897,n898,n902);
xnor (n898,n899,n12);
nor (n899,n900,n901);
and (n900,n124,n429);
and (n901,n101,n431);
xnor (n902,n903,n23);
nor (n903,n904,n905);
and (n904,n57,n17);
and (n905,n117,n22);
and (n906,n902,n907);
xnor (n907,n908,n39);
nor (n908,n909,n910);
and (n909,n72,n31);
and (n910,n48,n36);
and (n911,n898,n907);
xnor (n912,n913,n125);
nand (n913,n516,n122);
and (n914,n912,n915);
xor (n915,n916,n853);
xor (n916,n844,n848);
and (n917,n896,n915);
xor (n918,n919,n796);
xor (n919,n787,n791);
and (n920,n918,n921);
xor (n921,n922,n871);
xor (n922,n842,n858);
and (n923,n894,n921);
xor (n924,n925,n877);
xor (n925,n840,n874);
and (n926,n927,n928);
xor (n927,n889,n891);
or (n928,n929,n981);
and (n929,n930,n931);
xor (n930,n892,n924);
and (n931,n932,n979);
or (n932,n933,n975,n978);
and (n933,n934,n968);
or (n934,n935,n962,n967);
and (n935,n936,n950);
or (n936,n937,n946,n949);
and (n937,n938,n942);
xnor (n938,n939,n39);
nor (n939,n940,n941);
and (n940,n64,n31);
and (n941,n72,n36);
xnor (n942,n943,n95);
nor (n943,n944,n945);
and (n944,n360,n87);
and (n945,n78,n92);
and (n946,n942,n947);
xnor (n947,n948,n110);
nand (n948,n516,n107);
and (n949,n938,n947);
or (n950,n951,n960,n961);
and (n951,n952,n956);
xnor (n952,n953,n12);
nor (n953,n954,n955);
and (n954,n117,n429);
and (n955,n124,n431);
xnor (n956,n957,n23);
nor (n957,n958,n959);
and (n958,n48,n17);
and (n959,n57,n22);
and (n960,n956,n110);
and (n961,n952,n110);
and (n962,n950,n963);
xnor (n963,n964,n95);
nor (n964,n965,n966);
and (n965,n78,n87);
and (n966,n64,n92);
and (n967,n936,n963);
and (n968,n969,n973);
xnor (n969,n970,n110);
nor (n970,n971,n972);
and (n971,n516,n102);
and (n972,n360,n107);
xor (n973,n974,n907);
xor (n974,n898,n902);
and (n975,n968,n976);
xor (n976,n977,n125);
xor (n977,n860,n864);
and (n978,n934,n976);
xor (n979,n980,n921);
xor (n980,n894,n918);
and (n981,n982,n983);
xor (n982,n930,n931);
or (n983,n984,n991);
and (n984,n985,n986);
xor (n985,n932,n979);
and (n986,n987,n989);
xor (n987,n988,n915);
xor (n988,n896,n912);
xor (n989,n990,n976);
xor (n990,n934,n968);
and (n991,n992,n993);
xor (n992,n985,n986);
or (n993,n994,n1027);
and (n994,n995,n996);
xor (n995,n987,n989);
or (n996,n997,n1024,n1026);
and (n997,n998,n1022);
or (n998,n999,n1018,n1021);
and (n999,n1000,n1016);
or (n1000,n1001,n1010,n1015);
and (n1001,n1002,n1006);
xnor (n1002,n1003,n12);
nor (n1003,n1004,n1005);
and (n1004,n57,n429);
and (n1005,n117,n431);
xnor (n1006,n1007,n23);
nor (n1007,n1008,n1009);
and (n1008,n72,n17);
and (n1009,n48,n22);
and (n1010,n1006,n1011);
xnor (n1011,n1012,n39);
nor (n1012,n1013,n1014);
and (n1013,n78,n31);
and (n1014,n64,n36);
and (n1015,n1002,n1011);
xor (n1016,n1017,n947);
xor (n1017,n938,n942);
and (n1018,n1016,n1019);
xor (n1019,n1020,n110);
xor (n1020,n952,n956);
and (n1021,n1000,n1019);
xor (n1022,n1023,n963);
xor (n1023,n936,n950);
and (n1024,n1022,n1025);
xor (n1025,n969,n973);
and (n1026,n998,n1025);
and (n1027,n1028,n1029);
xor (n1028,n995,n996);
or (n1029,n1030,n1063);
and (n1030,n1031,n1033);
xor (n1031,n1032,n1025);
xor (n1032,n998,n1022);
and (n1033,n1034,n1061);
or (n1034,n1035,n1055,n1060);
and (n1035,n1036,n1048);
or (n1036,n1037,n1046,n1047);
and (n1037,n1038,n1042);
xnor (n1038,n1039,n12);
nor (n1039,n1040,n1041);
and (n1040,n48,n429);
and (n1041,n57,n431);
xnor (n1042,n1043,n23);
nor (n1043,n1044,n1045);
and (n1044,n64,n17);
and (n1045,n72,n22);
and (n1046,n1042,n95);
and (n1047,n1038,n95);
and (n1048,n1049,n1053);
xnor (n1049,n1050,n39);
nor (n1050,n1051,n1052);
and (n1051,n360,n31);
and (n1052,n78,n36);
xnor (n1053,n1054,n95);
nand (n1054,n516,n92);
and (n1055,n1048,n1056);
xnor (n1056,n1057,n95);
nor (n1057,n1058,n1059);
and (n1058,n516,n87);
and (n1059,n360,n92);
and (n1060,n1036,n1056);
xor (n1061,n1062,n1019);
xor (n1062,n1000,n1016);
and (n1063,n1064,n1065);
xor (n1064,n1031,n1033);
or (n1065,n1066,n1073);
and (n1066,n1067,n1068);
xor (n1067,n1034,n1061);
and (n1068,n1069,n1071);
xor (n1069,n1070,n1011);
xor (n1070,n1002,n1006);
xor (n1071,n1072,n1056);
xor (n1072,n1036,n1048);
and (n1073,n1074,n1075);
xor (n1074,n1067,n1068);
or (n1075,n1076,n1101);
and (n1076,n1077,n1078);
xor (n1077,n1069,n1071);
or (n1078,n1079,n1098,n1100);
and (n1079,n1080,n1096);
or (n1080,n1081,n1090,n1095);
and (n1081,n1082,n1086);
xnor (n1082,n1083,n12);
nor (n1083,n1084,n1085);
and (n1084,n72,n429);
and (n1085,n48,n431);
xnor (n1086,n1087,n23);
nor (n1087,n1088,n1089);
and (n1088,n78,n17);
and (n1089,n64,n22);
and (n1090,n1086,n1091);
xnor (n1091,n1092,n39);
nor (n1092,n1093,n1094);
and (n1093,n516,n31);
and (n1094,n360,n36);
and (n1095,n1082,n1091);
xor (n1096,n1097,n95);
xor (n1097,n1038,n1042);
and (n1098,n1096,n1099);
xor (n1099,n1049,n1053);
and (n1100,n1080,n1099);
and (n1101,n1102,n1103);
xor (n1102,n1077,n1078);
or (n1103,n1104,n1122);
and (n1104,n1105,n1107);
xor (n1105,n1106,n1099);
xor (n1106,n1080,n1096);
and (n1107,n1108,n1120);
or (n1108,n1109,n1118,n1119);
and (n1109,n1110,n1114);
xnor (n1110,n1111,n12);
nor (n1111,n1112,n1113);
and (n1112,n64,n429);
and (n1113,n72,n431);
xnor (n1114,n1115,n23);
nor (n1115,n1116,n1117);
and (n1116,n360,n17);
and (n1117,n78,n22);
and (n1118,n1114,n39);
and (n1119,n1110,n39);
xor (n1120,n1121,n1091);
xor (n1121,n1082,n1086);
and (n1122,n1123,n1124);
xor (n1123,n1105,n1107);
or (n1124,n1125,n1132);
and (n1125,n1126,n1127);
xor (n1126,n1108,n1120);
and (n1127,n1128,n1130);
xnor (n1128,n1129,n39);
nand (n1129,n516,n36);
xor (n1130,n1131,n39);
xor (n1131,n1110,n1114);
and (n1132,n1133,n1134);
xor (n1133,n1126,n1127);
or (n1134,n1135,n1146);
and (n1135,n1136,n1137);
xor (n1136,n1128,n1130);
and (n1137,n1138,n1142);
xnor (n1138,n1139,n12);
nor (n1139,n1140,n1141);
and (n1140,n78,n429);
and (n1141,n64,n431);
xnor (n1142,n1143,n23);
nor (n1143,n1144,n1145);
and (n1144,n516,n17);
and (n1145,n360,n22);
and (n1146,n1147,n1148);
xor (n1147,n1136,n1137);
or (n1148,n1149,n1156);
and (n1149,n1150,n1151);
xor (n1150,n1138,n1142);
and (n1151,n1152,n23);
xnor (n1152,n1153,n12);
nor (n1153,n1154,n1155);
and (n1154,n360,n429);
and (n1155,n78,n431);
and (n1156,n1157,n1158);
xor (n1157,n1150,n1151);
or (n1158,n1159,n1163);
and (n1159,n1160,n1162);
xnor (n1160,n1161,n23);
nand (n1161,n516,n22);
xor (n1162,n1152,n23);
and (n1163,n1164,n1165);
xor (n1164,n1160,n1162);
and (n1165,n1166,n1170);
xnor (n1166,n1167,n12);
nor (n1167,n1168,n1169);
and (n1168,n516,n429);
and (n1169,n360,n431);
and (n1170,n1171,n12);
xnor (n1171,n1172,n12);
nand (n1172,n516,n431);
xor (n1173,n1174,n1283);
xor (n1174,n1175,n1253);
xor (n1175,n1176,n1228);
or (n1176,n1177,n1212,n1227);
and (n1177,n1178,n1204);
or (n1178,n1179,n1195,n1203);
and (n1179,n1180,n1191);
or (n1180,n1181,n1188,n1190);
and (n1181,n1182,n1185);
or (n1182,n26,n1183,n1184);
and (n1183,n27,n83);
and (n1184,n13,n83);
or (n1185,n113,n1186,n1187);
and (n1186,n114,n45);
and (n1187,n98,n45);
and (n1188,n1185,n1189);
or (n1189,n61,n77);
and (n1190,n1182,n1189);
or (n1191,n1192,n1193,n1194);
and (n1192,n371,n142);
and (n1193,n142,n372);
and (n1194,n371,n372);
and (n1195,n1191,n1196);
xor (n1196,n1197,n1202);
xor (n1197,n1198,n1200);
xor (n1198,n1199,n179);
xor (n1199,n170,n173);
xor (n1200,n1201,n192);
xor (n1201,n183,n187);
not (n1202,n196);
and (n1203,n1180,n1196);
xor (n1204,n1205,n196);
xor (n1205,n1206,n1209);
or (n1206,n202,n1207,n1208);
and (n1207,n173,n179);
and (n1208,n170,n179);
or (n1209,n206,n1210,n1211);
and (n1210,n187,n192);
and (n1211,n183,n192);
and (n1212,n1204,n1213);
xor (n1213,n1214,n229);
xor (n1214,n1215,n1223);
or (n1215,n1216,n1220,n1222);
and (n1216,n1217,n218);
or (n1217,n1218,n216,n1219);
and (n1218,n169,n134);
and (n1219,n169,n138);
and (n1220,n218,n1221);
and (n1221,n158,n162);
and (n1222,n1217,n1221);
or (n1223,n1224,n1225,n1226);
and (n1224,n1198,n1200);
and (n1225,n1200,n1202);
and (n1226,n1198,n1202);
and (n1227,n1178,n1213);
xor (n1228,n1229,n1246);
xor (n1229,n1230,n1234);
or (n1230,n1231,n1232,n1233);
and (n1231,n1215,n1223);
and (n1232,n1223,n229);
and (n1233,n1215,n229);
xor (n1234,n1235,n1244);
xor (n1235,n1236,n1240);
or (n1236,n1237,n1238,n1239);
and (n1237,n1206,n1209);
and (n1238,n1209,n196);
and (n1239,n1206,n196);
or (n1240,n1241,n1242,n1243);
and (n1241,n231,n232);
and (n1242,n232,n243);
and (n1243,n231,n243);
xor (n1244,n1245,n287);
xor (n1245,n294,n298);
xor (n1246,n1247,n1249);
xor (n1247,n1248,n290);
xor (n1248,n305,n308);
xnor (n1249,n1250,n270);
or (n1250,n1251,n268,n1252);
and (n1251,n304,n235);
and (n1252,n304,n239);
and (n1253,n1254,n1281);
or (n1254,n1255,n1277,n1280);
and (n1255,n1256,n1275);
or (n1256,n1257,n1273,n1274);
and (n1257,n1258,n1264);
or (n1258,n1259,n1263,n362);
and (n1259,n319,n1260);
or (n1260,n1261,n341,n1262);
and (n1261,n11,n337);
and (n1262,n11,n342);
and (n1263,n1260,n348);
or (n1264,n1265,n1270,n1272);
and (n1265,n1266,n1268);
xor (n1266,n1267,n83);
xor (n1267,n13,n27);
xor (n1268,n1269,n45);
xor (n1269,n98,n114);
and (n1270,n1268,n1271);
xnor (n1271,n61,n77);
and (n1272,n1266,n1271);
and (n1273,n1264,n369);
and (n1274,n1258,n369);
xor (n1275,n1276,n1221);
xor (n1276,n1217,n218);
and (n1277,n1275,n1278);
xor (n1278,n1279,n1196);
xor (n1279,n1180,n1191);
and (n1280,n1256,n1278);
xor (n1281,n1282,n1213);
xor (n1282,n1178,n1204);
or (n1283,n1284,n1304);
and (n1284,n1285,n1286);
xor (n1285,n1254,n1281);
and (n1286,n1287,n1302);
or (n1287,n1288,n1298,n1301);
and (n1288,n1289,n1296);
or (n1289,n1290,n1292,n1295);
and (n1290,n390,n1291);
or (n1291,n440,n445);
and (n1292,n1291,n1293);
xor (n1293,n1294,n1271);
xor (n1294,n1266,n1268);
and (n1295,n390,n1293);
xor (n1296,n1297,n1189);
xor (n1297,n1182,n1185);
and (n1298,n1296,n1299);
xor (n1299,n1300,n369);
xor (n1300,n1258,n1264);
and (n1301,n1289,n1299);
xor (n1302,n1303,n1278);
xor (n1303,n1256,n1275);
and (n1304,n1305,n1306);
xor (n1305,n1285,n1286);
or (n1306,n1307,n1323);
and (n1307,n1308,n1309);
xor (n1308,n1287,n1302);
and (n1309,n1310,n1321);
or (n1310,n1311,n1317,n1320);
and (n1311,n1312,n1315);
or (n1312,n472,n1313,n1314);
and (n1313,n519,n641);
and (n1314,n473,n641);
xor (n1315,n1316,n348);
xor (n1316,n319,n1260);
and (n1317,n1315,n1318);
xor (n1318,n1319,n1293);
xor (n1319,n390,n1291);
and (n1320,n1312,n1318);
xor (n1321,n1322,n1299);
xor (n1322,n1289,n1296);
and (n1323,n1324,n1325);
xor (n1324,n1308,n1309);
or (n1325,n1326,n1334);
and (n1326,n1327,n1328);
xor (n1327,n1310,n1321);
and (n1328,n1329,n1332);
or (n1329,n552,n1330,n1331);
and (n1330,n613,n643);
and (n1331,n553,n643);
xor (n1332,n1333,n1318);
xor (n1333,n1312,n1315);
and (n1334,n1335,n1336);
xor (n1335,n1327,n1328);
or (n1336,n1337,n634);
and (n1337,n1338,n1339);
xor (n1338,n1329,n1332);
or (n1339,n1340,n1341,n1342);
and (n1340,n619,n640);
and (n1341,n640,n642);
and (n1342,n619,n642);
endmodule
