module top (out,n20,n22,n26,n32,n38,n47,n49,n54,n58
        ,n65,n75,n80,n84,n90,n100,n102,n109,n111,n121
        ,n128,n130,n136,n140,n146,n155,n156,n162,n166,n174
        ,n185,n194,n199,n208,n210,n218,n224,n234,n241,n247
        ,n260,n266,n274,n281,n312,n331,n333,n341,n356,n373
        ,n378,n386,n412,n429,n469,n565,n570,n574,n580,n712
        ,n753,n922,n942,n959,n1122);
output out;
input n20;
input n22;
input n26;
input n32;
input n38;
input n47;
input n49;
input n54;
input n58;
input n65;
input n75;
input n80;
input n84;
input n90;
input n100;
input n102;
input n109;
input n111;
input n121;
input n128;
input n130;
input n136;
input n140;
input n146;
input n155;
input n156;
input n162;
input n166;
input n174;
input n185;
input n194;
input n199;
input n208;
input n210;
input n218;
input n224;
input n234;
input n241;
input n247;
input n260;
input n266;
input n274;
input n281;
input n312;
input n331;
input n333;
input n341;
input n356;
input n373;
input n378;
input n386;
input n412;
input n429;
input n469;
input n565;
input n570;
input n574;
input n580;
input n712;
input n753;
input n922;
input n942;
input n959;
input n1122;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n332;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n374;
wire n375;
wire n376;
wire n377;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n566;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
xor (out,n0,n4242);
nand (n0,n1,n4241);
or (n1,n2,n1086);
not (n2,n3);
nand (n3,n4,n1085);
not (n4,n5);
nor (n5,n6,n1000);
xor (n6,n7,n891);
xor (n7,n8,n632);
xor (n8,n9,n551);
xor (n9,n10,n250);
xor (n10,n11,n176);
xor (n11,n12,n93);
xor (n12,n13,n68);
xor (n13,n14,n41);
nand (n14,n15,n35);
or (n15,n16,n29);
nand (n16,n17,n24);
not (n17,n18);
nand (n18,n19,n23);
or (n19,n20,n21);
not (n21,n22);
nand (n23,n21,n20);
nand (n24,n25,n28);
or (n25,n26,n27);
not (n27,n20);
nand (n28,n26,n27);
nor (n29,n30,n33);
and (n30,n31,n32);
not (n31,n26);
and (n33,n26,n34);
not (n34,n32);
or (n35,n17,n36);
nor (n36,n37,n39);
and (n37,n31,n38);
and (n39,n26,n40);
not (n40,n38);
nand (n41,n42,n61);
or (n42,n43,n56);
not (n43,n44);
nor (n44,n45,n51);
nand (n45,n46,n50);
or (n46,n47,n48);
not (n48,n49);
nand (n50,n47,n48);
nor (n51,n52,n55);
and (n52,n49,n53);
not (n53,n54);
and (n55,n54,n48);
nor (n56,n57,n59);
and (n57,n53,n58);
and (n59,n54,n60);
not (n60,n58);
or (n61,n62,n63);
not (n62,n45);
nor (n63,n64,n66);
and (n64,n53,n65);
and (n66,n54,n67);
not (n67,n65);
nand (n68,n69,n87);
or (n69,n70,n82);
not (n70,n71);
and (n71,n72,n77);
and (n72,n73,n76);
nand (n73,n54,n74);
not (n74,n75);
nand (n76,n75,n53);
nor (n77,n78,n81);
and (n78,n74,n79);
not (n79,n80);
and (n81,n75,n80);
nor (n82,n83,n85);
and (n83,n79,n84);
and (n85,n80,n86);
not (n86,n84);
or (n87,n72,n88);
nor (n88,n89,n91);
and (n89,n79,n90);
and (n91,n80,n92);
not (n92,n90);
xor (n93,n94,n149);
xor (n94,n95,n123);
nand (n95,n96,n117);
or (n96,n97,n105);
not (n97,n98);
nand (n98,n99,n103);
or (n99,n100,n101);
not (n101,n102);
or (n103,n104,n102);
not (n104,n100);
not (n105,n106);
nor (n106,n107,n113);
nand (n107,n108,n112);
or (n108,n109,n110);
not (n110,n111);
nand (n112,n109,n110);
nor (n113,n114,n115);
and (n114,n104,n109);
and (n115,n100,n116);
not (n116,n109);
nand (n117,n107,n118);
nand (n118,n119,n122);
or (n119,n100,n120);
not (n120,n121);
or (n122,n104,n121);
nand (n123,n124,n143);
or (n124,n125,n138);
nand (n125,n126,n133);
and (n126,n127,n131);
nand (n127,n128,n129);
not (n129,n130);
nand (n131,n130,n132);
not (n132,n128);
nand (n133,n134,n137);
or (n134,n130,n135);
not (n135,n136);
nand (n137,n130,n135);
nor (n138,n139,n141);
and (n139,n135,n140);
and (n141,n136,n142);
not (n142,n140);
or (n143,n126,n144);
nor (n144,n145,n147);
and (n145,n135,n146);
and (n147,n136,n148);
not (n148,n146);
nand (n149,n150,n169);
or (n150,n151,n164);
nand (n151,n152,n159);
nor (n152,n153,n157);
and (n153,n154,n156);
not (n154,n155);
and (n157,n155,n158);
not (n158,n156);
nor (n159,n160,n163);
and (n160,n158,n161);
not (n161,n162);
and (n163,n156,n162);
nor (n164,n165,n167);
and (n165,n166,n161);
and (n167,n168,n162);
not (n168,n166);
or (n169,n152,n170);
not (n170,n171);
nand (n171,n172,n175);
or (n172,n173,n162);
not (n173,n174);
or (n175,n161,n174);
xor (n176,n177,n228);
xor (n177,n178,n202);
nand (n178,n179,n196);
or (n179,n180,n191);
nand (n180,n181,n187);
not (n181,n182);
nor (n182,n183,n186);
and (n183,n184,n128);
not (n184,n185);
and (n186,n185,n132);
not (n187,n188);
nand (n188,n189,n190);
or (n189,n31,n185);
nand (n190,n185,n31);
nor (n191,n192,n195);
and (n192,n193,n128);
not (n193,n194);
and (n195,n194,n132);
or (n196,n187,n197);
nor (n197,n198,n200);
and (n198,n132,n199);
and (n200,n128,n201);
not (n201,n199);
nand (n202,n203,n221);
or (n203,n204,n215);
not (n204,n205);
nor (n205,n206,n212);
nor (n206,n207,n211);
and (n207,n208,n209);
not (n209,n210);
nor (n211,n208,n209);
nand (n212,n213,n214);
or (n213,n209,n80);
nand (n214,n80,n209);
nor (n215,n216,n219);
and (n216,n217,n218);
not (n217,n208);
and (n219,n208,n220);
not (n220,n218);
or (n221,n222,n227);
nor (n222,n223,n225);
and (n223,n217,n224);
and (n225,n208,n226);
not (n226,n224);
not (n227,n212);
nand (n228,n229,n244);
or (n229,n230,n239);
nand (n230,n231,n236);
nor (n231,n232,n235);
and (n232,n233,n208);
not (n233,n234);
and (n235,n234,n217);
nand (n236,n237,n238);
or (n237,n234,n154);
nand (n238,n154,n234);
nor (n239,n240,n242);
and (n240,n154,n241);
and (n242,n155,n243);
not (n243,n241);
or (n244,n231,n245);
nor (n245,n246,n248);
and (n246,n154,n247);
and (n248,n155,n249);
not (n249,n247);
or (n250,n251,n550);
and (n251,n252,n475);
xor (n252,n253,n320);
or (n253,n254,n319);
and (n254,n255,n284);
xor (n255,n256,n269);
nand (n256,n257,n263);
or (n257,n125,n258);
nor (n258,n259,n261);
and (n259,n135,n260);
and (n261,n136,n262);
not (n262,n260);
or (n263,n126,n264);
nor (n264,n265,n267);
and (n265,n135,n266);
and (n267,n136,n268);
not (n268,n266);
not (n269,n270);
nand (n270,n271,n277);
or (n271,n105,n272);
nor (n272,n273,n275);
and (n273,n104,n274);
and (n275,n100,n276);
not (n276,n274);
or (n277,n278,n279);
not (n278,n107);
nor (n279,n280,n282);
and (n280,n104,n281);
and (n282,n100,n283);
not (n283,n281);
or (n284,n285,n318);
and (n285,n286,n306);
xor (n286,n287,n296);
nand (n287,n288,n292);
or (n288,n16,n289);
nor (n289,n290,n291);
and (n290,n146,n31);
and (n291,n26,n148);
or (n292,n17,n293);
nor (n293,n294,n295);
and (n294,n193,n26);
and (n295,n194,n31);
nand (n296,n297,n302);
or (n297,n298,n204);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n173,n217);
and (n301,n174,n208);
nand (n302,n303,n212);
nor (n303,n304,n305);
and (n304,n243,n217);
and (n305,n241,n208);
nand (n306,n307,n314);
or (n307,n230,n308);
not (n308,n309);
nand (n309,n310,n313);
or (n310,n311,n155);
not (n311,n312);
or (n313,n154,n312);
or (n314,n231,n315);
nor (n315,n316,n317);
and (n316,n154,n166);
and (n317,n155,n168);
and (n318,n287,n296);
and (n319,n256,n269);
or (n320,n321,n474);
and (n321,n322,n444);
xor (n322,n323,n390);
or (n323,n324,n389);
and (n324,n325,n367);
xor (n325,n326,n346);
nand (n326,n327,n343);
or (n327,n328,n336);
not (n328,n329);
nor (n329,n330,n334);
and (n330,n331,n332);
not (n332,n333);
and (n334,n335,n333);
not (n335,n331);
not (n336,n337);
nand (n337,n329,n338);
nand (n338,n339,n342);
or (n339,n333,n340);
not (n340,n341);
nand (n342,n340,n333);
nor (n343,n344,n345);
and (n344,n121,n341);
and (n345,n120,n340);
nand (n346,n347,n362);
or (n347,n348,n352);
not (n348,n349);
nor (n349,n350,n351);
and (n350,n281,n111);
and (n351,n283,n110);
not (n352,n353);
nor (n353,n354,n359);
nand (n354,n355,n357);
or (n355,n356,n340);
or (n357,n341,n358);
not (n358,n356);
nor (n359,n360,n361);
and (n360,n110,n356);
and (n361,n111,n358);
nand (n362,n363,n354);
not (n363,n364);
nor (n364,n365,n366);
and (n365,n101,n111);
and (n366,n102,n110);
nand (n367,n368,n383);
or (n368,n369,n380);
nand (n369,n370,n375);
and (n370,n371,n374);
nand (n371,n100,n372);
not (n372,n373);
nand (n374,n373,n104);
nand (n375,n376,n379);
or (n376,n373,n377);
not (n377,n378);
nand (n379,n377,n373);
nor (n380,n381,n382);
and (n381,n377,n38);
and (n382,n378,n40);
or (n383,n370,n384);
nor (n384,n385,n387);
and (n385,n377,n386);
and (n387,n378,n388);
not (n388,n386);
and (n389,n326,n346);
or (n390,n391,n443);
and (n391,n392,n423);
xor (n392,n393,n401);
nand (n393,n394,n395);
or (n394,n126,n258);
nand (n395,n396,n400);
not (n396,n397);
nor (n397,n398,n399);
and (n398,n135,n65);
and (n399,n136,n67);
not (n400,n125);
nand (n401,n402,n418);
or (n402,n403,n408);
not (n403,n404);
nand (n404,n405,n406);
or (n405,n47,n92);
or (n406,n407,n90);
not (n407,n47);
nand (n408,n409,n415);
not (n409,n410);
nor (n410,n411,n413);
and (n411,n407,n412);
and (n413,n47,n414);
not (n414,n412);
and (n415,n416,n417);
nand (n416,n136,n414);
nand (n417,n135,n412);
nand (n418,n419,n420);
not (n419,n415);
nand (n420,n421,n422);
or (n421,n47,n60);
or (n422,n407,n58);
nand (n423,n424,n439);
or (n424,n425,n436);
not (n425,n426);
nor (n426,n427,n432);
nor (n427,n428,n430);
and (n428,n21,n429);
and (n430,n22,n431);
not (n431,n429);
not (n432,n433);
nor (n433,n434,n435);
and (n434,n377,n429);
and (n435,n378,n431);
nor (n436,n437,n438);
and (n437,n21,n199);
and (n438,n22,n201);
or (n439,n433,n440);
nor (n440,n441,n442);
and (n441,n21,n32);
and (n442,n22,n34);
and (n443,n393,n401);
or (n444,n445,n473);
and (n445,n446,n465);
xor (n446,n447,n456);
nand (n447,n448,n452);
or (n448,n43,n449);
nor (n449,n450,n451);
and (n450,n53,n224);
and (n451,n54,n226);
or (n452,n62,n453);
nor (n453,n454,n455);
and (n454,n53,n84);
and (n455,n54,n86);
nand (n456,n457,n461);
or (n457,n70,n458);
nor (n458,n459,n460);
and (n459,n247,n79);
and (n460,n80,n249);
or (n461,n72,n462);
nor (n462,n463,n464);
and (n463,n79,n218);
and (n464,n80,n220);
nand (n465,n466,n472);
or (n466,n105,n467);
nor (n467,n468,n470);
and (n468,n104,n469);
and (n470,n100,n471);
not (n471,n469);
or (n472,n278,n272);
and (n473,n447,n456);
and (n474,n323,n390);
xor (n475,n476,n524);
xor (n476,n477,n501);
or (n477,n478,n500);
and (n478,n479,n494);
xor (n479,n480,n486);
nand (n480,n481,n482);
or (n481,n425,n440);
or (n482,n433,n483);
nor (n483,n484,n485);
and (n484,n21,n38);
and (n485,n22,n40);
nand (n486,n487,n489);
or (n487,n488,n408);
not (n488,n420);
nand (n489,n490,n419);
not (n490,n491);
nor (n491,n492,n493);
and (n492,n407,n65);
and (n493,n47,n67);
nand (n494,n495,n496);
or (n495,n43,n453);
or (n496,n62,n497);
nor (n497,n498,n499);
and (n498,n53,n90);
and (n499,n54,n92);
and (n500,n480,n486);
or (n501,n502,n523);
and (n502,n503,n516);
xor (n503,n504,n510);
nand (n504,n505,n506);
or (n505,n16,n293);
or (n506,n17,n507);
nor (n507,n508,n509);
and (n508,n31,n199);
and (n509,n26,n201);
nand (n510,n511,n512);
or (n511,n70,n462);
or (n512,n72,n513);
nor (n513,n514,n515);
and (n514,n79,n224);
and (n515,n80,n226);
nand (n516,n517,n519);
or (n517,n204,n518);
not (n518,n303);
or (n519,n520,n227);
nor (n520,n521,n522);
and (n521,n217,n247);
and (n522,n208,n249);
and (n523,n504,n510);
or (n524,n525,n549);
and (n525,n526,n543);
xor (n526,n527,n534);
nand (n527,n528,n529);
or (n528,n352,n364);
or (n529,n530,n531);
not (n530,n354);
nor (n531,n532,n533);
and (n532,n110,n121);
and (n533,n111,n120);
nand (n534,n535,n539);
or (n535,n180,n536);
nor (n536,n537,n538);
and (n537,n132,n140);
and (n538,n128,n142);
or (n539,n187,n540);
nor (n540,n541,n542);
and (n541,n132,n146);
and (n542,n128,n148);
nand (n543,n544,n545);
or (n544,n230,n315);
or (n545,n231,n546);
nor (n546,n547,n548);
and (n547,n154,n174);
and (n548,n155,n173);
and (n549,n527,n534);
and (n550,n253,n320);
xor (n551,n552,n587);
xor (n552,n553,n584);
or (n553,n554,n583);
and (n554,n555,n270);
xor (n555,n556,n559);
nand (n556,n557,n558);
or (n557,n125,n264);
or (n558,n126,n138);
nand (n559,n560,n577);
or (n560,n561,n572);
nand (n561,n562,n567);
not (n562,n563);
nand (n563,n564,n566);
or (n564,n161,n565);
nand (n566,n565,n161);
nand (n567,n568,n571);
or (n568,n569,n565);
not (n569,n570);
nand (n571,n569,n565);
nor (n572,n573,n575);
and (n573,n569,n574);
and (n575,n576,n570);
not (n576,n574);
or (n577,n562,n578);
nor (n578,n579,n581);
and (n579,n580,n569);
and (n581,n582,n570);
not (n582,n580);
and (n583,n556,n559);
or (n584,n585,n586);
and (n585,n476,n524);
and (n586,n477,n501);
xor (n587,n588,n616);
xor (n588,n589,n600);
not (n589,n590);
nand (n590,n591,n596);
or (n591,n592,n369);
not (n592,n593);
nand (n593,n594,n595);
or (n594,n378,n276);
or (n595,n377,n274);
or (n596,n370,n597);
nor (n597,n598,n599);
and (n598,n377,n281);
and (n599,n378,n283);
or (n600,n601,n615);
and (n601,n602,n612);
xor (n602,n603,n609);
nand (n603,n604,n605);
or (n604,n408,n491);
or (n605,n415,n606);
nor (n606,n607,n608);
and (n607,n407,n260);
and (n608,n47,n262);
nand (n609,n610,n611);
or (n610,n43,n497);
or (n611,n62,n56);
nand (n612,n613,n614);
or (n613,n16,n507);
or (n614,n17,n29);
and (n615,n603,n609);
or (n616,n617,n631);
and (n617,n618,n625);
xor (n618,n619,n622);
nand (n619,n620,n621);
or (n620,n70,n513);
or (n621,n72,n82);
nand (n622,n623,n624);
or (n623,n204,n520);
or (n624,n227,n215);
nand (n625,n626,n627);
or (n626,n592,n370);
or (n627,n369,n628);
nor (n628,n629,n630);
and (n629,n377,n469);
and (n630,n378,n471);
and (n631,n619,n622);
xor (n632,n633,n764);
xor (n633,n634,n727);
xor (n634,n635,n720);
xor (n635,n636,n691);
xor (n636,n637,n671);
xor (n637,n638,n655);
or (n638,n639,n654);
and (n639,n640,n648);
xor (n640,n641,n645);
nand (n641,n642,n643);
or (n642,n540,n180);
nand (n643,n644,n188);
not (n644,n191);
nand (n645,n646,n647);
or (n646,n230,n546);
or (n647,n231,n239);
nand (n648,n649,n653);
or (n649,n151,n650);
nor (n650,n651,n652);
and (n651,n312,n161);
and (n652,n162,n311);
or (n653,n152,n164);
and (n654,n641,n645);
or (n655,n656,n670);
and (n656,n657,n664);
xor (n657,n658,n661);
nand (n658,n659,n660);
or (n659,n353,n354);
not (n660,n531);
nand (n661,n662,n663);
or (n662,n105,n279);
or (n663,n278,n97);
nand (n664,n665,n666);
or (n665,n425,n483);
or (n666,n433,n667);
nor (n667,n668,n669);
and (n668,n21,n386);
and (n669,n22,n388);
and (n670,n658,n661);
xor (n671,n672,n685);
xor (n672,n673,n679);
nand (n673,n674,n675);
or (n674,n561,n578);
or (n675,n562,n676);
nor (n676,n677,n678);
and (n677,n312,n569);
and (n678,n311,n570);
nand (n679,n680,n681);
or (n680,n425,n667);
or (n681,n433,n682);
nor (n682,n683,n684);
and (n683,n21,n469);
and (n684,n22,n471);
nand (n685,n686,n687);
or (n686,n408,n606);
or (n687,n415,n688);
nor (n688,n689,n690);
and (n689,n407,n266);
and (n690,n47,n268);
or (n691,n692,n719);
and (n692,n693,n718);
xor (n693,n694,n717);
or (n694,n695,n716);
and (n695,n696,n708);
xor (n696,n697,n703);
nand (n697,n698,n702);
or (n698,n151,n699);
nor (n699,n700,n701);
and (n700,n580,n161);
and (n701,n162,n582);
or (n702,n152,n650);
nand (n703,n704,n705);
or (n704,n384,n369);
nand (n705,n706,n707);
not (n706,n628);
not (n707,n370);
nand (n708,n709,n715);
or (n709,n561,n710);
nor (n710,n711,n713);
and (n711,n569,n712);
and (n713,n714,n570);
not (n714,n712);
or (n715,n562,n572);
and (n716,n697,n703);
xor (n717,n602,n612);
xor (n718,n657,n664);
and (n719,n694,n717);
or (n720,n721,n726);
and (n721,n722,n725);
xor (n722,n723,n724);
xor (n723,n640,n648);
xor (n724,n618,n625);
xor (n725,n555,n270);
and (n726,n723,n724);
or (n727,n728,n763);
and (n728,n729,n762);
xor (n729,n730,n761);
or (n730,n731,n760);
and (n731,n732,n759);
xor (n732,n733,n758);
or (n733,n734,n757);
and (n734,n735,n749);
xor (n735,n736,n743);
nand (n736,n737,n741);
or (n737,n738,n180);
nor (n738,n739,n740);
and (n739,n132,n266);
and (n740,n128,n268);
nand (n741,n742,n188);
not (n742,n536);
nand (n743,n744,n748);
or (n744,n151,n745);
nor (n745,n746,n747);
and (n746,n574,n161);
and (n747,n162,n576);
or (n748,n152,n699);
nand (n749,n750,n756);
or (n750,n561,n751);
nor (n751,n752,n754);
and (n752,n753,n569);
and (n754,n755,n570);
not (n755,n753);
or (n756,n562,n710);
and (n757,n736,n743);
xor (n758,n696,n708);
xor (n759,n479,n494);
and (n760,n733,n758);
xor (n761,n693,n718);
xor (n762,n722,n725);
and (n763,n730,n761);
or (n764,n765,n890);
and (n765,n766,n775);
xor (n766,n767,n774);
or (n767,n768,n773);
and (n768,n769,n772);
xor (n769,n770,n771);
xor (n770,n526,n543);
xor (n771,n503,n516);
xor (n772,n255,n284);
and (n773,n770,n771);
xor (n774,n252,n475);
or (n775,n776,n889);
and (n776,n777,n837);
xor (n777,n778,n836);
or (n778,n779,n835);
and (n779,n780,n813);
xor (n780,n781,n789);
not (n781,n782);
nor (n782,n783,n788);
and (n783,n336,n784);
not (n784,n785);
nor (n785,n786,n787);
and (n786,n340,n102);
and (n787,n341,n101);
and (n788,n328,n343);
or (n789,n790,n812);
and (n790,n791,n806);
xor (n791,n792,n799);
nand (n792,n793,n798);
or (n793,n794,n352);
not (n794,n795);
nand (n795,n796,n797);
or (n796,n111,n276);
or (n797,n110,n274);
nand (n798,n354,n349);
nand (n799,n800,n805);
or (n800,n801,n369);
not (n801,n802);
nand (n802,n803,n804);
or (n803,n378,n34);
or (n804,n377,n32);
or (n805,n370,n380);
nand (n806,n807,n811);
or (n807,n125,n808);
nor (n808,n809,n810);
and (n809,n135,n58);
and (n810,n136,n60);
or (n811,n126,n397);
and (n812,n792,n799);
or (n813,n814,n834);
and (n814,n815,n828);
xor (n815,n816,n822);
nand (n816,n817,n821);
or (n817,n818,n408);
nor (n818,n819,n820);
and (n819,n407,n84);
and (n820,n47,n86);
nand (n821,n419,n404);
nand (n822,n823,n827);
or (n823,n425,n824);
nor (n824,n825,n826);
and (n825,n21,n194);
and (n826,n22,n193);
or (n827,n433,n436);
nand (n828,n829,n833);
or (n829,n43,n830);
nor (n830,n831,n832);
and (n831,n53,n218);
and (n832,n54,n220);
or (n833,n62,n449);
and (n834,n816,n822);
and (n835,n781,n789);
xor (n836,n322,n444);
or (n837,n838,n888);
and (n838,n839,n887);
xor (n839,n840,n863);
or (n840,n841,n862);
and (n841,n842,n856);
xor (n842,n843,n849);
nand (n843,n844,n848);
or (n844,n70,n845);
nor (n845,n846,n847);
and (n846,n241,n79);
and (n847,n80,n243);
or (n848,n458,n72);
nand (n849,n850,n854);
or (n850,n851,n105);
nor (n851,n852,n853);
and (n852,n388,n100);
and (n853,n386,n104);
nand (n854,n855,n107);
not (n855,n467);
nand (n856,n857,n861);
or (n857,n16,n858);
nor (n858,n859,n860);
and (n859,n31,n140);
and (n860,n26,n142);
or (n861,n17,n289);
and (n862,n843,n849);
or (n863,n864,n886);
and (n864,n865,n880);
xor (n865,n866,n872);
nand (n866,n867,n868);
or (n867,n227,n298);
or (n868,n204,n869);
nor (n869,n870,n871);
and (n870,n217,n166);
and (n871,n208,n168);
nand (n872,n873,n878);
or (n873,n874,n230);
not (n874,n875);
nand (n875,n876,n877);
or (n876,n582,n155);
or (n877,n154,n580);
nand (n878,n309,n879);
not (n879,n231);
nand (n880,n881,n885);
or (n881,n180,n882);
nor (n882,n883,n884);
and (n883,n132,n260);
and (n884,n128,n262);
or (n885,n187,n738);
and (n886,n866,n872);
xor (n887,n392,n423);
and (n888,n840,n863);
and (n889,n778,n836);
and (n890,n767,n774);
or (n891,n892,n999);
and (n892,n893,n998);
xor (n893,n894,n997);
or (n894,n895,n996);
and (n895,n896,n905);
xor (n896,n897,n904);
or (n897,n898,n903);
and (n898,n899,n902);
xor (n899,n900,n901);
xor (n900,n735,n749);
xor (n901,n325,n367);
xor (n902,n286,n306);
and (n903,n900,n901);
xor (n904,n732,n759);
or (n905,n906,n995);
and (n906,n907,n927);
xor (n907,n908,n909);
xor (n908,n446,n465);
or (n909,n910,n926);
and (n910,n911,n782);
xor (n911,n912,n918);
nand (n912,n913,n917);
or (n913,n151,n914);
nor (n914,n915,n916);
and (n915,n712,n161);
and (n916,n714,n162);
or (n917,n152,n745);
nand (n918,n919,n925);
or (n919,n561,n920);
nor (n920,n921,n923);
and (n921,n922,n569);
and (n923,n570,n924);
not (n924,n922);
or (n925,n562,n751);
and (n926,n912,n918);
or (n927,n928,n994);
and (n928,n929,n970);
xor (n929,n930,n946);
or (n930,n931,n937);
nand (n931,n932,n936);
or (n932,n337,n933);
nor (n933,n934,n935);
and (n934,n283,n341);
and (n935,n281,n340);
or (n936,n329,n785);
nand (n937,n938,n943);
or (n938,n939,n942);
not (n939,n940);
nand (n940,n941,n331);
not (n941,n942);
nor (n943,n944,n945);
and (n944,n121,n331);
and (n945,n120,n335);
or (n946,n947,n969);
and (n947,n948,n963);
xor (n948,n949,n955);
nand (n949,n950,n954);
or (n950,n105,n951);
nor (n951,n952,n953);
and (n952,n40,n100);
and (n953,n38,n104);
or (n954,n278,n851);
nand (n955,n956,n962);
or (n956,n561,n957);
nor (n957,n958,n960);
and (n958,n959,n569);
and (n960,n570,n961);
not (n961,n959);
or (n962,n920,n562);
nand (n963,n964,n968);
or (n964,n180,n965);
nor (n965,n966,n967);
and (n966,n132,n65);
and (n967,n128,n67);
or (n968,n187,n882);
and (n969,n949,n955);
or (n970,n971,n993);
and (n971,n972,n987);
xor (n972,n973,n979);
nand (n973,n974,n978);
or (n974,n125,n975);
nor (n975,n976,n977);
and (n976,n135,n90);
and (n977,n136,n92);
or (n978,n126,n808);
nand (n979,n980,n981);
or (n980,n801,n370);
nand (n981,n982,n986);
not (n982,n983);
nor (n983,n984,n985);
and (n984,n377,n199);
and (n985,n378,n201);
not (n986,n369);
nand (n987,n988,n992);
or (n988,n408,n989);
nor (n989,n990,n991);
and (n990,n407,n224);
and (n991,n47,n226);
or (n992,n415,n818);
and (n993,n973,n979);
and (n994,n930,n946);
and (n995,n908,n909);
and (n996,n897,n904);
xor (n997,n729,n762);
xor (n998,n766,n775);
and (n999,n894,n997);
or (n1000,n1001,n1084);
and (n1001,n1002,n1065);
xor (n1002,n1003,n1064);
or (n1003,n1004,n1063);
and (n1004,n1005,n1062);
xor (n1005,n1006,n1007);
xor (n1006,n769,n772);
or (n1007,n1008,n1061);
and (n1008,n1009,n1012);
xor (n1009,n1010,n1011);
xor (n1010,n780,n813);
xor (n1011,n839,n887);
or (n1012,n1013,n1060);
and (n1013,n1014,n1059);
xor (n1014,n1015,n1037);
or (n1015,n1016,n1036);
and (n1016,n1017,n1030);
xor (n1017,n1018,n1024);
nand (n1018,n1019,n1023);
or (n1019,n1020,n43);
nor (n1020,n1021,n1022);
and (n1021,n249,n54);
and (n1022,n247,n53);
or (n1023,n62,n830);
nand (n1024,n1025,n1029);
or (n1025,n1026,n352);
nor (n1026,n1027,n1028);
and (n1027,n110,n469);
and (n1028,n111,n471);
nand (n1029,n354,n795);
nand (n1030,n1031,n1035);
or (n1031,n425,n1032);
nor (n1032,n1033,n1034);
and (n1033,n21,n146);
and (n1034,n22,n148);
or (n1035,n433,n824);
and (n1036,n1018,n1024);
or (n1037,n1038,n1058);
and (n1038,n1039,n1052);
xor (n1039,n1040,n1046);
nand (n1040,n1041,n1045);
or (n1041,n70,n1042);
nor (n1042,n1043,n1044);
and (n1043,n79,n174);
and (n1044,n80,n173);
or (n1045,n72,n845);
nand (n1046,n1047,n1051);
or (n1047,n204,n1048);
nor (n1048,n1049,n1050);
and (n1049,n217,n312);
and (n1050,n208,n311);
or (n1051,n227,n869);
nand (n1052,n1053,n1054);
or (n1053,n858,n17);
or (n1054,n16,n1055);
nor (n1055,n1056,n1057);
and (n1056,n31,n266);
and (n1057,n26,n268);
and (n1058,n1040,n1046);
xor (n1059,n791,n806);
and (n1060,n1015,n1037);
and (n1061,n1010,n1011);
xor (n1062,n777,n837);
and (n1063,n1006,n1007);
xor (n1064,n893,n998);
or (n1065,n1066,n1083);
and (n1066,n1067,n1082);
xor (n1067,n1068,n1069);
xor (n1068,n896,n905);
or (n1069,n1070,n1081);
and (n1070,n1071,n1080);
xor (n1071,n1072,n1079);
or (n1072,n1073,n1078);
and (n1073,n1074,n1077);
xor (n1074,n1075,n1076);
xor (n1075,n865,n880);
xor (n1076,n815,n828);
xor (n1077,n842,n856);
and (n1078,n1075,n1076);
xor (n1079,n899,n902);
xor (n1080,n907,n927);
and (n1081,n1072,n1079);
xor (n1082,n1005,n1062);
and (n1083,n1068,n1069);
and (n1084,n1003,n1064);
nand (n1085,n6,n1000);
not (n1086,n1087);
nand (n1087,n1088,n4240);
or (n1088,n1089,n1437);
nor (n1089,n1090,n1091);
xor (n1090,n1002,n1065);
or (n1091,n1092,n1436);
and (n1092,n1093,n1273);
xor (n1093,n1094,n1272);
or (n1094,n1095,n1271);
and (n1095,n1096,n1270);
xor (n1096,n1097,n1210);
or (n1097,n1098,n1209);
and (n1098,n1099,n1135);
xor (n1099,n1100,n1101);
xor (n1100,n911,n782);
or (n1101,n1102,n1134);
and (n1102,n1103,n1116);
xor (n1103,n1104,n1110);
nand (n1104,n1105,n1109);
or (n1105,n230,n1106);
nor (n1106,n1107,n1108);
and (n1107,n154,n574);
and (n1108,n155,n576);
or (n1109,n231,n874);
nand (n1110,n1111,n1115);
or (n1111,n151,n1112);
nor (n1112,n1113,n1114);
and (n1113,n753,n161);
and (n1114,n755,n162);
or (n1115,n152,n914);
and (n1116,n1117,n1126);
nor (n1117,n1118,n569);
nor (n1118,n1119,n1123);
and (n1119,n1120,n161);
not (n1120,n1121);
and (n1121,n1122,n565);
and (n1123,n1124,n1125);
not (n1124,n1122);
not (n1125,n565);
nand (n1126,n1127,n1129);
or (n1127,n941,n1128);
not (n1128,n943);
or (n1129,n940,n1130);
not (n1130,n1131);
nand (n1131,n1132,n1133);
or (n1132,n102,n335);
nand (n1133,n335,n102);
and (n1134,n1104,n1110);
or (n1135,n1136,n1208);
and (n1136,n1137,n1186);
xor (n1137,n1138,n1164);
or (n1138,n1139,n1163);
and (n1139,n1140,n1157);
xor (n1140,n1141,n1149);
nand (n1141,n1142,n1147);
or (n1142,n1143,n337);
not (n1143,n1144);
nor (n1144,n1145,n1146);
and (n1145,n274,n341);
and (n1146,n276,n340);
nand (n1147,n1148,n328);
not (n1148,n933);
nand (n1149,n1150,n1155);
or (n1150,n1151,n105);
not (n1151,n1152);
nand (n1152,n1153,n1154);
or (n1153,n100,n34);
or (n1154,n104,n32);
nand (n1155,n1156,n107);
not (n1156,n951);
nand (n1157,n1158,n1162);
or (n1158,n561,n1159);
nor (n1159,n1160,n1161);
and (n1160,n1124,n570);
and (n1161,n1122,n569);
or (n1162,n562,n957);
and (n1163,n1141,n1149);
or (n1164,n1165,n1185);
and (n1165,n1166,n1179);
xor (n1166,n1167,n1173);
nand (n1167,n1168,n1172);
or (n1168,n180,n1169);
nor (n1169,n1170,n1171);
and (n1170,n58,n132);
and (n1171,n60,n128);
or (n1172,n187,n965);
nand (n1173,n1174,n1178);
or (n1174,n125,n1175);
nor (n1175,n1176,n1177);
and (n1176,n135,n84);
and (n1177,n136,n86);
or (n1178,n126,n975);
nand (n1179,n1180,n1184);
or (n1180,n369,n1181);
nor (n1181,n1182,n1183);
and (n1182,n193,n378);
and (n1183,n194,n377);
or (n1184,n370,n983);
and (n1185,n1167,n1173);
or (n1186,n1187,n1207);
and (n1187,n1188,n1201);
xor (n1188,n1189,n1195);
nand (n1189,n1190,n1194);
or (n1190,n408,n1191);
nor (n1191,n1192,n1193);
and (n1192,n220,n47);
and (n1193,n218,n407);
or (n1194,n415,n989);
nand (n1195,n1196,n1200);
or (n1196,n43,n1197);
nor (n1197,n1198,n1199);
and (n1198,n53,n241);
and (n1199,n54,n243);
or (n1200,n62,n1020);
nand (n1201,n1202,n1206);
or (n1202,n352,n1203);
nor (n1203,n1204,n1205);
and (n1204,n110,n386);
and (n1205,n111,n388);
or (n1206,n530,n1026);
and (n1207,n1189,n1195);
and (n1208,n1138,n1164);
and (n1209,n1100,n1101);
or (n1210,n1211,n1269);
and (n1211,n1212,n1268);
xor (n1212,n1213,n1267);
or (n1213,n1214,n1266);
and (n1214,n1215,n1262);
xor (n1215,n1216,n1239);
or (n1216,n1217,n1238);
and (n1217,n1218,n1232);
xor (n1218,n1219,n1226);
nand (n1219,n1220,n1224);
or (n1220,n1221,n425);
nor (n1221,n1222,n1223);
and (n1222,n142,n22);
and (n1223,n140,n21);
nand (n1224,n1225,n432);
not (n1225,n1032);
nand (n1226,n1227,n1231);
or (n1227,n70,n1228);
nor (n1228,n1229,n1230);
and (n1229,n79,n166);
and (n1230,n80,n168);
or (n1231,n72,n1042);
nand (n1232,n1233,n1237);
or (n1233,n204,n1234);
nor (n1234,n1235,n1236);
and (n1235,n217,n580);
and (n1236,n208,n582);
or (n1237,n227,n1048);
and (n1238,n1219,n1226);
or (n1239,n1240,n1261);
and (n1240,n1241,n1255);
xor (n1241,n1242,n1249);
nand (n1242,n1243,n1248);
or (n1243,n1244,n16);
not (n1244,n1245);
nand (n1245,n1246,n1247);
or (n1246,n26,n262);
or (n1247,n31,n260);
or (n1248,n1055,n17);
nand (n1249,n1250,n1254);
or (n1250,n1251,n230);
nor (n1251,n1252,n1253);
and (n1252,n154,n712);
and (n1253,n155,n714);
or (n1254,n231,n1106);
nand (n1255,n1256,n1260);
or (n1256,n151,n1257);
nor (n1257,n1258,n1259);
and (n1258,n922,n161);
and (n1259,n924,n162);
or (n1260,n152,n1112);
and (n1261,n1242,n1249);
nand (n1262,n1263,n930);
or (n1263,n1264,n1265);
not (n1264,n937);
not (n1265,n931);
and (n1266,n1216,n1239);
xor (n1267,n929,n970);
xor (n1268,n1014,n1059);
and (n1269,n1213,n1267);
xor (n1270,n1009,n1012);
and (n1271,n1097,n1210);
xor (n1272,n1067,n1082);
or (n1273,n1274,n1435);
and (n1274,n1275,n1290);
xor (n1275,n1276,n1277);
xor (n1276,n1071,n1080);
or (n1277,n1278,n1289);
and (n1278,n1279,n1288);
xor (n1279,n1280,n1287);
or (n1280,n1281,n1286);
and (n1281,n1282,n1285);
xor (n1282,n1283,n1284);
xor (n1283,n972,n987);
xor (n1284,n1017,n1030);
xor (n1285,n1039,n1052);
and (n1286,n1283,n1284);
xor (n1287,n1074,n1077);
xor (n1288,n1099,n1135);
and (n1289,n1280,n1287);
or (n1290,n1291,n1434);
and (n1291,n1292,n1433);
xor (n1292,n1293,n1374);
or (n1293,n1294,n1373);
and (n1294,n1295,n1298);
xor (n1295,n1296,n1297);
xor (n1296,n948,n963);
xor (n1297,n1103,n1116);
or (n1298,n1299,n1372);
and (n1299,n1300,n1348);
xor (n1300,n1301,n1325);
or (n1301,n1302,n1324);
and (n1302,n1303,n1318);
xor (n1303,n1304,n1312);
nand (n1304,n1305,n1310);
or (n1305,n1306,n369);
not (n1306,n1307);
nor (n1307,n1308,n1309);
and (n1308,n146,n378);
and (n1309,n148,n377);
nand (n1310,n1311,n707);
not (n1311,n1181);
nand (n1312,n1313,n1317);
or (n1313,n408,n1314);
nor (n1314,n1315,n1316);
and (n1315,n407,n247);
and (n1316,n47,n249);
or (n1317,n415,n1191);
nand (n1318,n1319,n1323);
or (n1319,n43,n1320);
nor (n1320,n1321,n1322);
and (n1321,n53,n174);
and (n1322,n54,n173);
or (n1323,n62,n1197);
and (n1324,n1304,n1312);
or (n1325,n1326,n1347);
and (n1326,n1327,n1341);
xor (n1327,n1328,n1335);
nand (n1328,n1329,n1333);
or (n1329,n1330,n352);
nor (n1330,n1331,n1332);
and (n1331,n40,n111);
and (n1332,n38,n110);
nand (n1333,n1334,n354);
not (n1334,n1203);
nand (n1335,n1336,n1340);
or (n1336,n425,n1337);
nor (n1337,n1338,n1339);
and (n1338,n21,n266);
and (n1339,n22,n268);
or (n1340,n433,n1221);
nand (n1341,n1342,n1346);
or (n1342,n70,n1343);
nor (n1343,n1344,n1345);
and (n1344,n79,n312);
and (n1345,n80,n311);
or (n1346,n72,n1228);
and (n1347,n1328,n1335);
or (n1348,n1349,n1371);
and (n1349,n1350,n1365);
xor (n1350,n1351,n1358);
nand (n1351,n1352,n1357);
or (n1352,n1353,n204);
not (n1353,n1354);
nand (n1354,n1355,n1356);
or (n1355,n208,n576);
or (n1356,n217,n574);
or (n1357,n227,n1234);
nand (n1358,n1359,n1364);
or (n1359,n1360,n16);
not (n1360,n1361);
nand (n1361,n1362,n1363);
or (n1362,n26,n67);
or (n1363,n31,n65);
nand (n1364,n18,n1245);
nand (n1365,n1366,n1370);
or (n1366,n230,n1367);
nor (n1367,n1368,n1369);
and (n1368,n154,n753);
and (n1369,n155,n755);
or (n1370,n231,n1251);
and (n1371,n1351,n1358);
and (n1372,n1301,n1325);
and (n1373,n1296,n1297);
or (n1374,n1375,n1432);
and (n1375,n1376,n1431);
xor (n1376,n1377,n1424);
or (n1377,n1378,n1423);
and (n1378,n1379,n1400);
xor (n1379,n1380,n1381);
xor (n1380,n1117,n1126);
or (n1381,n1382,n1399);
and (n1382,n1383,n1392);
xor (n1383,n1384,n1385);
nor (n1384,n562,n1124);
nand (n1385,n1386,n1391);
or (n1386,n940,n1387);
not (n1387,n1388);
nor (n1388,n1389,n1390);
and (n1389,n283,n335);
and (n1390,n281,n331);
nand (n1391,n1131,n942);
nand (n1392,n1393,n1398);
or (n1393,n1394,n337);
not (n1394,n1395);
nand (n1395,n1396,n1397);
or (n1396,n341,n471);
or (n1397,n340,n469);
nand (n1398,n328,n1144);
and (n1399,n1384,n1385);
or (n1400,n1401,n1422);
and (n1401,n1402,n1416);
xor (n1402,n1403,n1410);
nand (n1403,n1404,n1409);
or (n1404,n1405,n105);
not (n1405,n1406);
nand (n1406,n1407,n1408);
or (n1407,n100,n201);
or (n1408,n104,n199);
nand (n1409,n107,n1152);
nand (n1410,n1411,n1415);
or (n1411,n180,n1412);
nor (n1412,n1413,n1414);
and (n1413,n132,n90);
and (n1414,n128,n92);
or (n1415,n187,n1169);
nand (n1416,n1417,n1421);
or (n1417,n125,n1418);
nor (n1418,n1419,n1420);
and (n1419,n135,n224);
and (n1420,n136,n226);
or (n1421,n126,n1175);
and (n1422,n1403,n1410);
and (n1423,n1380,n1381);
or (n1424,n1425,n1430);
and (n1425,n1426,n1429);
xor (n1426,n1427,n1428);
xor (n1427,n1241,n1255);
xor (n1428,n1140,n1157);
xor (n1429,n1166,n1179);
and (n1430,n1427,n1428);
xor (n1431,n1215,n1262);
and (n1432,n1377,n1424);
xor (n1433,n1212,n1268);
and (n1434,n1293,n1374);
and (n1435,n1276,n1277);
and (n1436,n1094,n1272);
not (n1437,n1438);
nand (n1438,n1439,n4225);
or (n1439,n1440,n2078);
nand (n1440,n1441,n1647);
nor (n1441,n1442,n1632);
nor (n1442,n1443,n1444);
xor (n1443,n1093,n1273);
or (n1444,n1445,n1631);
and (n1445,n1446,n1449);
xor (n1446,n1447,n1448);
xor (n1447,n1096,n1270);
xor (n1448,n1275,n1290);
or (n1449,n1450,n1630);
and (n1450,n1451,n1539);
xor (n1451,n1452,n1453);
xor (n1452,n1279,n1288);
or (n1453,n1454,n1538);
and (n1454,n1455,n1458);
xor (n1455,n1456,n1457);
xor (n1456,n1137,n1186);
xor (n1457,n1282,n1285);
or (n1458,n1459,n1537);
and (n1459,n1460,n1463);
xor (n1460,n1461,n1462);
xor (n1461,n1188,n1201);
xor (n1462,n1218,n1232);
or (n1463,n1464,n1536);
and (n1464,n1465,n1513);
xor (n1465,n1466,n1489);
or (n1466,n1467,n1488);
and (n1467,n1468,n1481);
xor (n1468,n1469,n1475);
nand (n1469,n1470,n1474);
or (n1470,n125,n1471);
nor (n1471,n1472,n1473);
and (n1472,n135,n218);
and (n1473,n136,n220);
or (n1474,n126,n1418);
nand (n1475,n1476,n1480);
or (n1476,n369,n1477);
nor (n1477,n1478,n1479);
and (n1478,n377,n140);
and (n1479,n378,n142);
or (n1480,n370,n1306);
nand (n1481,n1482,n1487);
or (n1482,n408,n1483);
not (n1483,n1484);
nor (n1484,n1485,n1486);
and (n1485,n241,n47);
and (n1486,n243,n407);
or (n1487,n415,n1314);
and (n1488,n1469,n1475);
or (n1489,n1490,n1512);
and (n1490,n1491,n1506);
xor (n1491,n1492,n1500);
nand (n1492,n1493,n1498);
or (n1493,n1494,n43);
not (n1494,n1495);
nand (n1495,n1496,n1497);
or (n1496,n54,n168);
or (n1497,n53,n166);
nand (n1498,n1499,n45);
not (n1499,n1320);
nand (n1500,n1501,n1505);
or (n1501,n352,n1502);
nor (n1502,n1503,n1504);
and (n1503,n110,n32);
and (n1504,n111,n34);
or (n1505,n530,n1330);
nand (n1506,n1507,n1511);
or (n1507,n425,n1508);
nor (n1508,n1509,n1510);
and (n1509,n21,n260);
and (n1510,n22,n262);
or (n1511,n433,n1337);
and (n1512,n1492,n1500);
or (n1513,n1514,n1535);
and (n1514,n1515,n1529);
xor (n1515,n1516,n1522);
nand (n1516,n1517,n1521);
or (n1517,n70,n1518);
nor (n1518,n1519,n1520);
and (n1519,n79,n580);
and (n1520,n80,n582);
or (n1521,n72,n1343);
nand (n1522,n1523,n1524);
or (n1523,n1353,n227);
nand (n1524,n1525,n205);
not (n1525,n1526);
nor (n1526,n1527,n1528);
and (n1527,n217,n712);
and (n1528,n714,n208);
nand (n1529,n1530,n1534);
or (n1530,n1531,n16);
nor (n1531,n1532,n1533);
and (n1532,n31,n58);
and (n1533,n26,n60);
or (n1534,n17,n1360);
and (n1535,n1516,n1522);
and (n1536,n1466,n1489);
and (n1537,n1461,n1462);
and (n1538,n1456,n1457);
or (n1539,n1540,n1629);
and (n1540,n1541,n1594);
xor (n1541,n1542,n1543);
xor (n1542,n1295,n1298);
or (n1543,n1544,n1593);
and (n1544,n1545,n1592);
xor (n1545,n1546,n1591);
or (n1546,n1547,n1590);
and (n1547,n1548,n1568);
xor (n1548,n1549,n1555);
nand (n1549,n1550,n1554);
or (n1550,n151,n1551);
nor (n1551,n1552,n1553);
and (n1552,n161,n959);
and (n1553,n961,n162);
or (n1554,n152,n1257);
and (n1555,n1556,n1562);
nor (n1556,n1557,n161);
nor (n1557,n1558,n1561);
and (n1558,n1559,n154);
not (n1559,n1560);
and (n1560,n1122,n156);
and (n1561,n1124,n158);
nand (n1562,n1563,n1564);
or (n1563,n941,n1387);
or (n1564,n940,n1565);
nor (n1565,n1566,n1567);
and (n1566,n335,n274);
and (n1567,n331,n276);
or (n1568,n1569,n1589);
and (n1569,n1570,n1583);
xor (n1570,n1571,n1577);
nand (n1571,n1572,n1573);
or (n1572,n1394,n329);
or (n1573,n337,n1574);
nor (n1574,n1575,n1576);
and (n1575,n388,n341);
and (n1576,n386,n340);
nand (n1577,n1578,n1579);
or (n1578,n1405,n278);
or (n1579,n105,n1580);
nor (n1580,n1581,n1582);
and (n1581,n104,n194);
and (n1582,n100,n193);
nand (n1583,n1584,n1588);
or (n1584,n180,n1585);
nor (n1585,n1586,n1587);
and (n1586,n132,n84);
and (n1587,n128,n86);
or (n1588,n187,n1412);
and (n1589,n1571,n1577);
and (n1590,n1549,n1555);
xor (n1591,n1300,n1348);
xor (n1592,n1379,n1400);
and (n1593,n1546,n1591);
or (n1594,n1595,n1628);
and (n1595,n1596,n1627);
xor (n1596,n1597,n1604);
or (n1597,n1598,n1603);
and (n1598,n1599,n1602);
xor (n1599,n1600,n1601);
xor (n1600,n1383,n1392);
xor (n1601,n1350,n1365);
xor (n1602,n1327,n1341);
and (n1603,n1600,n1601);
or (n1604,n1605,n1626);
and (n1605,n1606,n1609);
xor (n1606,n1607,n1608);
xor (n1607,n1303,n1318);
xor (n1608,n1402,n1416);
or (n1609,n1610,n1625);
and (n1610,n1611,n1624);
xor (n1611,n1612,n1618);
nand (n1612,n1613,n1617);
or (n1613,n230,n1614);
nor (n1614,n1615,n1616);
and (n1615,n154,n922);
and (n1616,n155,n924);
or (n1617,n231,n1367);
nand (n1618,n1619,n1623);
or (n1619,n151,n1620);
nor (n1620,n1621,n1622);
and (n1621,n1124,n162);
and (n1622,n1122,n161);
or (n1623,n152,n1551);
xor (n1624,n1556,n1562);
and (n1625,n1612,n1618);
and (n1626,n1607,n1608);
xor (n1627,n1426,n1429);
and (n1628,n1597,n1604);
and (n1629,n1542,n1543);
and (n1630,n1452,n1453);
and (n1631,n1447,n1448);
nor (n1632,n1633,n1646);
or (n1633,n1634,n1645);
and (n1634,n1635,n1638);
xor (n1635,n1636,n1637);
xor (n1636,n1292,n1433);
xor (n1637,n1451,n1539);
or (n1638,n1639,n1644);
and (n1639,n1640,n1643);
xor (n1640,n1641,n1642);
xor (n1641,n1376,n1431);
xor (n1642,n1455,n1458);
xor (n1643,n1541,n1594);
and (n1644,n1641,n1642);
and (n1645,n1636,n1637);
xor (n1646,n1446,n1449);
nor (n1647,n1648,n1940);
nor (n1648,n1649,n1650);
xor (n1649,n1635,n1638);
or (n1650,n1651,n1939);
and (n1651,n1652,n1938);
xor (n1652,n1653,n1795);
or (n1653,n1654,n1794);
and (n1654,n1655,n1738);
xor (n1655,n1656,n1657);
xor (n1656,n1460,n1463);
or (n1657,n1658,n1737);
and (n1658,n1659,n1730);
xor (n1659,n1660,n1661);
xor (n1660,n1548,n1568);
or (n1661,n1662,n1729);
and (n1662,n1663,n1706);
xor (n1663,n1664,n1687);
or (n1664,n1665,n1686);
and (n1665,n1666,n1680);
xor (n1666,n1667,n1674);
nand (n1667,n1668,n1673);
or (n1668,n1669,n408);
not (n1669,n1670);
nor (n1670,n1671,n1672);
and (n1671,n174,n47);
and (n1672,n173,n407);
nand (n1673,n1484,n419);
nand (n1674,n1675,n1679);
or (n1675,n1676,n43);
nor (n1676,n1677,n1678);
and (n1677,n311,n54);
and (n1678,n312,n53);
nand (n1679,n1495,n45);
nand (n1680,n1681,n1685);
or (n1681,n940,n1682);
nor (n1682,n1683,n1684);
and (n1683,n335,n469);
and (n1684,n331,n471);
or (n1685,n1565,n941);
and (n1686,n1667,n1674);
or (n1687,n1688,n1705);
and (n1688,n1689,n1699);
xor (n1689,n1690,n1691);
nor (n1690,n152,n1124);
nand (n1691,n1692,n1697);
or (n1692,n1693,n337);
not (n1693,n1694);
nand (n1694,n1695,n1696);
or (n1695,n341,n40);
or (n1696,n340,n38);
nand (n1697,n1698,n328);
not (n1698,n1574);
nand (n1699,n1700,n1704);
or (n1700,n105,n1701);
nor (n1701,n1702,n1703);
and (n1702,n104,n146);
and (n1703,n100,n148);
or (n1704,n278,n1580);
and (n1705,n1690,n1691);
or (n1706,n1707,n1728);
and (n1707,n1708,n1722);
xor (n1708,n1709,n1716);
nand (n1709,n1710,n1714);
or (n1710,n1711,n180);
nor (n1711,n1712,n1713);
and (n1712,n224,n132);
and (n1713,n226,n128);
nand (n1714,n1715,n188);
not (n1715,n1585);
nand (n1716,n1717,n1721);
or (n1717,n125,n1718);
nor (n1718,n1719,n1720);
and (n1719,n135,n247);
and (n1720,n136,n249);
or (n1721,n126,n1471);
nand (n1722,n1723,n1727);
or (n1723,n369,n1724);
nor (n1724,n1725,n1726);
and (n1725,n377,n266);
and (n1726,n378,n268);
or (n1727,n370,n1477);
and (n1728,n1709,n1716);
and (n1729,n1664,n1687);
or (n1730,n1731,n1736);
and (n1731,n1732,n1735);
xor (n1732,n1733,n1734);
xor (n1733,n1515,n1529);
xor (n1734,n1468,n1481);
xor (n1735,n1491,n1506);
and (n1736,n1733,n1734);
and (n1737,n1660,n1661);
or (n1738,n1739,n1793);
and (n1739,n1740,n1792);
xor (n1740,n1741,n1742);
xor (n1741,n1465,n1513);
or (n1742,n1743,n1791);
and (n1743,n1744,n1790);
xor (n1744,n1745,n1768);
or (n1745,n1746,n1767);
and (n1746,n1747,n1761);
xor (n1747,n1748,n1755);
nand (n1748,n1749,n1754);
or (n1749,n1750,n425);
not (n1750,n1751);
nor (n1751,n1752,n1753);
and (n1752,n65,n22);
and (n1753,n67,n21);
or (n1754,n433,n1508);
nand (n1755,n1756,n1760);
or (n1756,n70,n1757);
nor (n1757,n1758,n1759);
and (n1758,n79,n574);
and (n1759,n80,n576);
or (n1760,n72,n1518);
nand (n1761,n1762,n1766);
or (n1762,n204,n1763);
nor (n1763,n1764,n1765);
and (n1764,n753,n217);
and (n1765,n208,n755);
or (n1766,n1526,n227);
and (n1767,n1748,n1755);
or (n1768,n1769,n1789);
and (n1769,n1770,n1783);
xor (n1770,n1771,n1777);
nand (n1771,n1772,n1776);
or (n1772,n352,n1773);
nor (n1773,n1774,n1775);
and (n1774,n201,n111);
and (n1775,n199,n110);
or (n1776,n530,n1502);
nand (n1777,n1778,n1782);
or (n1778,n230,n1779);
nor (n1779,n1780,n1781);
and (n1780,n959,n154);
and (n1781,n155,n961);
or (n1782,n231,n1614);
nand (n1783,n1784,n1788);
or (n1784,n16,n1785);
nor (n1785,n1786,n1787);
and (n1786,n31,n90);
and (n1787,n26,n92);
or (n1788,n17,n1531);
and (n1789,n1771,n1777);
xor (n1790,n1570,n1583);
and (n1791,n1745,n1768);
xor (n1792,n1606,n1609);
and (n1793,n1741,n1742);
and (n1794,n1656,n1657);
or (n1795,n1796,n1937);
and (n1796,n1797,n1800);
xor (n1797,n1798,n1799);
xor (n1798,n1545,n1592);
xor (n1799,n1596,n1627);
or (n1800,n1801,n1936);
and (n1801,n1802,n1859);
xor (n1802,n1803,n1804);
xor (n1803,n1599,n1602);
or (n1804,n1805,n1858);
and (n1805,n1806,n1857);
xor (n1806,n1807,n1808);
xor (n1807,n1663,n1706);
or (n1808,n1809,n1856);
and (n1809,n1810,n1855);
xor (n1810,n1811,n1833);
or (n1811,n1812,n1832);
and (n1812,n1813,n1826);
xor (n1813,n1814,n1820);
nand (n1814,n1815,n1819);
or (n1815,n204,n1816);
nor (n1816,n1817,n1818);
and (n1817,n924,n208);
and (n1818,n922,n217);
or (n1819,n1763,n227);
nand (n1820,n1821,n1825);
or (n1821,n352,n1822);
nor (n1822,n1823,n1824);
and (n1823,n110,n194);
and (n1824,n111,n193);
or (n1825,n530,n1773);
nand (n1826,n1827,n1831);
or (n1827,n230,n1828);
nor (n1828,n1829,n1830);
and (n1829,n1124,n155);
and (n1830,n1122,n154);
or (n1831,n1779,n231);
and (n1832,n1814,n1820);
or (n1833,n1834,n1854);
and (n1834,n1835,n1848);
xor (n1835,n1836,n1842);
nand (n1836,n1837,n1841);
or (n1837,n940,n1838);
nor (n1838,n1839,n1840);
and (n1839,n388,n331);
and (n1840,n386,n335);
or (n1841,n1682,n941);
nand (n1842,n1843,n1847);
or (n1843,n1844,n425);
nor (n1844,n1845,n1846);
and (n1845,n21,n58);
and (n1846,n22,n60);
nand (n1847,n432,n1751);
nand (n1848,n1849,n1853);
or (n1849,n70,n1850);
nor (n1850,n1851,n1852);
and (n1851,n79,n712);
and (n1852,n80,n714);
or (n1853,n72,n1757);
and (n1854,n1836,n1842);
xor (n1855,n1708,n1722);
and (n1856,n1811,n1833);
xor (n1857,n1744,n1790);
and (n1858,n1807,n1808);
or (n1859,n1860,n1935);
and (n1860,n1861,n1928);
xor (n1861,n1862,n1863);
xor (n1862,n1611,n1624);
or (n1863,n1864,n1927);
and (n1864,n1865,n1903);
xor (n1865,n1866,n1880);
and (n1866,n1867,n1873);
nand (n1867,n1868,n1872);
or (n1868,n1869,n337);
nor (n1869,n1870,n1871);
and (n1870,n340,n32);
and (n1871,n341,n34);
nand (n1872,n328,n1694);
not (n1873,n1874);
nand (n1874,n1875,n155);
nand (n1875,n1876,n1877);
or (n1876,n1122,n234);
nand (n1877,n1878,n217);
not (n1878,n1879);
and (n1879,n1122,n234);
or (n1880,n1881,n1902);
and (n1881,n1882,n1896);
xor (n1882,n1883,n1890);
nand (n1883,n1884,n1888);
or (n1884,n1885,n105);
nor (n1885,n1886,n1887);
and (n1886,n104,n140);
and (n1887,n100,n142);
nand (n1888,n1889,n107);
not (n1889,n1701);
nand (n1890,n1891,n1895);
or (n1891,n180,n1892);
nor (n1892,n1893,n1894);
and (n1893,n132,n218);
and (n1894,n128,n220);
or (n1895,n187,n1711);
nand (n1896,n1897,n1901);
or (n1897,n125,n1898);
nor (n1898,n1899,n1900);
and (n1899,n241,n135);
and (n1900,n136,n243);
or (n1901,n126,n1718);
and (n1902,n1883,n1890);
or (n1903,n1904,n1926);
and (n1904,n1905,n1920);
xor (n1905,n1906,n1913);
nand (n1906,n1907,n1911);
or (n1907,n1908,n369);
nor (n1908,n1909,n1910);
and (n1909,n377,n260);
and (n1910,n378,n262);
nand (n1911,n1912,n707);
not (n1912,n1724);
nand (n1913,n1914,n1919);
or (n1914,n1915,n408);
not (n1915,n1916);
nand (n1916,n1917,n1918);
or (n1917,n47,n168);
or (n1918,n407,n166);
nand (n1919,n419,n1670);
nand (n1920,n1921,n1925);
or (n1921,n43,n1922);
nor (n1922,n1923,n1924);
and (n1923,n53,n580);
and (n1924,n54,n582);
or (n1925,n62,n1676);
and (n1926,n1906,n1913);
and (n1927,n1866,n1880);
or (n1928,n1929,n1934);
and (n1929,n1930,n1933);
xor (n1930,n1931,n1932);
xor (n1931,n1770,n1783);
xor (n1932,n1689,n1699);
xor (n1933,n1666,n1680);
and (n1934,n1931,n1932);
and (n1935,n1862,n1863);
and (n1936,n1803,n1804);
and (n1937,n1798,n1799);
xor (n1938,n1640,n1643);
and (n1939,n1653,n1795);
nor (n1940,n1941,n2077);
or (n1941,n1942,n2076);
and (n1942,n1943,n1946);
xor (n1943,n1944,n1945);
xor (n1944,n1655,n1738);
xor (n1945,n1797,n1800);
or (n1946,n1947,n2075);
and (n1947,n1948,n1951);
xor (n1948,n1949,n1950);
xor (n1949,n1659,n1730);
xor (n1950,n1740,n1792);
or (n1951,n1952,n2074);
and (n1952,n1953,n2061);
xor (n1953,n1954,n1955);
xor (n1954,n1732,n1735);
or (n1955,n1956,n2060);
and (n1956,n1957,n2030);
xor (n1957,n1958,n1959);
xor (n1958,n1747,n1761);
or (n1959,n1960,n2029);
and (n1960,n1961,n2007);
xor (n1961,n1962,n1984);
or (n1962,n1963,n1983);
and (n1963,n1964,n1977);
xor (n1964,n1965,n1971);
nand (n1965,n1966,n1970);
or (n1966,n180,n1967);
nor (n1967,n1968,n1969);
and (n1968,n249,n128);
and (n1969,n247,n132);
or (n1970,n1892,n187);
nand (n1971,n1972,n1976);
or (n1972,n125,n1973);
nor (n1973,n1974,n1975);
and (n1974,n174,n135);
and (n1975,n136,n173);
or (n1976,n126,n1898);
nand (n1977,n1978,n1982);
or (n1978,n369,n1979);
nor (n1979,n1980,n1981);
and (n1980,n377,n65);
and (n1981,n378,n67);
or (n1982,n370,n1908);
and (n1983,n1965,n1971);
or (n1984,n1985,n2006);
and (n1985,n1986,n2000);
xor (n1986,n1987,n1994);
nand (n1987,n1988,n1989);
or (n1988,n415,n1915);
nand (n1989,n1990,n1991);
not (n1990,n408);
nand (n1991,n1992,n1993);
or (n1992,n47,n311);
or (n1993,n407,n312);
nand (n1994,n1995,n1999);
or (n1995,n43,n1996);
nor (n1996,n1997,n1998);
and (n1997,n53,n574);
and (n1998,n54,n576);
or (n1999,n62,n1922);
nand (n2000,n2001,n2005);
or (n2001,n940,n2002);
nor (n2002,n2003,n2004);
and (n2003,n335,n38);
and (n2004,n331,n40);
or (n2005,n1838,n941);
and (n2006,n1987,n1994);
or (n2007,n2008,n2028);
and (n2008,n2009,n2022);
xor (n2009,n2010,n2016);
nand (n2010,n2011,n2015);
or (n2011,n425,n2012);
nor (n2012,n2013,n2014);
and (n2013,n21,n90);
and (n2014,n22,n92);
or (n2015,n433,n1844);
nand (n2016,n2017,n2021);
or (n2017,n70,n2018);
nor (n2018,n2019,n2020);
and (n2019,n79,n753);
and (n2020,n80,n755);
or (n2021,n72,n1850);
nand (n2022,n2023,n2027);
or (n2023,n204,n2024);
nor (n2024,n2025,n2026);
and (n2025,n217,n959);
and (n2026,n208,n961);
or (n2027,n227,n1816);
and (n2028,n2010,n2016);
and (n2029,n1962,n1984);
or (n2030,n2031,n2059);
and (n2031,n2032,n2042);
xor (n2032,n2033,n2039);
nand (n2033,n2034,n2038);
or (n2034,n16,n2035);
nor (n2035,n2036,n2037);
and (n2036,n31,n84);
and (n2037,n26,n86);
or (n2038,n17,n1785);
nor (n2039,n1866,n2040);
and (n2040,n2041,n1874);
not (n2041,n1867);
or (n2042,n2043,n2058);
and (n2043,n2044,n2052);
xor (n2044,n2045,n2046);
nor (n2045,n231,n1124);
nand (n2046,n2047,n2051);
or (n2047,n337,n2048);
nor (n2048,n2049,n2050);
and (n2049,n340,n199);
and (n2050,n341,n201);
or (n2051,n329,n1869);
nand (n2052,n2053,n2057);
or (n2053,n105,n2054);
nor (n2054,n2055,n2056);
and (n2055,n104,n266);
and (n2056,n100,n268);
or (n2057,n278,n1885);
and (n2058,n2045,n2046);
and (n2059,n2033,n2039);
and (n2060,n1958,n1959);
or (n2061,n2062,n2073);
and (n2062,n2063,n2066);
xor (n2063,n2064,n2065);
xor (n2064,n1865,n1903);
xor (n2065,n1810,n1855);
or (n2066,n2067,n2072);
and (n2067,n2068,n2071);
xor (n2068,n2069,n2070);
xor (n2069,n1813,n1826);
xor (n2070,n1882,n1896);
xor (n2071,n1835,n1848);
and (n2072,n2069,n2070);
and (n2073,n2064,n2065);
and (n2074,n1954,n1955);
and (n2075,n1949,n1950);
and (n2076,n1944,n1945);
xor (n2077,n1652,n1938);
not (n2078,n2079);
nand (n2079,n2080,n4202,n4215);
nand (n2080,n2081,n2268,n3981,n4185);
nor (n2081,n2082,n2097);
nor (n2082,n2083,n2084);
xor (n2083,n1943,n1946);
or (n2084,n2085,n2096);
and (n2085,n2086,n2089);
xor (n2086,n2087,n2088);
xor (n2087,n1802,n1859);
xor (n2088,n1948,n1951);
or (n2089,n2090,n2095);
and (n2090,n2091,n2094);
xor (n2091,n2092,n2093);
xor (n2092,n1861,n1928);
xor (n2093,n1806,n1857);
xor (n2094,n1953,n2061);
and (n2095,n2092,n2093);
and (n2096,n2087,n2088);
nor (n2097,n2098,n2099);
xor (n2098,n2086,n2089);
or (n2099,n2100,n2267);
and (n2100,n2101,n2266);
xor (n2101,n2102,n2247);
or (n2102,n2103,n2246);
and (n2103,n2104,n2141);
xor (n2104,n2105,n2106);
xor (n2105,n1930,n1933);
or (n2106,n2107,n2140);
and (n2107,n2108,n2139);
xor (n2108,n2109,n2110);
xor (n2109,n1905,n1920);
or (n2110,n2111,n2138);
and (n2111,n2112,n2125);
xor (n2112,n2113,n2119);
nand (n2113,n2114,n2118);
or (n2114,n352,n2115);
nor (n2115,n2116,n2117);
and (n2116,n110,n146);
and (n2117,n111,n148);
or (n2118,n530,n1822);
nand (n2119,n2120,n2124);
or (n2120,n16,n2121);
nor (n2121,n2122,n2123);
and (n2122,n31,n224);
and (n2123,n26,n226);
or (n2124,n17,n2035);
and (n2125,n2126,n2132);
nor (n2126,n2127,n217);
nor (n2127,n2128,n2131);
and (n2128,n2129,n79);
not (n2129,n2130);
and (n2130,n1122,n210);
and (n2131,n1124,n209);
nand (n2132,n2133,n2137);
or (n2133,n337,n2134);
nor (n2134,n2135,n2136);
and (n2135,n340,n194);
and (n2136,n341,n193);
or (n2137,n329,n2048);
and (n2138,n2113,n2119);
xor (n2139,n2032,n2042);
and (n2140,n2109,n2110);
or (n2141,n2142,n2245);
and (n2142,n2143,n2244);
xor (n2143,n2144,n2216);
or (n2144,n2145,n2215);
and (n2145,n2146,n2193);
xor (n2146,n2147,n2170);
or (n2147,n2148,n2169);
and (n2148,n2149,n2163);
xor (n2149,n2150,n2157);
nand (n2150,n2151,n2155);
or (n2151,n2152,n105);
nor (n2152,n2153,n2154);
and (n2153,n104,n260);
and (n2154,n100,n262);
nand (n2155,n2156,n107);
not (n2156,n2054);
nand (n2157,n2158,n2162);
or (n2158,n180,n2159);
nor (n2159,n2160,n2161);
and (n2160,n132,n241);
and (n2161,n128,n243);
or (n2162,n187,n1967);
nand (n2163,n2164,n2168);
or (n2164,n125,n2165);
nor (n2165,n2166,n2167);
and (n2166,n135,n166);
and (n2167,n136,n168);
or (n2168,n126,n1973);
and (n2169,n2150,n2157);
or (n2170,n2171,n2192);
and (n2171,n2172,n2186);
xor (n2172,n2173,n2179);
nand (n2173,n2174,n2178);
or (n2174,n369,n2175);
nor (n2175,n2176,n2177);
and (n2176,n377,n58);
and (n2177,n378,n60);
or (n2178,n370,n1979);
nand (n2179,n2180,n2184);
or (n2180,n408,n2181);
nor (n2181,n2182,n2183);
and (n2182,n407,n580);
and (n2183,n47,n582);
or (n2184,n415,n2185);
not (n2185,n1991);
nand (n2186,n2187,n2191);
or (n2187,n43,n2188);
nor (n2188,n2189,n2190);
and (n2189,n53,n712);
and (n2190,n54,n714);
or (n2191,n62,n1996);
and (n2192,n2173,n2179);
or (n2193,n2194,n2214);
and (n2194,n2195,n2208);
xor (n2195,n2196,n2202);
nand (n2196,n2197,n2201);
or (n2197,n940,n2198);
nor (n2198,n2199,n2200);
and (n2199,n335,n32);
and (n2200,n331,n34);
or (n2201,n2002,n941);
nand (n2202,n2203,n2207);
or (n2203,n425,n2204);
nor (n2204,n2205,n2206);
and (n2205,n21,n84);
and (n2206,n22,n86);
or (n2207,n433,n2012);
nand (n2208,n2209,n2210);
or (n2209,n2018,n72);
or (n2210,n70,n2211);
nor (n2211,n2212,n2213);
and (n2212,n922,n79);
and (n2213,n80,n924);
and (n2214,n2196,n2202);
and (n2215,n2147,n2170);
or (n2216,n2217,n2243);
and (n2217,n2218,n2242);
xor (n2218,n2219,n2241);
or (n2219,n2220,n2240);
and (n2220,n2221,n2234);
xor (n2221,n2222,n2228);
nand (n2222,n2223,n2227);
or (n2223,n204,n2224);
nor (n2224,n2225,n2226);
and (n2225,n1124,n208);
and (n2226,n1122,n217);
or (n2227,n2024,n227);
nand (n2228,n2229,n2233);
or (n2229,n352,n2230);
nor (n2230,n2231,n2232);
and (n2231,n110,n140);
and (n2232,n111,n142);
or (n2233,n530,n2115);
nand (n2234,n2235,n2239);
or (n2235,n16,n2236);
nor (n2236,n2237,n2238);
and (n2237,n31,n218);
and (n2238,n26,n220);
or (n2239,n17,n2121);
and (n2240,n2222,n2228);
xor (n2241,n2044,n2052);
xor (n2242,n1986,n2000);
and (n2243,n2219,n2241);
xor (n2244,n1961,n2007);
and (n2245,n2144,n2216);
and (n2246,n2105,n2106);
or (n2247,n2248,n2265);
and (n2248,n2249,n2252);
xor (n2249,n2250,n2251);
xor (n2250,n1957,n2030);
xor (n2251,n2063,n2066);
or (n2252,n2253,n2264);
and (n2253,n2254,n2263);
xor (n2254,n2255,n2262);
or (n2255,n2256,n2261);
and (n2256,n2257,n2260);
xor (n2257,n2258,n2259);
xor (n2258,n1964,n1977);
xor (n2259,n2009,n2022);
xor (n2260,n2112,n2125);
and (n2261,n2258,n2259);
xor (n2262,n2068,n2071);
xor (n2263,n2108,n2139);
and (n2264,n2255,n2262);
and (n2265,n2250,n2251);
xor (n2266,n2091,n2094);
and (n2267,n2102,n2247);
nand (n2268,n2269,n3462);
nor (n2269,n2270,n3448);
and (n2270,n2271,n2860,n3182);
nor (n2271,n2272,n2774);
nor (n2272,n2273,n2661);
xor (n2273,n2274,n2654);
xor (n2274,n2275,n2447);
or (n2275,n2276,n2446);
and (n2276,n2277,n2371);
xor (n2277,n2278,n2314);
xor (n2278,n2279,n2298);
xor (n2279,n2280,n2289);
nand (n2280,n2281,n2285);
or (n2281,n425,n2282);
nor (n2282,n2283,n2284);
and (n2283,n21,n174);
and (n2284,n22,n173);
or (n2285,n433,n2286);
nor (n2286,n2287,n2288);
and (n2287,n21,n241);
and (n2288,n22,n243);
nand (n2289,n2290,n2294);
or (n2290,n16,n2291);
nor (n2291,n2292,n2293);
and (n2292,n312,n31);
and (n2293,n26,n311);
or (n2294,n17,n2295);
nor (n2295,n2296,n2297);
and (n2296,n31,n166);
and (n2297,n26,n168);
and (n2298,n2299,n2305);
nor (n2299,n2300,n407);
nor (n2300,n2301,n2304);
and (n2301,n2302,n135);
not (n2302,n2303);
and (n2303,n1122,n412);
and (n2304,n1124,n414);
nand (n2305,n2306,n2310);
or (n2306,n940,n2307);
nor (n2307,n2308,n2309);
and (n2308,n335,n260);
and (n2309,n331,n262);
or (n2310,n2311,n941);
nor (n2311,n2312,n2313);
and (n2312,n335,n266);
and (n2313,n331,n268);
or (n2314,n2315,n2370);
and (n2315,n2316,n2339);
xor (n2316,n2317,n2318);
xor (n2317,n2299,n2305);
or (n2318,n2319,n2338);
and (n2319,n2320,n2328);
xor (n2320,n2321,n2322);
and (n2321,n419,n1122);
nand (n2322,n2323,n2327);
or (n2323,n940,n2324);
nor (n2324,n2325,n2326);
and (n2325,n335,n65);
and (n2326,n331,n67);
or (n2327,n2307,n941);
nand (n2328,n2329,n2333);
or (n2329,n105,n2330);
nor (n2330,n2331,n2332);
and (n2331,n104,n247);
and (n2332,n100,n249);
or (n2333,n278,n2334);
not (n2334,n2335);
nor (n2335,n2336,n2337);
and (n2336,n218,n100);
and (n2337,n220,n104);
and (n2338,n2321,n2322);
or (n2339,n2340,n2369);
and (n2340,n2341,n2360);
xor (n2341,n2342,n2351);
nand (n2342,n2343,n2347);
or (n2343,n180,n2344);
nor (n2344,n2345,n2346);
and (n2345,n132,n753);
and (n2346,n128,n755);
or (n2347,n187,n2348);
nor (n2348,n2349,n2350);
and (n2349,n712,n132);
and (n2350,n714,n128);
nand (n2351,n2352,n2356);
or (n2352,n125,n2353);
nor (n2353,n2354,n2355);
and (n2354,n135,n959);
and (n2355,n136,n961);
or (n2356,n126,n2357);
nor (n2357,n2358,n2359);
and (n2358,n135,n922);
and (n2359,n136,n924);
nand (n2360,n2361,n2365);
or (n2361,n337,n2362);
nor (n2362,n2363,n2364);
and (n2363,n340,n90);
and (n2364,n341,n92);
or (n2365,n329,n2366);
nor (n2366,n2367,n2368);
and (n2367,n58,n340);
and (n2368,n60,n341);
and (n2369,n2342,n2351);
and (n2370,n2317,n2318);
or (n2371,n2372,n2445);
and (n2372,n2373,n2425);
xor (n2373,n2374,n2406);
or (n2374,n2375,n2405);
and (n2375,n2376,n2396);
xor (n2376,n2377,n2387);
nand (n2377,n2378,n2383);
or (n2378,n2379,n369);
not (n2379,n2380);
nand (n2380,n2381,n2382);
or (n2381,n378,n173);
or (n2382,n377,n174);
nand (n2383,n707,n2384);
nor (n2384,n2385,n2386);
and (n2385,n243,n377);
and (n2386,n241,n378);
nand (n2387,n2388,n2392);
or (n2388,n2389,n352);
nor (n2389,n2390,n2391);
and (n2390,n110,n224);
and (n2391,n111,n226);
nand (n2392,n354,n2393);
nand (n2393,n2394,n2395);
or (n2394,n111,n86);
or (n2395,n110,n84);
nand (n2396,n2397,n2401);
or (n2397,n425,n2398);
nor (n2398,n2399,n2400);
and (n2399,n21,n312);
and (n2400,n22,n311);
or (n2401,n433,n2402);
nor (n2402,n2403,n2404);
and (n2403,n166,n21);
and (n2404,n22,n168);
and (n2405,n2377,n2387);
xor (n2406,n2407,n2419);
xor (n2407,n2408,n2416);
nand (n2408,n2409,n2411);
or (n2409,n2410,n352);
not (n2410,n2393);
nand (n2411,n2412,n354);
not (n2412,n2413);
nor (n2413,n2414,n2415);
and (n2414,n92,n111);
and (n2415,n90,n110);
nand (n2416,n2417,n2418);
or (n2417,n425,n2402);
or (n2418,n2282,n433);
nand (n2419,n2420,n2424);
or (n2420,n16,n2421);
nor (n2421,n2422,n2423);
and (n2422,n580,n31);
and (n2423,n26,n582);
or (n2424,n17,n2291);
xor (n2425,n2426,n2439);
xor (n2426,n2427,n2433);
nand (n2427,n2428,n2429);
or (n2428,n2334,n105);
nand (n2429,n2430,n107);
nor (n2430,n2431,n2432);
and (n2431,n226,n104);
and (n2432,n224,n100);
nand (n2433,n2434,n2435);
or (n2434,n2348,n180);
nand (n2435,n2436,n188);
nor (n2436,n2437,n2438);
and (n2437,n576,n132);
and (n2438,n574,n128);
nand (n2439,n2440,n2441);
or (n2440,n125,n2357);
or (n2441,n2442,n126);
nor (n2442,n2443,n2444);
and (n2443,n135,n753);
and (n2444,n136,n755);
and (n2445,n2374,n2406);
and (n2446,n2278,n2314);
xor (n2447,n2448,n2572);
xor (n2448,n2449,n2523);
or (n2449,n2450,n2522);
and (n2450,n2451,n2493);
xor (n2451,n2452,n2469);
xor (n2452,n2453,n2461);
xor (n2453,n2454,n2455);
and (n2454,n45,n1122);
nand (n2455,n2456,n2457);
or (n2456,n940,n2311);
or (n2457,n2458,n941);
nor (n2458,n2459,n2460);
and (n2459,n142,n331);
and (n2460,n140,n335);
nand (n2461,n2462,n2464);
or (n2462,n105,n2463);
not (n2463,n2430);
or (n2464,n278,n2465);
not (n2465,n2466);
nor (n2466,n2467,n2468);
and (n2467,n84,n100);
and (n2468,n86,n104);
xor (n2469,n2470,n2484);
xor (n2470,n2471,n2478);
nand (n2471,n2472,n2474);
or (n2472,n2473,n180);
not (n2473,n2436);
or (n2474,n187,n2475);
nor (n2475,n2476,n2477);
and (n2476,n582,n128);
and (n2477,n580,n132);
nand (n2478,n2479,n2480);
or (n2479,n125,n2442);
or (n2480,n126,n2481);
nor (n2481,n2482,n2483);
and (n2482,n135,n712);
and (n2483,n136,n714);
nand (n2484,n2485,n2489);
or (n2485,n337,n2486);
nor (n2486,n2487,n2488);
and (n2487,n340,n65);
and (n2488,n341,n67);
or (n2489,n329,n2490);
nor (n2490,n2491,n2492);
and (n2491,n340,n260);
and (n2492,n341,n262);
xor (n2493,n2494,n2516);
xor (n2494,n2495,n2505);
nand (n2495,n2496,n2501);
or (n2496,n2497,n408);
not (n2497,n2498);
nand (n2498,n2499,n2500);
or (n2499,n47,n961);
or (n2500,n407,n959);
or (n2501,n415,n2502);
nor (n2502,n2503,n2504);
and (n2503,n924,n47);
and (n2504,n922,n407);
nand (n2505,n2506,n2511);
or (n2506,n2507,n370);
not (n2507,n2508);
nand (n2508,n2509,n2510);
or (n2509,n378,n220);
or (n2510,n377,n218);
nand (n2511,n2512,n986);
not (n2512,n2513);
nor (n2513,n2514,n2515);
and (n2514,n377,n247);
and (n2515,n378,n249);
nand (n2516,n2517,n2518);
or (n2517,n352,n2413);
or (n2518,n530,n2519);
nor (n2519,n2520,n2521);
and (n2520,n110,n58);
and (n2521,n111,n60);
and (n2522,n2452,n2469);
xor (n2523,n2524,n2569);
xor (n2524,n2525,n2545);
xor (n2525,n2526,n2539);
xor (n2526,n2527,n2533);
nand (n2527,n2528,n2529);
or (n2528,n2465,n105);
nand (n2529,n107,n2530);
nor (n2530,n2531,n2532);
and (n2531,n90,n100);
and (n2532,n92,n104);
nand (n2533,n2534,n2535);
or (n2534,n2475,n180);
nand (n2535,n188,n2536);
nand (n2536,n2537,n2538);
or (n2537,n128,n311);
or (n2538,n132,n312);
nand (n2539,n2540,n2541);
or (n2540,n125,n2481);
or (n2541,n126,n2542);
nor (n2542,n2543,n2544);
and (n2543,n135,n574);
and (n2544,n136,n576);
xor (n2545,n2546,n2560);
xor (n2546,n2547,n2554);
nand (n2547,n2548,n2549);
or (n2548,n2507,n369);
nand (n2549,n2550,n707);
not (n2550,n2551);
nor (n2551,n2552,n2553);
and (n2552,n226,n378);
and (n2553,n224,n377);
nand (n2554,n2555,n2556);
or (n2555,n408,n2502);
nand (n2556,n419,n2557);
nor (n2557,n2558,n2559);
and (n2558,n755,n407);
and (n2559,n753,n47);
nand (n2560,n2561,n2565);
or (n2561,n43,n2562);
nor (n2562,n2563,n2564);
and (n2563,n1124,n54);
and (n2564,n53,n1122);
or (n2565,n62,n2566);
nor (n2566,n2567,n2568);
and (n2567,n53,n959);
and (n2568,n54,n961);
or (n2569,n2570,n2571);
and (n2570,n2279,n2298);
and (n2571,n2280,n2289);
xor (n2572,n2573,n2626);
xor (n2573,n2574,n2602);
or (n2574,n2575,n2601);
and (n2575,n2576,n2583);
xor (n2576,n2577,n2580);
or (n2577,n2578,n2579);
and (n2578,n2426,n2439);
and (n2579,n2427,n2433);
or (n2580,n2581,n2582);
and (n2581,n2407,n2419);
and (n2582,n2408,n2416);
or (n2583,n2584,n2600);
and (n2584,n2585,n2596);
xor (n2585,n2586,n2590);
nand (n2586,n2587,n2588);
or (n2587,n2366,n337);
nand (n2588,n2589,n328);
not (n2589,n2486);
nand (n2590,n2591,n2592);
or (n2591,n2497,n415);
or (n2592,n408,n2593);
nor (n2593,n2594,n2595);
and (n2594,n47,n1124);
and (n2595,n407,n1122);
nand (n2596,n2597,n2599);
or (n2597,n369,n2598);
not (n2598,n2384);
or (n2599,n370,n2513);
and (n2600,n2586,n2590);
and (n2601,n2577,n2580);
xor (n2602,n2603,n2623);
xor (n2603,n2604,n2610);
nand (n2604,n2605,n2606);
or (n2605,n16,n2295);
or (n2606,n17,n2607);
nor (n2607,n2608,n2609);
and (n2608,n31,n174);
and (n2609,n26,n173);
xor (n2610,n2611,n2617);
and (n2611,n2612,n54);
nand (n2612,n2613,n2614);
or (n2613,n1122,n49);
nand (n2614,n2615,n407);
not (n2615,n2616);
and (n2616,n1122,n49);
nand (n2617,n2618,n2619);
or (n2618,n2490,n337);
nand (n2619,n328,n2620);
nor (n2620,n2621,n2622);
and (n2621,n266,n341);
and (n2622,n268,n340);
or (n2623,n2624,n2625);
and (n2624,n2470,n2484);
and (n2625,n2471,n2478);
xor (n2626,n2627,n2634);
xor (n2627,n2628,n2631);
or (n2628,n2629,n2630);
and (n2629,n2453,n2461);
and (n2630,n2454,n2455);
or (n2631,n2632,n2633);
and (n2632,n2494,n2516);
and (n2633,n2495,n2505);
xor (n2634,n2635,n2648);
xor (n2635,n2636,n2642);
nand (n2636,n2637,n2638);
or (n2637,n940,n2458);
or (n2638,n2639,n941);
nor (n2639,n2640,n2641);
and (n2640,n335,n146);
and (n2641,n331,n148);
nand (n2642,n2643,n2644);
or (n2643,n352,n2519);
nand (n2644,n354,n2645);
nor (n2645,n2646,n2647);
and (n2646,n65,n111);
and (n2647,n67,n110);
nand (n2648,n2649,n2650);
or (n2649,n425,n2286);
or (n2650,n433,n2651);
nor (n2651,n2652,n2653);
and (n2652,n21,n247);
and (n2653,n22,n249);
or (n2654,n2655,n2660);
and (n2655,n2656,n2659);
xor (n2656,n2657,n2658);
xor (n2657,n2576,n2583);
xor (n2658,n2451,n2493);
xor (n2659,n2277,n2371);
and (n2660,n2657,n2658);
or (n2661,n2662,n2773);
and (n2662,n2663,n2772);
xor (n2663,n2664,n2716);
or (n2664,n2665,n2715);
and (n2665,n2666,n2714);
xor (n2666,n2667,n2668);
xor (n2667,n2585,n2596);
or (n2668,n2669,n2713);
and (n2669,n2670,n2690);
xor (n2670,n2671,n2677);
nand (n2671,n2672,n2676);
or (n2672,n16,n2673);
nor (n2673,n2674,n2675);
and (n2674,n31,n574);
and (n2675,n26,n576);
or (n2676,n17,n2421);
and (n2677,n2678,n2684);
nor (n2678,n2679,n135);
nor (n2679,n2680,n2683);
and (n2680,n2681,n132);
not (n2681,n2682);
and (n2682,n1122,n130);
and (n2683,n1124,n129);
nand (n2684,n2685,n2689);
or (n2685,n940,n2686);
nor (n2686,n2687,n2688);
and (n2687,n335,n58);
and (n2688,n331,n60);
or (n2689,n2324,n941);
or (n2690,n2691,n2712);
and (n2691,n2692,n2706);
xor (n2692,n2693,n2700);
nand (n2693,n2694,n2698);
or (n2694,n2695,n105);
nor (n2695,n2696,n2697);
and (n2696,n104,n241);
and (n2697,n100,n243);
nand (n2698,n2699,n107);
not (n2699,n2330);
nand (n2700,n2701,n2705);
or (n2701,n180,n2702);
nor (n2702,n2703,n2704);
and (n2703,n132,n922);
and (n2704,n128,n924);
or (n2705,n187,n2344);
nand (n2706,n2707,n2711);
or (n2707,n125,n2708);
nor (n2708,n2709,n2710);
and (n2709,n1124,n136);
and (n2710,n135,n1122);
or (n2711,n126,n2353);
and (n2712,n2693,n2700);
and (n2713,n2671,n2677);
xor (n2714,n2316,n2339);
and (n2715,n2667,n2668);
or (n2716,n2717,n2771);
and (n2717,n2718,n2748);
xor (n2718,n2719,n2747);
or (n2719,n2720,n2746);
and (n2720,n2721,n2745);
xor (n2721,n2722,n2744);
or (n2722,n2723,n2743);
and (n2723,n2724,n2737);
xor (n2724,n2725,n2731);
nand (n2725,n2726,n2730);
or (n2726,n337,n2727);
nor (n2727,n2728,n2729);
and (n2728,n340,n84);
and (n2729,n341,n86);
or (n2730,n329,n2362);
nand (n2731,n2732,n2736);
or (n2732,n369,n2733);
nor (n2733,n2734,n2735);
and (n2734,n377,n166);
and (n2735,n378,n168);
or (n2736,n370,n2379);
nand (n2737,n2738,n2742);
or (n2738,n352,n2739);
nor (n2739,n2740,n2741);
and (n2740,n110,n218);
and (n2741,n111,n220);
or (n2742,n530,n2389);
and (n2743,n2725,n2731);
xor (n2744,n2376,n2396);
xor (n2745,n2320,n2328);
and (n2746,n2722,n2744);
xor (n2747,n2373,n2425);
or (n2748,n2749,n2770);
and (n2749,n2750,n2769);
xor (n2750,n2751,n2752);
xor (n2751,n2341,n2360);
or (n2752,n2753,n2768);
and (n2753,n2754,n2767);
xor (n2754,n2755,n2761);
nand (n2755,n2756,n2760);
or (n2756,n425,n2757);
nor (n2757,n2758,n2759);
and (n2758,n21,n580);
and (n2759,n22,n582);
or (n2760,n433,n2398);
nand (n2761,n2762,n2766);
or (n2762,n16,n2763);
nor (n2763,n2764,n2765);
and (n2764,n31,n712);
and (n2765,n26,n714);
or (n2766,n17,n2673);
xor (n2767,n2678,n2684);
and (n2768,n2755,n2761);
xor (n2769,n2670,n2690);
and (n2770,n2751,n2752);
and (n2771,n2719,n2747);
xor (n2772,n2656,n2659);
and (n2773,n2664,n2716);
nor (n2774,n2775,n2776);
xor (n2775,n2663,n2772);
or (n2776,n2777,n2859);
and (n2777,n2778,n2858);
xor (n2778,n2779,n2780);
xor (n2779,n2666,n2714);
or (n2780,n2781,n2857);
and (n2781,n2782,n2856);
xor (n2782,n2783,n2849);
or (n2783,n2784,n2848);
and (n2784,n2785,n2826);
xor (n2785,n2786,n2804);
or (n2786,n2787,n2803);
and (n2787,n2788,n2797);
xor (n2788,n2789,n2791);
and (n2789,n2790,n1122);
not (n2790,n126);
nand (n2791,n2792,n2796);
or (n2792,n940,n2793);
nor (n2793,n2794,n2795);
and (n2794,n335,n90);
and (n2795,n331,n92);
or (n2796,n2686,n941);
nand (n2797,n2798,n2802);
or (n2798,n337,n2799);
nor (n2799,n2800,n2801);
and (n2800,n340,n224);
and (n2801,n341,n226);
or (n2802,n329,n2727);
and (n2803,n2789,n2791);
or (n2804,n2805,n2825);
and (n2805,n2806,n2819);
xor (n2806,n2807,n2813);
nand (n2807,n2808,n2812);
or (n2808,n352,n2809);
nor (n2809,n2810,n2811);
and (n2810,n110,n247);
and (n2811,n111,n249);
or (n2812,n530,n2739);
nand (n2813,n2814,n2818);
or (n2814,n425,n2815);
nor (n2815,n2816,n2817);
and (n2816,n21,n574);
and (n2817,n22,n576);
or (n2818,n433,n2757);
nand (n2819,n2820,n2824);
or (n2820,n16,n2821);
nor (n2821,n2822,n2823);
and (n2822,n31,n753);
and (n2823,n26,n755);
or (n2824,n17,n2763);
and (n2825,n2807,n2813);
or (n2826,n2827,n2847);
and (n2827,n2828,n2841);
xor (n2828,n2829,n2835);
nand (n2829,n2830,n2834);
or (n2830,n180,n2831);
nor (n2831,n2832,n2833);
and (n2832,n132,n959);
and (n2833,n128,n961);
or (n2834,n187,n2702);
nand (n2835,n2836,n2840);
or (n2836,n105,n2837);
nor (n2837,n2838,n2839);
and (n2838,n104,n174);
and (n2839,n100,n173);
or (n2840,n278,n2695);
nand (n2841,n2842,n2846);
or (n2842,n369,n2843);
nor (n2843,n2844,n2845);
and (n2844,n312,n377);
and (n2845,n378,n311);
or (n2846,n370,n2733);
and (n2847,n2829,n2835);
and (n2848,n2786,n2804);
or (n2849,n2850,n2855);
and (n2850,n2851,n2854);
xor (n2851,n2852,n2853);
xor (n2852,n2692,n2706);
xor (n2853,n2724,n2737);
xor (n2854,n2754,n2767);
and (n2855,n2852,n2853);
xor (n2856,n2721,n2745);
and (n2857,n2783,n2849);
xor (n2858,n2718,n2748);
and (n2859,n2779,n2780);
nand (n2860,n2861,n3181);
or (n2861,n2862,n3176);
nor (n2862,n2863,n3175);
and (n2863,n2864,n3163);
not (n2864,n2865);
nand (n2865,n2866,n3160);
or (n2866,n2867,n3140);
not (n2867,n2868);
nand (n2868,n2869,n3082);
xor (n2869,n2870,n3013);
xor (n2870,n2871,n2876);
xor (n2871,n2872,n2875);
xor (n2872,n2873,n2874);
xor (n2873,n2806,n2819);
xor (n2874,n2788,n2797);
xor (n2875,n2828,n2841);
or (n2876,n2877,n3012);
and (n2877,n2878,n2953);
xor (n2878,n2879,n2918);
or (n2879,n2880,n2917);
and (n2880,n2881,n2901);
xor (n2881,n2882,n2891);
nand (n2882,n2883,n2887);
or (n2883,n425,n2884);
nor (n2884,n2885,n2886);
and (n2885,n21,n753);
and (n2886,n22,n755);
or (n2887,n433,n2888);
nor (n2888,n2889,n2890);
and (n2889,n21,n712);
and (n2890,n22,n714);
nand (n2891,n2892,n2897);
or (n2892,n2893,n16);
not (n2893,n2894);
nand (n2894,n2895,n2896);
or (n2895,n961,n26);
or (n2896,n31,n959);
or (n2897,n17,n2898);
nor (n2898,n2899,n2900);
and (n2899,n31,n922);
and (n2900,n26,n924);
and (n2901,n2902,n2908);
nor (n2902,n2903,n31);
nor (n2903,n2904,n2907);
and (n2904,n2905,n21);
not (n2905,n2906);
and (n2906,n1122,n20);
and (n2907,n1124,n27);
nand (n2908,n2909,n2913);
or (n2909,n2910,n940);
nor (n2910,n2911,n2912);
and (n2911,n335,n218);
and (n2912,n331,n220);
or (n2913,n2914,n941);
nor (n2914,n2915,n2916);
and (n2915,n335,n224);
and (n2916,n331,n226);
and (n2917,n2882,n2891);
xor (n2918,n2919,n2936);
xor (n2919,n2920,n2923);
nand (n2920,n2921,n2922);
or (n2921,n16,n2898);
or (n2922,n17,n2821);
xor (n2923,n2924,n2930);
nor (n2924,n2925,n132);
nor (n2925,n2926,n2929);
and (n2926,n2927,n31);
not (n2927,n2928);
and (n2928,n1122,n185);
and (n2929,n1124,n184);
nand (n2930,n2931,n2935);
or (n2931,n940,n2932);
nor (n2932,n2933,n2934);
and (n2933,n335,n84);
and (n2934,n331,n86);
or (n2935,n2793,n941);
or (n2936,n2937,n2952);
and (n2937,n2938,n2943);
xor (n2938,n2939,n2940);
nor (n2939,n187,n1124);
nand (n2940,n2941,n2942);
or (n2941,n940,n2914);
or (n2942,n2932,n941);
nand (n2943,n2944,n2948);
or (n2944,n337,n2945);
nor (n2945,n2946,n2947);
and (n2946,n340,n247);
and (n2947,n341,n249);
or (n2948,n329,n2949);
nor (n2949,n2950,n2951);
and (n2950,n340,n218);
and (n2951,n341,n220);
and (n2952,n2939,n2940);
or (n2953,n2954,n3011);
and (n2954,n2955,n3010);
xor (n2955,n2956,n2985);
or (n2956,n2957,n2984);
and (n2957,n2958,n2975);
xor (n2958,n2959,n2965);
nand (n2959,n2960,n2964);
or (n2960,n337,n2961);
nor (n2961,n2962,n2963);
and (n2962,n340,n241);
and (n2963,n341,n243);
or (n2964,n329,n2945);
nand (n2965,n2966,n2970);
or (n2966,n105,n2967);
nor (n2967,n2968,n2969);
and (n2968,n104,n580);
and (n2969,n100,n582);
or (n2970,n278,n2971);
not (n2971,n2972);
nor (n2972,n2973,n2974);
and (n2973,n312,n100);
and (n2974,n311,n104);
nand (n2975,n2976,n2980);
or (n2976,n369,n2977);
nor (n2977,n2978,n2979);
and (n2978,n377,n712);
and (n2979,n378,n714);
or (n2980,n370,n2981);
nor (n2981,n2982,n2983);
and (n2982,n377,n574);
and (n2983,n378,n576);
and (n2984,n2959,n2965);
or (n2985,n2986,n3009);
and (n2986,n2987,n3003);
xor (n2987,n2988,n2997);
nand (n2988,n2989,n2993);
or (n2989,n352,n2990);
nor (n2990,n2991,n2992);
and (n2991,n110,n166);
and (n2992,n111,n168);
or (n2993,n530,n2994);
nor (n2994,n2995,n2996);
and (n2995,n110,n174);
and (n2996,n111,n173);
nand (n2997,n2998,n3002);
or (n2998,n425,n2999);
nor (n2999,n3000,n3001);
and (n3000,n21,n922);
and (n3001,n22,n924);
or (n3002,n433,n2884);
nand (n3003,n3004,n3005);
or (n3004,n2893,n17);
or (n3005,n16,n3006);
nor (n3006,n3007,n3008);
and (n3007,n1124,n26);
and (n3008,n1122,n31);
and (n3009,n2988,n2997);
xor (n3010,n2938,n2943);
and (n3011,n2956,n2985);
and (n3012,n2879,n2918);
xor (n3013,n3014,n3062);
xor (n3014,n3015,n3018);
or (n3015,n3016,n3017);
and (n3016,n2919,n2936);
and (n3017,n2920,n2923);
xor (n3018,n3019,n3041);
xor (n3019,n3020,n3021);
and (n3020,n2924,n2930);
or (n3021,n3022,n3040);
and (n3022,n3023,n3034);
xor (n3023,n3024,n3028);
nand (n3024,n3025,n3026);
or (n3025,n2799,n329);
nand (n3026,n3027,n336);
not (n3027,n2949);
nand (n3028,n3029,n3033);
or (n3029,n180,n3030);
nor (n3030,n3031,n3032);
and (n3031,n128,n1124);
and (n3032,n132,n1122);
or (n3033,n187,n2831);
nand (n3034,n3035,n3039);
or (n3035,n105,n3036);
nor (n3036,n3037,n3038);
and (n3037,n104,n166);
and (n3038,n100,n168);
or (n3039,n278,n2837);
and (n3040,n3024,n3028);
or (n3041,n3042,n3061);
and (n3042,n3043,n3058);
xor (n3043,n3044,n3051);
nand (n3044,n3045,n3049);
or (n3045,n3046,n369);
nor (n3046,n3047,n3048);
and (n3047,n582,n378);
and (n3048,n580,n377);
nand (n3049,n3050,n707);
not (n3050,n2843);
nand (n3051,n3052,n3056);
or (n3052,n3053,n352);
nor (n3053,n3054,n3055);
and (n3054,n110,n241);
and (n3055,n111,n243);
nand (n3056,n3057,n354);
not (n3057,n2809);
nand (n3058,n3059,n3060);
or (n3059,n425,n2888);
or (n3060,n433,n2815);
and (n3061,n3044,n3051);
or (n3062,n3063,n3081);
and (n3063,n3064,n3080);
xor (n3064,n3065,n3079);
or (n3065,n3066,n3078);
and (n3066,n3067,n3075);
xor (n3067,n3068,n3072);
nand (n3068,n3069,n3070);
or (n3069,n2971,n105);
nand (n3070,n3071,n107);
not (n3071,n3036);
nand (n3072,n3073,n3074);
or (n3073,n369,n2981);
or (n3074,n370,n3046);
nand (n3075,n3076,n3077);
or (n3076,n352,n2994);
or (n3077,n530,n3053);
and (n3078,n3068,n3072);
xor (n3079,n3043,n3058);
xor (n3080,n3023,n3034);
and (n3081,n3065,n3079);
or (n3082,n3083,n3139);
and (n3083,n3084,n3138);
xor (n3084,n3085,n3086);
xor (n3085,n3064,n3080);
or (n3086,n3087,n3137);
and (n3087,n3088,n3091);
xor (n3088,n3089,n3090);
xor (n3089,n3067,n3075);
xor (n3090,n2881,n2901);
or (n3091,n3092,n3136);
and (n3092,n3093,n3113);
xor (n3093,n3094,n3095);
xor (n3094,n2902,n2908);
or (n3095,n3096,n3112);
and (n3096,n3097,n3106);
xor (n3097,n3098,n3099);
nor (n3098,n17,n1124);
nand (n3099,n3100,n3105);
or (n3100,n3101,n337);
not (n3101,n3102);
nand (n3102,n3103,n3104);
or (n3103,n341,n173);
or (n3104,n340,n174);
or (n3105,n329,n2961);
nand (n3106,n3107,n3111);
or (n3107,n105,n3108);
nor (n3108,n3109,n3110);
and (n3109,n104,n574);
and (n3110,n100,n576);
or (n3111,n278,n2967);
and (n3112,n3098,n3099);
or (n3113,n3114,n3135);
and (n3114,n3115,n3129);
xor (n3115,n3116,n3122);
nand (n3116,n3117,n3121);
or (n3117,n369,n3118);
nor (n3118,n3119,n3120);
and (n3119,n377,n753);
and (n3120,n378,n755);
or (n3121,n370,n2977);
nand (n3122,n3123,n3128);
or (n3123,n940,n3124);
not (n3124,n3125);
nor (n3125,n3126,n3127);
and (n3126,n247,n331);
and (n3127,n249,n335);
or (n3128,n2910,n941);
nand (n3129,n3130,n3134);
or (n3130,n425,n3131);
nor (n3131,n3132,n3133);
and (n3132,n21,n959);
and (n3133,n22,n961);
or (n3134,n433,n2999);
and (n3135,n3116,n3122);
and (n3136,n3094,n3095);
and (n3137,n3089,n3090);
xor (n3138,n2878,n2953);
and (n3139,n3085,n3086);
not (n3140,n3141);
nand (n3141,n3142,n3157);
xor (n3142,n3143,n3148);
xor (n3143,n3144,n3145);
xor (n3144,n2851,n2854);
or (n3145,n3146,n3147);
and (n3146,n3014,n3062);
and (n3147,n3015,n3018);
xor (n3148,n3149,n3154);
xor (n3149,n3150,n3153);
or (n3150,n3151,n3152);
and (n3151,n3019,n3041);
and (n3152,n3020,n3021);
xor (n3153,n2785,n2826);
or (n3154,n3155,n3156);
and (n3155,n2872,n2875);
and (n3156,n2873,n2874);
or (n3157,n3158,n3159);
and (n3158,n2870,n3013);
and (n3159,n2871,n2876);
nand (n3160,n3161,n3162);
not (n3161,n3142);
not (n3162,n3157);
not (n3163,n3164);
nor (n3164,n3165,n3172);
xor (n3165,n3166,n3171);
xor (n3166,n3167,n3168);
xor (n3167,n2750,n2769);
or (n3168,n3169,n3170);
and (n3169,n3149,n3154);
and (n3170,n3150,n3153);
xor (n3171,n2782,n2856);
or (n3172,n3173,n3174);
and (n3173,n3143,n3148);
and (n3174,n3144,n3145);
and (n3175,n3165,n3172);
nor (n3176,n3177,n3178);
xor (n3177,n2778,n2858);
or (n3178,n3179,n3180);
and (n3179,n3166,n3171);
and (n3180,n3167,n3168);
nand (n3181,n3177,n3178);
nor (n3182,n3183,n3308);
nor (n3183,n3184,n3305);
xor (n3184,n3185,n3302);
xor (n3185,n3186,n3203);
xor (n3186,n3187,n3200);
xor (n3187,n3188,n3191);
or (n3188,n3189,n3190);
and (n3189,n2627,n2634);
and (n3190,n2628,n2631);
xor (n3191,n3192,n3197);
xor (n3192,n3193,n3194);
and (n3193,n2611,n2617);
or (n3194,n3195,n3196);
and (n3195,n2635,n2648);
and (n3196,n2636,n2642);
or (n3197,n3198,n3199);
and (n3198,n2546,n2560);
and (n3199,n2547,n2554);
or (n3200,n3201,n3202);
and (n3201,n2524,n2569);
and (n3202,n2525,n2545);
xor (n3203,n3204,n3299);
xor (n3204,n3205,n3253);
xor (n3205,n3206,n3231);
xor (n3206,n3207,n3210);
or (n3207,n3208,n3209);
and (n3208,n2526,n2539);
and (n3209,n2527,n2533);
xor (n3210,n3211,n3225);
xor (n3211,n3212,n3219);
nand (n3212,n3213,n3215);
or (n3213,n3214,n352);
not (n3214,n2645);
nand (n3215,n354,n3216);
nor (n3216,n3217,n3218);
and (n3217,n260,n111);
and (n3218,n262,n110);
nand (n3219,n3220,n3221);
or (n3220,n425,n2651);
or (n3221,n3222,n433);
nor (n3222,n3223,n3224);
and (n3223,n21,n218);
and (n3224,n22,n220);
nand (n3225,n3226,n3227);
or (n3226,n16,n2607);
or (n3227,n17,n3228);
nor (n3228,n3229,n3230);
and (n3229,n31,n241);
and (n3230,n26,n243);
xor (n3231,n3232,n3246);
xor (n3232,n3233,n3240);
nand (n3233,n3234,n3236);
or (n3234,n3235,n180);
not (n3235,n2536);
nand (n3236,n3237,n188);
nor (n3237,n3238,n3239);
and (n3238,n166,n128);
and (n3239,n168,n132);
nand (n3240,n3241,n3242);
or (n3241,n125,n2542);
or (n3242,n126,n3243);
nor (n3243,n3244,n3245);
and (n3244,n135,n580);
and (n3245,n136,n582);
nand (n3246,n3247,n3248);
or (n3247,n369,n2551);
or (n3248,n370,n3249);
not (n3249,n3250);
nand (n3250,n3251,n3252);
or (n3251,n378,n86);
or (n3252,n377,n84);
xor (n3253,n3254,n3296);
xor (n3254,n3255,n3278);
xor (n3255,n3256,n3272);
xor (n3256,n3257,n3264);
nand (n3257,n3258,n3260);
or (n3258,n3259,n408);
not (n3259,n2557);
nand (n3260,n3261,n419);
nor (n3261,n3262,n3263);
and (n3262,n714,n407);
and (n3263,n712,n47);
nand (n3264,n3265,n3270);
or (n3265,n3266,n62);
not (n3266,n3267);
nand (n3267,n3268,n3269);
or (n3268,n54,n924);
or (n3269,n53,n922);
nand (n3270,n3271,n44);
not (n3271,n2566);
nand (n3272,n3273,n3274);
or (n3273,n940,n2639);
or (n3274,n3275,n941);
nor (n3275,n3276,n3277);
and (n3276,n193,n331);
and (n3277,n194,n335);
xor (n3278,n3279,n3289);
xor (n3279,n3280,n3281);
nor (n3280,n72,n1124);
nand (n3281,n3282,n3284);
or (n3282,n3283,n337);
not (n3283,n2620);
nand (n3284,n3285,n328);
not (n3285,n3286);
nor (n3286,n3287,n3288);
and (n3287,n142,n341);
and (n3288,n140,n340);
nand (n3289,n3290,n3292);
or (n3290,n3291,n105);
not (n3291,n2530);
nand (n3292,n107,n3293);
nand (n3293,n3294,n3295);
or (n3294,n100,n60);
or (n3295,n104,n58);
or (n3296,n3297,n3298);
and (n3297,n2603,n2623);
and (n3298,n2604,n2610);
or (n3299,n3300,n3301);
and (n3300,n2573,n2626);
and (n3301,n2574,n2602);
or (n3302,n3303,n3304);
and (n3303,n2448,n2572);
and (n3304,n2449,n2523);
or (n3305,n3306,n3307);
and (n3306,n2274,n2654);
and (n3307,n2275,n2447);
nor (n3308,n3309,n3312);
or (n3309,n3310,n3311);
and (n3310,n3185,n3302);
and (n3311,n3186,n3203);
xor (n3312,n3313,n3320);
xor (n3313,n3314,n3317);
or (n3314,n3315,n3316);
and (n3315,n3187,n3200);
and (n3316,n3188,n3191);
or (n3317,n3318,n3319);
and (n3318,n3204,n3299);
and (n3319,n3205,n3253);
xor (n3320,n3321,n3381);
xor (n3321,n3322,n3378);
xor (n3322,n3323,n3375);
xor (n3323,n3324,n3347);
xor (n3324,n3325,n3341);
xor (n3325,n3326,n3334);
nand (n3326,n3327,n3329);
or (n3327,n3328,n105);
not (n3328,n3293);
nand (n3329,n3330,n107);
not (n3330,n3331);
nor (n3331,n3332,n3333);
and (n3332,n104,n65);
and (n3333,n100,n67);
nand (n3334,n3335,n3337);
or (n3335,n180,n3336);
not (n3336,n3237);
or (n3337,n187,n3338);
nor (n3338,n3339,n3340);
and (n3339,n132,n174);
and (n3340,n128,n173);
nand (n3341,n3342,n3343);
or (n3342,n125,n3243);
or (n3343,n126,n3344);
nor (n3344,n3345,n3346);
and (n3345,n135,n312);
and (n3346,n136,n311);
xor (n3347,n3348,n3361);
xor (n3348,n3349,n3355);
nand (n3349,n3350,n3351);
or (n3350,n425,n3222);
or (n3351,n433,n3352);
nor (n3352,n3353,n3354);
and (n3353,n21,n224);
and (n3354,n22,n226);
nand (n3355,n3356,n3357);
or (n3356,n16,n3228);
or (n3357,n17,n3358);
nor (n3358,n3359,n3360);
and (n3359,n31,n247);
and (n3360,n26,n249);
xor (n3361,n3362,n3368);
nor (n3362,n3363,n79);
nor (n3363,n3364,n3367);
and (n3364,n3365,n53);
not (n3365,n3366);
and (n3366,n1122,n75);
and (n3367,n1124,n74);
nand (n3368,n3369,n3374);
or (n3369,n3370,n329);
not (n3370,n3371);
nand (n3371,n3372,n3373);
or (n3372,n341,n148);
or (n3373,n340,n146);
or (n3374,n337,n3286);
or (n3375,n3376,n3377);
and (n3376,n3192,n3197);
and (n3377,n3193,n3194);
or (n3378,n3379,n3380);
and (n3379,n3254,n3296);
and (n3380,n3255,n3278);
xor (n3381,n3382,n3397);
xor (n3382,n3383,n3394);
xor (n3383,n3384,n3391);
xor (n3384,n3385,n3388);
or (n3385,n3386,n3387);
and (n3386,n3256,n3272);
and (n3387,n3257,n3264);
or (n3388,n3389,n3390);
and (n3389,n3211,n3225);
and (n3390,n3212,n3219);
or (n3391,n3392,n3393);
and (n3392,n3279,n3289);
and (n3393,n3280,n3281);
or (n3394,n3395,n3396);
and (n3395,n3206,n3231);
and (n3396,n3207,n3210);
xor (n3397,n3398,n3426);
xor (n3398,n3399,n3402);
or (n3399,n3400,n3401);
and (n3400,n3232,n3246);
and (n3401,n3233,n3240);
xor (n3402,n3403,n3417);
xor (n3403,n3404,n3410);
nand (n3404,n3405,n3406);
or (n3405,n940,n3275);
or (n3406,n3407,n941);
nor (n3407,n3408,n3409);
and (n3408,n199,n335);
and (n3409,n201,n331);
nand (n3410,n3411,n3413);
or (n3411,n3412,n352);
not (n3412,n3216);
nand (n3413,n354,n3414);
nand (n3414,n3415,n3416);
or (n3415,n111,n268);
or (n3416,n110,n266);
nand (n3417,n3418,n3422);
or (n3418,n70,n3419);
nor (n3419,n3420,n3421);
and (n3420,n1124,n80);
and (n3421,n1122,n79);
or (n3422,n72,n3423);
nor (n3423,n3424,n3425);
and (n3424,n959,n79);
and (n3425,n80,n961);
xor (n3426,n3427,n3442);
xor (n3427,n3428,n3435);
nand (n3428,n3429,n3434);
or (n3429,n3430,n370);
not (n3430,n3431);
nand (n3431,n3432,n3433);
or (n3432,n378,n92);
or (n3433,n377,n90);
nand (n3434,n986,n3250);
nand (n3435,n3436,n3438);
or (n3436,n408,n3437);
not (n3437,n3261);
or (n3438,n415,n3439);
nor (n3439,n3440,n3441);
and (n3440,n407,n574);
and (n3441,n47,n576);
nand (n3442,n3443,n3444);
or (n3443,n43,n3266);
or (n3444,n62,n3445);
nor (n3445,n3446,n3447);
and (n3446,n53,n753);
and (n3447,n54,n755);
nand (n3448,n3449,n3456);
or (n3449,n3450,n3451);
not (n3450,n3182);
not (n3451,n3452);
nand (n3452,n3453,n3455);
or (n3453,n2272,n3454);
nand (n3454,n2775,n2776);
nand (n3455,n2273,n2661);
nor (n3456,n3457,n3461);
and (n3457,n3458,n3460);
not (n3458,n3459);
nand (n3459,n3184,n3305);
not (n3460,n3308);
and (n3461,n3309,n3312);
nand (n3462,n2271,n3182,n3463,n3467);
and (n3463,n3464,n3465,n3163);
not (n3464,n3176);
and (n3465,n3160,n3466);
or (n3466,n3082,n2869);
nand (n3467,n3468,n3971,n3980);
nand (n3468,n3469,n3905,n3964);
or (n3469,n3470,n3904);
and (n3470,n3471,n3647);
xor (n3471,n3472,n3595);
or (n3472,n3473,n3594);
and (n3473,n3474,n3555);
xor (n3474,n3475,n3504);
xor (n3475,n3476,n3495);
xor (n3476,n3477,n3486);
nand (n3477,n3478,n3482);
or (n3478,n369,n3479);
nor (n3479,n3480,n3481);
and (n3480,n377,n959);
and (n3481,n378,n961);
or (n3482,n370,n3483);
nor (n3483,n3484,n3485);
and (n3484,n377,n922);
and (n3485,n378,n924);
nand (n3486,n3487,n3491);
or (n3487,n3488,n940);
nor (n3488,n3489,n3490);
and (n3489,n335,n174);
and (n3490,n331,n173);
or (n3491,n3492,n941);
nor (n3492,n3493,n3494);
and (n3493,n335,n241);
and (n3494,n331,n243);
nand (n3495,n3496,n3500);
or (n3496,n352,n3497);
nor (n3497,n3498,n3499);
and (n3498,n110,n574);
and (n3499,n111,n576);
or (n3500,n530,n3501);
nor (n3501,n3502,n3503);
and (n3502,n110,n580);
and (n3503,n111,n582);
or (n3504,n3505,n3554);
and (n3505,n3506,n3529);
xor (n3506,n3507,n3513);
nand (n3507,n3508,n3512);
or (n3508,n352,n3509);
nor (n3509,n3510,n3511);
and (n3510,n110,n712);
and (n3511,n111,n714);
or (n3512,n530,n3497);
xor (n3513,n3514,n3520);
and (n3514,n3515,n378);
nand (n3515,n3516,n3517);
or (n3516,n1122,n373);
nand (n3517,n3518,n104);
not (n3518,n3519);
and (n3519,n1122,n373);
nand (n3520,n3521,n3525);
or (n3521,n337,n3522);
nor (n3522,n3523,n3524);
and (n3523,n340,n580);
and (n3524,n341,n582);
or (n3525,n329,n3526);
nor (n3526,n3527,n3528);
and (n3527,n340,n312);
and (n3528,n341,n311);
or (n3529,n3530,n3553);
and (n3530,n3531,n3542);
xor (n3531,n3532,n3533);
and (n3532,n707,n1122);
nand (n3533,n3534,n3538);
or (n3534,n940,n3535);
nor (n3535,n3536,n3537);
and (n3536,n335,n312);
and (n3537,n331,n311);
or (n3538,n3539,n941);
nor (n3539,n3540,n3541);
and (n3540,n335,n166);
and (n3541,n331,n168);
nand (n3542,n3543,n3548);
or (n3543,n3544,n105);
not (n3544,n3545);
nor (n3545,n3546,n3547);
and (n3546,n959,n100);
and (n3547,n961,n104);
nand (n3548,n3549,n107);
not (n3549,n3550);
nor (n3550,n3551,n3552);
and (n3551,n104,n922);
and (n3552,n100,n924);
and (n3553,n3532,n3533);
and (n3554,n3507,n3513);
xor (n3555,n3556,n3579);
xor (n3556,n3557,n3558);
and (n3557,n3514,n3520);
or (n3558,n3559,n3578);
and (n3559,n3560,n3575);
xor (n3560,n3561,n3567);
nand (n3561,n3562,n3563);
or (n3562,n105,n3550);
or (n3563,n278,n3564);
nor (n3564,n3565,n3566);
and (n3565,n104,n753);
and (n3566,n100,n755);
nand (n3567,n3568,n3573);
or (n3568,n3569,n369);
not (n3569,n3570);
nand (n3570,n3571,n3572);
or (n3571,n377,n1122);
or (n3572,n1124,n378);
nand (n3573,n3574,n707);
not (n3574,n3479);
nand (n3575,n3576,n3577);
or (n3576,n940,n3539);
or (n3577,n3488,n941);
and (n3578,n3561,n3567);
xor (n3579,n3580,n3588);
xor (n3580,n3581,n3582);
nor (n3581,n433,n1124);
nand (n3582,n3583,n3584);
or (n3583,n337,n3526);
or (n3584,n329,n3585);
nor (n3585,n3586,n3587);
and (n3586,n340,n166);
and (n3587,n341,n168);
nand (n3588,n3589,n3590);
or (n3589,n105,n3564);
or (n3590,n278,n3591);
nor (n3591,n3592,n3593);
and (n3592,n104,n712);
and (n3593,n100,n714);
and (n3594,n3475,n3504);
xor (n3595,n3596,n3644);
xor (n3596,n3597,n3625);
xor (n3597,n3598,n3611);
xor (n3598,n3599,n3605);
nand (n3599,n3600,n3604);
or (n3600,n425,n3601);
nor (n3601,n3602,n3603);
and (n3602,n1124,n22);
and (n3603,n21,n1122);
or (n3604,n433,n3131);
nand (n3605,n3606,n3607);
or (n3606,n352,n3501);
or (n3607,n530,n3608);
nor (n3608,n3609,n3610);
and (n3609,n110,n312);
and (n3610,n111,n311);
nand (n3611,n3612,n3624);
or (n3612,n3613,n3620);
not (n3613,n3614);
nand (n3614,n3615,n22);
nand (n3615,n3616,n3617);
or (n3616,n1122,n429);
nand (n3617,n3618,n377);
not (n3618,n3619);
and (n3619,n1122,n429);
not (n3620,n3621);
nand (n3621,n3622,n3623);
or (n3622,n337,n3585);
or (n3623,n329,n3101);
or (n3624,n3621,n3614);
xor (n3625,n3626,n3633);
xor (n3626,n3627,n3630);
or (n3627,n3628,n3629);
and (n3628,n3580,n3588);
and (n3629,n3581,n3582);
or (n3630,n3631,n3632);
and (n3631,n3476,n3495);
and (n3632,n3477,n3486);
xor (n3633,n3634,n3641);
xor (n3634,n3635,n3638);
nand (n3635,n3636,n3637);
or (n3636,n105,n3591);
or (n3637,n278,n3108);
nand (n3638,n3639,n3640);
or (n3639,n369,n3483);
or (n3640,n370,n3118);
nand (n3641,n3642,n3643);
or (n3642,n941,n3124);
or (n3643,n3492,n940);
or (n3644,n3645,n3646);
and (n3645,n3556,n3579);
and (n3646,n3557,n3558);
or (n3647,n3648,n3903);
and (n3648,n3649,n3689);
xor (n3649,n3650,n3688);
or (n3650,n3651,n3687);
and (n3651,n3652,n3686);
xor (n3652,n3653,n3654);
xor (n3653,n3560,n3575);
or (n3654,n3655,n3685);
and (n3655,n3656,n3671);
xor (n3656,n3657,n3663);
nand (n3657,n3658,n3662);
or (n3658,n337,n3659);
nor (n3659,n3660,n3661);
and (n3660,n576,n341);
and (n3661,n574,n340);
or (n3662,n329,n3522);
nand (n3663,n3664,n3669);
or (n3664,n3665,n352);
not (n3665,n3666);
nand (n3666,n3667,n3668);
or (n3667,n111,n755);
or (n3668,n110,n753);
nand (n3669,n3670,n354);
not (n3670,n3509);
and (n3671,n3672,n3678);
nor (n3672,n3673,n104);
nor (n3673,n3674,n3677);
and (n3674,n3675,n110);
not (n3675,n3676);
and (n3676,n1122,n109);
and (n3677,n1124,n116);
nand (n3678,n3679,n3684);
or (n3679,n940,n3680);
not (n3680,n3681);
nor (n3681,n3682,n3683);
and (n3682,n582,n335);
and (n3683,n580,n331);
or (n3684,n3535,n941);
and (n3685,n3657,n3663);
xor (n3686,n3506,n3529);
and (n3687,n3653,n3654);
xor (n3688,n3474,n3555);
or (n3689,n3690,n3902);
and (n3690,n3691,n3725);
xor (n3691,n3692,n3724);
or (n3692,n3693,n3723);
and (n3693,n3694,n3722);
xor (n3694,n3695,n3721);
or (n3695,n3696,n3720);
and (n3696,n3697,n3713);
xor (n3697,n3698,n3705);
nand (n3698,n3699,n3704);
or (n3699,n3700,n105);
not (n3700,n3701);
nand (n3701,n3702,n3703);
or (n3702,n104,n1122);
or (n3703,n1124,n100);
nand (n3704,n107,n3545);
nand (n3705,n3706,n3711);
or (n3706,n3707,n337);
not (n3707,n3708);
nor (n3708,n3709,n3710);
and (n3709,n714,n340);
and (n3710,n712,n341);
nand (n3711,n3712,n328);
not (n3712,n3659);
nand (n3713,n3714,n3719);
or (n3714,n3715,n352);
not (n3715,n3716);
nor (n3716,n3717,n3718);
and (n3717,n922,n111);
and (n3718,n924,n110);
nand (n3719,n354,n3666);
and (n3720,n3698,n3705);
xor (n3721,n3531,n3542);
xor (n3722,n3656,n3671);
and (n3723,n3695,n3721);
xor (n3724,n3652,n3686);
nand (n3725,n3726,n3901);
or (n3726,n3727,n3757);
not (n3727,n3728);
nand (n3728,n3729,n3731);
not (n3729,n3730);
xor (n3730,n3694,n3722);
not (n3731,n3732);
or (n3732,n3733,n3756);
and (n3733,n3734,n3755);
xor (n3734,n3735,n3736);
xor (n3735,n3672,n3678);
or (n3736,n3737,n3754);
and (n3737,n3738,n3747);
xor (n3738,n3739,n3740);
and (n3739,n107,n1122);
nand (n3740,n3741,n3746);
or (n3741,n940,n3742);
not (n3742,n3743);
nor (n3743,n3744,n3745);
and (n3744,n574,n331);
and (n3745,n576,n335);
nand (n3746,n3681,n942);
nand (n3747,n3748,n3753);
or (n3748,n3749,n337);
not (n3749,n3750);
nor (n3750,n3751,n3752);
and (n3751,n755,n340);
and (n3752,n753,n341);
nand (n3753,n328,n3708);
and (n3754,n3739,n3740);
xor (n3755,n3697,n3713);
and (n3756,n3735,n3736);
not (n3757,n3758);
nand (n3758,n3759,n3900);
or (n3759,n3760,n3790);
not (n3760,n3761);
nand (n3761,n3762,n3764);
not (n3762,n3763);
xor (n3763,n3734,n3755);
not (n3764,n3765);
or (n3765,n3766,n3789);
and (n3766,n3767,n3788);
xor (n3767,n3768,n3775);
nand (n3768,n3769,n3774);
or (n3769,n3770,n352);
not (n3770,n3771);
nor (n3771,n3772,n3773);
and (n3772,n959,n111);
and (n3773,n961,n110);
nand (n3774,n354,n3716);
and (n3775,n3776,n3781);
and (n3776,n3777,n111);
nand (n3777,n3778,n3780);
or (n3778,n3779,n341);
and (n3779,n1122,n356);
or (n3780,n1122,n356);
nand (n3781,n3782,n3783);
or (n3782,n941,n3742);
nand (n3783,n3784,n939);
not (n3784,n3785);
nor (n3785,n3786,n3787);
and (n3786,n712,n335);
and (n3787,n714,n331);
xor (n3788,n3738,n3747);
and (n3789,n3768,n3775);
not (n3790,n3791);
nand (n3791,n3792,n3899);
or (n3792,n3793,n3817);
not (n3793,n3794);
nand (n3794,n3795,n3797);
not (n3795,n3796);
xor (n3796,n3767,n3788);
not (n3797,n3798);
or (n3798,n3799,n3816);
and (n3799,n3800,n3815);
xor (n3800,n3801,n3808);
nand (n3801,n3802,n3807);
or (n3802,n3803,n337);
not (n3803,n3804);
nor (n3804,n3805,n3806);
and (n3805,n924,n340);
and (n3806,n922,n341);
nand (n3807,n328,n3750);
nand (n3808,n3809,n3814);
or (n3809,n3810,n352);
not (n3810,n3811);
nand (n3811,n3812,n3813);
or (n3812,n110,n1122);
or (n3813,n111,n1124);
nand (n3814,n354,n3771);
xor (n3815,n3776,n3781);
and (n3816,n3801,n3808);
not (n3817,n3818);
nand (n3818,n3819,n3898);
or (n3819,n3820,n3844);
not (n3820,n3821);
nand (n3821,n3822,n3824);
not (n3822,n3823);
xor (n3823,n3800,n3815);
not (n3824,n3825);
or (n3825,n3826,n3843);
and (n3826,n3827,n3836);
xor (n3827,n3828,n3829);
and (n3828,n354,n1122);
nand (n3829,n3830,n3835);
or (n3830,n3831,n337);
not (n3831,n3832);
nor (n3832,n3833,n3834);
and (n3833,n959,n341);
and (n3834,n961,n340);
nand (n3835,n328,n3804);
nand (n3836,n3837,n3842);
or (n3837,n940,n3838);
not (n3838,n3839);
nor (n3839,n3840,n3841);
and (n3840,n755,n335);
and (n3841,n753,n331);
or (n3842,n3785,n941);
and (n3843,n3828,n3829);
not (n3844,n3845);
nand (n3845,n3846,n3897);
or (n3846,n3847,n3863);
nor (n3847,n3848,n3849);
xor (n3848,n3827,n3836);
and (n3849,n3850,n3856);
nor (n3850,n3851,n340);
nor (n3851,n3852,n3853);
and (n3852,n332,n1124);
and (n3853,n3854,n335);
not (n3854,n3855);
and (n3855,n1122,n333);
nand (n3856,n3857,n3858);
or (n3857,n941,n3838);
nand (n3858,n3859,n939);
not (n3859,n3860);
nor (n3860,n3861,n3862);
and (n3861,n335,n922);
and (n3862,n331,n924);
not (n3863,n3864);
or (n3864,n3865,n3896);
and (n3865,n3866,n3875);
xor (n3866,n3867,n3874);
nand (n3867,n3868,n3873);
or (n3868,n3869,n337);
not (n3869,n3870);
nand (n3870,n3871,n3872);
or (n3871,n340,n1122);
or (n3872,n341,n1124);
nand (n3873,n328,n3832);
xor (n3874,n3850,n3856);
or (n3875,n3876,n3895);
and (n3876,n3877,n3885);
xor (n3877,n3878,n3879);
nor (n3878,n329,n1124);
nand (n3879,n3880,n3884);
or (n3880,n3881,n940);
nor (n3881,n3882,n3883);
and (n3882,n335,n959);
and (n3883,n331,n961);
or (n3884,n3860,n941);
nor (n3885,n3886,n3893);
nor (n3886,n3887,n3889);
and (n3887,n3888,n942);
not (n3888,n3881);
nor (n3889,n3890,n940);
nor (n3890,n3891,n3892);
and (n3891,n1122,n335);
and (n3892,n1124,n331);
or (n3893,n3894,n335);
and (n3894,n1122,n942);
and (n3895,n3878,n3879);
and (n3896,n3867,n3874);
nand (n3897,n3848,n3849);
nand (n3898,n3823,n3825);
nand (n3899,n3796,n3798);
nand (n3900,n3763,n3765);
nand (n3901,n3730,n3732);
and (n3902,n3692,n3724);
and (n3903,n3650,n3688);
and (n3904,n3472,n3595);
nor (n3905,n3906,n3946);
not (n3906,n3907);
nand (n3907,n3908,n3930);
not (n3908,n3909);
xor (n3909,n3910,n3913);
xor (n3910,n3911,n3912);
xor (n3911,n2955,n3010);
xor (n3912,n3088,n3091);
or (n3913,n3914,n3929);
and (n3914,n3915,n3918);
xor (n3915,n3916,n3917);
xor (n3916,n2987,n3003);
xor (n3917,n2958,n2975);
or (n3918,n3919,n3928);
and (n3919,n3920,n3925);
xor (n3920,n3921,n3924);
nand (n3921,n3922,n3923);
or (n3922,n352,n3608);
or (n3923,n530,n2990);
and (n3924,n3621,n3613);
or (n3925,n3926,n3927);
and (n3926,n3634,n3641);
and (n3927,n3635,n3638);
and (n3928,n3921,n3924);
and (n3929,n3916,n3917);
not (n3930,n3931);
or (n3931,n3932,n3945);
and (n3932,n3933,n3944);
xor (n3933,n3934,n3935);
xor (n3934,n3093,n3113);
or (n3935,n3936,n3943);
and (n3936,n3937,n3940);
xor (n3937,n3938,n3939);
xor (n3938,n3115,n3129);
xor (n3939,n3097,n3106);
or (n3940,n3941,n3942);
and (n3941,n3598,n3611);
and (n3942,n3599,n3605);
and (n3943,n3938,n3939);
xor (n3944,n3915,n3918);
and (n3945,n3934,n3935);
nand (n3946,n3947,n3959);
not (n3947,n3948);
nor (n3948,n3949,n3950);
xor (n3949,n3933,n3944);
or (n3950,n3951,n3958);
and (n3951,n3952,n3957);
xor (n3952,n3953,n3954);
xor (n3953,n3920,n3925);
or (n3954,n3955,n3956);
and (n3955,n3626,n3633);
and (n3956,n3627,n3630);
xor (n3957,n3937,n3940);
and (n3958,n3953,n3954);
or (n3959,n3960,n3963);
or (n3960,n3961,n3962);
and (n3961,n3596,n3644);
and (n3962,n3597,n3625);
xor (n3963,n3952,n3957);
nand (n3964,n3965,n3967);
not (n3965,n3966);
xor (n3966,n3084,n3138);
not (n3967,n3968);
or (n3968,n3969,n3970);
and (n3969,n3910,n3913);
and (n3970,n3911,n3912);
nand (n3971,n3972,n3964);
nand (n3972,n3973,n3979);
or (n3973,n3906,n3974);
not (n3974,n3975);
nand (n3975,n3976,n3978);
or (n3976,n3948,n3977);
nand (n3977,n3960,n3963);
nand (n3978,n3949,n3950);
nand (n3979,n3909,n3931);
nand (n3980,n3966,n3968);
and (n3981,n3982,n4148,n4179);
nand (n3982,n3983,n4116);
not (n3983,n3984);
xor (n3984,n3985,n4103);
xor (n3985,n3986,n3987);
xor (n3986,n2254,n2263);
or (n3987,n3988,n4102);
and (n3988,n3989,n4085);
xor (n3989,n3990,n4062);
or (n3990,n3991,n4061);
and (n3991,n3992,n4033);
xor (n3992,n3993,n4004);
or (n3993,n3994,n4003);
and (n3994,n3995,n4000);
xor (n3995,n3996,n3999);
nand (n3996,n3997,n3998);
or (n3997,n16,n3358);
or (n3998,n17,n2236);
and (n3999,n3362,n3368);
or (n4000,n4001,n4002);
and (n4001,n3427,n3442);
and (n4002,n3428,n3435);
and (n4003,n3996,n3999);
xor (n4004,n4005,n4032);
xor (n4005,n4006,n4021);
or (n4006,n4007,n4020);
and (n4007,n4008,n4017);
xor (n4008,n4009,n4014);
nand (n4009,n4010,n4012);
or (n4010,n4011,n352);
not (n4011,n3414);
nand (n4012,n4013,n354);
not (n4013,n2230);
nand (n4014,n4015,n4016);
or (n4015,n70,n3423);
or (n4016,n72,n2211);
nand (n4017,n4018,n4019);
or (n4018,n425,n3352);
or (n4019,n433,n2204);
and (n4020,n4009,n4014);
or (n4021,n4022,n4031);
and (n4022,n4023,n4028);
xor (n4023,n4024,n4025);
nor (n4024,n227,n1124);
nand (n4025,n4026,n4027);
or (n4026,n3370,n337);
or (n4027,n329,n2134);
nand (n4028,n4029,n4030);
or (n4029,n105,n3331);
or (n4030,n278,n2152);
and (n4031,n4024,n4025);
xor (n4032,n2221,n2234);
or (n4033,n4034,n4060);
and (n4034,n4035,n4049);
xor (n4035,n4036,n4048);
xor (n4036,n4037,n4045);
xor (n4037,n4038,n4042);
nand (n4038,n4039,n4040);
or (n4039,n3439,n408);
nand (n4040,n4041,n419);
not (n4041,n2181);
nand (n4042,n4043,n4044);
or (n4043,n43,n3445);
or (n4044,n62,n2188);
nand (n4045,n4046,n4047);
or (n4046,n940,n3407);
or (n4047,n2198,n941);
xor (n4048,n4023,n4028);
xor (n4049,n4050,n4057);
xor (n4050,n4051,n4054);
nand (n4051,n4052,n4053);
or (n4052,n180,n3338);
or (n4053,n187,n2159);
nand (n4054,n4055,n4056);
or (n4055,n125,n3344);
or (n4056,n126,n2165);
nand (n4057,n4058,n4059);
or (n4058,n369,n3430);
or (n4059,n370,n2175);
and (n4060,n4036,n4048);
and (n4061,n3993,n4004);
xor (n4062,n4063,n4078);
xor (n4063,n4064,n4075);
or (n4064,n4065,n4074);
and (n4065,n4066,n4071);
xor (n4066,n4067,n4068);
xor (n4067,n2126,n2132);
or (n4068,n4069,n4070);
and (n4069,n4050,n4057);
and (n4070,n4051,n4054);
or (n4071,n4072,n4073);
and (n4072,n4037,n4045);
and (n4073,n4038,n4042);
and (n4074,n4067,n4068);
or (n4075,n4076,n4077);
and (n4076,n4005,n4032);
and (n4077,n4006,n4021);
or (n4078,n4079,n4084);
and (n4079,n4080,n4083);
xor (n4080,n4081,n4082);
xor (n4081,n2149,n2163);
xor (n4082,n2172,n2186);
xor (n4083,n2195,n2208);
and (n4084,n4081,n4082);
or (n4085,n4086,n4101);
and (n4086,n4087,n4100);
xor (n4087,n4088,n4099);
or (n4088,n4089,n4098);
and (n4089,n4090,n4097);
xor (n4090,n4091,n4094);
or (n4091,n4092,n4093);
and (n4092,n3403,n3417);
and (n4093,n3404,n3410);
or (n4094,n4095,n4096);
and (n4095,n3325,n3341);
and (n4096,n3326,n3334);
xor (n4097,n4008,n4017);
and (n4098,n4091,n4094);
xor (n4099,n4066,n4071);
xor (n4100,n4080,n4083);
and (n4101,n4088,n4099);
and (n4102,n3990,n4062);
xor (n4103,n4104,n4115);
xor (n4104,n4105,n4108);
or (n4105,n4106,n4107);
and (n4106,n4063,n4078);
and (n4107,n4064,n4075);
or (n4108,n4109,n4114);
and (n4109,n4110,n4113);
xor (n4110,n4111,n4112);
xor (n4111,n2146,n2193);
xor (n4112,n2257,n2260);
xor (n4113,n2218,n2242);
and (n4114,n4111,n4112);
xor (n4115,n2143,n2244);
not (n4116,n4117);
or (n4117,n4118,n4147);
and (n4118,n4119,n4146);
xor (n4119,n4120,n4121);
xor (n4120,n4110,n4113);
or (n4121,n4122,n4145);
and (n4122,n4123,n4144);
xor (n4123,n4124,n4135);
or (n4124,n4125,n4134);
and (n4125,n4126,n4133);
xor (n4126,n4127,n4130);
or (n4127,n4128,n4129);
and (n4128,n3348,n3361);
and (n4129,n3349,n3355);
or (n4130,n4131,n4132);
and (n4131,n3384,n3391);
and (n4132,n3385,n3388);
xor (n4133,n3995,n4000);
and (n4134,n4127,n4130);
or (n4135,n4136,n4143);
and (n4136,n4137,n4142);
xor (n4137,n4138,n4139);
xor (n4138,n4090,n4097);
or (n4139,n4140,n4141);
and (n4140,n3398,n3426);
and (n4141,n3399,n3402);
xor (n4142,n4035,n4049);
and (n4143,n4138,n4139);
xor (n4144,n3992,n4033);
and (n4145,n4124,n4135);
xor (n4146,n3989,n4085);
and (n4147,n4120,n4121);
nor (n4148,n4149,n4168);
nor (n4149,n4150,n4165);
xor (n4150,n4151,n4162);
xor (n4151,n4152,n4153);
xor (n4152,n4137,n4142);
xor (n4153,n4154,n4159);
xor (n4154,n4155,n4158);
or (n4155,n4156,n4157);
and (n4156,n3323,n3375);
and (n4157,n3324,n3347);
xor (n4158,n4126,n4133);
or (n4159,n4160,n4161);
and (n4160,n3382,n3397);
and (n4161,n3383,n3394);
or (n4162,n4163,n4164);
and (n4163,n3321,n3381);
and (n4164,n3322,n3378);
or (n4165,n4166,n4167);
and (n4166,n3313,n3320);
and (n4167,n3314,n3317);
nor (n4168,n4169,n4172);
or (n4169,n4170,n4171);
and (n4170,n4151,n4162);
and (n4171,n4152,n4153);
xor (n4172,n4173,n4178);
xor (n4173,n4174,n4175);
xor (n4174,n4087,n4100);
or (n4175,n4176,n4177);
and (n4176,n4154,n4159);
and (n4177,n4155,n4158);
xor (n4178,n4123,n4144);
not (n4179,n4180);
nor (n4180,n4181,n4182);
xor (n4181,n4119,n4146);
or (n4182,n4183,n4184);
and (n4183,n4173,n4178);
and (n4184,n4174,n4175);
nor (n4185,n4186,n4197);
nor (n4186,n4187,n4188);
xor (n4187,n2101,n2266);
or (n4188,n4189,n4196);
and (n4189,n4190,n4195);
xor (n4190,n4191,n4192);
xor (n4191,n2104,n2141);
or (n4192,n4193,n4194);
and (n4193,n4104,n4115);
and (n4194,n4105,n4108);
xor (n4195,n2249,n2252);
and (n4196,n4191,n4192);
nor (n4197,n4198,n4199);
xor (n4198,n4190,n4195);
or (n4199,n4200,n4201);
and (n4200,n3985,n4103);
and (n4201,n3986,n3987);
nand (n4202,n4203,n2081,n4185);
nand (n4203,n4204,n4214);
or (n4204,n4205,n4206);
not (n4205,n3982);
not (n4206,n4207);
nand (n4207,n4208,n4213);
or (n4208,n4209,n4180);
nor (n4209,n4210,n4212);
nor (n4210,n4168,n4211);
nand (n4211,n4150,n4165);
and (n4212,n4169,n4172);
nand (n4213,n4181,n4182);
nand (n4214,n3984,n4117);
nor (n4215,n4216,n4221);
and (n4216,n2081,n4217);
nand (n4217,n4218,n4220);
or (n4218,n4186,n4219);
nand (n4219,n4198,n4199);
nand (n4220,n4187,n4188);
nand (n4221,n4222,n4224);
or (n4222,n2082,n4223);
nand (n4223,n2098,n2099);
nand (n4224,n2083,n2084);
not (n4225,n4226);
nand (n4226,n4227,n4234);
or (n4227,n4228,n4233);
not (n4228,n4229);
nand (n4229,n4230,n4232);
or (n4230,n1648,n4231);
nand (n4231,n1941,n2077);
nand (n4232,n1649,n1650);
not (n4233,n1441);
nor (n4234,n4235,n4239);
and (n4235,n4236,n4237);
not (n4236,n1442);
not (n4237,n4238);
nand (n4238,n1633,n1646);
and (n4239,n1443,n1444);
nand (n4240,n1090,n1091);
or (n4241,n1087,n3);
xor (n4242,n4243,n8031);
xor (n4243,n4244,n8090);
xor (n4244,n4245,n8026);
xor (n4245,n4246,n8083);
xor (n4246,n4247,n8020);
xor (n4247,n4248,n8071);
xor (n4248,n4249,n8014);
xor (n4249,n4250,n8054);
xor (n4250,n4251,n8008);
xor (n4251,n4252,n8032);
xor (n4252,n4253,n8002);
xor (n4253,n4254,n7999);
xor (n4254,n4255,n7998);
xor (n4255,n4256,n7960);
xor (n4256,n4257,n7959);
xor (n4257,n4258,n7914);
xor (n4258,n4259,n7913);
xor (n4259,n4260,n7863);
xor (n4260,n4261,n7862);
xor (n4261,n4262,n7805);
xor (n4262,n4263,n7804);
xor (n4263,n4264,n7742);
xor (n4264,n4265,n7741);
xor (n4265,n4266,n7674);
xor (n4266,n4267,n7673);
xor (n4267,n4268,n7599);
xor (n4268,n4269,n7598);
xor (n4269,n4270,n7517);
xor (n4270,n4271,n7516);
xor (n4271,n4272,n7430);
xor (n4272,n4273,n7429);
xor (n4273,n4274,n7336);
xor (n4274,n4275,n7335);
xor (n4275,n4276,n7237);
xor (n4276,n4277,n7236);
xor (n4277,n4278,n7135);
xor (n4278,n4279,n7134);
xor (n4279,n4280,n7024);
xor (n4280,n4281,n7023);
xor (n4281,n4282,n6906);
xor (n4282,n4283,n6905);
xor (n4283,n4284,n6783);
xor (n4284,n4285,n6782);
xor (n4285,n4286,n6655);
xor (n4286,n4287,n6654);
xor (n4287,n4288,n6520);
xor (n4288,n4289,n6519);
xor (n4289,n4290,n6378);
xor (n4290,n4291,n6377);
xor (n4291,n4292,n6231);
xor (n4292,n4293,n6230);
xor (n4293,n4294,n6078);
xor (n4294,n4295,n6077);
xor (n4295,n4296,n5919);
xor (n4296,n4297,n5918);
xor (n4297,n4298,n5755);
xor (n4298,n4299,n5754);
xor (n4299,n4300,n5584);
xor (n4300,n4301,n5583);
xor (n4301,n4302,n5412);
xor (n4302,n4303,n5411);
xor (n4303,n4304,n5229);
xor (n4304,n4305,n5228);
xor (n4305,n4306,n5047);
xor (n4306,n4307,n5046);
xor (n4307,n4308,n4861);
xor (n4308,n4309,n4860);
xor (n4309,n4310,n4680);
xor (n4310,n4311,n344);
xor (n4311,n4312,n4318);
xor (n4312,n4313,n4317);
xor (n4313,n4314,n4316);
xor (n4314,n4315,n944);
and (n4315,n121,n942);
and (n4316,n4315,n944);
and (n4317,n121,n333);
or (n4318,n4319,n4320);
and (n4319,n4313,n4317);
and (n4320,n4312,n4321);
or (n4321,n4322,n4502);
and (n4322,n4323,n4501);
xor (n4323,n4314,n4324);
or (n4324,n4325,n4327);
and (n4325,n4315,n4326);
and (n4326,n102,n331);
and (n4327,n4328,n4329);
xor (n4328,n4315,n4326);
or (n4329,n4330,n4332);
and (n4330,n4331,n1390);
and (n4331,n102,n942);
and (n4332,n4333,n4334);
xor (n4333,n4331,n1390);
or (n4334,n4335,n4338);
and (n4335,n4336,n4337);
and (n4336,n281,n942);
and (n4337,n274,n331);
and (n4338,n4339,n4340);
xor (n4339,n4336,n4337);
or (n4340,n4341,n4344);
and (n4341,n4342,n4343);
and (n4342,n274,n942);
and (n4343,n469,n331);
and (n4344,n4345,n4346);
xor (n4345,n4342,n4343);
or (n4346,n4347,n4350);
and (n4347,n4348,n4349);
and (n4348,n469,n942);
and (n4349,n386,n331);
and (n4350,n4351,n4352);
xor (n4351,n4348,n4349);
or (n4352,n4353,n4356);
and (n4353,n4354,n4355);
and (n4354,n386,n942);
and (n4355,n38,n331);
and (n4356,n4357,n4358);
xor (n4357,n4354,n4355);
or (n4358,n4359,n4362);
and (n4359,n4360,n4361);
and (n4360,n38,n942);
and (n4361,n32,n331);
and (n4362,n4363,n4364);
xor (n4363,n4360,n4361);
or (n4364,n4365,n4368);
and (n4365,n4366,n4367);
and (n4366,n32,n942);
and (n4367,n199,n331);
and (n4368,n4369,n4370);
xor (n4369,n4366,n4367);
or (n4370,n4371,n4374);
and (n4371,n4372,n4373);
and (n4372,n199,n942);
and (n4373,n194,n331);
and (n4374,n4375,n4376);
xor (n4375,n4372,n4373);
or (n4376,n4377,n4380);
and (n4377,n4378,n4379);
and (n4378,n194,n942);
and (n4379,n146,n331);
and (n4380,n4381,n4382);
xor (n4381,n4378,n4379);
or (n4382,n4383,n4386);
and (n4383,n4384,n4385);
and (n4384,n146,n942);
and (n4385,n140,n331);
and (n4386,n4387,n4388);
xor (n4387,n4384,n4385);
or (n4388,n4389,n4392);
and (n4389,n4390,n4391);
and (n4390,n140,n942);
and (n4391,n266,n331);
and (n4392,n4393,n4394);
xor (n4393,n4390,n4391);
or (n4394,n4395,n4398);
and (n4395,n4396,n4397);
and (n4396,n266,n942);
and (n4397,n260,n331);
and (n4398,n4399,n4400);
xor (n4399,n4396,n4397);
or (n4400,n4401,n4404);
and (n4401,n4402,n4403);
and (n4402,n260,n942);
and (n4403,n65,n331);
and (n4404,n4405,n4406);
xor (n4405,n4402,n4403);
or (n4406,n4407,n4410);
and (n4407,n4408,n4409);
and (n4408,n65,n942);
and (n4409,n58,n331);
and (n4410,n4411,n4412);
xor (n4411,n4408,n4409);
or (n4412,n4413,n4416);
and (n4413,n4414,n4415);
and (n4414,n58,n942);
and (n4415,n90,n331);
and (n4416,n4417,n4418);
xor (n4417,n4414,n4415);
or (n4418,n4419,n4422);
and (n4419,n4420,n4421);
and (n4420,n90,n942);
and (n4421,n84,n331);
and (n4422,n4423,n4424);
xor (n4423,n4420,n4421);
or (n4424,n4425,n4428);
and (n4425,n4426,n4427);
and (n4426,n84,n942);
and (n4427,n224,n331);
and (n4428,n4429,n4430);
xor (n4429,n4426,n4427);
or (n4430,n4431,n4434);
and (n4431,n4432,n4433);
and (n4432,n224,n942);
and (n4433,n218,n331);
and (n4434,n4435,n4436);
xor (n4435,n4432,n4433);
or (n4436,n4437,n4439);
and (n4437,n4438,n3126);
and (n4438,n218,n942);
and (n4439,n4440,n4441);
xor (n4440,n4438,n3126);
or (n4441,n4442,n4445);
and (n4442,n4443,n4444);
and (n4443,n247,n942);
and (n4444,n241,n331);
and (n4445,n4446,n4447);
xor (n4446,n4443,n4444);
or (n4447,n4448,n4451);
and (n4448,n4449,n4450);
and (n4449,n241,n942);
and (n4450,n174,n331);
and (n4451,n4452,n4453);
xor (n4452,n4449,n4450);
or (n4453,n4454,n4457);
and (n4454,n4455,n4456);
and (n4455,n174,n942);
and (n4456,n166,n331);
and (n4457,n4458,n4459);
xor (n4458,n4455,n4456);
or (n4459,n4460,n4463);
and (n4460,n4461,n4462);
and (n4461,n166,n942);
and (n4462,n312,n331);
and (n4463,n4464,n4465);
xor (n4464,n4461,n4462);
or (n4465,n4466,n4468);
and (n4466,n4467,n3683);
and (n4467,n312,n942);
and (n4468,n4469,n4470);
xor (n4469,n4467,n3683);
or (n4470,n4471,n4473);
and (n4471,n4472,n3744);
and (n4472,n580,n942);
and (n4473,n4474,n4475);
xor (n4474,n4472,n3744);
or (n4475,n4476,n4479);
and (n4476,n4477,n4478);
and (n4477,n574,n942);
and (n4478,n712,n331);
and (n4479,n4480,n4481);
xor (n4480,n4477,n4478);
or (n4481,n4482,n4484);
and (n4482,n4483,n3841);
and (n4483,n712,n942);
and (n4484,n4485,n4486);
xor (n4485,n4483,n3841);
or (n4486,n4487,n4490);
and (n4487,n4488,n4489);
and (n4488,n753,n942);
and (n4489,n922,n331);
and (n4490,n4491,n4492);
xor (n4491,n4488,n4489);
or (n4492,n4493,n4496);
and (n4493,n4494,n4495);
and (n4494,n922,n942);
and (n4495,n959,n331);
and (n4496,n4497,n4498);
xor (n4497,n4494,n4495);
and (n4498,n4499,n4500);
and (n4499,n959,n942);
and (n4500,n1122,n331);
and (n4501,n102,n333);
and (n4502,n4503,n4504);
xor (n4503,n4323,n4501);
or (n4504,n4505,n4508);
and (n4505,n4506,n4507);
xor (n4506,n4328,n4329);
and (n4507,n281,n333);
and (n4508,n4509,n4510);
xor (n4509,n4506,n4507);
or (n4510,n4511,n4514);
and (n4511,n4512,n4513);
xor (n4512,n4333,n4334);
and (n4513,n274,n333);
and (n4514,n4515,n4516);
xor (n4515,n4512,n4513);
or (n4516,n4517,n4520);
and (n4517,n4518,n4519);
xor (n4518,n4339,n4340);
and (n4519,n469,n333);
and (n4520,n4521,n4522);
xor (n4521,n4518,n4519);
or (n4522,n4523,n4526);
and (n4523,n4524,n4525);
xor (n4524,n4345,n4346);
and (n4525,n386,n333);
and (n4526,n4527,n4528);
xor (n4527,n4524,n4525);
or (n4528,n4529,n4532);
and (n4529,n4530,n4531);
xor (n4530,n4351,n4352);
and (n4531,n38,n333);
and (n4532,n4533,n4534);
xor (n4533,n4530,n4531);
or (n4534,n4535,n4538);
and (n4535,n4536,n4537);
xor (n4536,n4357,n4358);
and (n4537,n32,n333);
and (n4538,n4539,n4540);
xor (n4539,n4536,n4537);
or (n4540,n4541,n4544);
and (n4541,n4542,n4543);
xor (n4542,n4363,n4364);
and (n4543,n199,n333);
and (n4544,n4545,n4546);
xor (n4545,n4542,n4543);
or (n4546,n4547,n4550);
and (n4547,n4548,n4549);
xor (n4548,n4369,n4370);
and (n4549,n194,n333);
and (n4550,n4551,n4552);
xor (n4551,n4548,n4549);
or (n4552,n4553,n4556);
and (n4553,n4554,n4555);
xor (n4554,n4375,n4376);
and (n4555,n146,n333);
and (n4556,n4557,n4558);
xor (n4557,n4554,n4555);
or (n4558,n4559,n4562);
and (n4559,n4560,n4561);
xor (n4560,n4381,n4382);
and (n4561,n140,n333);
and (n4562,n4563,n4564);
xor (n4563,n4560,n4561);
or (n4564,n4565,n4568);
and (n4565,n4566,n4567);
xor (n4566,n4387,n4388);
and (n4567,n266,n333);
and (n4568,n4569,n4570);
xor (n4569,n4566,n4567);
or (n4570,n4571,n4574);
and (n4571,n4572,n4573);
xor (n4572,n4393,n4394);
and (n4573,n260,n333);
and (n4574,n4575,n4576);
xor (n4575,n4572,n4573);
or (n4576,n4577,n4580);
and (n4577,n4578,n4579);
xor (n4578,n4399,n4400);
and (n4579,n65,n333);
and (n4580,n4581,n4582);
xor (n4581,n4578,n4579);
or (n4582,n4583,n4586);
and (n4583,n4584,n4585);
xor (n4584,n4405,n4406);
and (n4585,n58,n333);
and (n4586,n4587,n4588);
xor (n4587,n4584,n4585);
or (n4588,n4589,n4592);
and (n4589,n4590,n4591);
xor (n4590,n4411,n4412);
and (n4591,n90,n333);
and (n4592,n4593,n4594);
xor (n4593,n4590,n4591);
or (n4594,n4595,n4598);
and (n4595,n4596,n4597);
xor (n4596,n4417,n4418);
and (n4597,n84,n333);
and (n4598,n4599,n4600);
xor (n4599,n4596,n4597);
or (n4600,n4601,n4604);
and (n4601,n4602,n4603);
xor (n4602,n4423,n4424);
and (n4603,n224,n333);
and (n4604,n4605,n4606);
xor (n4605,n4602,n4603);
or (n4606,n4607,n4610);
and (n4607,n4608,n4609);
xor (n4608,n4429,n4430);
and (n4609,n218,n333);
and (n4610,n4611,n4612);
xor (n4611,n4608,n4609);
or (n4612,n4613,n4616);
and (n4613,n4614,n4615);
xor (n4614,n4435,n4436);
and (n4615,n247,n333);
and (n4616,n4617,n4618);
xor (n4617,n4614,n4615);
or (n4618,n4619,n4622);
and (n4619,n4620,n4621);
xor (n4620,n4440,n4441);
and (n4621,n241,n333);
and (n4622,n4623,n4624);
xor (n4623,n4620,n4621);
or (n4624,n4625,n4628);
and (n4625,n4626,n4627);
xor (n4626,n4446,n4447);
and (n4627,n174,n333);
and (n4628,n4629,n4630);
xor (n4629,n4626,n4627);
or (n4630,n4631,n4634);
and (n4631,n4632,n4633);
xor (n4632,n4452,n4453);
and (n4633,n166,n333);
and (n4634,n4635,n4636);
xor (n4635,n4632,n4633);
or (n4636,n4637,n4640);
and (n4637,n4638,n4639);
xor (n4638,n4458,n4459);
and (n4639,n312,n333);
and (n4640,n4641,n4642);
xor (n4641,n4638,n4639);
or (n4642,n4643,n4646);
and (n4643,n4644,n4645);
xor (n4644,n4464,n4465);
and (n4645,n580,n333);
and (n4646,n4647,n4648);
xor (n4647,n4644,n4645);
or (n4648,n4649,n4652);
and (n4649,n4650,n4651);
xor (n4650,n4469,n4470);
and (n4651,n574,n333);
and (n4652,n4653,n4654);
xor (n4653,n4650,n4651);
or (n4654,n4655,n4658);
and (n4655,n4656,n4657);
xor (n4656,n4474,n4475);
and (n4657,n712,n333);
and (n4658,n4659,n4660);
xor (n4659,n4656,n4657);
or (n4660,n4661,n4664);
and (n4661,n4662,n4663);
xor (n4662,n4480,n4481);
and (n4663,n753,n333);
and (n4664,n4665,n4666);
xor (n4665,n4662,n4663);
or (n4666,n4667,n4670);
and (n4667,n4668,n4669);
xor (n4668,n4485,n4486);
and (n4669,n922,n333);
and (n4670,n4671,n4672);
xor (n4671,n4668,n4669);
or (n4672,n4673,n4676);
and (n4673,n4674,n4675);
xor (n4674,n4491,n4492);
and (n4675,n959,n333);
and (n4676,n4677,n4678);
xor (n4677,n4674,n4675);
and (n4678,n4679,n3855);
xor (n4679,n4497,n4498);
or (n4680,n4681,n4682);
and (n4681,n4311,n344);
and (n4682,n4310,n4683);
or (n4683,n4684,n4687);
and (n4684,n4685,n4686);
xor (n4685,n4312,n4321);
and (n4686,n102,n341);
and (n4687,n4688,n4689);
xor (n4688,n4685,n4686);
or (n4689,n4690,n4693);
and (n4690,n4691,n4692);
xor (n4691,n4503,n4504);
and (n4692,n281,n341);
and (n4693,n4694,n4695);
xor (n4694,n4691,n4692);
or (n4695,n4696,n4698);
and (n4696,n4697,n1145);
xor (n4697,n4509,n4510);
and (n4698,n4699,n4700);
xor (n4699,n4697,n1145);
or (n4700,n4701,n4704);
and (n4701,n4702,n4703);
xor (n4702,n4515,n4516);
and (n4703,n469,n341);
and (n4704,n4705,n4706);
xor (n4705,n4702,n4703);
or (n4706,n4707,n4710);
and (n4707,n4708,n4709);
xor (n4708,n4521,n4522);
and (n4709,n386,n341);
and (n4710,n4711,n4712);
xor (n4711,n4708,n4709);
or (n4712,n4713,n4716);
and (n4713,n4714,n4715);
xor (n4714,n4527,n4528);
and (n4715,n38,n341);
and (n4716,n4717,n4718);
xor (n4717,n4714,n4715);
or (n4718,n4719,n4722);
and (n4719,n4720,n4721);
xor (n4720,n4533,n4534);
and (n4721,n32,n341);
and (n4722,n4723,n4724);
xor (n4723,n4720,n4721);
or (n4724,n4725,n4728);
and (n4725,n4726,n4727);
xor (n4726,n4539,n4540);
and (n4727,n199,n341);
and (n4728,n4729,n4730);
xor (n4729,n4726,n4727);
or (n4730,n4731,n4734);
and (n4731,n4732,n4733);
xor (n4732,n4545,n4546);
and (n4733,n194,n341);
and (n4734,n4735,n4736);
xor (n4735,n4732,n4733);
or (n4736,n4737,n4740);
and (n4737,n4738,n4739);
xor (n4738,n4551,n4552);
and (n4739,n146,n341);
and (n4740,n4741,n4742);
xor (n4741,n4738,n4739);
or (n4742,n4743,n4746);
and (n4743,n4744,n4745);
xor (n4744,n4557,n4558);
and (n4745,n140,n341);
and (n4746,n4747,n4748);
xor (n4747,n4744,n4745);
or (n4748,n4749,n4751);
and (n4749,n4750,n2621);
xor (n4750,n4563,n4564);
and (n4751,n4752,n4753);
xor (n4752,n4750,n2621);
or (n4753,n4754,n4757);
and (n4754,n4755,n4756);
xor (n4755,n4569,n4570);
and (n4756,n260,n341);
and (n4757,n4758,n4759);
xor (n4758,n4755,n4756);
or (n4759,n4760,n4763);
and (n4760,n4761,n4762);
xor (n4761,n4575,n4576);
and (n4762,n65,n341);
and (n4763,n4764,n4765);
xor (n4764,n4761,n4762);
or (n4765,n4766,n4769);
and (n4766,n4767,n4768);
xor (n4767,n4581,n4582);
and (n4768,n58,n341);
and (n4769,n4770,n4771);
xor (n4770,n4767,n4768);
or (n4771,n4772,n4775);
and (n4772,n4773,n4774);
xor (n4773,n4587,n4588);
and (n4774,n90,n341);
and (n4775,n4776,n4777);
xor (n4776,n4773,n4774);
or (n4777,n4778,n4781);
and (n4778,n4779,n4780);
xor (n4779,n4593,n4594);
and (n4780,n84,n341);
and (n4781,n4782,n4783);
xor (n4782,n4779,n4780);
or (n4783,n4784,n4787);
and (n4784,n4785,n4786);
xor (n4785,n4599,n4600);
and (n4786,n224,n341);
and (n4787,n4788,n4789);
xor (n4788,n4785,n4786);
or (n4789,n4790,n4793);
and (n4790,n4791,n4792);
xor (n4791,n4605,n4606);
and (n4792,n218,n341);
and (n4793,n4794,n4795);
xor (n4794,n4791,n4792);
or (n4795,n4796,n4799);
and (n4796,n4797,n4798);
xor (n4797,n4611,n4612);
and (n4798,n247,n341);
and (n4799,n4800,n4801);
xor (n4800,n4797,n4798);
or (n4801,n4802,n4805);
and (n4802,n4803,n4804);
xor (n4803,n4617,n4618);
and (n4804,n241,n341);
and (n4805,n4806,n4807);
xor (n4806,n4803,n4804);
or (n4807,n4808,n4811);
and (n4808,n4809,n4810);
xor (n4809,n4623,n4624);
and (n4810,n174,n341);
and (n4811,n4812,n4813);
xor (n4812,n4809,n4810);
or (n4813,n4814,n4817);
and (n4814,n4815,n4816);
xor (n4815,n4629,n4630);
and (n4816,n166,n341);
and (n4817,n4818,n4819);
xor (n4818,n4815,n4816);
or (n4819,n4820,n4823);
and (n4820,n4821,n4822);
xor (n4821,n4635,n4636);
and (n4822,n312,n341);
and (n4823,n4824,n4825);
xor (n4824,n4821,n4822);
or (n4825,n4826,n4829);
and (n4826,n4827,n4828);
xor (n4827,n4641,n4642);
and (n4828,n580,n341);
and (n4829,n4830,n4831);
xor (n4830,n4827,n4828);
or (n4831,n4832,n4835);
and (n4832,n4833,n4834);
xor (n4833,n4647,n4648);
and (n4834,n574,n341);
and (n4835,n4836,n4837);
xor (n4836,n4833,n4834);
or (n4837,n4838,n4840);
and (n4838,n4839,n3710);
xor (n4839,n4653,n4654);
and (n4840,n4841,n4842);
xor (n4841,n4839,n3710);
or (n4842,n4843,n4845);
and (n4843,n4844,n3752);
xor (n4844,n4659,n4660);
and (n4845,n4846,n4847);
xor (n4846,n4844,n3752);
or (n4847,n4848,n4850);
and (n4848,n4849,n3806);
xor (n4849,n4665,n4666);
and (n4850,n4851,n4852);
xor (n4851,n4849,n3806);
or (n4852,n4853,n4855);
and (n4853,n4854,n3833);
xor (n4854,n4671,n4672);
and (n4855,n4856,n4857);
xor (n4856,n4854,n3833);
and (n4857,n4858,n4859);
xor (n4858,n4677,n4678);
and (n4859,n1122,n341);
and (n4860,n121,n356);
or (n4861,n4862,n4863);
and (n4862,n4309,n4860);
and (n4863,n4308,n4864);
or (n4864,n4865,n4868);
and (n4865,n4866,n4867);
xor (n4866,n4310,n4683);
and (n4867,n102,n356);
and (n4868,n4869,n4870);
xor (n4869,n4866,n4867);
or (n4870,n4871,n4874);
and (n4871,n4872,n4873);
xor (n4872,n4688,n4689);
and (n4873,n281,n356);
and (n4874,n4875,n4876);
xor (n4875,n4872,n4873);
or (n4876,n4877,n4880);
and (n4877,n4878,n4879);
xor (n4878,n4694,n4695);
and (n4879,n274,n356);
and (n4880,n4881,n4882);
xor (n4881,n4878,n4879);
or (n4882,n4883,n4886);
and (n4883,n4884,n4885);
xor (n4884,n4699,n4700);
and (n4885,n469,n356);
and (n4886,n4887,n4888);
xor (n4887,n4884,n4885);
or (n4888,n4889,n4892);
and (n4889,n4890,n4891);
xor (n4890,n4705,n4706);
and (n4891,n386,n356);
and (n4892,n4893,n4894);
xor (n4893,n4890,n4891);
or (n4894,n4895,n4898);
and (n4895,n4896,n4897);
xor (n4896,n4711,n4712);
and (n4897,n38,n356);
and (n4898,n4899,n4900);
xor (n4899,n4896,n4897);
or (n4900,n4901,n4904);
and (n4901,n4902,n4903);
xor (n4902,n4717,n4718);
and (n4903,n32,n356);
and (n4904,n4905,n4906);
xor (n4905,n4902,n4903);
or (n4906,n4907,n4910);
and (n4907,n4908,n4909);
xor (n4908,n4723,n4724);
and (n4909,n199,n356);
and (n4910,n4911,n4912);
xor (n4911,n4908,n4909);
or (n4912,n4913,n4916);
and (n4913,n4914,n4915);
xor (n4914,n4729,n4730);
and (n4915,n194,n356);
and (n4916,n4917,n4918);
xor (n4917,n4914,n4915);
or (n4918,n4919,n4922);
and (n4919,n4920,n4921);
xor (n4920,n4735,n4736);
and (n4921,n146,n356);
and (n4922,n4923,n4924);
xor (n4923,n4920,n4921);
or (n4924,n4925,n4928);
and (n4925,n4926,n4927);
xor (n4926,n4741,n4742);
and (n4927,n140,n356);
and (n4928,n4929,n4930);
xor (n4929,n4926,n4927);
or (n4930,n4931,n4934);
and (n4931,n4932,n4933);
xor (n4932,n4747,n4748);
and (n4933,n266,n356);
and (n4934,n4935,n4936);
xor (n4935,n4932,n4933);
or (n4936,n4937,n4940);
and (n4937,n4938,n4939);
xor (n4938,n4752,n4753);
and (n4939,n260,n356);
and (n4940,n4941,n4942);
xor (n4941,n4938,n4939);
or (n4942,n4943,n4946);
and (n4943,n4944,n4945);
xor (n4944,n4758,n4759);
and (n4945,n65,n356);
and (n4946,n4947,n4948);
xor (n4947,n4944,n4945);
or (n4948,n4949,n4952);
and (n4949,n4950,n4951);
xor (n4950,n4764,n4765);
and (n4951,n58,n356);
and (n4952,n4953,n4954);
xor (n4953,n4950,n4951);
or (n4954,n4955,n4958);
and (n4955,n4956,n4957);
xor (n4956,n4770,n4771);
and (n4957,n90,n356);
and (n4958,n4959,n4960);
xor (n4959,n4956,n4957);
or (n4960,n4961,n4964);
and (n4961,n4962,n4963);
xor (n4962,n4776,n4777);
and (n4963,n84,n356);
and (n4964,n4965,n4966);
xor (n4965,n4962,n4963);
or (n4966,n4967,n4970);
and (n4967,n4968,n4969);
xor (n4968,n4782,n4783);
and (n4969,n224,n356);
and (n4970,n4971,n4972);
xor (n4971,n4968,n4969);
or (n4972,n4973,n4976);
and (n4973,n4974,n4975);
xor (n4974,n4788,n4789);
and (n4975,n218,n356);
and (n4976,n4977,n4978);
xor (n4977,n4974,n4975);
or (n4978,n4979,n4982);
and (n4979,n4980,n4981);
xor (n4980,n4794,n4795);
and (n4981,n247,n356);
and (n4982,n4983,n4984);
xor (n4983,n4980,n4981);
or (n4984,n4985,n4988);
and (n4985,n4986,n4987);
xor (n4986,n4800,n4801);
and (n4987,n241,n356);
and (n4988,n4989,n4990);
xor (n4989,n4986,n4987);
or (n4990,n4991,n4994);
and (n4991,n4992,n4993);
xor (n4992,n4806,n4807);
and (n4993,n174,n356);
and (n4994,n4995,n4996);
xor (n4995,n4992,n4993);
or (n4996,n4997,n5000);
and (n4997,n4998,n4999);
xor (n4998,n4812,n4813);
and (n4999,n166,n356);
and (n5000,n5001,n5002);
xor (n5001,n4998,n4999);
or (n5002,n5003,n5006);
and (n5003,n5004,n5005);
xor (n5004,n4818,n4819);
and (n5005,n312,n356);
and (n5006,n5007,n5008);
xor (n5007,n5004,n5005);
or (n5008,n5009,n5012);
and (n5009,n5010,n5011);
xor (n5010,n4824,n4825);
and (n5011,n580,n356);
and (n5012,n5013,n5014);
xor (n5013,n5010,n5011);
or (n5014,n5015,n5018);
and (n5015,n5016,n5017);
xor (n5016,n4830,n4831);
and (n5017,n574,n356);
and (n5018,n5019,n5020);
xor (n5019,n5016,n5017);
or (n5020,n5021,n5024);
and (n5021,n5022,n5023);
xor (n5022,n4836,n4837);
and (n5023,n712,n356);
and (n5024,n5025,n5026);
xor (n5025,n5022,n5023);
or (n5026,n5027,n5030);
and (n5027,n5028,n5029);
xor (n5028,n4841,n4842);
and (n5029,n753,n356);
and (n5030,n5031,n5032);
xor (n5031,n5028,n5029);
or (n5032,n5033,n5036);
and (n5033,n5034,n5035);
xor (n5034,n4846,n4847);
and (n5035,n922,n356);
and (n5036,n5037,n5038);
xor (n5037,n5034,n5035);
or (n5038,n5039,n5042);
and (n5039,n5040,n5041);
xor (n5040,n4851,n4852);
and (n5041,n959,n356);
and (n5042,n5043,n5044);
xor (n5043,n5040,n5041);
and (n5044,n5045,n3779);
xor (n5045,n4856,n4857);
and (n5046,n121,n111);
or (n5047,n5048,n5049);
and (n5048,n4307,n5046);
and (n5049,n4306,n5050);
or (n5050,n5051,n5054);
and (n5051,n5052,n5053);
xor (n5052,n4308,n4864);
and (n5053,n102,n111);
and (n5054,n5055,n5056);
xor (n5055,n5052,n5053);
or (n5056,n5057,n5059);
and (n5057,n5058,n350);
xor (n5058,n4869,n4870);
and (n5059,n5060,n5061);
xor (n5060,n5058,n350);
or (n5061,n5062,n5065);
and (n5062,n5063,n5064);
xor (n5063,n4875,n4876);
and (n5064,n274,n111);
and (n5065,n5066,n5067);
xor (n5066,n5063,n5064);
or (n5067,n5068,n5071);
and (n5068,n5069,n5070);
xor (n5069,n4881,n4882);
and (n5070,n469,n111);
and (n5071,n5072,n5073);
xor (n5072,n5069,n5070);
or (n5073,n5074,n5077);
and (n5074,n5075,n5076);
xor (n5075,n4887,n4888);
and (n5076,n386,n111);
and (n5077,n5078,n5079);
xor (n5078,n5075,n5076);
or (n5079,n5080,n5083);
and (n5080,n5081,n5082);
xor (n5081,n4893,n4894);
and (n5082,n38,n111);
and (n5083,n5084,n5085);
xor (n5084,n5081,n5082);
or (n5085,n5086,n5089);
and (n5086,n5087,n5088);
xor (n5087,n4899,n4900);
and (n5088,n32,n111);
and (n5089,n5090,n5091);
xor (n5090,n5087,n5088);
or (n5091,n5092,n5095);
and (n5092,n5093,n5094);
xor (n5093,n4905,n4906);
and (n5094,n199,n111);
and (n5095,n5096,n5097);
xor (n5096,n5093,n5094);
or (n5097,n5098,n5101);
and (n5098,n5099,n5100);
xor (n5099,n4911,n4912);
and (n5100,n194,n111);
and (n5101,n5102,n5103);
xor (n5102,n5099,n5100);
or (n5103,n5104,n5107);
and (n5104,n5105,n5106);
xor (n5105,n4917,n4918);
and (n5106,n146,n111);
and (n5107,n5108,n5109);
xor (n5108,n5105,n5106);
or (n5109,n5110,n5113);
and (n5110,n5111,n5112);
xor (n5111,n4923,n4924);
and (n5112,n140,n111);
and (n5113,n5114,n5115);
xor (n5114,n5111,n5112);
or (n5115,n5116,n5119);
and (n5116,n5117,n5118);
xor (n5117,n4929,n4930);
and (n5118,n266,n111);
and (n5119,n5120,n5121);
xor (n5120,n5117,n5118);
or (n5121,n5122,n5124);
and (n5122,n5123,n3217);
xor (n5123,n4935,n4936);
and (n5124,n5125,n5126);
xor (n5125,n5123,n3217);
or (n5126,n5127,n5129);
and (n5127,n5128,n2646);
xor (n5128,n4941,n4942);
and (n5129,n5130,n5131);
xor (n5130,n5128,n2646);
or (n5131,n5132,n5135);
and (n5132,n5133,n5134);
xor (n5133,n4947,n4948);
and (n5134,n58,n111);
and (n5135,n5136,n5137);
xor (n5136,n5133,n5134);
or (n5137,n5138,n5141);
and (n5138,n5139,n5140);
xor (n5139,n4953,n4954);
and (n5140,n90,n111);
and (n5141,n5142,n5143);
xor (n5142,n5139,n5140);
or (n5143,n5144,n5147);
and (n5144,n5145,n5146);
xor (n5145,n4959,n4960);
and (n5146,n84,n111);
and (n5147,n5148,n5149);
xor (n5148,n5145,n5146);
or (n5149,n5150,n5153);
and (n5150,n5151,n5152);
xor (n5151,n4965,n4966);
and (n5152,n224,n111);
and (n5153,n5154,n5155);
xor (n5154,n5151,n5152);
or (n5155,n5156,n5159);
and (n5156,n5157,n5158);
xor (n5157,n4971,n4972);
and (n5158,n218,n111);
and (n5159,n5160,n5161);
xor (n5160,n5157,n5158);
or (n5161,n5162,n5165);
and (n5162,n5163,n5164);
xor (n5163,n4977,n4978);
and (n5164,n247,n111);
and (n5165,n5166,n5167);
xor (n5166,n5163,n5164);
or (n5167,n5168,n5171);
and (n5168,n5169,n5170);
xor (n5169,n4983,n4984);
and (n5170,n241,n111);
and (n5171,n5172,n5173);
xor (n5172,n5169,n5170);
or (n5173,n5174,n5177);
and (n5174,n5175,n5176);
xor (n5175,n4989,n4990);
and (n5176,n174,n111);
and (n5177,n5178,n5179);
xor (n5178,n5175,n5176);
or (n5179,n5180,n5183);
and (n5180,n5181,n5182);
xor (n5181,n4995,n4996);
and (n5182,n166,n111);
and (n5183,n5184,n5185);
xor (n5184,n5181,n5182);
or (n5185,n5186,n5189);
and (n5186,n5187,n5188);
xor (n5187,n5001,n5002);
and (n5188,n312,n111);
and (n5189,n5190,n5191);
xor (n5190,n5187,n5188);
or (n5191,n5192,n5195);
and (n5192,n5193,n5194);
xor (n5193,n5007,n5008);
and (n5194,n580,n111);
and (n5195,n5196,n5197);
xor (n5196,n5193,n5194);
or (n5197,n5198,n5201);
and (n5198,n5199,n5200);
xor (n5199,n5013,n5014);
and (n5200,n574,n111);
and (n5201,n5202,n5203);
xor (n5202,n5199,n5200);
or (n5203,n5204,n5207);
and (n5204,n5205,n5206);
xor (n5205,n5019,n5020);
and (n5206,n712,n111);
and (n5207,n5208,n5209);
xor (n5208,n5205,n5206);
or (n5209,n5210,n5213);
and (n5210,n5211,n5212);
xor (n5211,n5025,n5026);
and (n5212,n753,n111);
and (n5213,n5214,n5215);
xor (n5214,n5211,n5212);
or (n5215,n5216,n5218);
and (n5216,n5217,n3717);
xor (n5217,n5031,n5032);
and (n5218,n5219,n5220);
xor (n5219,n5217,n3717);
or (n5220,n5221,n5223);
and (n5221,n5222,n3772);
xor (n5222,n5037,n5038);
and (n5223,n5224,n5225);
xor (n5224,n5222,n3772);
and (n5225,n5226,n5227);
xor (n5226,n5043,n5044);
and (n5227,n1122,n111);
and (n5228,n121,n109);
or (n5229,n5230,n5233);
and (n5230,n5231,n5232);
xor (n5231,n4306,n5050);
and (n5232,n102,n109);
and (n5233,n5234,n5235);
xor (n5234,n5231,n5232);
or (n5235,n5236,n5239);
and (n5236,n5237,n5238);
xor (n5237,n5055,n5056);
and (n5238,n281,n109);
and (n5239,n5240,n5241);
xor (n5240,n5237,n5238);
or (n5241,n5242,n5245);
and (n5242,n5243,n5244);
xor (n5243,n5060,n5061);
and (n5244,n274,n109);
and (n5245,n5246,n5247);
xor (n5246,n5243,n5244);
or (n5247,n5248,n5251);
and (n5248,n5249,n5250);
xor (n5249,n5066,n5067);
and (n5250,n469,n109);
and (n5251,n5252,n5253);
xor (n5252,n5249,n5250);
or (n5253,n5254,n5257);
and (n5254,n5255,n5256);
xor (n5255,n5072,n5073);
and (n5256,n386,n109);
and (n5257,n5258,n5259);
xor (n5258,n5255,n5256);
or (n5259,n5260,n5263);
and (n5260,n5261,n5262);
xor (n5261,n5078,n5079);
and (n5262,n38,n109);
and (n5263,n5264,n5265);
xor (n5264,n5261,n5262);
or (n5265,n5266,n5269);
and (n5266,n5267,n5268);
xor (n5267,n5084,n5085);
and (n5268,n32,n109);
and (n5269,n5270,n5271);
xor (n5270,n5267,n5268);
or (n5271,n5272,n5275);
and (n5272,n5273,n5274);
xor (n5273,n5090,n5091);
and (n5274,n199,n109);
and (n5275,n5276,n5277);
xor (n5276,n5273,n5274);
or (n5277,n5278,n5281);
and (n5278,n5279,n5280);
xor (n5279,n5096,n5097);
and (n5280,n194,n109);
and (n5281,n5282,n5283);
xor (n5282,n5279,n5280);
or (n5283,n5284,n5287);
and (n5284,n5285,n5286);
xor (n5285,n5102,n5103);
and (n5286,n146,n109);
and (n5287,n5288,n5289);
xor (n5288,n5285,n5286);
or (n5289,n5290,n5293);
and (n5290,n5291,n5292);
xor (n5291,n5108,n5109);
and (n5292,n140,n109);
and (n5293,n5294,n5295);
xor (n5294,n5291,n5292);
or (n5295,n5296,n5299);
and (n5296,n5297,n5298);
xor (n5297,n5114,n5115);
and (n5298,n266,n109);
and (n5299,n5300,n5301);
xor (n5300,n5297,n5298);
or (n5301,n5302,n5305);
and (n5302,n5303,n5304);
xor (n5303,n5120,n5121);
and (n5304,n260,n109);
and (n5305,n5306,n5307);
xor (n5306,n5303,n5304);
or (n5307,n5308,n5311);
and (n5308,n5309,n5310);
xor (n5309,n5125,n5126);
and (n5310,n65,n109);
and (n5311,n5312,n5313);
xor (n5312,n5309,n5310);
or (n5313,n5314,n5317);
and (n5314,n5315,n5316);
xor (n5315,n5130,n5131);
and (n5316,n58,n109);
and (n5317,n5318,n5319);
xor (n5318,n5315,n5316);
or (n5319,n5320,n5323);
and (n5320,n5321,n5322);
xor (n5321,n5136,n5137);
and (n5322,n90,n109);
and (n5323,n5324,n5325);
xor (n5324,n5321,n5322);
or (n5325,n5326,n5329);
and (n5326,n5327,n5328);
xor (n5327,n5142,n5143);
and (n5328,n84,n109);
and (n5329,n5330,n5331);
xor (n5330,n5327,n5328);
or (n5331,n5332,n5335);
and (n5332,n5333,n5334);
xor (n5333,n5148,n5149);
and (n5334,n224,n109);
and (n5335,n5336,n5337);
xor (n5336,n5333,n5334);
or (n5337,n5338,n5341);
and (n5338,n5339,n5340);
xor (n5339,n5154,n5155);
and (n5340,n218,n109);
and (n5341,n5342,n5343);
xor (n5342,n5339,n5340);
or (n5343,n5344,n5347);
and (n5344,n5345,n5346);
xor (n5345,n5160,n5161);
and (n5346,n247,n109);
and (n5347,n5348,n5349);
xor (n5348,n5345,n5346);
or (n5349,n5350,n5353);
and (n5350,n5351,n5352);
xor (n5351,n5166,n5167);
and (n5352,n241,n109);
and (n5353,n5354,n5355);
xor (n5354,n5351,n5352);
or (n5355,n5356,n5359);
and (n5356,n5357,n5358);
xor (n5357,n5172,n5173);
and (n5358,n174,n109);
and (n5359,n5360,n5361);
xor (n5360,n5357,n5358);
or (n5361,n5362,n5365);
and (n5362,n5363,n5364);
xor (n5363,n5178,n5179);
and (n5364,n166,n109);
and (n5365,n5366,n5367);
xor (n5366,n5363,n5364);
or (n5367,n5368,n5371);
and (n5368,n5369,n5370);
xor (n5369,n5184,n5185);
and (n5370,n312,n109);
and (n5371,n5372,n5373);
xor (n5372,n5369,n5370);
or (n5373,n5374,n5377);
and (n5374,n5375,n5376);
xor (n5375,n5190,n5191);
and (n5376,n580,n109);
and (n5377,n5378,n5379);
xor (n5378,n5375,n5376);
or (n5379,n5380,n5383);
and (n5380,n5381,n5382);
xor (n5381,n5196,n5197);
and (n5382,n574,n109);
and (n5383,n5384,n5385);
xor (n5384,n5381,n5382);
or (n5385,n5386,n5389);
and (n5386,n5387,n5388);
xor (n5387,n5202,n5203);
and (n5388,n712,n109);
and (n5389,n5390,n5391);
xor (n5390,n5387,n5388);
or (n5391,n5392,n5395);
and (n5392,n5393,n5394);
xor (n5393,n5208,n5209);
and (n5394,n753,n109);
and (n5395,n5396,n5397);
xor (n5396,n5393,n5394);
or (n5397,n5398,n5401);
and (n5398,n5399,n5400);
xor (n5399,n5214,n5215);
and (n5400,n922,n109);
and (n5401,n5402,n5403);
xor (n5402,n5399,n5400);
or (n5403,n5404,n5407);
and (n5404,n5405,n5406);
xor (n5405,n5219,n5220);
and (n5406,n959,n109);
and (n5407,n5408,n5409);
xor (n5408,n5405,n5406);
and (n5409,n5410,n3676);
xor (n5410,n5224,n5225);
and (n5411,n102,n100);
or (n5412,n5413,n5416);
and (n5413,n5414,n5415);
xor (n5414,n5234,n5235);
and (n5415,n281,n100);
and (n5416,n5417,n5418);
xor (n5417,n5414,n5415);
or (n5418,n5419,n5422);
and (n5419,n5420,n5421);
xor (n5420,n5240,n5241);
and (n5421,n274,n100);
and (n5422,n5423,n5424);
xor (n5423,n5420,n5421);
or (n5424,n5425,n5428);
and (n5425,n5426,n5427);
xor (n5426,n5246,n5247);
and (n5427,n469,n100);
and (n5428,n5429,n5430);
xor (n5429,n5426,n5427);
or (n5430,n5431,n5434);
and (n5431,n5432,n5433);
xor (n5432,n5252,n5253);
and (n5433,n386,n100);
and (n5434,n5435,n5436);
xor (n5435,n5432,n5433);
or (n5436,n5437,n5440);
and (n5437,n5438,n5439);
xor (n5438,n5258,n5259);
and (n5439,n38,n100);
and (n5440,n5441,n5442);
xor (n5441,n5438,n5439);
or (n5442,n5443,n5446);
and (n5443,n5444,n5445);
xor (n5444,n5264,n5265);
and (n5445,n32,n100);
and (n5446,n5447,n5448);
xor (n5447,n5444,n5445);
or (n5448,n5449,n5452);
and (n5449,n5450,n5451);
xor (n5450,n5270,n5271);
and (n5451,n199,n100);
and (n5452,n5453,n5454);
xor (n5453,n5450,n5451);
or (n5454,n5455,n5458);
and (n5455,n5456,n5457);
xor (n5456,n5276,n5277);
and (n5457,n194,n100);
and (n5458,n5459,n5460);
xor (n5459,n5456,n5457);
or (n5460,n5461,n5464);
and (n5461,n5462,n5463);
xor (n5462,n5282,n5283);
and (n5463,n146,n100);
and (n5464,n5465,n5466);
xor (n5465,n5462,n5463);
or (n5466,n5467,n5470);
and (n5467,n5468,n5469);
xor (n5468,n5288,n5289);
and (n5469,n140,n100);
and (n5470,n5471,n5472);
xor (n5471,n5468,n5469);
or (n5472,n5473,n5476);
and (n5473,n5474,n5475);
xor (n5474,n5294,n5295);
and (n5475,n266,n100);
and (n5476,n5477,n5478);
xor (n5477,n5474,n5475);
or (n5478,n5479,n5482);
and (n5479,n5480,n5481);
xor (n5480,n5300,n5301);
and (n5481,n260,n100);
and (n5482,n5483,n5484);
xor (n5483,n5480,n5481);
or (n5484,n5485,n5488);
and (n5485,n5486,n5487);
xor (n5486,n5306,n5307);
and (n5487,n65,n100);
and (n5488,n5489,n5490);
xor (n5489,n5486,n5487);
or (n5490,n5491,n5494);
and (n5491,n5492,n5493);
xor (n5492,n5312,n5313);
and (n5493,n58,n100);
and (n5494,n5495,n5496);
xor (n5495,n5492,n5493);
or (n5496,n5497,n5499);
and (n5497,n5498,n2531);
xor (n5498,n5318,n5319);
and (n5499,n5500,n5501);
xor (n5500,n5498,n2531);
or (n5501,n5502,n5504);
and (n5502,n5503,n2467);
xor (n5503,n5324,n5325);
and (n5504,n5505,n5506);
xor (n5505,n5503,n2467);
or (n5506,n5507,n5509);
and (n5507,n5508,n2432);
xor (n5508,n5330,n5331);
and (n5509,n5510,n5511);
xor (n5510,n5508,n2432);
or (n5511,n5512,n5514);
and (n5512,n5513,n2336);
xor (n5513,n5336,n5337);
and (n5514,n5515,n5516);
xor (n5515,n5513,n2336);
or (n5516,n5517,n5520);
and (n5517,n5518,n5519);
xor (n5518,n5342,n5343);
and (n5519,n247,n100);
and (n5520,n5521,n5522);
xor (n5521,n5518,n5519);
or (n5522,n5523,n5526);
and (n5523,n5524,n5525);
xor (n5524,n5348,n5349);
and (n5525,n241,n100);
and (n5526,n5527,n5528);
xor (n5527,n5524,n5525);
or (n5528,n5529,n5532);
and (n5529,n5530,n5531);
xor (n5530,n5354,n5355);
and (n5531,n174,n100);
and (n5532,n5533,n5534);
xor (n5533,n5530,n5531);
or (n5534,n5535,n5538);
and (n5535,n5536,n5537);
xor (n5536,n5360,n5361);
and (n5537,n166,n100);
and (n5538,n5539,n5540);
xor (n5539,n5536,n5537);
or (n5540,n5541,n5543);
and (n5541,n5542,n2973);
xor (n5542,n5366,n5367);
and (n5543,n5544,n5545);
xor (n5544,n5542,n2973);
or (n5545,n5546,n5549);
and (n5546,n5547,n5548);
xor (n5547,n5372,n5373);
and (n5548,n580,n100);
and (n5549,n5550,n5551);
xor (n5550,n5547,n5548);
or (n5551,n5552,n5555);
and (n5552,n5553,n5554);
xor (n5553,n5378,n5379);
and (n5554,n574,n100);
and (n5555,n5556,n5557);
xor (n5556,n5553,n5554);
or (n5557,n5558,n5561);
and (n5558,n5559,n5560);
xor (n5559,n5384,n5385);
and (n5560,n712,n100);
and (n5561,n5562,n5563);
xor (n5562,n5559,n5560);
or (n5563,n5564,n5567);
and (n5564,n5565,n5566);
xor (n5565,n5390,n5391);
and (n5566,n753,n100);
and (n5567,n5568,n5569);
xor (n5568,n5565,n5566);
or (n5569,n5570,n5573);
and (n5570,n5571,n5572);
xor (n5571,n5396,n5397);
and (n5572,n922,n100);
and (n5573,n5574,n5575);
xor (n5574,n5571,n5572);
or (n5575,n5576,n5578);
and (n5576,n5577,n3546);
xor (n5577,n5402,n5403);
and (n5578,n5579,n5580);
xor (n5579,n5577,n3546);
and (n5580,n5581,n5582);
xor (n5581,n5408,n5409);
and (n5582,n1122,n100);
and (n5583,n281,n373);
or (n5584,n5585,n5588);
and (n5585,n5586,n5587);
xor (n5586,n5417,n5418);
and (n5587,n274,n373);
and (n5588,n5589,n5590);
xor (n5589,n5586,n5587);
or (n5590,n5591,n5594);
and (n5591,n5592,n5593);
xor (n5592,n5423,n5424);
and (n5593,n469,n373);
and (n5594,n5595,n5596);
xor (n5595,n5592,n5593);
or (n5596,n5597,n5600);
and (n5597,n5598,n5599);
xor (n5598,n5429,n5430);
and (n5599,n386,n373);
and (n5600,n5601,n5602);
xor (n5601,n5598,n5599);
or (n5602,n5603,n5606);
and (n5603,n5604,n5605);
xor (n5604,n5435,n5436);
and (n5605,n38,n373);
and (n5606,n5607,n5608);
xor (n5607,n5604,n5605);
or (n5608,n5609,n5612);
and (n5609,n5610,n5611);
xor (n5610,n5441,n5442);
and (n5611,n32,n373);
and (n5612,n5613,n5614);
xor (n5613,n5610,n5611);
or (n5614,n5615,n5618);
and (n5615,n5616,n5617);
xor (n5616,n5447,n5448);
and (n5617,n199,n373);
and (n5618,n5619,n5620);
xor (n5619,n5616,n5617);
or (n5620,n5621,n5624);
and (n5621,n5622,n5623);
xor (n5622,n5453,n5454);
and (n5623,n194,n373);
and (n5624,n5625,n5626);
xor (n5625,n5622,n5623);
or (n5626,n5627,n5630);
and (n5627,n5628,n5629);
xor (n5628,n5459,n5460);
and (n5629,n146,n373);
and (n5630,n5631,n5632);
xor (n5631,n5628,n5629);
or (n5632,n5633,n5636);
and (n5633,n5634,n5635);
xor (n5634,n5465,n5466);
and (n5635,n140,n373);
and (n5636,n5637,n5638);
xor (n5637,n5634,n5635);
or (n5638,n5639,n5642);
and (n5639,n5640,n5641);
xor (n5640,n5471,n5472);
and (n5641,n266,n373);
and (n5642,n5643,n5644);
xor (n5643,n5640,n5641);
or (n5644,n5645,n5648);
and (n5645,n5646,n5647);
xor (n5646,n5477,n5478);
and (n5647,n260,n373);
and (n5648,n5649,n5650);
xor (n5649,n5646,n5647);
or (n5650,n5651,n5654);
and (n5651,n5652,n5653);
xor (n5652,n5483,n5484);
and (n5653,n65,n373);
and (n5654,n5655,n5656);
xor (n5655,n5652,n5653);
or (n5656,n5657,n5660);
and (n5657,n5658,n5659);
xor (n5658,n5489,n5490);
and (n5659,n58,n373);
and (n5660,n5661,n5662);
xor (n5661,n5658,n5659);
or (n5662,n5663,n5666);
and (n5663,n5664,n5665);
xor (n5664,n5495,n5496);
and (n5665,n90,n373);
and (n5666,n5667,n5668);
xor (n5667,n5664,n5665);
or (n5668,n5669,n5672);
and (n5669,n5670,n5671);
xor (n5670,n5500,n5501);
and (n5671,n84,n373);
and (n5672,n5673,n5674);
xor (n5673,n5670,n5671);
or (n5674,n5675,n5678);
and (n5675,n5676,n5677);
xor (n5676,n5505,n5506);
and (n5677,n224,n373);
and (n5678,n5679,n5680);
xor (n5679,n5676,n5677);
or (n5680,n5681,n5684);
and (n5681,n5682,n5683);
xor (n5682,n5510,n5511);
and (n5683,n218,n373);
and (n5684,n5685,n5686);
xor (n5685,n5682,n5683);
or (n5686,n5687,n5690);
and (n5687,n5688,n5689);
xor (n5688,n5515,n5516);
and (n5689,n247,n373);
and (n5690,n5691,n5692);
xor (n5691,n5688,n5689);
or (n5692,n5693,n5696);
and (n5693,n5694,n5695);
xor (n5694,n5521,n5522);
and (n5695,n241,n373);
and (n5696,n5697,n5698);
xor (n5697,n5694,n5695);
or (n5698,n5699,n5702);
and (n5699,n5700,n5701);
xor (n5700,n5527,n5528);
and (n5701,n174,n373);
and (n5702,n5703,n5704);
xor (n5703,n5700,n5701);
or (n5704,n5705,n5708);
and (n5705,n5706,n5707);
xor (n5706,n5533,n5534);
and (n5707,n166,n373);
and (n5708,n5709,n5710);
xor (n5709,n5706,n5707);
or (n5710,n5711,n5714);
and (n5711,n5712,n5713);
xor (n5712,n5539,n5540);
and (n5713,n312,n373);
and (n5714,n5715,n5716);
xor (n5715,n5712,n5713);
or (n5716,n5717,n5720);
and (n5717,n5718,n5719);
xor (n5718,n5544,n5545);
and (n5719,n580,n373);
and (n5720,n5721,n5722);
xor (n5721,n5718,n5719);
or (n5722,n5723,n5726);
and (n5723,n5724,n5725);
xor (n5724,n5550,n5551);
and (n5725,n574,n373);
and (n5726,n5727,n5728);
xor (n5727,n5724,n5725);
or (n5728,n5729,n5732);
and (n5729,n5730,n5731);
xor (n5730,n5556,n5557);
and (n5731,n712,n373);
and (n5732,n5733,n5734);
xor (n5733,n5730,n5731);
or (n5734,n5735,n5738);
and (n5735,n5736,n5737);
xor (n5736,n5562,n5563);
and (n5737,n753,n373);
and (n5738,n5739,n5740);
xor (n5739,n5736,n5737);
or (n5740,n5741,n5744);
and (n5741,n5742,n5743);
xor (n5742,n5568,n5569);
and (n5743,n922,n373);
and (n5744,n5745,n5746);
xor (n5745,n5742,n5743);
or (n5746,n5747,n5750);
and (n5747,n5748,n5749);
xor (n5748,n5574,n5575);
and (n5749,n959,n373);
and (n5750,n5751,n5752);
xor (n5751,n5748,n5749);
and (n5752,n5753,n3519);
xor (n5753,n5579,n5580);
and (n5754,n274,n378);
or (n5755,n5756,n5759);
and (n5756,n5757,n5758);
xor (n5757,n5589,n5590);
and (n5758,n469,n378);
and (n5759,n5760,n5761);
xor (n5760,n5757,n5758);
or (n5761,n5762,n5765);
and (n5762,n5763,n5764);
xor (n5763,n5595,n5596);
and (n5764,n386,n378);
and (n5765,n5766,n5767);
xor (n5766,n5763,n5764);
or (n5767,n5768,n5771);
and (n5768,n5769,n5770);
xor (n5769,n5601,n5602);
and (n5770,n38,n378);
and (n5771,n5772,n5773);
xor (n5772,n5769,n5770);
or (n5773,n5774,n5777);
and (n5774,n5775,n5776);
xor (n5775,n5607,n5608);
and (n5776,n32,n378);
and (n5777,n5778,n5779);
xor (n5778,n5775,n5776);
or (n5779,n5780,n5783);
and (n5780,n5781,n5782);
xor (n5781,n5613,n5614);
and (n5782,n199,n378);
and (n5783,n5784,n5785);
xor (n5784,n5781,n5782);
or (n5785,n5786,n5789);
and (n5786,n5787,n5788);
xor (n5787,n5619,n5620);
and (n5788,n194,n378);
and (n5789,n5790,n5791);
xor (n5790,n5787,n5788);
or (n5791,n5792,n5794);
and (n5792,n5793,n1308);
xor (n5793,n5625,n5626);
and (n5794,n5795,n5796);
xor (n5795,n5793,n1308);
or (n5796,n5797,n5800);
and (n5797,n5798,n5799);
xor (n5798,n5631,n5632);
and (n5799,n140,n378);
and (n5800,n5801,n5802);
xor (n5801,n5798,n5799);
or (n5802,n5803,n5806);
and (n5803,n5804,n5805);
xor (n5804,n5637,n5638);
and (n5805,n266,n378);
and (n5806,n5807,n5808);
xor (n5807,n5804,n5805);
or (n5808,n5809,n5812);
and (n5809,n5810,n5811);
xor (n5810,n5643,n5644);
and (n5811,n260,n378);
and (n5812,n5813,n5814);
xor (n5813,n5810,n5811);
or (n5814,n5815,n5818);
and (n5815,n5816,n5817);
xor (n5816,n5649,n5650);
and (n5817,n65,n378);
and (n5818,n5819,n5820);
xor (n5819,n5816,n5817);
or (n5820,n5821,n5824);
and (n5821,n5822,n5823);
xor (n5822,n5655,n5656);
and (n5823,n58,n378);
and (n5824,n5825,n5826);
xor (n5825,n5822,n5823);
or (n5826,n5827,n5830);
and (n5827,n5828,n5829);
xor (n5828,n5661,n5662);
and (n5829,n90,n378);
and (n5830,n5831,n5832);
xor (n5831,n5828,n5829);
or (n5832,n5833,n5836);
and (n5833,n5834,n5835);
xor (n5834,n5667,n5668);
and (n5835,n84,n378);
and (n5836,n5837,n5838);
xor (n5837,n5834,n5835);
or (n5838,n5839,n5842);
and (n5839,n5840,n5841);
xor (n5840,n5673,n5674);
and (n5841,n224,n378);
and (n5842,n5843,n5844);
xor (n5843,n5840,n5841);
or (n5844,n5845,n5848);
and (n5845,n5846,n5847);
xor (n5846,n5679,n5680);
and (n5847,n218,n378);
and (n5848,n5849,n5850);
xor (n5849,n5846,n5847);
or (n5850,n5851,n5854);
and (n5851,n5852,n5853);
xor (n5852,n5685,n5686);
and (n5853,n247,n378);
and (n5854,n5855,n5856);
xor (n5855,n5852,n5853);
or (n5856,n5857,n5859);
and (n5857,n5858,n2386);
xor (n5858,n5691,n5692);
and (n5859,n5860,n5861);
xor (n5860,n5858,n2386);
or (n5861,n5862,n5865);
and (n5862,n5863,n5864);
xor (n5863,n5697,n5698);
and (n5864,n174,n378);
and (n5865,n5866,n5867);
xor (n5866,n5863,n5864);
or (n5867,n5868,n5871);
and (n5868,n5869,n5870);
xor (n5869,n5703,n5704);
and (n5870,n166,n378);
and (n5871,n5872,n5873);
xor (n5872,n5869,n5870);
or (n5873,n5874,n5877);
and (n5874,n5875,n5876);
xor (n5875,n5709,n5710);
and (n5876,n312,n378);
and (n5877,n5878,n5879);
xor (n5878,n5875,n5876);
or (n5879,n5880,n5883);
and (n5880,n5881,n5882);
xor (n5881,n5715,n5716);
and (n5882,n580,n378);
and (n5883,n5884,n5885);
xor (n5884,n5881,n5882);
or (n5885,n5886,n5889);
and (n5886,n5887,n5888);
xor (n5887,n5721,n5722);
and (n5888,n574,n378);
and (n5889,n5890,n5891);
xor (n5890,n5887,n5888);
or (n5891,n5892,n5895);
and (n5892,n5893,n5894);
xor (n5893,n5727,n5728);
and (n5894,n712,n378);
and (n5895,n5896,n5897);
xor (n5896,n5893,n5894);
or (n5897,n5898,n5901);
and (n5898,n5899,n5900);
xor (n5899,n5733,n5734);
and (n5900,n753,n378);
and (n5901,n5902,n5903);
xor (n5902,n5899,n5900);
or (n5903,n5904,n5907);
and (n5904,n5905,n5906);
xor (n5905,n5739,n5740);
and (n5906,n922,n378);
and (n5907,n5908,n5909);
xor (n5908,n5905,n5906);
or (n5909,n5910,n5913);
and (n5910,n5911,n5912);
xor (n5911,n5745,n5746);
and (n5912,n959,n378);
and (n5913,n5914,n5915);
xor (n5914,n5911,n5912);
and (n5915,n5916,n5917);
xor (n5916,n5751,n5752);
and (n5917,n1122,n378);
and (n5918,n469,n429);
or (n5919,n5920,n5923);
and (n5920,n5921,n5922);
xor (n5921,n5760,n5761);
and (n5922,n386,n429);
and (n5923,n5924,n5925);
xor (n5924,n5921,n5922);
or (n5925,n5926,n5929);
and (n5926,n5927,n5928);
xor (n5927,n5766,n5767);
and (n5928,n38,n429);
and (n5929,n5930,n5931);
xor (n5930,n5927,n5928);
or (n5931,n5932,n5935);
and (n5932,n5933,n5934);
xor (n5933,n5772,n5773);
and (n5934,n32,n429);
and (n5935,n5936,n5937);
xor (n5936,n5933,n5934);
or (n5937,n5938,n5941);
and (n5938,n5939,n5940);
xor (n5939,n5778,n5779);
and (n5940,n199,n429);
and (n5941,n5942,n5943);
xor (n5942,n5939,n5940);
or (n5943,n5944,n5947);
and (n5944,n5945,n5946);
xor (n5945,n5784,n5785);
and (n5946,n194,n429);
and (n5947,n5948,n5949);
xor (n5948,n5945,n5946);
or (n5949,n5950,n5953);
and (n5950,n5951,n5952);
xor (n5951,n5790,n5791);
and (n5952,n146,n429);
and (n5953,n5954,n5955);
xor (n5954,n5951,n5952);
or (n5955,n5956,n5959);
and (n5956,n5957,n5958);
xor (n5957,n5795,n5796);
and (n5958,n140,n429);
and (n5959,n5960,n5961);
xor (n5960,n5957,n5958);
or (n5961,n5962,n5965);
and (n5962,n5963,n5964);
xor (n5963,n5801,n5802);
and (n5964,n266,n429);
and (n5965,n5966,n5967);
xor (n5966,n5963,n5964);
or (n5967,n5968,n5971);
and (n5968,n5969,n5970);
xor (n5969,n5807,n5808);
and (n5970,n260,n429);
and (n5971,n5972,n5973);
xor (n5972,n5969,n5970);
or (n5973,n5974,n5977);
and (n5974,n5975,n5976);
xor (n5975,n5813,n5814);
and (n5976,n65,n429);
and (n5977,n5978,n5979);
xor (n5978,n5975,n5976);
or (n5979,n5980,n5983);
and (n5980,n5981,n5982);
xor (n5981,n5819,n5820);
and (n5982,n58,n429);
and (n5983,n5984,n5985);
xor (n5984,n5981,n5982);
or (n5985,n5986,n5989);
and (n5986,n5987,n5988);
xor (n5987,n5825,n5826);
and (n5988,n90,n429);
and (n5989,n5990,n5991);
xor (n5990,n5987,n5988);
or (n5991,n5992,n5995);
and (n5992,n5993,n5994);
xor (n5993,n5831,n5832);
and (n5994,n84,n429);
and (n5995,n5996,n5997);
xor (n5996,n5993,n5994);
or (n5997,n5998,n6001);
and (n5998,n5999,n6000);
xor (n5999,n5837,n5838);
and (n6000,n224,n429);
and (n6001,n6002,n6003);
xor (n6002,n5999,n6000);
or (n6003,n6004,n6007);
and (n6004,n6005,n6006);
xor (n6005,n5843,n5844);
and (n6006,n218,n429);
and (n6007,n6008,n6009);
xor (n6008,n6005,n6006);
or (n6009,n6010,n6013);
and (n6010,n6011,n6012);
xor (n6011,n5849,n5850);
and (n6012,n247,n429);
and (n6013,n6014,n6015);
xor (n6014,n6011,n6012);
or (n6015,n6016,n6019);
and (n6016,n6017,n6018);
xor (n6017,n5855,n5856);
and (n6018,n241,n429);
and (n6019,n6020,n6021);
xor (n6020,n6017,n6018);
or (n6021,n6022,n6025);
and (n6022,n6023,n6024);
xor (n6023,n5860,n5861);
and (n6024,n174,n429);
and (n6025,n6026,n6027);
xor (n6026,n6023,n6024);
or (n6027,n6028,n6031);
and (n6028,n6029,n6030);
xor (n6029,n5866,n5867);
and (n6030,n166,n429);
and (n6031,n6032,n6033);
xor (n6032,n6029,n6030);
or (n6033,n6034,n6037);
and (n6034,n6035,n6036);
xor (n6035,n5872,n5873);
and (n6036,n312,n429);
and (n6037,n6038,n6039);
xor (n6038,n6035,n6036);
or (n6039,n6040,n6043);
and (n6040,n6041,n6042);
xor (n6041,n5878,n5879);
and (n6042,n580,n429);
and (n6043,n6044,n6045);
xor (n6044,n6041,n6042);
or (n6045,n6046,n6049);
and (n6046,n6047,n6048);
xor (n6047,n5884,n5885);
and (n6048,n574,n429);
and (n6049,n6050,n6051);
xor (n6050,n6047,n6048);
or (n6051,n6052,n6055);
and (n6052,n6053,n6054);
xor (n6053,n5890,n5891);
and (n6054,n712,n429);
and (n6055,n6056,n6057);
xor (n6056,n6053,n6054);
or (n6057,n6058,n6061);
and (n6058,n6059,n6060);
xor (n6059,n5896,n5897);
and (n6060,n753,n429);
and (n6061,n6062,n6063);
xor (n6062,n6059,n6060);
or (n6063,n6064,n6067);
and (n6064,n6065,n6066);
xor (n6065,n5902,n5903);
and (n6066,n922,n429);
and (n6067,n6068,n6069);
xor (n6068,n6065,n6066);
or (n6069,n6070,n6073);
and (n6070,n6071,n6072);
xor (n6071,n5908,n5909);
and (n6072,n959,n429);
and (n6073,n6074,n6075);
xor (n6074,n6071,n6072);
and (n6075,n6076,n3619);
xor (n6076,n5914,n5915);
and (n6077,n386,n22);
or (n6078,n6079,n6082);
and (n6079,n6080,n6081);
xor (n6080,n5924,n5925);
and (n6081,n38,n22);
and (n6082,n6083,n6084);
xor (n6083,n6080,n6081);
or (n6084,n6085,n6088);
and (n6085,n6086,n6087);
xor (n6086,n5930,n5931);
and (n6087,n32,n22);
and (n6088,n6089,n6090);
xor (n6089,n6086,n6087);
or (n6090,n6091,n6094);
and (n6091,n6092,n6093);
xor (n6092,n5936,n5937);
and (n6093,n199,n22);
and (n6094,n6095,n6096);
xor (n6095,n6092,n6093);
or (n6096,n6097,n6100);
and (n6097,n6098,n6099);
xor (n6098,n5942,n5943);
and (n6099,n194,n22);
and (n6100,n6101,n6102);
xor (n6101,n6098,n6099);
or (n6102,n6103,n6106);
and (n6103,n6104,n6105);
xor (n6104,n5948,n5949);
and (n6105,n146,n22);
and (n6106,n6107,n6108);
xor (n6107,n6104,n6105);
or (n6108,n6109,n6112);
and (n6109,n6110,n6111);
xor (n6110,n5954,n5955);
and (n6111,n140,n22);
and (n6112,n6113,n6114);
xor (n6113,n6110,n6111);
or (n6114,n6115,n6118);
and (n6115,n6116,n6117);
xor (n6116,n5960,n5961);
and (n6117,n266,n22);
and (n6118,n6119,n6120);
xor (n6119,n6116,n6117);
or (n6120,n6121,n6124);
and (n6121,n6122,n6123);
xor (n6122,n5966,n5967);
and (n6123,n260,n22);
and (n6124,n6125,n6126);
xor (n6125,n6122,n6123);
or (n6126,n6127,n6129);
and (n6127,n6128,n1752);
xor (n6128,n5972,n5973);
and (n6129,n6130,n6131);
xor (n6130,n6128,n1752);
or (n6131,n6132,n6135);
and (n6132,n6133,n6134);
xor (n6133,n5978,n5979);
and (n6134,n58,n22);
and (n6135,n6136,n6137);
xor (n6136,n6133,n6134);
or (n6137,n6138,n6141);
and (n6138,n6139,n6140);
xor (n6139,n5984,n5985);
and (n6140,n90,n22);
and (n6141,n6142,n6143);
xor (n6142,n6139,n6140);
or (n6143,n6144,n6147);
and (n6144,n6145,n6146);
xor (n6145,n5990,n5991);
and (n6146,n84,n22);
and (n6147,n6148,n6149);
xor (n6148,n6145,n6146);
or (n6149,n6150,n6153);
and (n6150,n6151,n6152);
xor (n6151,n5996,n5997);
and (n6152,n224,n22);
and (n6153,n6154,n6155);
xor (n6154,n6151,n6152);
or (n6155,n6156,n6159);
and (n6156,n6157,n6158);
xor (n6157,n6002,n6003);
and (n6158,n218,n22);
and (n6159,n6160,n6161);
xor (n6160,n6157,n6158);
or (n6161,n6162,n6165);
and (n6162,n6163,n6164);
xor (n6163,n6008,n6009);
and (n6164,n247,n22);
and (n6165,n6166,n6167);
xor (n6166,n6163,n6164);
or (n6167,n6168,n6171);
and (n6168,n6169,n6170);
xor (n6169,n6014,n6015);
and (n6170,n241,n22);
and (n6171,n6172,n6173);
xor (n6172,n6169,n6170);
or (n6173,n6174,n6177);
and (n6174,n6175,n6176);
xor (n6175,n6020,n6021);
and (n6176,n174,n22);
and (n6177,n6178,n6179);
xor (n6178,n6175,n6176);
or (n6179,n6180,n6183);
and (n6180,n6181,n6182);
xor (n6181,n6026,n6027);
and (n6182,n166,n22);
and (n6183,n6184,n6185);
xor (n6184,n6181,n6182);
or (n6185,n6186,n6189);
and (n6186,n6187,n6188);
xor (n6187,n6032,n6033);
and (n6188,n312,n22);
and (n6189,n6190,n6191);
xor (n6190,n6187,n6188);
or (n6191,n6192,n6195);
and (n6192,n6193,n6194);
xor (n6193,n6038,n6039);
and (n6194,n580,n22);
and (n6195,n6196,n6197);
xor (n6196,n6193,n6194);
or (n6197,n6198,n6201);
and (n6198,n6199,n6200);
xor (n6199,n6044,n6045);
and (n6200,n574,n22);
and (n6201,n6202,n6203);
xor (n6202,n6199,n6200);
or (n6203,n6204,n6207);
and (n6204,n6205,n6206);
xor (n6205,n6050,n6051);
and (n6206,n712,n22);
and (n6207,n6208,n6209);
xor (n6208,n6205,n6206);
or (n6209,n6210,n6213);
and (n6210,n6211,n6212);
xor (n6211,n6056,n6057);
and (n6212,n753,n22);
and (n6213,n6214,n6215);
xor (n6214,n6211,n6212);
or (n6215,n6216,n6219);
and (n6216,n6217,n6218);
xor (n6217,n6062,n6063);
and (n6218,n922,n22);
and (n6219,n6220,n6221);
xor (n6220,n6217,n6218);
or (n6221,n6222,n6225);
and (n6222,n6223,n6224);
xor (n6223,n6068,n6069);
and (n6224,n959,n22);
and (n6225,n6226,n6227);
xor (n6226,n6223,n6224);
and (n6227,n6228,n6229);
xor (n6228,n6074,n6075);
and (n6229,n1122,n22);
and (n6230,n38,n20);
or (n6231,n6232,n6235);
and (n6232,n6233,n6234);
xor (n6233,n6083,n6084);
and (n6234,n32,n20);
and (n6235,n6236,n6237);
xor (n6236,n6233,n6234);
or (n6237,n6238,n6241);
and (n6238,n6239,n6240);
xor (n6239,n6089,n6090);
and (n6240,n199,n20);
and (n6241,n6242,n6243);
xor (n6242,n6239,n6240);
or (n6243,n6244,n6247);
and (n6244,n6245,n6246);
xor (n6245,n6095,n6096);
and (n6246,n194,n20);
and (n6247,n6248,n6249);
xor (n6248,n6245,n6246);
or (n6249,n6250,n6253);
and (n6250,n6251,n6252);
xor (n6251,n6101,n6102);
and (n6252,n146,n20);
and (n6253,n6254,n6255);
xor (n6254,n6251,n6252);
or (n6255,n6256,n6259);
and (n6256,n6257,n6258);
xor (n6257,n6107,n6108);
and (n6258,n140,n20);
and (n6259,n6260,n6261);
xor (n6260,n6257,n6258);
or (n6261,n6262,n6265);
and (n6262,n6263,n6264);
xor (n6263,n6113,n6114);
and (n6264,n266,n20);
and (n6265,n6266,n6267);
xor (n6266,n6263,n6264);
or (n6267,n6268,n6271);
and (n6268,n6269,n6270);
xor (n6269,n6119,n6120);
and (n6270,n260,n20);
and (n6271,n6272,n6273);
xor (n6272,n6269,n6270);
or (n6273,n6274,n6277);
and (n6274,n6275,n6276);
xor (n6275,n6125,n6126);
and (n6276,n65,n20);
and (n6277,n6278,n6279);
xor (n6278,n6275,n6276);
or (n6279,n6280,n6283);
and (n6280,n6281,n6282);
xor (n6281,n6130,n6131);
and (n6282,n58,n20);
and (n6283,n6284,n6285);
xor (n6284,n6281,n6282);
or (n6285,n6286,n6289);
and (n6286,n6287,n6288);
xor (n6287,n6136,n6137);
and (n6288,n90,n20);
and (n6289,n6290,n6291);
xor (n6290,n6287,n6288);
or (n6291,n6292,n6295);
and (n6292,n6293,n6294);
xor (n6293,n6142,n6143);
and (n6294,n84,n20);
and (n6295,n6296,n6297);
xor (n6296,n6293,n6294);
or (n6297,n6298,n6301);
and (n6298,n6299,n6300);
xor (n6299,n6148,n6149);
and (n6300,n224,n20);
and (n6301,n6302,n6303);
xor (n6302,n6299,n6300);
or (n6303,n6304,n6307);
and (n6304,n6305,n6306);
xor (n6305,n6154,n6155);
and (n6306,n218,n20);
and (n6307,n6308,n6309);
xor (n6308,n6305,n6306);
or (n6309,n6310,n6313);
and (n6310,n6311,n6312);
xor (n6311,n6160,n6161);
and (n6312,n247,n20);
and (n6313,n6314,n6315);
xor (n6314,n6311,n6312);
or (n6315,n6316,n6319);
and (n6316,n6317,n6318);
xor (n6317,n6166,n6167);
and (n6318,n241,n20);
and (n6319,n6320,n6321);
xor (n6320,n6317,n6318);
or (n6321,n6322,n6325);
and (n6322,n6323,n6324);
xor (n6323,n6172,n6173);
and (n6324,n174,n20);
and (n6325,n6326,n6327);
xor (n6326,n6323,n6324);
or (n6327,n6328,n6331);
and (n6328,n6329,n6330);
xor (n6329,n6178,n6179);
and (n6330,n166,n20);
and (n6331,n6332,n6333);
xor (n6332,n6329,n6330);
or (n6333,n6334,n6337);
and (n6334,n6335,n6336);
xor (n6335,n6184,n6185);
and (n6336,n312,n20);
and (n6337,n6338,n6339);
xor (n6338,n6335,n6336);
or (n6339,n6340,n6343);
and (n6340,n6341,n6342);
xor (n6341,n6190,n6191);
and (n6342,n580,n20);
and (n6343,n6344,n6345);
xor (n6344,n6341,n6342);
or (n6345,n6346,n6349);
and (n6346,n6347,n6348);
xor (n6347,n6196,n6197);
and (n6348,n574,n20);
and (n6349,n6350,n6351);
xor (n6350,n6347,n6348);
or (n6351,n6352,n6355);
and (n6352,n6353,n6354);
xor (n6353,n6202,n6203);
and (n6354,n712,n20);
and (n6355,n6356,n6357);
xor (n6356,n6353,n6354);
or (n6357,n6358,n6361);
and (n6358,n6359,n6360);
xor (n6359,n6208,n6209);
and (n6360,n753,n20);
and (n6361,n6362,n6363);
xor (n6362,n6359,n6360);
or (n6363,n6364,n6367);
and (n6364,n6365,n6366);
xor (n6365,n6214,n6215);
and (n6366,n922,n20);
and (n6367,n6368,n6369);
xor (n6368,n6365,n6366);
or (n6369,n6370,n6373);
and (n6370,n6371,n6372);
xor (n6371,n6220,n6221);
and (n6372,n959,n20);
and (n6373,n6374,n6375);
xor (n6374,n6371,n6372);
and (n6375,n6376,n2906);
xor (n6376,n6226,n6227);
and (n6377,n32,n26);
or (n6378,n6379,n6382);
and (n6379,n6380,n6381);
xor (n6380,n6236,n6237);
and (n6381,n199,n26);
and (n6382,n6383,n6384);
xor (n6383,n6380,n6381);
or (n6384,n6385,n6388);
and (n6385,n6386,n6387);
xor (n6386,n6242,n6243);
and (n6387,n194,n26);
and (n6388,n6389,n6390);
xor (n6389,n6386,n6387);
or (n6390,n6391,n6394);
and (n6391,n6392,n6393);
xor (n6392,n6248,n6249);
and (n6393,n146,n26);
and (n6394,n6395,n6396);
xor (n6395,n6392,n6393);
or (n6396,n6397,n6400);
and (n6397,n6398,n6399);
xor (n6398,n6254,n6255);
and (n6399,n140,n26);
and (n6400,n6401,n6402);
xor (n6401,n6398,n6399);
or (n6402,n6403,n6406);
and (n6403,n6404,n6405);
xor (n6404,n6260,n6261);
and (n6405,n266,n26);
and (n6406,n6407,n6408);
xor (n6407,n6404,n6405);
or (n6408,n6409,n6412);
and (n6409,n6410,n6411);
xor (n6410,n6266,n6267);
and (n6411,n260,n26);
and (n6412,n6413,n6414);
xor (n6413,n6410,n6411);
or (n6414,n6415,n6418);
and (n6415,n6416,n6417);
xor (n6416,n6272,n6273);
and (n6417,n65,n26);
and (n6418,n6419,n6420);
xor (n6419,n6416,n6417);
or (n6420,n6421,n6424);
and (n6421,n6422,n6423);
xor (n6422,n6278,n6279);
and (n6423,n58,n26);
and (n6424,n6425,n6426);
xor (n6425,n6422,n6423);
or (n6426,n6427,n6430);
and (n6427,n6428,n6429);
xor (n6428,n6284,n6285);
and (n6429,n90,n26);
and (n6430,n6431,n6432);
xor (n6431,n6428,n6429);
or (n6432,n6433,n6436);
and (n6433,n6434,n6435);
xor (n6434,n6290,n6291);
and (n6435,n84,n26);
and (n6436,n6437,n6438);
xor (n6437,n6434,n6435);
or (n6438,n6439,n6442);
and (n6439,n6440,n6441);
xor (n6440,n6296,n6297);
and (n6441,n224,n26);
and (n6442,n6443,n6444);
xor (n6443,n6440,n6441);
or (n6444,n6445,n6448);
and (n6445,n6446,n6447);
xor (n6446,n6302,n6303);
and (n6447,n218,n26);
and (n6448,n6449,n6450);
xor (n6449,n6446,n6447);
or (n6450,n6451,n6454);
and (n6451,n6452,n6453);
xor (n6452,n6308,n6309);
and (n6453,n247,n26);
and (n6454,n6455,n6456);
xor (n6455,n6452,n6453);
or (n6456,n6457,n6460);
and (n6457,n6458,n6459);
xor (n6458,n6314,n6315);
and (n6459,n241,n26);
and (n6460,n6461,n6462);
xor (n6461,n6458,n6459);
or (n6462,n6463,n6466);
and (n6463,n6464,n6465);
xor (n6464,n6320,n6321);
and (n6465,n174,n26);
and (n6466,n6467,n6468);
xor (n6467,n6464,n6465);
or (n6468,n6469,n6472);
and (n6469,n6470,n6471);
xor (n6470,n6326,n6327);
and (n6471,n166,n26);
and (n6472,n6473,n6474);
xor (n6473,n6470,n6471);
or (n6474,n6475,n6478);
and (n6475,n6476,n6477);
xor (n6476,n6332,n6333);
and (n6477,n312,n26);
and (n6478,n6479,n6480);
xor (n6479,n6476,n6477);
or (n6480,n6481,n6484);
and (n6481,n6482,n6483);
xor (n6482,n6338,n6339);
and (n6483,n580,n26);
and (n6484,n6485,n6486);
xor (n6485,n6482,n6483);
or (n6486,n6487,n6490);
and (n6487,n6488,n6489);
xor (n6488,n6344,n6345);
and (n6489,n574,n26);
and (n6490,n6491,n6492);
xor (n6491,n6488,n6489);
or (n6492,n6493,n6496);
and (n6493,n6494,n6495);
xor (n6494,n6350,n6351);
and (n6495,n712,n26);
and (n6496,n6497,n6498);
xor (n6497,n6494,n6495);
or (n6498,n6499,n6502);
and (n6499,n6500,n6501);
xor (n6500,n6356,n6357);
and (n6501,n753,n26);
and (n6502,n6503,n6504);
xor (n6503,n6500,n6501);
or (n6504,n6505,n6508);
and (n6505,n6506,n6507);
xor (n6506,n6362,n6363);
and (n6507,n922,n26);
and (n6508,n6509,n6510);
xor (n6509,n6506,n6507);
or (n6510,n6511,n6514);
and (n6511,n6512,n6513);
xor (n6512,n6368,n6369);
and (n6513,n959,n26);
and (n6514,n6515,n6516);
xor (n6515,n6512,n6513);
and (n6516,n6517,n6518);
xor (n6517,n6374,n6375);
and (n6518,n1122,n26);
and (n6519,n199,n185);
or (n6520,n6521,n6524);
and (n6521,n6522,n6523);
xor (n6522,n6383,n6384);
and (n6523,n194,n185);
and (n6524,n6525,n6526);
xor (n6525,n6522,n6523);
or (n6526,n6527,n6530);
and (n6527,n6528,n6529);
xor (n6528,n6389,n6390);
and (n6529,n146,n185);
and (n6530,n6531,n6532);
xor (n6531,n6528,n6529);
or (n6532,n6533,n6536);
and (n6533,n6534,n6535);
xor (n6534,n6395,n6396);
and (n6535,n140,n185);
and (n6536,n6537,n6538);
xor (n6537,n6534,n6535);
or (n6538,n6539,n6542);
and (n6539,n6540,n6541);
xor (n6540,n6401,n6402);
and (n6541,n266,n185);
and (n6542,n6543,n6544);
xor (n6543,n6540,n6541);
or (n6544,n6545,n6548);
and (n6545,n6546,n6547);
xor (n6546,n6407,n6408);
and (n6547,n260,n185);
and (n6548,n6549,n6550);
xor (n6549,n6546,n6547);
or (n6550,n6551,n6554);
and (n6551,n6552,n6553);
xor (n6552,n6413,n6414);
and (n6553,n65,n185);
and (n6554,n6555,n6556);
xor (n6555,n6552,n6553);
or (n6556,n6557,n6560);
and (n6557,n6558,n6559);
xor (n6558,n6419,n6420);
and (n6559,n58,n185);
and (n6560,n6561,n6562);
xor (n6561,n6558,n6559);
or (n6562,n6563,n6566);
and (n6563,n6564,n6565);
xor (n6564,n6425,n6426);
and (n6565,n90,n185);
and (n6566,n6567,n6568);
xor (n6567,n6564,n6565);
or (n6568,n6569,n6572);
and (n6569,n6570,n6571);
xor (n6570,n6431,n6432);
and (n6571,n84,n185);
and (n6572,n6573,n6574);
xor (n6573,n6570,n6571);
or (n6574,n6575,n6578);
and (n6575,n6576,n6577);
xor (n6576,n6437,n6438);
and (n6577,n224,n185);
and (n6578,n6579,n6580);
xor (n6579,n6576,n6577);
or (n6580,n6581,n6584);
and (n6581,n6582,n6583);
xor (n6582,n6443,n6444);
and (n6583,n218,n185);
and (n6584,n6585,n6586);
xor (n6585,n6582,n6583);
or (n6586,n6587,n6590);
and (n6587,n6588,n6589);
xor (n6588,n6449,n6450);
and (n6589,n247,n185);
and (n6590,n6591,n6592);
xor (n6591,n6588,n6589);
or (n6592,n6593,n6596);
and (n6593,n6594,n6595);
xor (n6594,n6455,n6456);
and (n6595,n241,n185);
and (n6596,n6597,n6598);
xor (n6597,n6594,n6595);
or (n6598,n6599,n6602);
and (n6599,n6600,n6601);
xor (n6600,n6461,n6462);
and (n6601,n174,n185);
and (n6602,n6603,n6604);
xor (n6603,n6600,n6601);
or (n6604,n6605,n6608);
and (n6605,n6606,n6607);
xor (n6606,n6467,n6468);
and (n6607,n166,n185);
and (n6608,n6609,n6610);
xor (n6609,n6606,n6607);
or (n6610,n6611,n6614);
and (n6611,n6612,n6613);
xor (n6612,n6473,n6474);
and (n6613,n312,n185);
and (n6614,n6615,n6616);
xor (n6615,n6612,n6613);
or (n6616,n6617,n6620);
and (n6617,n6618,n6619);
xor (n6618,n6479,n6480);
and (n6619,n580,n185);
and (n6620,n6621,n6622);
xor (n6621,n6618,n6619);
or (n6622,n6623,n6626);
and (n6623,n6624,n6625);
xor (n6624,n6485,n6486);
and (n6625,n574,n185);
and (n6626,n6627,n6628);
xor (n6627,n6624,n6625);
or (n6628,n6629,n6632);
and (n6629,n6630,n6631);
xor (n6630,n6491,n6492);
and (n6631,n712,n185);
and (n6632,n6633,n6634);
xor (n6633,n6630,n6631);
or (n6634,n6635,n6638);
and (n6635,n6636,n6637);
xor (n6636,n6497,n6498);
and (n6637,n753,n185);
and (n6638,n6639,n6640);
xor (n6639,n6636,n6637);
or (n6640,n6641,n6644);
and (n6641,n6642,n6643);
xor (n6642,n6503,n6504);
and (n6643,n922,n185);
and (n6644,n6645,n6646);
xor (n6645,n6642,n6643);
or (n6646,n6647,n6650);
and (n6647,n6648,n6649);
xor (n6648,n6509,n6510);
and (n6649,n959,n185);
and (n6650,n6651,n6652);
xor (n6651,n6648,n6649);
and (n6652,n6653,n2928);
xor (n6653,n6515,n6516);
and (n6654,n194,n128);
or (n6655,n6656,n6659);
and (n6656,n6657,n6658);
xor (n6657,n6525,n6526);
and (n6658,n146,n128);
and (n6659,n6660,n6661);
xor (n6660,n6657,n6658);
or (n6661,n6662,n6665);
and (n6662,n6663,n6664);
xor (n6663,n6531,n6532);
and (n6664,n140,n128);
and (n6665,n6666,n6667);
xor (n6666,n6663,n6664);
or (n6667,n6668,n6671);
and (n6668,n6669,n6670);
xor (n6669,n6537,n6538);
and (n6670,n266,n128);
and (n6671,n6672,n6673);
xor (n6672,n6669,n6670);
or (n6673,n6674,n6677);
and (n6674,n6675,n6676);
xor (n6675,n6543,n6544);
and (n6676,n260,n128);
and (n6677,n6678,n6679);
xor (n6678,n6675,n6676);
or (n6679,n6680,n6683);
and (n6680,n6681,n6682);
xor (n6681,n6549,n6550);
and (n6682,n65,n128);
and (n6683,n6684,n6685);
xor (n6684,n6681,n6682);
or (n6685,n6686,n6689);
and (n6686,n6687,n6688);
xor (n6687,n6555,n6556);
and (n6688,n58,n128);
and (n6689,n6690,n6691);
xor (n6690,n6687,n6688);
or (n6691,n6692,n6695);
and (n6692,n6693,n6694);
xor (n6693,n6561,n6562);
and (n6694,n90,n128);
and (n6695,n6696,n6697);
xor (n6696,n6693,n6694);
or (n6697,n6698,n6701);
and (n6698,n6699,n6700);
xor (n6699,n6567,n6568);
and (n6700,n84,n128);
and (n6701,n6702,n6703);
xor (n6702,n6699,n6700);
or (n6703,n6704,n6707);
and (n6704,n6705,n6706);
xor (n6705,n6573,n6574);
and (n6706,n224,n128);
and (n6707,n6708,n6709);
xor (n6708,n6705,n6706);
or (n6709,n6710,n6713);
and (n6710,n6711,n6712);
xor (n6711,n6579,n6580);
and (n6712,n218,n128);
and (n6713,n6714,n6715);
xor (n6714,n6711,n6712);
or (n6715,n6716,n6719);
and (n6716,n6717,n6718);
xor (n6717,n6585,n6586);
and (n6718,n247,n128);
and (n6719,n6720,n6721);
xor (n6720,n6717,n6718);
or (n6721,n6722,n6725);
and (n6722,n6723,n6724);
xor (n6723,n6591,n6592);
and (n6724,n241,n128);
and (n6725,n6726,n6727);
xor (n6726,n6723,n6724);
or (n6727,n6728,n6731);
and (n6728,n6729,n6730);
xor (n6729,n6597,n6598);
and (n6730,n174,n128);
and (n6731,n6732,n6733);
xor (n6732,n6729,n6730);
or (n6733,n6734,n6736);
and (n6734,n6735,n3238);
xor (n6735,n6603,n6604);
and (n6736,n6737,n6738);
xor (n6737,n6735,n3238);
or (n6738,n6739,n6742);
and (n6739,n6740,n6741);
xor (n6740,n6609,n6610);
and (n6741,n312,n128);
and (n6742,n6743,n6744);
xor (n6743,n6740,n6741);
or (n6744,n6745,n6748);
and (n6745,n6746,n6747);
xor (n6746,n6615,n6616);
and (n6747,n580,n128);
and (n6748,n6749,n6750);
xor (n6749,n6746,n6747);
or (n6750,n6751,n6753);
and (n6751,n6752,n2438);
xor (n6752,n6621,n6622);
and (n6753,n6754,n6755);
xor (n6754,n6752,n2438);
or (n6755,n6756,n6759);
and (n6756,n6757,n6758);
xor (n6757,n6627,n6628);
and (n6758,n712,n128);
and (n6759,n6760,n6761);
xor (n6760,n6757,n6758);
or (n6761,n6762,n6765);
and (n6762,n6763,n6764);
xor (n6763,n6633,n6634);
and (n6764,n753,n128);
and (n6765,n6766,n6767);
xor (n6766,n6763,n6764);
or (n6767,n6768,n6771);
and (n6768,n6769,n6770);
xor (n6769,n6639,n6640);
and (n6770,n922,n128);
and (n6771,n6772,n6773);
xor (n6772,n6769,n6770);
or (n6773,n6774,n6777);
and (n6774,n6775,n6776);
xor (n6775,n6645,n6646);
and (n6776,n959,n128);
and (n6777,n6778,n6779);
xor (n6778,n6775,n6776);
and (n6779,n6780,n6781);
xor (n6780,n6651,n6652);
and (n6781,n1122,n128);
and (n6782,n146,n130);
or (n6783,n6784,n6787);
and (n6784,n6785,n6786);
xor (n6785,n6660,n6661);
and (n6786,n140,n130);
and (n6787,n6788,n6789);
xor (n6788,n6785,n6786);
or (n6789,n6790,n6793);
and (n6790,n6791,n6792);
xor (n6791,n6666,n6667);
and (n6792,n266,n130);
and (n6793,n6794,n6795);
xor (n6794,n6791,n6792);
or (n6795,n6796,n6799);
and (n6796,n6797,n6798);
xor (n6797,n6672,n6673);
and (n6798,n260,n130);
and (n6799,n6800,n6801);
xor (n6800,n6797,n6798);
or (n6801,n6802,n6805);
and (n6802,n6803,n6804);
xor (n6803,n6678,n6679);
and (n6804,n65,n130);
and (n6805,n6806,n6807);
xor (n6806,n6803,n6804);
or (n6807,n6808,n6811);
and (n6808,n6809,n6810);
xor (n6809,n6684,n6685);
and (n6810,n58,n130);
and (n6811,n6812,n6813);
xor (n6812,n6809,n6810);
or (n6813,n6814,n6817);
and (n6814,n6815,n6816);
xor (n6815,n6690,n6691);
and (n6816,n90,n130);
and (n6817,n6818,n6819);
xor (n6818,n6815,n6816);
or (n6819,n6820,n6823);
and (n6820,n6821,n6822);
xor (n6821,n6696,n6697);
and (n6822,n84,n130);
and (n6823,n6824,n6825);
xor (n6824,n6821,n6822);
or (n6825,n6826,n6829);
and (n6826,n6827,n6828);
xor (n6827,n6702,n6703);
and (n6828,n224,n130);
and (n6829,n6830,n6831);
xor (n6830,n6827,n6828);
or (n6831,n6832,n6835);
and (n6832,n6833,n6834);
xor (n6833,n6708,n6709);
and (n6834,n218,n130);
and (n6835,n6836,n6837);
xor (n6836,n6833,n6834);
or (n6837,n6838,n6841);
and (n6838,n6839,n6840);
xor (n6839,n6714,n6715);
and (n6840,n247,n130);
and (n6841,n6842,n6843);
xor (n6842,n6839,n6840);
or (n6843,n6844,n6847);
and (n6844,n6845,n6846);
xor (n6845,n6720,n6721);
and (n6846,n241,n130);
and (n6847,n6848,n6849);
xor (n6848,n6845,n6846);
or (n6849,n6850,n6853);
and (n6850,n6851,n6852);
xor (n6851,n6726,n6727);
and (n6852,n174,n130);
and (n6853,n6854,n6855);
xor (n6854,n6851,n6852);
or (n6855,n6856,n6859);
and (n6856,n6857,n6858);
xor (n6857,n6732,n6733);
and (n6858,n166,n130);
and (n6859,n6860,n6861);
xor (n6860,n6857,n6858);
or (n6861,n6862,n6865);
and (n6862,n6863,n6864);
xor (n6863,n6737,n6738);
and (n6864,n312,n130);
and (n6865,n6866,n6867);
xor (n6866,n6863,n6864);
or (n6867,n6868,n6871);
and (n6868,n6869,n6870);
xor (n6869,n6743,n6744);
and (n6870,n580,n130);
and (n6871,n6872,n6873);
xor (n6872,n6869,n6870);
or (n6873,n6874,n6877);
and (n6874,n6875,n6876);
xor (n6875,n6749,n6750);
and (n6876,n574,n130);
and (n6877,n6878,n6879);
xor (n6878,n6875,n6876);
or (n6879,n6880,n6883);
and (n6880,n6881,n6882);
xor (n6881,n6754,n6755);
and (n6882,n712,n130);
and (n6883,n6884,n6885);
xor (n6884,n6881,n6882);
or (n6885,n6886,n6889);
and (n6886,n6887,n6888);
xor (n6887,n6760,n6761);
and (n6888,n753,n130);
and (n6889,n6890,n6891);
xor (n6890,n6887,n6888);
or (n6891,n6892,n6895);
and (n6892,n6893,n6894);
xor (n6893,n6766,n6767);
and (n6894,n922,n130);
and (n6895,n6896,n6897);
xor (n6896,n6893,n6894);
or (n6897,n6898,n6901);
and (n6898,n6899,n6900);
xor (n6899,n6772,n6773);
and (n6900,n959,n130);
and (n6901,n6902,n6903);
xor (n6902,n6899,n6900);
and (n6903,n6904,n2682);
xor (n6904,n6778,n6779);
and (n6905,n140,n136);
or (n6906,n6907,n6910);
and (n6907,n6908,n6909);
xor (n6908,n6788,n6789);
and (n6909,n266,n136);
and (n6910,n6911,n6912);
xor (n6911,n6908,n6909);
or (n6912,n6913,n6916);
and (n6913,n6914,n6915);
xor (n6914,n6794,n6795);
and (n6915,n260,n136);
and (n6916,n6917,n6918);
xor (n6917,n6914,n6915);
or (n6918,n6919,n6922);
and (n6919,n6920,n6921);
xor (n6920,n6800,n6801);
and (n6921,n65,n136);
and (n6922,n6923,n6924);
xor (n6923,n6920,n6921);
or (n6924,n6925,n6928);
and (n6925,n6926,n6927);
xor (n6926,n6806,n6807);
and (n6927,n58,n136);
and (n6928,n6929,n6930);
xor (n6929,n6926,n6927);
or (n6930,n6931,n6934);
and (n6931,n6932,n6933);
xor (n6932,n6812,n6813);
and (n6933,n90,n136);
and (n6934,n6935,n6936);
xor (n6935,n6932,n6933);
or (n6936,n6937,n6940);
and (n6937,n6938,n6939);
xor (n6938,n6818,n6819);
and (n6939,n84,n136);
and (n6940,n6941,n6942);
xor (n6941,n6938,n6939);
or (n6942,n6943,n6946);
and (n6943,n6944,n6945);
xor (n6944,n6824,n6825);
and (n6945,n224,n136);
and (n6946,n6947,n6948);
xor (n6947,n6944,n6945);
or (n6948,n6949,n6952);
and (n6949,n6950,n6951);
xor (n6950,n6830,n6831);
and (n6951,n218,n136);
and (n6952,n6953,n6954);
xor (n6953,n6950,n6951);
or (n6954,n6955,n6958);
and (n6955,n6956,n6957);
xor (n6956,n6836,n6837);
and (n6957,n247,n136);
and (n6958,n6959,n6960);
xor (n6959,n6956,n6957);
or (n6960,n6961,n6964);
and (n6961,n6962,n6963);
xor (n6962,n6842,n6843);
and (n6963,n241,n136);
and (n6964,n6965,n6966);
xor (n6965,n6962,n6963);
or (n6966,n6967,n6970);
and (n6967,n6968,n6969);
xor (n6968,n6848,n6849);
and (n6969,n174,n136);
and (n6970,n6971,n6972);
xor (n6971,n6968,n6969);
or (n6972,n6973,n6976);
and (n6973,n6974,n6975);
xor (n6974,n6854,n6855);
and (n6975,n166,n136);
and (n6976,n6977,n6978);
xor (n6977,n6974,n6975);
or (n6978,n6979,n6982);
and (n6979,n6980,n6981);
xor (n6980,n6860,n6861);
and (n6981,n312,n136);
and (n6982,n6983,n6984);
xor (n6983,n6980,n6981);
or (n6984,n6985,n6988);
and (n6985,n6986,n6987);
xor (n6986,n6866,n6867);
and (n6987,n580,n136);
and (n6988,n6989,n6990);
xor (n6989,n6986,n6987);
or (n6990,n6991,n6994);
and (n6991,n6992,n6993);
xor (n6992,n6872,n6873);
and (n6993,n574,n136);
and (n6994,n6995,n6996);
xor (n6995,n6992,n6993);
or (n6996,n6997,n7000);
and (n6997,n6998,n6999);
xor (n6998,n6878,n6879);
and (n6999,n712,n136);
and (n7000,n7001,n7002);
xor (n7001,n6998,n6999);
or (n7002,n7003,n7006);
and (n7003,n7004,n7005);
xor (n7004,n6884,n6885);
and (n7005,n753,n136);
and (n7006,n7007,n7008);
xor (n7007,n7004,n7005);
or (n7008,n7009,n7012);
and (n7009,n7010,n7011);
xor (n7010,n6890,n6891);
and (n7011,n922,n136);
and (n7012,n7013,n7014);
xor (n7013,n7010,n7011);
or (n7014,n7015,n7018);
and (n7015,n7016,n7017);
xor (n7016,n6896,n6897);
and (n7017,n959,n136);
and (n7018,n7019,n7020);
xor (n7019,n7016,n7017);
and (n7020,n7021,n7022);
xor (n7021,n6902,n6903);
and (n7022,n1122,n136);
and (n7023,n266,n412);
or (n7024,n7025,n7028);
and (n7025,n7026,n7027);
xor (n7026,n6911,n6912);
and (n7027,n260,n412);
and (n7028,n7029,n7030);
xor (n7029,n7026,n7027);
or (n7030,n7031,n7034);
and (n7031,n7032,n7033);
xor (n7032,n6917,n6918);
and (n7033,n65,n412);
and (n7034,n7035,n7036);
xor (n7035,n7032,n7033);
or (n7036,n7037,n7040);
and (n7037,n7038,n7039);
xor (n7038,n6923,n6924);
and (n7039,n58,n412);
and (n7040,n7041,n7042);
xor (n7041,n7038,n7039);
or (n7042,n7043,n7046);
and (n7043,n7044,n7045);
xor (n7044,n6929,n6930);
and (n7045,n90,n412);
and (n7046,n7047,n7048);
xor (n7047,n7044,n7045);
or (n7048,n7049,n7052);
and (n7049,n7050,n7051);
xor (n7050,n6935,n6936);
and (n7051,n84,n412);
and (n7052,n7053,n7054);
xor (n7053,n7050,n7051);
or (n7054,n7055,n7058);
and (n7055,n7056,n7057);
xor (n7056,n6941,n6942);
and (n7057,n224,n412);
and (n7058,n7059,n7060);
xor (n7059,n7056,n7057);
or (n7060,n7061,n7064);
and (n7061,n7062,n7063);
xor (n7062,n6947,n6948);
and (n7063,n218,n412);
and (n7064,n7065,n7066);
xor (n7065,n7062,n7063);
or (n7066,n7067,n7070);
and (n7067,n7068,n7069);
xor (n7068,n6953,n6954);
and (n7069,n247,n412);
and (n7070,n7071,n7072);
xor (n7071,n7068,n7069);
or (n7072,n7073,n7076);
and (n7073,n7074,n7075);
xor (n7074,n6959,n6960);
and (n7075,n241,n412);
and (n7076,n7077,n7078);
xor (n7077,n7074,n7075);
or (n7078,n7079,n7082);
and (n7079,n7080,n7081);
xor (n7080,n6965,n6966);
and (n7081,n174,n412);
and (n7082,n7083,n7084);
xor (n7083,n7080,n7081);
or (n7084,n7085,n7088);
and (n7085,n7086,n7087);
xor (n7086,n6971,n6972);
and (n7087,n166,n412);
and (n7088,n7089,n7090);
xor (n7089,n7086,n7087);
or (n7090,n7091,n7094);
and (n7091,n7092,n7093);
xor (n7092,n6977,n6978);
and (n7093,n312,n412);
and (n7094,n7095,n7096);
xor (n7095,n7092,n7093);
or (n7096,n7097,n7100);
and (n7097,n7098,n7099);
xor (n7098,n6983,n6984);
and (n7099,n580,n412);
and (n7100,n7101,n7102);
xor (n7101,n7098,n7099);
or (n7102,n7103,n7106);
and (n7103,n7104,n7105);
xor (n7104,n6989,n6990);
and (n7105,n574,n412);
and (n7106,n7107,n7108);
xor (n7107,n7104,n7105);
or (n7108,n7109,n7112);
and (n7109,n7110,n7111);
xor (n7110,n6995,n6996);
and (n7111,n712,n412);
and (n7112,n7113,n7114);
xor (n7113,n7110,n7111);
or (n7114,n7115,n7118);
and (n7115,n7116,n7117);
xor (n7116,n7001,n7002);
and (n7117,n753,n412);
and (n7118,n7119,n7120);
xor (n7119,n7116,n7117);
or (n7120,n7121,n7124);
and (n7121,n7122,n7123);
xor (n7122,n7007,n7008);
and (n7123,n922,n412);
and (n7124,n7125,n7126);
xor (n7125,n7122,n7123);
or (n7126,n7127,n7130);
and (n7127,n7128,n7129);
xor (n7128,n7013,n7014);
and (n7129,n959,n412);
and (n7130,n7131,n7132);
xor (n7131,n7128,n7129);
and (n7132,n7133,n2303);
xor (n7133,n7019,n7020);
and (n7134,n260,n47);
or (n7135,n7136,n7139);
and (n7136,n7137,n7138);
xor (n7137,n7029,n7030);
and (n7138,n65,n47);
and (n7139,n7140,n7141);
xor (n7140,n7137,n7138);
or (n7141,n7142,n7145);
and (n7142,n7143,n7144);
xor (n7143,n7035,n7036);
and (n7144,n58,n47);
and (n7145,n7146,n7147);
xor (n7146,n7143,n7144);
or (n7147,n7148,n7151);
and (n7148,n7149,n7150);
xor (n7149,n7041,n7042);
and (n7150,n90,n47);
and (n7151,n7152,n7153);
xor (n7152,n7149,n7150);
or (n7153,n7154,n7157);
and (n7154,n7155,n7156);
xor (n7155,n7047,n7048);
and (n7156,n84,n47);
and (n7157,n7158,n7159);
xor (n7158,n7155,n7156);
or (n7159,n7160,n7163);
and (n7160,n7161,n7162);
xor (n7161,n7053,n7054);
and (n7162,n224,n47);
and (n7163,n7164,n7165);
xor (n7164,n7161,n7162);
or (n7165,n7166,n7169);
and (n7166,n7167,n7168);
xor (n7167,n7059,n7060);
and (n7168,n218,n47);
and (n7169,n7170,n7171);
xor (n7170,n7167,n7168);
or (n7171,n7172,n7175);
and (n7172,n7173,n7174);
xor (n7173,n7065,n7066);
and (n7174,n247,n47);
and (n7175,n7176,n7177);
xor (n7176,n7173,n7174);
or (n7177,n7178,n7180);
and (n7178,n7179,n1485);
xor (n7179,n7071,n7072);
and (n7180,n7181,n7182);
xor (n7181,n7179,n1485);
or (n7182,n7183,n7185);
and (n7183,n7184,n1671);
xor (n7184,n7077,n7078);
and (n7185,n7186,n7187);
xor (n7186,n7184,n1671);
or (n7187,n7188,n7191);
and (n7188,n7189,n7190);
xor (n7189,n7083,n7084);
and (n7190,n166,n47);
and (n7191,n7192,n7193);
xor (n7192,n7189,n7190);
or (n7193,n7194,n7197);
and (n7194,n7195,n7196);
xor (n7195,n7089,n7090);
and (n7196,n312,n47);
and (n7197,n7198,n7199);
xor (n7198,n7195,n7196);
or (n7199,n7200,n7203);
and (n7200,n7201,n7202);
xor (n7201,n7095,n7096);
and (n7202,n580,n47);
and (n7203,n7204,n7205);
xor (n7204,n7201,n7202);
or (n7205,n7206,n7209);
and (n7206,n7207,n7208);
xor (n7207,n7101,n7102);
and (n7208,n574,n47);
and (n7209,n7210,n7211);
xor (n7210,n7207,n7208);
or (n7211,n7212,n7214);
and (n7212,n7213,n3263);
xor (n7213,n7107,n7108);
and (n7214,n7215,n7216);
xor (n7215,n7213,n3263);
or (n7216,n7217,n7219);
and (n7217,n7218,n2559);
xor (n7218,n7113,n7114);
and (n7219,n7220,n7221);
xor (n7220,n7218,n2559);
or (n7221,n7222,n7225);
and (n7222,n7223,n7224);
xor (n7223,n7119,n7120);
and (n7224,n922,n47);
and (n7225,n7226,n7227);
xor (n7226,n7223,n7224);
or (n7227,n7228,n7231);
and (n7228,n7229,n7230);
xor (n7229,n7125,n7126);
and (n7230,n959,n47);
and (n7231,n7232,n7233);
xor (n7232,n7229,n7230);
and (n7233,n7234,n7235);
xor (n7234,n7131,n7132);
and (n7235,n1122,n47);
and (n7236,n65,n49);
or (n7237,n7238,n7241);
and (n7238,n7239,n7240);
xor (n7239,n7140,n7141);
and (n7240,n58,n49);
and (n7241,n7242,n7243);
xor (n7242,n7239,n7240);
or (n7243,n7244,n7247);
and (n7244,n7245,n7246);
xor (n7245,n7146,n7147);
and (n7246,n90,n49);
and (n7247,n7248,n7249);
xor (n7248,n7245,n7246);
or (n7249,n7250,n7253);
and (n7250,n7251,n7252);
xor (n7251,n7152,n7153);
and (n7252,n84,n49);
and (n7253,n7254,n7255);
xor (n7254,n7251,n7252);
or (n7255,n7256,n7259);
and (n7256,n7257,n7258);
xor (n7257,n7158,n7159);
and (n7258,n224,n49);
and (n7259,n7260,n7261);
xor (n7260,n7257,n7258);
or (n7261,n7262,n7265);
and (n7262,n7263,n7264);
xor (n7263,n7164,n7165);
and (n7264,n218,n49);
and (n7265,n7266,n7267);
xor (n7266,n7263,n7264);
or (n7267,n7268,n7271);
and (n7268,n7269,n7270);
xor (n7269,n7170,n7171);
and (n7270,n247,n49);
and (n7271,n7272,n7273);
xor (n7272,n7269,n7270);
or (n7273,n7274,n7277);
and (n7274,n7275,n7276);
xor (n7275,n7176,n7177);
and (n7276,n241,n49);
and (n7277,n7278,n7279);
xor (n7278,n7275,n7276);
or (n7279,n7280,n7283);
and (n7280,n7281,n7282);
xor (n7281,n7181,n7182);
and (n7282,n174,n49);
and (n7283,n7284,n7285);
xor (n7284,n7281,n7282);
or (n7285,n7286,n7289);
and (n7286,n7287,n7288);
xor (n7287,n7186,n7187);
and (n7288,n166,n49);
and (n7289,n7290,n7291);
xor (n7290,n7287,n7288);
or (n7291,n7292,n7295);
and (n7292,n7293,n7294);
xor (n7293,n7192,n7193);
and (n7294,n312,n49);
and (n7295,n7296,n7297);
xor (n7296,n7293,n7294);
or (n7297,n7298,n7301);
and (n7298,n7299,n7300);
xor (n7299,n7198,n7199);
and (n7300,n580,n49);
and (n7301,n7302,n7303);
xor (n7302,n7299,n7300);
or (n7303,n7304,n7307);
and (n7304,n7305,n7306);
xor (n7305,n7204,n7205);
and (n7306,n574,n49);
and (n7307,n7308,n7309);
xor (n7308,n7305,n7306);
or (n7309,n7310,n7313);
and (n7310,n7311,n7312);
xor (n7311,n7210,n7211);
and (n7312,n712,n49);
and (n7313,n7314,n7315);
xor (n7314,n7311,n7312);
or (n7315,n7316,n7319);
and (n7316,n7317,n7318);
xor (n7317,n7215,n7216);
and (n7318,n753,n49);
and (n7319,n7320,n7321);
xor (n7320,n7317,n7318);
or (n7321,n7322,n7325);
and (n7322,n7323,n7324);
xor (n7323,n7220,n7221);
and (n7324,n922,n49);
and (n7325,n7326,n7327);
xor (n7326,n7323,n7324);
or (n7327,n7328,n7331);
and (n7328,n7329,n7330);
xor (n7329,n7226,n7227);
and (n7330,n959,n49);
and (n7331,n7332,n7333);
xor (n7332,n7329,n7330);
and (n7333,n7334,n2616);
xor (n7334,n7232,n7233);
and (n7335,n58,n54);
or (n7336,n7337,n7340);
and (n7337,n7338,n7339);
xor (n7338,n7242,n7243);
and (n7339,n90,n54);
and (n7340,n7341,n7342);
xor (n7341,n7338,n7339);
or (n7342,n7343,n7346);
and (n7343,n7344,n7345);
xor (n7344,n7248,n7249);
and (n7345,n84,n54);
and (n7346,n7347,n7348);
xor (n7347,n7344,n7345);
or (n7348,n7349,n7352);
and (n7349,n7350,n7351);
xor (n7350,n7254,n7255);
and (n7351,n224,n54);
and (n7352,n7353,n7354);
xor (n7353,n7350,n7351);
or (n7354,n7355,n7358);
and (n7355,n7356,n7357);
xor (n7356,n7260,n7261);
and (n7357,n218,n54);
and (n7358,n7359,n7360);
xor (n7359,n7356,n7357);
or (n7360,n7361,n7364);
and (n7361,n7362,n7363);
xor (n7362,n7266,n7267);
and (n7363,n247,n54);
and (n7364,n7365,n7366);
xor (n7365,n7362,n7363);
or (n7366,n7367,n7370);
and (n7367,n7368,n7369);
xor (n7368,n7272,n7273);
and (n7369,n241,n54);
and (n7370,n7371,n7372);
xor (n7371,n7368,n7369);
or (n7372,n7373,n7376);
and (n7373,n7374,n7375);
xor (n7374,n7278,n7279);
and (n7375,n174,n54);
and (n7376,n7377,n7378);
xor (n7377,n7374,n7375);
or (n7378,n7379,n7382);
and (n7379,n7380,n7381);
xor (n7380,n7284,n7285);
and (n7381,n166,n54);
and (n7382,n7383,n7384);
xor (n7383,n7380,n7381);
or (n7384,n7385,n7388);
and (n7385,n7386,n7387);
xor (n7386,n7290,n7291);
and (n7387,n312,n54);
and (n7388,n7389,n7390);
xor (n7389,n7386,n7387);
or (n7390,n7391,n7394);
and (n7391,n7392,n7393);
xor (n7392,n7296,n7297);
and (n7393,n580,n54);
and (n7394,n7395,n7396);
xor (n7395,n7392,n7393);
or (n7396,n7397,n7400);
and (n7397,n7398,n7399);
xor (n7398,n7302,n7303);
and (n7399,n574,n54);
and (n7400,n7401,n7402);
xor (n7401,n7398,n7399);
or (n7402,n7403,n7406);
and (n7403,n7404,n7405);
xor (n7404,n7308,n7309);
and (n7405,n712,n54);
and (n7406,n7407,n7408);
xor (n7407,n7404,n7405);
or (n7408,n7409,n7412);
and (n7409,n7410,n7411);
xor (n7410,n7314,n7315);
and (n7411,n753,n54);
and (n7412,n7413,n7414);
xor (n7413,n7410,n7411);
or (n7414,n7415,n7418);
and (n7415,n7416,n7417);
xor (n7416,n7320,n7321);
and (n7417,n922,n54);
and (n7418,n7419,n7420);
xor (n7419,n7416,n7417);
or (n7420,n7421,n7424);
and (n7421,n7422,n7423);
xor (n7422,n7326,n7327);
and (n7423,n959,n54);
and (n7424,n7425,n7426);
xor (n7425,n7422,n7423);
and (n7426,n7427,n7428);
xor (n7427,n7332,n7333);
and (n7428,n1122,n54);
and (n7429,n90,n75);
or (n7430,n7431,n7434);
and (n7431,n7432,n7433);
xor (n7432,n7341,n7342);
and (n7433,n84,n75);
and (n7434,n7435,n7436);
xor (n7435,n7432,n7433);
or (n7436,n7437,n7440);
and (n7437,n7438,n7439);
xor (n7438,n7347,n7348);
and (n7439,n224,n75);
and (n7440,n7441,n7442);
xor (n7441,n7438,n7439);
or (n7442,n7443,n7446);
and (n7443,n7444,n7445);
xor (n7444,n7353,n7354);
and (n7445,n218,n75);
and (n7446,n7447,n7448);
xor (n7447,n7444,n7445);
or (n7448,n7449,n7452);
and (n7449,n7450,n7451);
xor (n7450,n7359,n7360);
and (n7451,n247,n75);
and (n7452,n7453,n7454);
xor (n7453,n7450,n7451);
or (n7454,n7455,n7458);
and (n7455,n7456,n7457);
xor (n7456,n7365,n7366);
and (n7457,n241,n75);
and (n7458,n7459,n7460);
xor (n7459,n7456,n7457);
or (n7460,n7461,n7464);
and (n7461,n7462,n7463);
xor (n7462,n7371,n7372);
and (n7463,n174,n75);
and (n7464,n7465,n7466);
xor (n7465,n7462,n7463);
or (n7466,n7467,n7470);
and (n7467,n7468,n7469);
xor (n7468,n7377,n7378);
and (n7469,n166,n75);
and (n7470,n7471,n7472);
xor (n7471,n7468,n7469);
or (n7472,n7473,n7476);
and (n7473,n7474,n7475);
xor (n7474,n7383,n7384);
and (n7475,n312,n75);
and (n7476,n7477,n7478);
xor (n7477,n7474,n7475);
or (n7478,n7479,n7482);
and (n7479,n7480,n7481);
xor (n7480,n7389,n7390);
and (n7481,n580,n75);
and (n7482,n7483,n7484);
xor (n7483,n7480,n7481);
or (n7484,n7485,n7488);
and (n7485,n7486,n7487);
xor (n7486,n7395,n7396);
and (n7487,n574,n75);
and (n7488,n7489,n7490);
xor (n7489,n7486,n7487);
or (n7490,n7491,n7494);
and (n7491,n7492,n7493);
xor (n7492,n7401,n7402);
and (n7493,n712,n75);
and (n7494,n7495,n7496);
xor (n7495,n7492,n7493);
or (n7496,n7497,n7500);
and (n7497,n7498,n7499);
xor (n7498,n7407,n7408);
and (n7499,n753,n75);
and (n7500,n7501,n7502);
xor (n7501,n7498,n7499);
or (n7502,n7503,n7506);
and (n7503,n7504,n7505);
xor (n7504,n7413,n7414);
and (n7505,n922,n75);
and (n7506,n7507,n7508);
xor (n7507,n7504,n7505);
or (n7508,n7509,n7512);
and (n7509,n7510,n7511);
xor (n7510,n7419,n7420);
and (n7511,n959,n75);
and (n7512,n7513,n7514);
xor (n7513,n7510,n7511);
and (n7514,n7515,n3366);
xor (n7515,n7425,n7426);
and (n7516,n84,n80);
or (n7517,n7518,n7521);
and (n7518,n7519,n7520);
xor (n7519,n7435,n7436);
and (n7520,n224,n80);
and (n7521,n7522,n7523);
xor (n7522,n7519,n7520);
or (n7523,n7524,n7527);
and (n7524,n7525,n7526);
xor (n7525,n7441,n7442);
and (n7526,n218,n80);
and (n7527,n7528,n7529);
xor (n7528,n7525,n7526);
or (n7529,n7530,n7533);
and (n7530,n7531,n7532);
xor (n7531,n7447,n7448);
and (n7532,n247,n80);
and (n7533,n7534,n7535);
xor (n7534,n7531,n7532);
or (n7535,n7536,n7539);
and (n7536,n7537,n7538);
xor (n7537,n7453,n7454);
and (n7538,n241,n80);
and (n7539,n7540,n7541);
xor (n7540,n7537,n7538);
or (n7541,n7542,n7545);
and (n7542,n7543,n7544);
xor (n7543,n7459,n7460);
and (n7544,n174,n80);
and (n7545,n7546,n7547);
xor (n7546,n7543,n7544);
or (n7547,n7548,n7551);
and (n7548,n7549,n7550);
xor (n7549,n7465,n7466);
and (n7550,n166,n80);
and (n7551,n7552,n7553);
xor (n7552,n7549,n7550);
or (n7553,n7554,n7557);
and (n7554,n7555,n7556);
xor (n7555,n7471,n7472);
and (n7556,n312,n80);
and (n7557,n7558,n7559);
xor (n7558,n7555,n7556);
or (n7559,n7560,n7563);
and (n7560,n7561,n7562);
xor (n7561,n7477,n7478);
and (n7562,n580,n80);
and (n7563,n7564,n7565);
xor (n7564,n7561,n7562);
or (n7565,n7566,n7569);
and (n7566,n7567,n7568);
xor (n7567,n7483,n7484);
and (n7568,n574,n80);
and (n7569,n7570,n7571);
xor (n7570,n7567,n7568);
or (n7571,n7572,n7575);
and (n7572,n7573,n7574);
xor (n7573,n7489,n7490);
and (n7574,n712,n80);
and (n7575,n7576,n7577);
xor (n7576,n7573,n7574);
or (n7577,n7578,n7581);
and (n7578,n7579,n7580);
xor (n7579,n7495,n7496);
and (n7580,n753,n80);
and (n7581,n7582,n7583);
xor (n7582,n7579,n7580);
or (n7583,n7584,n7587);
and (n7584,n7585,n7586);
xor (n7585,n7501,n7502);
and (n7586,n922,n80);
and (n7587,n7588,n7589);
xor (n7588,n7585,n7586);
or (n7589,n7590,n7593);
and (n7590,n7591,n7592);
xor (n7591,n7507,n7508);
and (n7592,n959,n80);
and (n7593,n7594,n7595);
xor (n7594,n7591,n7592);
and (n7595,n7596,n7597);
xor (n7596,n7513,n7514);
and (n7597,n1122,n80);
and (n7598,n224,n210);
or (n7599,n7600,n7603);
and (n7600,n7601,n7602);
xor (n7601,n7522,n7523);
and (n7602,n218,n210);
and (n7603,n7604,n7605);
xor (n7604,n7601,n7602);
or (n7605,n7606,n7609);
and (n7606,n7607,n7608);
xor (n7607,n7528,n7529);
and (n7608,n247,n210);
and (n7609,n7610,n7611);
xor (n7610,n7607,n7608);
or (n7611,n7612,n7615);
and (n7612,n7613,n7614);
xor (n7613,n7534,n7535);
and (n7614,n241,n210);
and (n7615,n7616,n7617);
xor (n7616,n7613,n7614);
or (n7617,n7618,n7621);
and (n7618,n7619,n7620);
xor (n7619,n7540,n7541);
and (n7620,n174,n210);
and (n7621,n7622,n7623);
xor (n7622,n7619,n7620);
or (n7623,n7624,n7627);
and (n7624,n7625,n7626);
xor (n7625,n7546,n7547);
and (n7626,n166,n210);
and (n7627,n7628,n7629);
xor (n7628,n7625,n7626);
or (n7629,n7630,n7633);
and (n7630,n7631,n7632);
xor (n7631,n7552,n7553);
and (n7632,n312,n210);
and (n7633,n7634,n7635);
xor (n7634,n7631,n7632);
or (n7635,n7636,n7639);
and (n7636,n7637,n7638);
xor (n7637,n7558,n7559);
and (n7638,n580,n210);
and (n7639,n7640,n7641);
xor (n7640,n7637,n7638);
or (n7641,n7642,n7645);
and (n7642,n7643,n7644);
xor (n7643,n7564,n7565);
and (n7644,n574,n210);
and (n7645,n7646,n7647);
xor (n7646,n7643,n7644);
or (n7647,n7648,n7651);
and (n7648,n7649,n7650);
xor (n7649,n7570,n7571);
and (n7650,n712,n210);
and (n7651,n7652,n7653);
xor (n7652,n7649,n7650);
or (n7653,n7654,n7657);
and (n7654,n7655,n7656);
xor (n7655,n7576,n7577);
and (n7656,n753,n210);
and (n7657,n7658,n7659);
xor (n7658,n7655,n7656);
or (n7659,n7660,n7663);
and (n7660,n7661,n7662);
xor (n7661,n7582,n7583);
and (n7662,n922,n210);
and (n7663,n7664,n7665);
xor (n7664,n7661,n7662);
or (n7665,n7666,n7669);
and (n7666,n7667,n7668);
xor (n7667,n7588,n7589);
and (n7668,n959,n210);
and (n7669,n7670,n7671);
xor (n7670,n7667,n7668);
and (n7671,n7672,n2130);
xor (n7672,n7594,n7595);
and (n7673,n218,n208);
or (n7674,n7675,n7678);
and (n7675,n7676,n7677);
xor (n7676,n7604,n7605);
and (n7677,n247,n208);
and (n7678,n7679,n7680);
xor (n7679,n7676,n7677);
or (n7680,n7681,n7683);
and (n7681,n7682,n305);
xor (n7682,n7610,n7611);
and (n7683,n7684,n7685);
xor (n7684,n7682,n305);
or (n7685,n7686,n7688);
and (n7686,n7687,n301);
xor (n7687,n7616,n7617);
and (n7688,n7689,n7690);
xor (n7689,n7687,n301);
or (n7690,n7691,n7694);
and (n7691,n7692,n7693);
xor (n7692,n7622,n7623);
and (n7693,n166,n208);
and (n7694,n7695,n7696);
xor (n7695,n7692,n7693);
or (n7696,n7697,n7700);
and (n7697,n7698,n7699);
xor (n7698,n7628,n7629);
and (n7699,n312,n208);
and (n7700,n7701,n7702);
xor (n7701,n7698,n7699);
or (n7702,n7703,n7706);
and (n7703,n7704,n7705);
xor (n7704,n7634,n7635);
and (n7705,n580,n208);
and (n7706,n7707,n7708);
xor (n7707,n7704,n7705);
or (n7708,n7709,n7712);
and (n7709,n7710,n7711);
xor (n7710,n7640,n7641);
and (n7711,n574,n208);
and (n7712,n7713,n7714);
xor (n7713,n7710,n7711);
or (n7714,n7715,n7718);
and (n7715,n7716,n7717);
xor (n7716,n7646,n7647);
and (n7717,n712,n208);
and (n7718,n7719,n7720);
xor (n7719,n7716,n7717);
or (n7720,n7721,n7724);
and (n7721,n7722,n7723);
xor (n7722,n7652,n7653);
and (n7723,n753,n208);
and (n7724,n7725,n7726);
xor (n7725,n7722,n7723);
or (n7726,n7727,n7730);
and (n7727,n7728,n7729);
xor (n7728,n7658,n7659);
and (n7729,n922,n208);
and (n7730,n7731,n7732);
xor (n7731,n7728,n7729);
or (n7732,n7733,n7736);
and (n7733,n7734,n7735);
xor (n7734,n7664,n7665);
and (n7735,n959,n208);
and (n7736,n7737,n7738);
xor (n7737,n7734,n7735);
and (n7738,n7739,n7740);
xor (n7739,n7670,n7671);
and (n7740,n1122,n208);
and (n7741,n247,n234);
or (n7742,n7743,n7746);
and (n7743,n7744,n7745);
xor (n7744,n7679,n7680);
and (n7745,n241,n234);
and (n7746,n7747,n7748);
xor (n7747,n7744,n7745);
or (n7748,n7749,n7752);
and (n7749,n7750,n7751);
xor (n7750,n7684,n7685);
and (n7751,n174,n234);
and (n7752,n7753,n7754);
xor (n7753,n7750,n7751);
or (n7754,n7755,n7758);
and (n7755,n7756,n7757);
xor (n7756,n7689,n7690);
and (n7757,n166,n234);
and (n7758,n7759,n7760);
xor (n7759,n7756,n7757);
or (n7760,n7761,n7764);
and (n7761,n7762,n7763);
xor (n7762,n7695,n7696);
and (n7763,n312,n234);
and (n7764,n7765,n7766);
xor (n7765,n7762,n7763);
or (n7766,n7767,n7770);
and (n7767,n7768,n7769);
xor (n7768,n7701,n7702);
and (n7769,n580,n234);
and (n7770,n7771,n7772);
xor (n7771,n7768,n7769);
or (n7772,n7773,n7776);
and (n7773,n7774,n7775);
xor (n7774,n7707,n7708);
and (n7775,n574,n234);
and (n7776,n7777,n7778);
xor (n7777,n7774,n7775);
or (n7778,n7779,n7782);
and (n7779,n7780,n7781);
xor (n7780,n7713,n7714);
and (n7781,n712,n234);
and (n7782,n7783,n7784);
xor (n7783,n7780,n7781);
or (n7784,n7785,n7788);
and (n7785,n7786,n7787);
xor (n7786,n7719,n7720);
and (n7787,n753,n234);
and (n7788,n7789,n7790);
xor (n7789,n7786,n7787);
or (n7790,n7791,n7794);
and (n7791,n7792,n7793);
xor (n7792,n7725,n7726);
and (n7793,n922,n234);
and (n7794,n7795,n7796);
xor (n7795,n7792,n7793);
or (n7796,n7797,n7800);
and (n7797,n7798,n7799);
xor (n7798,n7731,n7732);
and (n7799,n959,n234);
and (n7800,n7801,n7802);
xor (n7801,n7798,n7799);
and (n7802,n7803,n1879);
xor (n7803,n7737,n7738);
and (n7804,n241,n155);
or (n7805,n7806,n7809);
and (n7806,n7807,n7808);
xor (n7807,n7747,n7748);
and (n7808,n174,n155);
and (n7809,n7810,n7811);
xor (n7810,n7807,n7808);
or (n7811,n7812,n7815);
and (n7812,n7813,n7814);
xor (n7813,n7753,n7754);
and (n7814,n166,n155);
and (n7815,n7816,n7817);
xor (n7816,n7813,n7814);
or (n7817,n7818,n7821);
and (n7818,n7819,n7820);
xor (n7819,n7759,n7760);
and (n7820,n312,n155);
and (n7821,n7822,n7823);
xor (n7822,n7819,n7820);
or (n7823,n7824,n7827);
and (n7824,n7825,n7826);
xor (n7825,n7765,n7766);
and (n7826,n580,n155);
and (n7827,n7828,n7829);
xor (n7828,n7825,n7826);
or (n7829,n7830,n7833);
and (n7830,n7831,n7832);
xor (n7831,n7771,n7772);
and (n7832,n574,n155);
and (n7833,n7834,n7835);
xor (n7834,n7831,n7832);
or (n7835,n7836,n7839);
and (n7836,n7837,n7838);
xor (n7837,n7777,n7778);
and (n7838,n712,n155);
and (n7839,n7840,n7841);
xor (n7840,n7837,n7838);
or (n7841,n7842,n7845);
and (n7842,n7843,n7844);
xor (n7843,n7783,n7784);
and (n7844,n753,n155);
and (n7845,n7846,n7847);
xor (n7846,n7843,n7844);
or (n7847,n7848,n7851);
and (n7848,n7849,n7850);
xor (n7849,n7789,n7790);
and (n7850,n922,n155);
and (n7851,n7852,n7853);
xor (n7852,n7849,n7850);
or (n7853,n7854,n7857);
and (n7854,n7855,n7856);
xor (n7855,n7795,n7796);
and (n7856,n959,n155);
and (n7857,n7858,n7859);
xor (n7858,n7855,n7856);
and (n7859,n7860,n7861);
xor (n7860,n7801,n7802);
and (n7861,n1122,n155);
and (n7862,n174,n156);
or (n7863,n7864,n7867);
and (n7864,n7865,n7866);
xor (n7865,n7810,n7811);
and (n7866,n166,n156);
and (n7867,n7868,n7869);
xor (n7868,n7865,n7866);
or (n7869,n7870,n7873);
and (n7870,n7871,n7872);
xor (n7871,n7816,n7817);
and (n7872,n312,n156);
and (n7873,n7874,n7875);
xor (n7874,n7871,n7872);
or (n7875,n7876,n7879);
and (n7876,n7877,n7878);
xor (n7877,n7822,n7823);
and (n7878,n580,n156);
and (n7879,n7880,n7881);
xor (n7880,n7877,n7878);
or (n7881,n7882,n7885);
and (n7882,n7883,n7884);
xor (n7883,n7828,n7829);
and (n7884,n574,n156);
and (n7885,n7886,n7887);
xor (n7886,n7883,n7884);
or (n7887,n7888,n7891);
and (n7888,n7889,n7890);
xor (n7889,n7834,n7835);
and (n7890,n712,n156);
and (n7891,n7892,n7893);
xor (n7892,n7889,n7890);
or (n7893,n7894,n7897);
and (n7894,n7895,n7896);
xor (n7895,n7840,n7841);
and (n7896,n753,n156);
and (n7897,n7898,n7899);
xor (n7898,n7895,n7896);
or (n7899,n7900,n7903);
and (n7900,n7901,n7902);
xor (n7901,n7846,n7847);
and (n7902,n922,n156);
and (n7903,n7904,n7905);
xor (n7904,n7901,n7902);
or (n7905,n7906,n7909);
and (n7906,n7907,n7908);
xor (n7907,n7852,n7853);
and (n7908,n959,n156);
and (n7909,n7910,n7911);
xor (n7910,n7907,n7908);
and (n7911,n7912,n1560);
xor (n7912,n7858,n7859);
and (n7913,n166,n162);
or (n7914,n7915,n7918);
and (n7915,n7916,n7917);
xor (n7916,n7868,n7869);
and (n7917,n312,n162);
and (n7918,n7919,n7920);
xor (n7919,n7916,n7917);
or (n7920,n7921,n7924);
and (n7921,n7922,n7923);
xor (n7922,n7874,n7875);
and (n7923,n580,n162);
and (n7924,n7925,n7926);
xor (n7925,n7922,n7923);
or (n7926,n7927,n7930);
and (n7927,n7928,n7929);
xor (n7928,n7880,n7881);
and (n7929,n574,n162);
and (n7930,n7931,n7932);
xor (n7931,n7928,n7929);
or (n7932,n7933,n7936);
and (n7933,n7934,n7935);
xor (n7934,n7886,n7887);
and (n7935,n712,n162);
and (n7936,n7937,n7938);
xor (n7937,n7934,n7935);
or (n7938,n7939,n7942);
and (n7939,n7940,n7941);
xor (n7940,n7892,n7893);
and (n7941,n753,n162);
and (n7942,n7943,n7944);
xor (n7943,n7940,n7941);
or (n7944,n7945,n7948);
and (n7945,n7946,n7947);
xor (n7946,n7898,n7899);
and (n7947,n922,n162);
and (n7948,n7949,n7950);
xor (n7949,n7946,n7947);
or (n7950,n7951,n7954);
and (n7951,n7952,n7953);
xor (n7952,n7904,n7905);
and (n7953,n959,n162);
and (n7954,n7955,n7956);
xor (n7955,n7952,n7953);
and (n7956,n7957,n7958);
xor (n7957,n7910,n7911);
and (n7958,n1122,n162);
and (n7959,n312,n565);
or (n7960,n7961,n7964);
and (n7961,n7962,n7963);
xor (n7962,n7919,n7920);
and (n7963,n580,n565);
and (n7964,n7965,n7966);
xor (n7965,n7962,n7963);
or (n7966,n7967,n7970);
and (n7967,n7968,n7969);
xor (n7968,n7925,n7926);
and (n7969,n574,n565);
and (n7970,n7971,n7972);
xor (n7971,n7968,n7969);
or (n7972,n7973,n7976);
and (n7973,n7974,n7975);
xor (n7974,n7931,n7932);
and (n7975,n712,n565);
and (n7976,n7977,n7978);
xor (n7977,n7974,n7975);
or (n7978,n7979,n7982);
and (n7979,n7980,n7981);
xor (n7980,n7937,n7938);
and (n7981,n753,n565);
and (n7982,n7983,n7984);
xor (n7983,n7980,n7981);
or (n7984,n7985,n7988);
and (n7985,n7986,n7987);
xor (n7986,n7943,n7944);
and (n7987,n922,n565);
and (n7988,n7989,n7990);
xor (n7989,n7986,n7987);
or (n7990,n7991,n7994);
and (n7991,n7992,n7993);
xor (n7992,n7949,n7950);
and (n7993,n959,n565);
and (n7994,n7995,n7996);
xor (n7995,n7992,n7993);
and (n7996,n7997,n1121);
xor (n7997,n7955,n7956);
and (n7998,n580,n570);
or (n7999,n8000,n8003);
and (n8000,n8001,n8002);
xor (n8001,n7965,n7966);
and (n8002,n574,n570);
and (n8003,n8004,n8005);
xor (n8004,n8001,n8002);
or (n8005,n8006,n8009);
and (n8006,n8007,n8008);
xor (n8007,n7971,n7972);
and (n8008,n712,n570);
and (n8009,n8010,n8011);
xor (n8010,n8007,n8008);
or (n8011,n8012,n8015);
and (n8012,n8013,n8014);
xor (n8013,n7977,n7978);
and (n8014,n753,n570);
and (n8015,n8016,n8017);
xor (n8016,n8013,n8014);
or (n8017,n8018,n8021);
and (n8018,n8019,n8020);
xor (n8019,n7983,n7984);
and (n8020,n922,n570);
and (n8021,n8022,n8023);
xor (n8022,n8019,n8020);
or (n8023,n8024,n8027);
and (n8024,n8025,n8026);
xor (n8025,n7989,n7990);
and (n8026,n959,n570);
and (n8027,n8028,n8029);
xor (n8028,n8025,n8026);
and (n8029,n8030,n8031);
xor (n8030,n7995,n7996);
and (n8031,n1122,n570);
or (n8032,n8033,n8035);
and (n8033,n8034,n8008);
xor (n8034,n8004,n8005);
and (n8035,n8036,n8037);
xor (n8036,n8034,n8008);
or (n8037,n8038,n8040);
and (n8038,n8039,n8014);
xor (n8039,n8010,n8011);
and (n8040,n8041,n8042);
xor (n8041,n8039,n8014);
or (n8042,n8043,n8045);
and (n8043,n8044,n8020);
xor (n8044,n8016,n8017);
and (n8045,n8046,n8047);
xor (n8046,n8044,n8020);
or (n8047,n8048,n8050);
and (n8048,n8049,n8026);
xor (n8049,n8022,n8023);
and (n8050,n8051,n8052);
xor (n8051,n8049,n8026);
and (n8052,n8053,n8031);
xor (n8053,n8028,n8029);
or (n8054,n8055,n8057);
and (n8055,n8056,n8014);
xor (n8056,n8036,n8037);
and (n8057,n8058,n8059);
xor (n8058,n8056,n8014);
or (n8059,n8060,n8062);
and (n8060,n8061,n8020);
xor (n8061,n8041,n8042);
and (n8062,n8063,n8064);
xor (n8063,n8061,n8020);
or (n8064,n8065,n8067);
and (n8065,n8066,n8026);
xor (n8066,n8046,n8047);
and (n8067,n8068,n8069);
xor (n8068,n8066,n8026);
and (n8069,n8070,n8031);
xor (n8070,n8051,n8052);
or (n8071,n8072,n8074);
and (n8072,n8073,n8020);
xor (n8073,n8058,n8059);
and (n8074,n8075,n8076);
xor (n8075,n8073,n8020);
or (n8076,n8077,n8079);
and (n8077,n8078,n8026);
xor (n8078,n8063,n8064);
and (n8079,n8080,n8081);
xor (n8080,n8078,n8026);
and (n8081,n8082,n8031);
xor (n8082,n8068,n8069);
or (n8083,n8084,n8086);
and (n8084,n8085,n8026);
xor (n8085,n8075,n8076);
and (n8086,n8087,n8088);
xor (n8087,n8085,n8026);
and (n8088,n8089,n8031);
xor (n8089,n8080,n8081);
and (n8090,n8091,n8031);
xor (n8091,n8087,n8088);
endmodule
