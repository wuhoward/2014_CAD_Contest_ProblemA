module top (out,n13,n15,n16,n20,n25,n27,n30,n35,n37
        ,n39,n42,n49,n51,n53,n56,n61,n63,n65,n68
        ,n84,n86,n89,n144,n176,n252,n266,n267,n339,n348
        ,n349,n385,n457,n487,n488,n678,n682,n684,n710,n711
        ,n818,n835,n836,n1022,n1026,n1028,n1039,n1051,n1065);
output out;
input n13;
input n15;
input n16;
input n20;
input n25;
input n27;
input n30;
input n35;
input n37;
input n39;
input n42;
input n49;
input n51;
input n53;
input n56;
input n61;
input n63;
input n65;
input n68;
input n84;
input n86;
input n89;
input n144;
input n176;
input n252;
input n266;
input n267;
input n339;
input n348;
input n349;
input n385;
input n457;
input n487;
input n488;
input n678;
input n682;
input n684;
input n710;
input n711;
input n818;
input n835;
input n836;
input n1022;
input n1026;
input n1028;
input n1039;
input n1051;
input n1065;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n17;
wire n18;
wire n19;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n38;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n64;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n679;
wire n680;
wire n681;
wire n683;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1023;
wire n1024;
wire n1025;
wire n1027;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
xor (out,n0,n3003);
xnor (n0,n1,n2963);
nand (n1,n2,n227);
nand (n2,n3,n187);
nand (n3,n4,n133,n186);
nand (n4,n5,n91);
nand (n5,n6,n70,n90);
nand (n6,n7,n44);
nand (n7,n8,n31,n43);
nand (n8,n9,n21);
not (n9,n10);
xor (n10,n11,n20);
or (n11,n12,n17);
and (n12,n13,n14);
xor (n14,n15,n16);
and (n17,n13,n18);
nor (n18,n14,n19);
xnor (n19,n20,n15);
xor (n21,n22,n30);
or (n22,n23,n26);
and (n23,n13,n24);
xor (n24,n25,n20);
and (n26,n27,n28);
nor (n28,n24,n29);
xnor (n29,n30,n25);
nand (n31,n32,n21);
xor (n32,n33,n42);
or (n33,n34,n38);
and (n34,n35,n36);
xor (n36,n37,n30);
and (n38,n39,n40);
nor (n40,n36,n41);
xnor (n41,n42,n37);
nand (n43,n9,n32);
nand (n44,n45,n57,n69);
nand (n45,n46,n10);
xor (n46,n47,n56);
or (n47,n48,n52);
and (n48,n49,n50);
xor (n50,n51,n42);
and (n52,n53,n54);
nor (n54,n50,n55);
xnor (n55,n56,n51);
nand (n57,n58,n10);
xor (n58,n59,n68);
or (n59,n60,n64);
and (n60,n61,n62);
xor (n62,n63,n56);
and (n64,n65,n66);
nor (n66,n62,n67);
xnor (n67,n68,n63);
nand (n69,n46,n58);
nand (n70,n71,n44);
xor (n71,n72,n80);
xor (n72,n73,n76);
xor (n73,n74,n30);
or (n74,n23,n75);
and (n75,n13,n28);
xor (n76,n77,n68);
or (n77,n78,n79);
and (n78,n53,n62);
and (n79,n61,n66);
xor (n80,n81,n89);
or (n81,n82,n85);
and (n82,n65,n83);
xor (n83,n84,n68);
and (n85,n86,n87);
nor (n87,n83,n88);
xnor (n88,n89,n84);
nand (n90,n7,n71);
xor (n91,n92,n116);
xor (n92,n93,n106);
nand (n93,n94,n104,n105);
nand (n94,n95,n99);
xor (n95,n96,n56);
or (n96,n97,n98);
and (n97,n39,n50);
and (n98,n49,n54);
not (n99,n100);
xor (n100,n101,n42);
or (n101,n102,n103);
and (n102,n27,n36);
and (n103,n35,n40);
nand (n104,n89,n99);
nand (n105,n95,n89);
xor (n106,n107,n89);
xor (n107,n108,n112);
xor (n108,n109,n89);
or (n109,n110,n111);
and (n110,n61,n83);
and (n111,n65,n87);
xor (n112,n113,n56);
or (n113,n114,n115);
and (n114,n35,n50);
and (n115,n39,n54);
xor (n116,n117,n122);
xor (n117,n100,n118);
nand (n118,n119,n120,n121);
nand (n119,n73,n76);
nand (n120,n80,n76);
nand (n121,n73,n80);
xor (n122,n123,n129);
xor (n123,n124,n125);
not (n124,n73);
xor (n125,n126,n42);
or (n126,n127,n128);
and (n127,n13,n36);
and (n128,n27,n40);
xor (n129,n130,n68);
or (n130,n131,n132);
and (n131,n49,n62);
and (n132,n53,n66);
nand (n133,n134,n91);
nand (n134,n135,n163,n185);
nand (n135,n136,n138);
xor (n136,n137,n89);
xor (n137,n95,n99);
nand (n138,n139,n145,n162);
nand (n139,n140,n89);
xor (n140,n141,n89);
or (n141,n142,n143);
and (n142,n86,n83);
and (n143,n144,n87);
nand (n145,n146,n89);
nand (n146,n147,n156,n161);
nand (n147,n148,n152);
xor (n148,n149,n30);
or (n149,n150,n151);
and (n150,n27,n24);
and (n151,n35,n28);
xor (n152,n153,n42);
or (n153,n154,n155);
and (n154,n39,n36);
and (n155,n49,n40);
nand (n156,n157,n152);
xor (n157,n158,n56);
or (n158,n159,n160);
and (n159,n53,n50);
and (n160,n61,n54);
nand (n161,n148,n157);
nand (n162,n140,n146);
nand (n163,n164,n138);
nand (n164,n165,n181,n184);
nand (n165,n166,n179);
nand (n166,n167,n177,n178);
nand (n167,n168,n172);
xor (n168,n169,n68);
or (n169,n170,n171);
and (n170,n65,n62);
and (n171,n86,n66);
xor (n172,n173,n89);
or (n173,n174,n175);
and (n174,n144,n83);
and (n175,n176,n87);
nand (n177,n9,n172);
nand (n178,n168,n9);
xor (n179,n180,n32);
xor (n180,n9,n21);
nand (n181,n182,n179);
xor (n182,n183,n58);
xor (n183,n46,n10);
nand (n184,n166,n182);
nand (n185,n136,n164);
nand (n186,n5,n134);
xor (n187,n188,n223);
xor (n188,n189,n193);
nand (n189,n190,n191,n192);
nand (n190,n100,n118);
nand (n191,n122,n118);
nand (n192,n100,n122);
xor (n193,n194,n213);
xor (n194,n195,n209);
xor (n195,n196,n205);
xor (n196,n197,n201);
xor (n197,n198,n56);
or (n198,n199,n200);
and (n199,n27,n50);
and (n200,n35,n54);
xor (n201,n202,n89);
or (n202,n203,n204);
and (n203,n53,n83);
and (n204,n61,n87);
xor (n205,n206,n68);
or (n206,n207,n208);
and (n207,n39,n62);
and (n208,n49,n66);
nand (n209,n210,n211,n212);
nand (n210,n108,n112);
nand (n211,n89,n112);
nand (n212,n108,n89);
xor (n213,n214,n219);
xor (n214,n215,n89);
not (n215,n216);
xor (n216,n217,n42);
or (n217,n127,n218);
and (n218,n13,n40);
nand (n219,n220,n221,n222);
nand (n220,n124,n125);
nand (n221,n129,n125);
nand (n222,n124,n129);
nand (n223,n224,n225,n226);
nand (n224,n93,n106);
nand (n225,n116,n106);
nand (n226,n93,n116);
nand (n227,n228,n2961);
nand (n228,n229,n999);
nor (n229,n230,n984);
nor (n230,n231,n577);
nand (n231,n232,n554);
nor (n232,n233,n530);
nor (n233,n234,n407);
xor (n234,n235,n364);
xor (n235,n236,n255);
xor (n236,n237,n242);
xor (n237,n238,n240);
xor (n238,n239,n157);
xor (n239,n148,n152);
xor (n240,n241,n9);
xor (n241,n168,n172);
nand (n242,n243,n253,n254);
nand (n243,n244,n248);
xor (n244,n245,n68);
or (n245,n246,n247);
and (n246,n86,n62);
and (n247,n144,n66);
xor (n248,n249,n89);
or (n249,n250,n251);
and (n250,n176,n83);
and (n251,n252,n87);
nand (n253,n89,n248);
nand (n254,n244,n89);
xor (n255,n256,n326);
xor (n256,n257,n292);
xor (n257,n258,n280);
xor (n258,n89,n259);
nand (n259,n260,n274,n279);
nand (n260,n261,n271);
not (n261,n262);
xor (n262,n263,n16);
or (n263,n264,n268);
and (n264,n13,n265);
xor (n265,n266,n267);
and (n268,n13,n269);
nor (n269,n265,n270);
xnor (n270,n16,n266);
xor (n271,n272,n20);
or (n272,n12,n273);
and (n273,n27,n18);
nand (n274,n275,n271);
xor (n275,n276,n42);
or (n276,n277,n278);
and (n277,n49,n36);
and (n278,n53,n40);
nand (n279,n261,n275);
nand (n280,n281,n286,n291);
nand (n281,n282,n262);
xor (n282,n283,n30);
or (n283,n284,n285);
and (n284,n35,n24);
and (n285,n39,n28);
nand (n286,n287,n262);
xor (n287,n288,n56);
or (n288,n289,n290);
and (n289,n61,n50);
and (n290,n65,n54);
nand (n291,n282,n287);
nand (n292,n293,n312,n325);
nand (n293,n294,n296);
xor (n294,n295,n275);
xor (n295,n261,n271);
nand (n296,n297,n306,n311);
nand (n297,n298,n302);
xor (n298,n299,n20);
or (n299,n300,n301);
and (n300,n27,n14);
and (n301,n35,n18);
xor (n302,n303,n42);
or (n303,n304,n305);
and (n304,n53,n36);
and (n305,n61,n40);
nand (n306,n307,n302);
xor (n307,n308,n30);
or (n308,n309,n310);
and (n309,n39,n24);
and (n310,n49,n28);
nand (n311,n298,n307);
nand (n312,n313,n296);
nand (n313,n314,n319,n324);
nand (n314,n261,n315);
xor (n315,n316,n56);
or (n316,n317,n318);
and (n317,n65,n50);
and (n318,n86,n54);
nand (n319,n320,n315);
xor (n320,n321,n68);
or (n321,n322,n323);
and (n322,n144,n62);
and (n323,n176,n66);
nand (n324,n261,n320);
nand (n325,n294,n313);
nand (n326,n327,n332,n363);
nand (n327,n328,n330);
xor (n328,n329,n89);
xor (n329,n244,n248);
xor (n330,n331,n287);
xor (n331,n282,n262);
nand (n332,n333,n330);
nand (n333,n334,n340,n362);
nand (n334,n335,n89);
xor (n335,n336,n89);
or (n336,n337,n338);
and (n337,n252,n83);
and (n338,n339,n87);
nand (n340,n341,n89);
nand (n341,n342,n356,n361);
nand (n342,n343,n353);
not (n343,n344);
xor (n344,n345,n267);
or (n345,n346,n350);
and (n346,n13,n347);
xor (n347,n348,n349);
and (n350,n13,n351);
nor (n351,n347,n352);
xnor (n352,n267,n348);
xor (n353,n354,n16);
or (n354,n264,n355);
and (n355,n27,n269);
nand (n356,n357,n353);
xor (n357,n358,n20);
or (n358,n359,n360);
and (n359,n35,n14);
and (n360,n39,n18);
nand (n361,n343,n357);
nand (n362,n335,n341);
nand (n363,n328,n333);
nand (n364,n365,n403,n406);
nand (n365,n366,n401);
nand (n366,n367,n387,n400);
nand (n367,n368,n370);
xor (n368,n369,n307);
xor (n369,n298,n302);
nand (n370,n371,n380,n386);
nand (n371,n372,n376);
xor (n372,n373,n30);
or (n373,n374,n375);
and (n374,n49,n24);
and (n375,n53,n28);
xor (n376,n377,n42);
or (n377,n378,n379);
and (n378,n61,n36);
and (n379,n65,n40);
nand (n380,n381,n376);
xor (n381,n382,n89);
or (n382,n383,n384);
and (n383,n339,n83);
and (n384,n385,n87);
nand (n386,n372,n381);
nand (n387,n388,n370);
nand (n388,n389,n394,n399);
nand (n389,n344,n390);
xor (n390,n391,n56);
or (n391,n392,n393);
and (n392,n86,n50);
and (n393,n144,n54);
nand (n394,n395,n390);
xor (n395,n396,n68);
or (n396,n397,n398);
and (n397,n176,n62);
and (n398,n252,n66);
nand (n399,n344,n395);
nand (n400,n368,n388);
xor (n401,n402,n313);
xor (n402,n294,n296);
nand (n403,n404,n401);
xor (n404,n405,n333);
xor (n405,n328,n330);
nand (n406,n366,n404);
nand (n407,n408,n440,n529);
nand (n408,n409,n438);
nand (n409,n410,n414,n437);
nand (n410,n411,n413);
xor (n411,n412,n320);
xor (n412,n261,n315);
xor (n413,n336,n341);
nand (n414,n415,n413);
nand (n415,n416,n419,n436);
nand (n416,n89,n417);
xor (n417,n418,n357);
xor (n418,n343,n353);
nand (n419,n420,n417);
nand (n420,n421,n430,n435);
nand (n421,n422,n426);
xor (n422,n423,n16);
or (n423,n424,n425);
and (n424,n27,n265);
and (n425,n35,n269);
xor (n426,n427,n20);
or (n427,n428,n429);
and (n428,n39,n14);
and (n429,n49,n18);
nand (n430,n431,n426);
xor (n431,n432,n30);
or (n432,n433,n434);
and (n433,n53,n24);
and (n434,n61,n28);
nand (n435,n422,n431);
nand (n436,n89,n420);
nand (n437,n411,n415);
xor (n438,n439,n404);
xor (n439,n366,n401);
nand (n440,n441,n438);
nand (n441,n442,n466,n528);
nand (n442,n443,n445);
xor (n443,n444,n388);
xor (n444,n368,n370);
nand (n445,n446,n462,n465);
nand (n446,n447,n460);
nand (n447,n448,n458,n459);
nand (n448,n449,n453);
xor (n449,n450,n42);
or (n450,n451,n452);
and (n451,n65,n36);
and (n452,n86,n40);
xor (n453,n454,n89);
or (n454,n455,n456);
and (n455,n385,n83);
and (n456,n457,n87);
nand (n458,n343,n453);
nand (n459,n449,n343);
xor (n460,n461,n381);
xor (n461,n372,n376);
nand (n462,n463,n460);
xor (n463,n464,n395);
xor (n464,n344,n390);
nand (n465,n447,n463);
nand (n466,n467,n445);
nand (n467,n468,n524,n527);
nand (n468,n469,n502);
nand (n469,n470,n479,n501);
nand (n470,n471,n475);
xor (n471,n472,n56);
or (n472,n473,n474);
and (n473,n144,n50);
and (n474,n176,n54);
xor (n475,n476,n68);
or (n476,n477,n478);
and (n477,n252,n62);
and (n478,n339,n66);
nand (n479,n480,n475);
nand (n480,n481,n495,n500);
nand (n481,n482,n492);
not (n482,n483);
xor (n483,n484,n349);
or (n484,n485,n489);
and (n485,n13,n486);
xor (n486,n487,n488);
and (n489,n13,n490);
nor (n490,n486,n491);
xnor (n491,n349,n487);
xor (n492,n493,n267);
or (n493,n346,n494);
and (n494,n27,n351);
nand (n495,n496,n492);
xor (n496,n497,n20);
or (n497,n498,n499);
and (n498,n49,n14);
and (n499,n53,n18);
nand (n500,n482,n496);
nand (n501,n471,n480);
nand (n502,n503,n506,n523);
nand (n503,n89,n504);
xor (n504,n505,n431);
xor (n505,n422,n426);
nand (n506,n507,n504);
nand (n507,n508,n517,n522);
nand (n508,n509,n513);
xor (n509,n510,n16);
or (n510,n511,n512);
and (n511,n35,n265);
and (n512,n39,n269);
xor (n513,n514,n30);
or (n514,n515,n516);
and (n515,n61,n24);
and (n516,n65,n28);
nand (n517,n518,n513);
xor (n518,n519,n42);
or (n519,n520,n521);
and (n520,n86,n36);
and (n521,n144,n40);
nand (n522,n509,n518);
nand (n523,n89,n507);
nand (n524,n525,n502);
xor (n525,n526,n420);
xor (n526,n89,n417);
nand (n527,n469,n525);
nand (n528,n443,n467);
nand (n529,n409,n441);
nor (n530,n531,n535);
nand (n531,n532,n533,n534);
nand (n532,n236,n255);
nand (n533,n364,n255);
nand (n534,n236,n364);
xor (n535,n536,n550);
xor (n536,n537,n541);
nand (n537,n538,n539,n540);
nand (n538,n238,n240);
nand (n539,n242,n240);
nand (n540,n238,n242);
xor (n541,n542,n548);
xor (n542,n543,n547);
nand (n543,n544,n545,n546);
nand (n544,n89,n259);
nand (n545,n280,n259);
nand (n546,n89,n280);
xor (n547,n141,n146);
xor (n548,n549,n182);
xor (n549,n166,n179);
nand (n550,n551,n552,n553);
nand (n551,n257,n292);
nand (n552,n326,n292);
nand (n553,n257,n326);
nor (n554,n555,n570);
nor (n555,n556,n560);
nand (n556,n557,n558,n559);
nand (n557,n537,n541);
nand (n558,n550,n541);
nand (n559,n537,n550);
xor (n560,n561,n566);
xor (n561,n562,n564);
xor (n562,n563,n71);
xor (n563,n7,n44);
xor (n564,n565,n164);
xor (n565,n136,n138);
nand (n566,n567,n568,n569);
nand (n567,n543,n547);
nand (n568,n548,n547);
nand (n569,n543,n548);
nor (n570,n571,n575);
nand (n571,n572,n573,n574);
nand (n572,n562,n564);
nand (n573,n566,n564);
nand (n574,n562,n566);
xor (n575,n576,n134);
xor (n576,n5,n91);
nor (n577,n578,n978);
nor (n578,n579,n954);
nor (n579,n580,n952);
nor (n580,n581,n927);
nand (n581,n582,n889);
nand (n582,n583,n805,n888);
nand (n583,n584,n668);
xor (n584,n585,n658);
xor (n585,n586,n608);
xor (n586,n587,n592);
xor (n587,n588,n89);
xor (n588,n589,n56);
or (n589,n590,n591);
and (n590,n176,n50);
and (n591,n252,n54);
nand (n592,n593,n602,n607);
nand (n593,n594,n598);
xor (n594,n595,n20);
or (n595,n596,n597);
and (n596,n53,n14);
and (n597,n61,n18);
xor (n598,n599,n267);
or (n599,n600,n601);
and (n600,n27,n347);
and (n601,n35,n351);
nand (n602,n603,n598);
xor (n603,n604,n16);
or (n604,n605,n606);
and (n605,n39,n265);
and (n606,n49,n269);
nand (n607,n594,n603);
nand (n608,n609,n640,n657);
nand (n609,n610,n626);
nand (n610,n611,n620,n625);
nand (n611,n612,n616);
xor (n612,n613,n20);
or (n613,n614,n615);
and (n614,n61,n14);
and (n615,n65,n18);
xor (n616,n617,n267);
or (n617,n618,n619);
and (n618,n35,n347);
and (n619,n39,n351);
nand (n620,n621,n616);
xor (n621,n622,n30);
or (n622,n623,n624);
and (n623,n86,n24);
and (n624,n144,n28);
nand (n625,n612,n621);
xor (n626,n627,n636);
xor (n627,n628,n632);
xor (n628,n629,n30);
or (n629,n630,n631);
and (n630,n65,n24);
and (n631,n86,n28);
xor (n632,n633,n42);
or (n633,n634,n635);
and (n634,n144,n36);
and (n635,n176,n40);
xor (n636,n637,n68);
or (n637,n638,n639);
and (n638,n385,n62);
and (n639,n457,n66);
nand (n640,n641,n626);
nand (n641,n642,n651,n656);
nand (n642,n643,n647);
xor (n643,n644,n349);
or (n644,n645,n646);
and (n645,n27,n486);
and (n646,n35,n490);
xor (n647,n648,n42);
or (n648,n649,n650);
and (n649,n176,n36);
and (n650,n252,n40);
nand (n651,n652,n647);
xor (n652,n653,n56);
or (n653,n654,n655);
and (n654,n339,n50);
and (n655,n385,n54);
nand (n656,n643,n652);
nand (n657,n610,n641);
xor (n658,n659,n664);
xor (n659,n660,n662);
xor (n660,n661,n496);
xor (n661,n482,n492);
xor (n662,n663,n518);
xor (n663,n509,n513);
nand (n664,n665,n666,n667);
nand (n665,n628,n632);
nand (n666,n636,n632);
nand (n667,n628,n636);
xor (n668,n669,n744);
xor (n669,n670,n724);
nand (n670,n671,n697,n723);
nand (n671,n672,n687);
nand (n672,n673,n685,n686);
nand (n673,n674,n679);
xor (n674,n675,n68);
or (n675,n676,n677);
and (n676,n457,n62);
and (n677,n678,n66);
xor (n679,n680,n89);
or (n680,n681,n683);
and (n681,n682,n83);
and (n683,n684,n87);
nand (n685,n89,n679);
nand (n686,n674,n89);
xor (n687,n688,n693);
xor (n688,n689,n482);
xor (n689,n690,n89);
or (n690,n691,n692);
and (n691,n678,n83);
and (n692,n682,n87);
xor (n693,n694,n56);
or (n694,n695,n696);
and (n695,n252,n50);
and (n696,n339,n54);
nand (n697,n698,n687);
xor (n698,n699,n721);
xor (n699,n89,n700);
nand (n700,n701,n715,n720);
nand (n701,n702,n705);
xor (n702,n703,n349);
or (n703,n485,n704);
and (n704,n27,n490);
not (n705,n706);
xor (n706,n707,n488);
or (n707,n708,n712);
and (n708,n13,n709);
xor (n709,n710,n711);
and (n712,n13,n713);
nor (n713,n709,n714);
xnor (n714,n488,n710);
nand (n715,n716,n705);
xor (n716,n717,n16);
or (n717,n718,n719);
and (n718,n49,n265);
and (n719,n53,n269);
nand (n720,n702,n716);
xor (n721,n722,n603);
xor (n722,n594,n598);
nand (n723,n672,n698);
xor (n724,n725,n740);
xor (n725,n726,n730);
nand (n726,n727,n728,n729);
nand (n727,n689,n482);
nand (n728,n693,n482);
nand (n729,n689,n693);
xor (n730,n731,n483);
xor (n731,n732,n736);
xor (n732,n733,n68);
or (n733,n734,n735);
and (n734,n339,n62);
and (n735,n385,n66);
xor (n736,n737,n89);
or (n737,n738,n739);
and (n738,n457,n83);
and (n739,n678,n87);
nand (n740,n741,n742,n743);
nand (n741,n89,n700);
nand (n742,n721,n700);
nand (n743,n89,n721);
nand (n744,n745,n801,n804);
nand (n745,n746,n766);
nand (n746,n747,n762,n765);
nand (n747,n748,n760);
nand (n748,n749,n754,n759);
nand (n749,n706,n750);
xor (n750,n751,n16);
or (n751,n752,n753);
and (n752,n53,n265);
and (n753,n61,n269);
nand (n754,n755,n750);
xor (n755,n756,n20);
or (n756,n757,n758);
and (n757,n65,n14);
and (n758,n86,n18);
nand (n759,n706,n755);
xor (n760,n761,n621);
xor (n761,n612,n616);
nand (n762,n763,n760);
xor (n763,n764,n716);
xor (n764,n702,n705);
nand (n765,n748,n763);
nand (n766,n767,n797,n800);
nand (n767,n768,n781);
nand (n768,n769,n775,n780);
nand (n769,n770,n774);
xor (n770,n771,n267);
or (n771,n772,n773);
and (n772,n39,n347);
and (n773,n49,n351);
not (n774,n643);
nand (n775,n776,n774);
xor (n776,n777,n30);
or (n777,n778,n779);
and (n778,n144,n24);
and (n779,n176,n28);
nand (n780,n770,n776);
nand (n781,n782,n791,n796);
nand (n782,n783,n787);
xor (n783,n784,n42);
or (n784,n785,n786);
and (n785,n252,n36);
and (n786,n339,n40);
xor (n787,n788,n56);
or (n788,n789,n790);
and (n789,n385,n50);
and (n790,n457,n54);
nand (n791,n792,n787);
xor (n792,n793,n68);
or (n793,n794,n795);
and (n794,n678,n62);
and (n795,n682,n66);
nand (n796,n783,n792);
nand (n797,n798,n781);
xor (n798,n799,n652);
xor (n799,n643,n647);
nand (n800,n768,n798);
nand (n801,n802,n766);
xor (n802,n803,n641);
xor (n803,n610,n626);
nand (n804,n746,n802);
nand (n805,n806,n668);
nand (n806,n807,n884,n887);
nand (n807,n808,n810);
xor (n808,n809,n698);
xor (n809,n672,n687);
nand (n810,n811,n844,n883);
nand (n811,n812,n842);
nand (n812,n813,n819,n841);
nand (n813,n814,n89);
xor (n814,n815,n89);
or (n815,n816,n817);
and (n816,n684,n83);
and (n817,n818,n87);
nand (n819,n820,n89);
nand (n820,n821,n829,n840);
nand (n821,n822,n825);
xor (n822,n823,n488);
or (n823,n708,n824);
and (n824,n27,n713);
xor (n825,n826,n349);
or (n826,n827,n828);
and (n827,n35,n486);
and (n828,n39,n490);
nand (n829,n830,n825);
not (n830,n831);
xor (n831,n832,n711);
or (n832,n833,n837);
and (n833,n13,n834);
xor (n834,n835,n836);
and (n837,n13,n838);
nor (n838,n834,n839);
xnor (n839,n711,n835);
nand (n840,n822,n830);
nand (n841,n814,n820);
xor (n842,n843,n89);
xor (n843,n674,n679);
nand (n844,n845,n842);
nand (n845,n846,n865,n882);
nand (n846,n847,n863);
nand (n847,n848,n857,n862);
nand (n848,n849,n853);
xor (n849,n850,n267);
or (n850,n851,n852);
and (n851,n49,n347);
and (n852,n53,n351);
xor (n853,n854,n16);
or (n854,n855,n856);
and (n855,n61,n265);
and (n856,n65,n269);
nand (n857,n858,n853);
xor (n858,n859,n20);
or (n859,n860,n861);
and (n860,n86,n14);
and (n861,n144,n18);
nand (n862,n849,n858);
xor (n863,n864,n755);
xor (n864,n706,n750);
nand (n865,n866,n863);
nand (n866,n867,n876,n881);
nand (n867,n868,n872);
xor (n868,n869,n42);
or (n869,n870,n871);
and (n870,n339,n36);
and (n871,n385,n40);
xor (n872,n873,n488);
or (n873,n874,n875);
and (n874,n27,n709);
and (n875,n35,n713);
nand (n876,n877,n872);
xor (n877,n878,n30);
or (n878,n879,n880);
and (n879,n176,n24);
and (n880,n252,n28);
nand (n881,n868,n877);
nand (n882,n847,n866);
nand (n883,n812,n845);
nand (n884,n885,n810);
xor (n885,n886,n802);
xor (n886,n746,n766);
nand (n887,n808,n885);
nand (n888,n584,n806);
xor (n889,n890,n923);
xor (n890,n891,n895);
nand (n891,n892,n893,n894);
nand (n892,n586,n608);
nand (n893,n658,n608);
nand (n894,n586,n658);
xor (n895,n896,n911);
xor (n896,n897,n901);
nand (n897,n898,n899,n900);
nand (n898,n726,n730);
nand (n899,n740,n730);
nand (n900,n726,n740);
xor (n901,n902,n909);
xor (n902,n903,n907);
nand (n903,n904,n905,n906);
nand (n904,n732,n736);
nand (n905,n483,n736);
nand (n906,n732,n483);
xor (n907,n908,n480);
xor (n908,n471,n475);
xor (n909,n910,n343);
xor (n910,n449,n453);
xor (n911,n912,n919);
xor (n912,n913,n917);
nand (n913,n914,n915,n916);
nand (n914,n588,n89);
nand (n915,n592,n89);
nand (n916,n588,n592);
xor (n917,n918,n507);
xor (n918,n89,n504);
nand (n919,n920,n921,n922);
nand (n920,n660,n662);
nand (n921,n664,n662);
nand (n922,n660,n664);
nand (n923,n924,n925,n926);
nand (n924,n670,n724);
nand (n925,n744,n724);
nand (n926,n670,n744);
nor (n927,n928,n932);
nand (n928,n929,n930,n931);
nand (n929,n891,n895);
nand (n930,n923,n895);
nand (n931,n891,n923);
xor (n932,n933,n948);
xor (n933,n934,n936);
xor (n934,n935,n525);
xor (n935,n469,n502);
xor (n936,n937,n944);
xor (n937,n938,n940);
xor (n938,n939,n463);
xor (n939,n447,n460);
nand (n940,n941,n942,n943);
nand (n941,n903,n907);
nand (n942,n909,n907);
nand (n943,n903,n909);
nand (n944,n945,n946,n947);
nand (n945,n913,n917);
nand (n946,n919,n917);
nand (n947,n913,n919);
nand (n948,n949,n950,n951);
nand (n949,n897,n901);
nand (n950,n911,n901);
nand (n951,n897,n911);
not (n952,n953);
nand (n953,n928,n932);
not (n954,n955);
nor (n955,n956,n971);
nor (n956,n957,n961);
nand (n957,n958,n959,n960);
nand (n958,n934,n936);
nand (n959,n948,n936);
nand (n960,n934,n948);
xor (n961,n962,n967);
xor (n962,n963,n965);
xor (n963,n964,n415);
xor (n964,n411,n413);
xor (n965,n966,n467);
xor (n966,n443,n445);
nand (n967,n968,n969,n970);
nand (n968,n938,n940);
nand (n969,n944,n940);
nand (n970,n938,n944);
nor (n971,n972,n976);
nand (n972,n973,n974,n975);
nand (n973,n963,n965);
nand (n974,n967,n965);
nand (n975,n963,n967);
xor (n976,n977,n441);
xor (n977,n409,n438);
not (n978,n979);
nor (n979,n980,n982);
nor (n980,n981,n971);
nand (n981,n957,n961);
not (n982,n983);
nand (n983,n972,n976);
not (n984,n985);
nor (n985,n986,n993);
nor (n986,n987,n992);
nor (n987,n988,n990);
nor (n988,n989,n530);
nand (n989,n234,n407);
not (n990,n991);
nand (n991,n531,n535);
not (n992,n554);
not (n993,n994);
nor (n994,n995,n997);
nor (n995,n996,n570);
nand (n996,n556,n560);
not (n997,n998);
nand (n998,n571,n575);
nand (n999,n1000,n1004);
nor (n1000,n1001,n231);
nand (n1001,n1002,n955);
nor (n1002,n1003,n927);
nor (n1003,n582,n889);
nand (n1004,n1005,n2535);
nor (n1005,n1006,n2503);
nor (n1006,n1007,n1976);
nor (n1007,n1008,n1961);
nor (n1008,n1009,n1682);
nand (n1009,n1010,n1465);
nor (n1010,n1011,n1364);
nor (n1011,n1012,n1274);
nand (n1012,n1013,n1189,n1273);
nand (n1013,n1014,n1091);
xor (n1014,n1015,n1067);
xor (n1015,n1016,n1041);
xor (n1016,n1017,n1029);
xor (n1017,n1018,n1023);
xor (n1018,n1019,n30);
or (n1019,n1020,n1021);
and (n1020,n818,n24);
and (n1021,n1022,n28);
xor (n1023,n1024,n42);
or (n1024,n1025,n1027);
and (n1025,n1026,n36);
and (n1027,n1028,n40);
xor (n1029,n1030,n1034);
xor (n1030,n1031,n711);
or (n1031,n1032,n1033);
and (n1032,n61,n834);
and (n1033,n65,n838);
xnor (n1034,n1035,n836);
nor (n1035,n1036,n1040);
and (n1036,n53,n1037);
and (n1037,n1038,n836);
not (n1038,n1039);
and (n1040,n49,n1039);
nand (n1041,n1042,n1052,n1066);
nand (n1042,n1043,n1047);
xor (n1043,n1044,n30);
or (n1044,n1045,n1046);
and (n1045,n1022,n24);
and (n1046,n1026,n28);
xor (n1047,n1048,n42);
or (n1048,n1049,n1050);
and (n1049,n1028,n36);
and (n1050,n1051,n40);
nand (n1052,n1053,n1047);
xor (n1053,n1054,n1063);
xor (n1054,n1055,n1059);
xor (n1055,n1056,n711);
or (n1056,n1057,n1058);
and (n1057,n65,n834);
and (n1058,n86,n838);
xor (n1059,n1060,n349);
or (n1060,n1061,n1062);
and (n1061,n252,n486);
and (n1062,n339,n490);
xnor (n1063,n1064,n56);
nand (n1064,n1065,n50);
nand (n1066,n1043,n1053);
xor (n1067,n1068,n1077);
xor (n1068,n1069,n1073);
xor (n1069,n1070,n56);
or (n1070,n1071,n1072);
and (n1071,n1051,n50);
and (n1072,n1065,n54);
nand (n1073,n1074,n1075,n1076);
nand (n1074,n1055,n1059);
nand (n1075,n1063,n1059);
nand (n1076,n1055,n1063);
xor (n1077,n1078,n1087);
xor (n1078,n1079,n1083);
xor (n1079,n1080,n349);
or (n1080,n1081,n1082);
and (n1081,n176,n486);
and (n1082,n252,n490);
xor (n1083,n1084,n488);
or (n1084,n1085,n1086);
and (n1085,n86,n709);
and (n1086,n144,n713);
xor (n1087,n1088,n267);
or (n1088,n1089,n1090);
and (n1089,n339,n347);
and (n1090,n385,n351);
nand (n1091,n1092,n1146,n1188);
nand (n1092,n1093,n1095);
xor (n1093,n1094,n1053);
xor (n1094,n1043,n1047);
xor (n1095,n1096,n1135);
xor (n1096,n1097,n1113);
nand (n1097,n1098,n1107,n1112);
nand (n1098,n1099,n1103);
xor (n1099,n1100,n349);
or (n1100,n1101,n1102);
and (n1101,n339,n486);
and (n1102,n385,n490);
xor (n1103,n1104,n488);
or (n1104,n1105,n1106);
and (n1105,n176,n709);
and (n1106,n252,n713);
nand (n1107,n1108,n1103);
xor (n1108,n1109,n267);
or (n1109,n1110,n1111);
and (n1110,n457,n347);
and (n1111,n678,n351);
nand (n1112,n1099,n1108);
nand (n1113,n1114,n1129,n1134);
nand (n1114,n1115,n1124);
xor (n1115,n1116,n1120);
xnor (n1116,n1117,n836);
nor (n1117,n1118,n1119);
and (n1118,n65,n1037);
and (n1119,n61,n1039);
xor (n1120,n1121,n711);
or (n1121,n1122,n1123);
and (n1122,n86,n834);
and (n1123,n144,n838);
and (n1124,n1125,n42);
xnor (n1125,n1126,n836);
nor (n1126,n1127,n1128);
and (n1127,n86,n1037);
and (n1128,n65,n1039);
nand (n1129,n1130,n1124);
xor (n1130,n1131,n16);
or (n1131,n1132,n1133);
and (n1132,n682,n265);
and (n1133,n684,n269);
nand (n1134,n1115,n1130);
xor (n1135,n1136,n1142);
xor (n1136,n1137,n1141);
xor (n1137,n1138,n16);
or (n1138,n1139,n1140);
and (n1139,n678,n265);
and (n1140,n682,n269);
and (n1141,n1116,n1120);
xor (n1142,n1143,n20);
or (n1143,n1144,n1145);
and (n1144,n684,n14);
and (n1145,n818,n18);
nand (n1146,n1147,n1095);
nand (n1147,n1148,n1172,n1187);
nand (n1148,n1149,n1170);
nand (n1149,n1150,n1164,n1169);
nand (n1150,n1151,n1160);
and (n1151,n1152,n1156);
xnor (n1152,n1153,n836);
nor (n1153,n1154,n1155);
and (n1154,n144,n1037);
and (n1155,n86,n1039);
xor (n1156,n1157,n711);
or (n1157,n1158,n1159);
and (n1158,n176,n834);
and (n1159,n252,n838);
xor (n1160,n1161,n16);
or (n1161,n1162,n1163);
and (n1162,n684,n265);
and (n1163,n818,n269);
nand (n1164,n1165,n1160);
xor (n1165,n1166,n20);
or (n1166,n1167,n1168);
and (n1167,n1022,n14);
and (n1168,n1026,n18);
nand (n1169,n1151,n1165);
xor (n1170,n1171,n1130);
xor (n1171,n1115,n1124);
nand (n1172,n1173,n1170);
xor (n1173,n1174,n1183);
xor (n1174,n1175,n1179);
xor (n1175,n1176,n20);
or (n1176,n1177,n1178);
and (n1177,n818,n14);
and (n1178,n1022,n18);
xor (n1179,n1180,n30);
or (n1180,n1181,n1182);
and (n1181,n1026,n24);
and (n1182,n1028,n28);
xor (n1183,n1184,n42);
or (n1184,n1185,n1186);
and (n1185,n1051,n36);
and (n1186,n1065,n40);
nand (n1187,n1149,n1173);
nand (n1188,n1093,n1147);
nand (n1189,n1190,n1091);
xor (n1190,n1191,n1230);
xor (n1191,n1192,n1196);
nand (n1192,n1193,n1194,n1195);
nand (n1193,n1097,n1113);
nand (n1194,n1135,n1113);
nand (n1195,n1097,n1135);
xor (n1196,n1197,n1219);
xor (n1197,n1198,n1215);
nand (n1198,n1199,n1209,n1214);
nand (n1199,n1200,n1204);
xor (n1200,n1201,n488);
or (n1201,n1202,n1203);
and (n1202,n144,n709);
and (n1203,n176,n713);
xor (n1204,n1205,n56);
xnor (n1205,n1206,n836);
nor (n1206,n1207,n1208);
and (n1207,n61,n1037);
and (n1208,n53,n1039);
nand (n1209,n1210,n1204);
xor (n1210,n1211,n267);
or (n1211,n1212,n1213);
and (n1212,n385,n347);
and (n1213,n457,n351);
nand (n1214,n1200,n1210);
nand (n1215,n1216,n1217,n1218);
nand (n1216,n1137,n1141);
nand (n1217,n1142,n1141);
nand (n1218,n1137,n1142);
xor (n1219,n1220,n1226);
xor (n1220,n1221,n1222);
and (n1221,n1205,n56);
xor (n1222,n1223,n16);
or (n1223,n1224,n1225);
and (n1224,n457,n265);
and (n1225,n678,n269);
xor (n1226,n1227,n20);
or (n1227,n1228,n1229);
and (n1228,n682,n14);
and (n1229,n684,n18);
nand (n1230,n1231,n1238,n1272);
nand (n1231,n1232,n1236);
nand (n1232,n1233,n1234,n1235);
nand (n1233,n1175,n1179);
nand (n1234,n1183,n1179);
nand (n1235,n1175,n1183);
xor (n1236,n1237,n1210);
xor (n1237,n1200,n1204);
nand (n1238,n1239,n1236);
nand (n1239,n1240,n1257,n1271);
nand (n1240,n1241,n1255);
nand (n1241,n1242,n1251,n1254);
nand (n1242,n1243,n1247);
xor (n1243,n1244,n711);
or (n1244,n1245,n1246);
and (n1245,n144,n834);
and (n1246,n176,n838);
xor (n1247,n1248,n349);
or (n1248,n1249,n1250);
and (n1249,n385,n486);
and (n1250,n457,n490);
nand (n1251,n1252,n1247);
xnor (n1252,n1253,n42);
nand (n1253,n1065,n36);
nand (n1254,n1243,n1252);
xor (n1255,n1256,n1108);
xor (n1256,n1099,n1103);
nand (n1257,n1258,n1255);
nand (n1258,n1259,n1265,n1270);
nand (n1259,n1260,n1264);
xor (n1260,n1261,n488);
or (n1261,n1262,n1263);
and (n1262,n252,n709);
and (n1263,n339,n713);
xor (n1264,n1125,n42);
nand (n1265,n1266,n1264);
xor (n1266,n1267,n267);
or (n1267,n1268,n1269);
and (n1268,n678,n347);
and (n1269,n682,n351);
nand (n1270,n1260,n1266);
nand (n1271,n1241,n1258);
nand (n1272,n1232,n1239);
nand (n1273,n1014,n1190);
xor (n1274,n1275,n1360);
xor (n1275,n1276,n1297);
xor (n1276,n1277,n1293);
xor (n1277,n1278,n1289);
xor (n1278,n1279,n1285);
xor (n1279,n1280,n1284);
xor (n1280,n1281,n42);
or (n1281,n1282,n1283);
and (n1282,n1022,n36);
and (n1283,n1026,n40);
and (n1284,n1030,n1034);
xor (n1285,n1286,n56);
or (n1286,n1287,n1288);
and (n1287,n1028,n50);
and (n1288,n1051,n54);
nand (n1289,n1290,n1291,n1292);
nand (n1290,n1069,n1073);
nand (n1291,n1077,n1073);
nand (n1292,n1069,n1077);
nand (n1293,n1294,n1295,n1296);
nand (n1294,n1198,n1215);
nand (n1295,n1219,n1215);
nand (n1296,n1198,n1219);
xor (n1297,n1298,n1356);
xor (n1298,n1299,n1323);
xor (n1299,n1300,n1319);
xor (n1300,n1301,n1305);
nand (n1301,n1302,n1303,n1304);
nand (n1302,n1221,n1222);
nand (n1303,n1226,n1222);
nand (n1304,n1221,n1226);
xor (n1305,n1306,n1315);
xor (n1306,n1307,n1311);
xnor (n1307,n1308,n836);
nor (n1308,n1309,n1310);
and (n1309,n49,n1037);
and (n1310,n39,n1039);
xor (n1311,n1312,n349);
or (n1312,n1313,n1314);
and (n1313,n144,n486);
and (n1314,n176,n490);
xor (n1315,n1316,n488);
or (n1316,n1317,n1318);
and (n1317,n65,n709);
and (n1318,n86,n713);
nand (n1319,n1320,n1321,n1322);
nand (n1320,n1079,n1083);
nand (n1321,n1087,n1083);
nand (n1322,n1079,n1087);
xor (n1323,n1324,n1342);
xor (n1324,n1325,n1329);
nand (n1325,n1326,n1327,n1328);
nand (n1326,n1018,n1023);
nand (n1327,n1029,n1023);
nand (n1328,n1018,n1029);
xor (n1329,n1330,n1340);
xor (n1330,n1331,n1335);
xor (n1331,n1332,n267);
or (n1332,n1333,n1334);
and (n1333,n252,n347);
and (n1334,n339,n351);
xor (n1335,n68,n1336);
xor (n1336,n1337,n711);
or (n1337,n1338,n1339);
and (n1338,n53,n834);
and (n1339,n61,n838);
xnor (n1340,n1341,n68);
nand (n1341,n1065,n62);
xor (n1342,n1343,n1352);
xor (n1343,n1344,n1348);
xor (n1344,n1345,n16);
or (n1345,n1346,n1347);
and (n1346,n385,n265);
and (n1347,n457,n269);
xor (n1348,n1349,n20);
or (n1349,n1350,n1351);
and (n1350,n678,n14);
and (n1351,n682,n18);
xor (n1352,n1353,n30);
or (n1353,n1354,n1355);
and (n1354,n684,n24);
and (n1355,n818,n28);
nand (n1356,n1357,n1358,n1359);
nand (n1357,n1016,n1041);
nand (n1358,n1067,n1041);
nand (n1359,n1016,n1067);
nand (n1360,n1361,n1362,n1363);
nand (n1361,n1192,n1196);
nand (n1362,n1230,n1196);
nand (n1363,n1192,n1230);
nor (n1364,n1365,n1369);
nand (n1365,n1366,n1367,n1368);
nand (n1366,n1276,n1297);
nand (n1367,n1360,n1297);
nand (n1368,n1276,n1360);
xor (n1369,n1370,n1379);
xor (n1370,n1371,n1375);
nand (n1371,n1372,n1373,n1374);
nand (n1372,n1278,n1289);
nand (n1373,n1293,n1289);
nand (n1374,n1278,n1293);
nand (n1375,n1376,n1377,n1378);
nand (n1376,n1299,n1323);
nand (n1377,n1356,n1323);
nand (n1378,n1299,n1356);
xor (n1379,n1380,n1441);
xor (n1380,n1381,n1412);
xor (n1381,n1382,n1401);
xor (n1382,n1383,n1397);
xor (n1383,n1384,n1393);
xor (n1384,n1385,n1389);
xor (n1385,n1386,n349);
or (n1386,n1387,n1388);
and (n1387,n86,n486);
and (n1388,n144,n490);
xor (n1389,n1390,n488);
or (n1390,n1391,n1392);
and (n1391,n61,n709);
and (n1392,n65,n713);
xor (n1393,n1394,n267);
or (n1394,n1395,n1396);
and (n1395,n176,n347);
and (n1396,n252,n351);
nand (n1397,n1398,n1399,n1400);
nand (n1398,n1331,n1335);
nand (n1399,n1340,n1335);
nand (n1400,n1331,n1340);
xor (n1401,n1402,n1408);
xor (n1402,n1403,n1407);
xor (n1403,n1404,n16);
or (n1404,n1405,n1406);
and (n1405,n339,n265);
and (n1406,n385,n269);
and (n1407,n68,n1336);
xor (n1408,n1409,n20);
or (n1409,n1410,n1411);
and (n1410,n457,n14);
and (n1411,n678,n18);
xor (n1412,n1413,n1437);
xor (n1413,n1414,n1418);
nand (n1414,n1415,n1416,n1417);
nand (n1415,n1344,n1348);
nand (n1416,n1352,n1348);
nand (n1417,n1344,n1352);
xor (n1418,n1419,n1428);
xor (n1419,n1420,n1424);
xor (n1420,n1421,n30);
or (n1421,n1422,n1423);
and (n1422,n682,n24);
and (n1423,n684,n28);
xor (n1424,n1425,n42);
or (n1425,n1426,n1427);
and (n1426,n818,n36);
and (n1427,n1022,n40);
xor (n1428,n1429,n1433);
xnor (n1429,n1430,n836);
nor (n1430,n1431,n1432);
and (n1431,n39,n1037);
and (n1432,n35,n1039);
xor (n1433,n1434,n711);
or (n1434,n1435,n1436);
and (n1435,n49,n834);
and (n1436,n53,n838);
nand (n1437,n1438,n1439,n1440);
nand (n1438,n1280,n1284);
nand (n1439,n1285,n1284);
nand (n1440,n1280,n1285);
xor (n1441,n1442,n1461);
xor (n1442,n1443,n1457);
xor (n1443,n1444,n1453);
xor (n1444,n1445,n1449);
xor (n1445,n1446,n56);
or (n1446,n1447,n1448);
and (n1447,n1026,n50);
and (n1448,n1028,n54);
xor (n1449,n1450,n68);
or (n1450,n1451,n1452);
and (n1451,n1051,n62);
and (n1452,n1065,n66);
nand (n1453,n1454,n1455,n1456);
nand (n1454,n1307,n1311);
nand (n1455,n1315,n1311);
nand (n1456,n1307,n1315);
nand (n1457,n1458,n1459,n1460);
nand (n1458,n1301,n1305);
nand (n1459,n1319,n1305);
nand (n1460,n1301,n1319);
nand (n1461,n1462,n1463,n1464);
nand (n1462,n1325,n1329);
nand (n1463,n1342,n1329);
nand (n1464,n1325,n1342);
nor (n1465,n1466,n1571);
nor (n1466,n1467,n1471);
nand (n1467,n1468,n1469,n1470);
nand (n1468,n1371,n1375);
nand (n1469,n1379,n1375);
nand (n1470,n1371,n1379);
xor (n1471,n1472,n1567);
xor (n1472,n1473,n1507);
xor (n1473,n1474,n1503);
xor (n1474,n1475,n1479);
nand (n1475,n1476,n1477,n1478);
nand (n1476,n1383,n1397);
nand (n1477,n1401,n1397);
nand (n1478,n1383,n1401);
xor (n1479,n1480,n1489);
xor (n1480,n1481,n1485);
xor (n1481,n1482,n68);
or (n1482,n1483,n1484);
and (n1483,n1028,n62);
and (n1484,n1051,n66);
nand (n1485,n1486,n1487,n1488);
nand (n1486,n1403,n1407);
nand (n1487,n1408,n1407);
nand (n1488,n1403,n1408);
xor (n1489,n1490,n1499);
xor (n1490,n1491,n1495);
xor (n1491,n1492,n349);
or (n1492,n1493,n1494);
and (n1493,n65,n486);
and (n1494,n86,n490);
xnor (n1495,n1496,n836);
nor (n1496,n1497,n1498);
and (n1497,n35,n1037);
and (n1498,n27,n1039);
xor (n1499,n1500,n488);
or (n1500,n1501,n1502);
and (n1501,n53,n709);
and (n1502,n61,n713);
nand (n1503,n1504,n1505,n1506);
nand (n1504,n1414,n1418);
nand (n1505,n1437,n1418);
nand (n1506,n1414,n1437);
xor (n1507,n1508,n1563);
xor (n1508,n1509,n1531);
xor (n1509,n1510,n1519);
xor (n1510,n1511,n1515);
nand (n1511,n1512,n1513,n1514);
nand (n1512,n1385,n1389);
nand (n1513,n1393,n1389);
nand (n1514,n1385,n1393);
nand (n1515,n1516,n1517,n1518);
nand (n1516,n1420,n1424);
nand (n1517,n1428,n1424);
nand (n1518,n1420,n1428);
xor (n1519,n1520,n1527);
xor (n1520,n1521,n1525);
xor (n1521,n1522,n267);
or (n1522,n1523,n1524);
and (n1523,n144,n347);
and (n1524,n176,n351);
xnor (n1525,n1526,n89);
nand (n1526,n1065,n83);
xor (n1527,n1528,n16);
or (n1528,n1529,n1530);
and (n1529,n252,n265);
and (n1530,n339,n269);
xor (n1531,n1532,n1551);
xor (n1532,n1533,n1537);
nand (n1533,n1534,n1535,n1536);
nand (n1534,n1445,n1449);
nand (n1535,n1453,n1449);
nand (n1536,n1445,n1453);
xor (n1537,n1538,n1547);
xor (n1538,n1539,n1543);
xor (n1539,n1540,n20);
or (n1540,n1541,n1542);
and (n1541,n385,n14);
and (n1542,n457,n18);
xor (n1543,n1544,n30);
or (n1544,n1545,n1546);
and (n1545,n678,n24);
and (n1546,n682,n28);
xor (n1547,n1548,n42);
or (n1548,n1549,n1550);
and (n1549,n684,n36);
and (n1550,n818,n40);
xor (n1551,n1552,n1559);
xor (n1552,n1553,n1558);
xor (n1553,n89,n1554);
xor (n1554,n1555,n711);
or (n1555,n1556,n1557);
and (n1556,n39,n834);
and (n1557,n49,n838);
and (n1558,n1429,n1433);
xor (n1559,n1560,n56);
or (n1560,n1561,n1562);
and (n1561,n1022,n50);
and (n1562,n1026,n54);
nand (n1563,n1564,n1565,n1566);
nand (n1564,n1443,n1457);
nand (n1565,n1461,n1457);
nand (n1566,n1443,n1461);
nand (n1567,n1568,n1569,n1570);
nand (n1568,n1381,n1412);
nand (n1569,n1441,n1412);
nand (n1570,n1381,n1441);
nor (n1571,n1572,n1576);
nand (n1572,n1573,n1574,n1575);
nand (n1573,n1473,n1507);
nand (n1574,n1567,n1507);
nand (n1575,n1473,n1567);
xor (n1576,n1577,n1586);
xor (n1577,n1578,n1582);
nand (n1578,n1579,n1580,n1581);
nand (n1579,n1475,n1479);
nand (n1580,n1503,n1479);
nand (n1581,n1475,n1503);
nand (n1582,n1583,n1584,n1585);
nand (n1583,n1509,n1531);
nand (n1584,n1563,n1531);
nand (n1585,n1509,n1563);
xor (n1586,n1587,n1648);
xor (n1587,n1588,n1612);
xor (n1588,n1589,n1608);
xor (n1589,n1590,n1594);
nand (n1590,n1591,n1592,n1593);
nand (n1591,n1539,n1543);
nand (n1592,n1547,n1543);
nand (n1593,n1539,n1547);
xor (n1594,n1595,n1604);
xor (n1595,n1596,n1600);
xor (n1596,n1597,n16);
or (n1597,n1598,n1599);
and (n1598,n176,n265);
and (n1599,n252,n269);
xor (n1600,n1601,n20);
or (n1601,n1602,n1603);
and (n1602,n339,n14);
and (n1603,n385,n18);
xor (n1604,n1605,n30);
or (n1605,n1606,n1607);
and (n1606,n457,n24);
and (n1607,n678,n28);
nand (n1608,n1609,n1610,n1611);
nand (n1609,n1553,n1558);
nand (n1610,n1559,n1558);
nand (n1611,n1553,n1559);
xor (n1612,n1613,n1634);
xor (n1613,n1614,n1630);
xor (n1614,n1615,n1629);
xor (n1615,n1616,n1620);
xor (n1616,n1617,n42);
or (n1617,n1618,n1619);
and (n1618,n682,n36);
and (n1619,n684,n40);
xor (n1620,n1621,n1625);
xnor (n1621,n1622,n836);
nor (n1622,n1623,n1624);
and (n1623,n27,n1037);
and (n1624,n13,n1039);
xor (n1625,n1626,n711);
or (n1626,n1627,n1628);
and (n1627,n35,n834);
and (n1628,n39,n838);
and (n1629,n89,n1554);
nand (n1630,n1631,n1632,n1633);
nand (n1631,n1481,n1485);
nand (n1632,n1489,n1485);
nand (n1633,n1481,n1489);
xor (n1634,n1635,n1644);
xor (n1635,n1636,n1640);
xor (n1636,n1637,n56);
or (n1637,n1638,n1639);
and (n1638,n818,n50);
and (n1639,n1022,n54);
xor (n1640,n1641,n89);
or (n1641,n1642,n1643);
and (n1642,n1051,n83);
and (n1643,n1065,n87);
xor (n1644,n1645,n68);
or (n1645,n1646,n1647);
and (n1646,n1026,n62);
and (n1647,n1028,n66);
xor (n1648,n1649,n1678);
xor (n1649,n1650,n1674);
xor (n1650,n1651,n1670);
xor (n1651,n1652,n1656);
nand (n1652,n1653,n1654,n1655);
nand (n1653,n1491,n1495);
nand (n1654,n1499,n1495);
nand (n1655,n1491,n1499);
xor (n1656,n1657,n1666);
xor (n1657,n1658,n1662);
xor (n1658,n1659,n349);
or (n1659,n1660,n1661);
and (n1660,n61,n486);
and (n1661,n65,n490);
xor (n1662,n1663,n488);
or (n1663,n1664,n1665);
and (n1664,n49,n709);
and (n1665,n53,n713);
xor (n1666,n1667,n267);
or (n1667,n1668,n1669);
and (n1668,n86,n347);
and (n1669,n144,n351);
nand (n1670,n1671,n1672,n1673);
nand (n1671,n1521,n1525);
nand (n1672,n1527,n1525);
nand (n1673,n1521,n1527);
nand (n1674,n1675,n1676,n1677);
nand (n1675,n1511,n1515);
nand (n1676,n1519,n1515);
nand (n1677,n1511,n1519);
nand (n1678,n1679,n1680,n1681);
nand (n1679,n1533,n1537);
nand (n1680,n1551,n1537);
nand (n1681,n1533,n1551);
nor (n1682,n1683,n1955);
nor (n1683,n1684,n1931);
nor (n1684,n1685,n1929);
nor (n1685,n1686,n1904);
nand (n1686,n1687,n1866);
nand (n1687,n1688,n1813,n1865);
nand (n1688,n1689,n1740);
xor (n1689,n1690,n1727);
xor (n1690,n1691,n1712);
nand (n1691,n1692,n1706,n1711);
nand (n1692,n1693,n1702);
and (n1693,n1694,n1698);
xnor (n1694,n1695,n836);
nor (n1695,n1696,n1697);
and (n1696,n252,n1037);
and (n1697,n176,n1039);
xor (n1698,n1699,n711);
or (n1699,n1700,n1701);
and (n1700,n339,n834);
and (n1701,n385,n838);
xor (n1702,n1703,n16);
or (n1703,n1704,n1705);
and (n1704,n1022,n265);
and (n1705,n1026,n269);
nand (n1706,n1707,n1702);
xor (n1707,n1708,n20);
or (n1708,n1709,n1710);
and (n1709,n1028,n14);
and (n1710,n1051,n18);
nand (n1711,n1693,n1707);
xor (n1712,n1713,n1722);
xor (n1713,n1714,n1718);
xor (n1714,n1715,n349);
or (n1715,n1716,n1717);
and (n1716,n457,n486);
and (n1717,n678,n490);
xor (n1718,n1719,n488);
or (n1719,n1720,n1721);
and (n1720,n339,n709);
and (n1721,n385,n713);
and (n1722,n1723,n30);
xnor (n1723,n1724,n836);
nor (n1724,n1725,n1726);
and (n1725,n176,n1037);
and (n1726,n144,n1039);
nand (n1727,n1728,n1734,n1739);
nand (n1728,n1729,n1733);
xor (n1729,n1730,n488);
or (n1730,n1731,n1732);
and (n1731,n385,n709);
and (n1732,n457,n713);
xor (n1733,n1723,n30);
nand (n1734,n1735,n1733);
xor (n1735,n1736,n267);
or (n1736,n1737,n1738);
and (n1737,n684,n347);
and (n1738,n818,n351);
nand (n1739,n1729,n1735);
xor (n1740,n1741,n1777);
xor (n1741,n1742,n1753);
xor (n1742,n1743,n1749);
xor (n1743,n1744,n1748);
xor (n1744,n1745,n267);
or (n1745,n1746,n1747);
and (n1746,n682,n347);
and (n1747,n684,n351);
xor (n1748,n1152,n1156);
xor (n1749,n1750,n16);
or (n1750,n1751,n1752);
and (n1751,n818,n265);
and (n1752,n1022,n269);
xor (n1753,n1754,n1763);
xor (n1754,n1755,n1759);
xor (n1755,n1756,n20);
or (n1756,n1757,n1758);
and (n1757,n1026,n14);
and (n1758,n1028,n18);
xor (n1759,n1760,n30);
or (n1760,n1761,n1762);
and (n1761,n1051,n24);
and (n1762,n1065,n28);
nand (n1763,n1764,n1771,n1776);
nand (n1764,n1765,n1769);
xor (n1765,n1766,n711);
or (n1766,n1767,n1768);
and (n1767,n252,n834);
and (n1768,n339,n838);
xnor (n1769,n1770,n30);
nand (n1770,n1065,n24);
nand (n1771,n1772,n1769);
xor (n1772,n1773,n349);
or (n1773,n1774,n1775);
and (n1774,n678,n486);
and (n1775,n682,n490);
nand (n1776,n1765,n1772);
nand (n1777,n1778,n1798,n1812);
nand (n1778,n1779,n1781);
xor (n1779,n1780,n1772);
xor (n1780,n1765,n1769);
nand (n1781,n1782,n1791,n1797);
nand (n1782,n1783,n1787);
xor (n1783,n1784,n349);
or (n1784,n1785,n1786);
and (n1785,n682,n486);
and (n1786,n684,n490);
xor (n1787,n1788,n488);
or (n1788,n1789,n1790);
and (n1789,n457,n709);
and (n1790,n678,n713);
nand (n1791,n1792,n1787);
and (n1792,n1793,n20);
xnor (n1793,n1794,n836);
nor (n1794,n1795,n1796);
and (n1795,n339,n1037);
and (n1796,n252,n1039);
nand (n1797,n1783,n1792);
nand (n1798,n1799,n1781);
nand (n1799,n1800,n1806,n1811);
nand (n1800,n1801,n1805);
xor (n1801,n1802,n267);
or (n1802,n1803,n1804);
and (n1803,n818,n347);
and (n1804,n1022,n351);
xor (n1805,n1694,n1698);
nand (n1806,n1807,n1805);
xor (n1807,n1808,n16);
or (n1808,n1809,n1810);
and (n1809,n1026,n265);
and (n1810,n1028,n269);
nand (n1811,n1801,n1807);
nand (n1812,n1779,n1799);
nand (n1813,n1814,n1740);
nand (n1814,n1815,n1820,n1864);
nand (n1815,n1816,n1818);
xor (n1816,n1817,n1707);
xor (n1817,n1693,n1702);
xor (n1818,n1819,n1735);
xor (n1819,n1729,n1733);
nand (n1820,n1821,n1818);
nand (n1821,n1822,n1841,n1863);
nand (n1822,n1823,n1827);
xor (n1823,n1824,n20);
or (n1824,n1825,n1826);
and (n1825,n1051,n14);
and (n1826,n1065,n18);
nand (n1827,n1828,n1835,n1840);
nand (n1828,n1829,n1833);
xor (n1829,n1830,n711);
or (n1830,n1831,n1832);
and (n1831,n385,n834);
and (n1832,n457,n838);
xnor (n1833,n1834,n20);
nand (n1834,n1065,n14);
nand (n1835,n1836,n1833);
xor (n1836,n1837,n349);
or (n1837,n1838,n1839);
and (n1838,n684,n486);
and (n1839,n818,n490);
nand (n1840,n1829,n1836);
nand (n1841,n1842,n1827);
nand (n1842,n1843,n1857,n1862);
nand (n1843,n1844,n1848);
xor (n1844,n1845,n488);
or (n1845,n1846,n1847);
and (n1846,n678,n709);
and (n1847,n682,n713);
and (n1848,n1849,n1853);
xnor (n1849,n1850,n836);
nor (n1850,n1851,n1852);
and (n1851,n385,n1037);
and (n1852,n339,n1039);
xor (n1853,n1854,n711);
or (n1854,n1855,n1856);
and (n1855,n457,n834);
and (n1856,n678,n838);
nand (n1857,n1858,n1848);
xor (n1858,n1859,n267);
or (n1859,n1860,n1861);
and (n1860,n1022,n347);
and (n1861,n1026,n351);
nand (n1862,n1844,n1858);
nand (n1863,n1823,n1842);
nand (n1864,n1816,n1821);
nand (n1865,n1689,n1814);
xor (n1866,n1867,n1882);
xor (n1867,n1868,n1878);
xor (n1868,n1869,n1876);
xor (n1869,n1870,n1874);
nand (n1870,n1871,n1872,n1873);
nand (n1871,n1714,n1718);
nand (n1872,n1722,n1718);
nand (n1873,n1714,n1722);
xor (n1874,n1875,n1165);
xor (n1875,n1151,n1160);
xor (n1876,n1877,n1266);
xor (n1877,n1260,n1264);
nand (n1878,n1879,n1880,n1881);
nand (n1879,n1742,n1753);
nand (n1880,n1777,n1753);
nand (n1881,n1742,n1777);
xor (n1882,n1883,n1892);
xor (n1883,n1884,n1888);
nand (n1884,n1885,n1886,n1887);
nand (n1885,n1755,n1759);
nand (n1886,n1763,n1759);
nand (n1887,n1755,n1763);
nand (n1888,n1889,n1890,n1891);
nand (n1889,n1691,n1712);
nand (n1890,n1727,n1712);
nand (n1891,n1691,n1727);
xor (n1892,n1893,n1902);
xor (n1893,n1894,n1898);
xor (n1894,n1895,n30);
or (n1895,n1896,n1897);
and (n1896,n1028,n24);
and (n1897,n1051,n28);
nand (n1898,n1899,n1900,n1901);
nand (n1899,n1744,n1748);
nand (n1900,n1749,n1748);
nand (n1901,n1744,n1749);
xor (n1902,n1903,n1252);
xor (n1903,n1243,n1247);
nor (n1904,n1905,n1909);
nand (n1905,n1906,n1907,n1908);
nand (n1906,n1868,n1878);
nand (n1907,n1882,n1878);
nand (n1908,n1868,n1882);
xor (n1909,n1910,n1917);
xor (n1910,n1911,n1913);
xor (n1911,n1912,n1173);
xor (n1912,n1149,n1170);
nand (n1913,n1914,n1915,n1916);
nand (n1914,n1884,n1888);
nand (n1915,n1892,n1888);
nand (n1916,n1884,n1892);
xor (n1917,n1918,n1927);
xor (n1918,n1919,n1923);
nand (n1919,n1920,n1921,n1922);
nand (n1920,n1894,n1898);
nand (n1921,n1902,n1898);
nand (n1922,n1894,n1902);
nand (n1923,n1924,n1925,n1926);
nand (n1924,n1870,n1874);
nand (n1925,n1876,n1874);
nand (n1926,n1870,n1876);
xor (n1927,n1928,n1258);
xor (n1928,n1241,n1255);
not (n1929,n1930);
nand (n1930,n1905,n1909);
not (n1931,n1932);
nor (n1932,n1933,n1948);
nor (n1933,n1934,n1938);
nand (n1934,n1935,n1936,n1937);
nand (n1935,n1911,n1913);
nand (n1936,n1917,n1913);
nand (n1937,n1911,n1917);
xor (n1938,n1939,n1946);
xor (n1939,n1940,n1942);
xor (n1940,n1941,n1239);
xor (n1941,n1232,n1236);
nand (n1942,n1943,n1944,n1945);
nand (n1943,n1919,n1923);
nand (n1944,n1927,n1923);
nand (n1945,n1919,n1927);
xor (n1946,n1947,n1147);
xor (n1947,n1093,n1095);
nor (n1948,n1949,n1953);
nand (n1949,n1950,n1951,n1952);
nand (n1950,n1940,n1942);
nand (n1951,n1946,n1942);
nand (n1952,n1940,n1946);
xor (n1953,n1954,n1190);
xor (n1954,n1014,n1091);
not (n1955,n1956);
nor (n1956,n1957,n1959);
nor (n1957,n1958,n1948);
nand (n1958,n1934,n1938);
not (n1959,n1960);
nand (n1960,n1949,n1953);
not (n1961,n1962);
nor (n1962,n1963,n1970);
nor (n1963,n1964,n1969);
nor (n1964,n1965,n1967);
nor (n1965,n1966,n1364);
nand (n1966,n1012,n1274);
not (n1967,n1968);
nand (n1968,n1365,n1369);
not (n1969,n1465);
not (n1970,n1971);
nor (n1971,n1972,n1974);
nor (n1972,n1973,n1571);
nand (n1973,n1467,n1471);
not (n1974,n1975);
nand (n1975,n1572,n1576);
not (n1976,n1977);
nor (n1977,n1978,n2393);
nand (n1978,n1979,n2206);
nor (n1979,n1980,n2092);
nor (n1980,n1981,n1985);
nand (n1981,n1982,n1983,n1984);
nand (n1982,n1578,n1582);
nand (n1983,n1586,n1582);
nand (n1984,n1578,n1586);
xor (n1985,n1986,n2088);
xor (n1986,n1987,n2020);
xor (n1987,n1988,n2016);
xor (n1988,n1989,n2012);
xor (n1989,n1990,n2008);
xor (n1990,n1991,n2004);
xor (n1991,n1992,n2001);
xor (n1992,n1993,n1997);
xor (n1993,n1994,n711);
or (n1994,n1995,n1996);
and (n1995,n27,n834);
and (n1996,n35,n838);
xor (n1997,n1998,n488);
or (n1998,n1999,n2000);
and (n1999,n39,n709);
and (n2000,n49,n713);
xnor (n2001,n2002,n836);
nor (n2002,n2003,n1624);
and (n2003,n13,n1037);
nand (n2004,n2005,n2006,n2007);
nand (n2005,n1596,n1600);
nand (n2006,n1604,n1600);
nand (n2007,n1596,n1604);
nand (n2008,n2009,n2010,n2011);
nand (n2009,n1616,n1620);
nand (n2010,n1629,n1620);
nand (n2011,n1616,n1629);
nand (n2012,n2013,n2014,n2015);
nand (n2013,n1590,n1594);
nand (n2014,n1608,n1594);
nand (n2015,n1590,n1608);
nand (n2016,n2017,n2018,n2019);
nand (n2017,n1614,n1630);
nand (n2018,n1634,n1630);
nand (n2019,n1614,n1634);
xor (n2020,n2021,n2084);
xor (n2021,n2022,n2060);
xor (n2022,n2023,n2045);
xor (n2023,n2024,n2038);
xor (n2024,n2025,n2034);
xor (n2025,n2026,n2030);
xor (n2026,n2027,n267);
or (n2027,n2028,n2029);
and (n2028,n65,n347);
and (n2029,n86,n351);
xor (n2030,n2031,n16);
or (n2031,n2032,n2033);
and (n2032,n144,n265);
and (n2033,n176,n269);
xor (n2034,n2035,n20);
or (n2035,n2036,n2037);
and (n2036,n252,n14);
and (n2037,n339,n18);
xor (n2038,n2039,n2041);
xor (n2039,n89,n2040);
and (n2040,n1621,n1625);
xor (n2041,n2042,n56);
or (n2042,n2043,n2044);
and (n2043,n684,n50);
and (n2044,n818,n54);
xor (n2045,n2046,n2055);
xor (n2046,n2047,n2051);
xor (n2047,n2048,n30);
or (n2048,n2049,n2050);
and (n2049,n385,n24);
and (n2050,n457,n28);
xor (n2051,n2052,n42);
or (n2052,n2053,n2054);
and (n2053,n678,n36);
and (n2054,n682,n40);
xor (n2055,n89,n2056);
xor (n2056,n2057,n349);
or (n2057,n2058,n2059);
and (n2058,n53,n486);
and (n2059,n61,n490);
xor (n2060,n2061,n2070);
xor (n2061,n2062,n2066);
nand (n2062,n2063,n2064,n2065);
nand (n2063,n1636,n1640);
nand (n2064,n1644,n1640);
nand (n2065,n1636,n1644);
nand (n2066,n2067,n2068,n2069);
nand (n2067,n1652,n1656);
nand (n2068,n1670,n1656);
nand (n2069,n1652,n1670);
xor (n2070,n2071,n2080);
xor (n2071,n2072,n2076);
xor (n2072,n2073,n68);
or (n2073,n2074,n2075);
and (n2074,n1022,n62);
and (n2075,n1026,n66);
xor (n2076,n2077,n89);
or (n2077,n2078,n2079);
and (n2078,n1028,n83);
and (n2079,n1051,n87);
nand (n2080,n2081,n2082,n2083);
nand (n2081,n1658,n1662);
nand (n2082,n1666,n1662);
nand (n2083,n1658,n1666);
nand (n2084,n2085,n2086,n2087);
nand (n2085,n1650,n1674);
nand (n2086,n1678,n1674);
nand (n2087,n1650,n1678);
nand (n2088,n2089,n2090,n2091);
nand (n2089,n1588,n1612);
nand (n2090,n1648,n1612);
nand (n2091,n1588,n1648);
nor (n2092,n2093,n2097);
nand (n2093,n2094,n2095,n2096);
nand (n2094,n1987,n2020);
nand (n2095,n2088,n2020);
nand (n2096,n1987,n2088);
xor (n2097,n2098,n2107);
xor (n2098,n2099,n2103);
nand (n2099,n2100,n2101,n2102);
nand (n2100,n1989,n2012);
nand (n2101,n2016,n2012);
nand (n2102,n1989,n2016);
nand (n2103,n2104,n2105,n2106);
nand (n2104,n2022,n2060);
nand (n2105,n2084,n2060);
nand (n2106,n2022,n2084);
xor (n2107,n2108,n2165);
xor (n2108,n2109,n2140);
xor (n2109,n2110,n2126);
xor (n2110,n2111,n2115);
nand (n2111,n2112,n2113,n2114);
nand (n2112,n89,n2040);
nand (n2113,n2041,n2040);
nand (n2114,n89,n2041);
xor (n2115,n2116,n2122);
xor (n2116,n2117,n2121);
xor (n2117,n2118,n42);
or (n2118,n2119,n2120);
and (n2119,n457,n36);
and (n2120,n678,n40);
and (n2121,n89,n2056);
xor (n2122,n2123,n56);
or (n2123,n2124,n2125);
and (n2124,n682,n50);
and (n2125,n684,n54);
xor (n2126,n2127,n2136);
xor (n2127,n2128,n2132);
xor (n2128,n2129,n68);
or (n2129,n2130,n2131);
and (n2130,n818,n62);
and (n2131,n1022,n66);
xor (n2132,n2133,n89);
or (n2133,n2134,n2135);
and (n2134,n1026,n83);
and (n2135,n1028,n87);
nand (n2136,n2137,n2138,n2139);
nand (n2137,n1993,n1997);
nand (n2138,n2001,n1997);
nand (n2139,n1993,n2001);
xor (n2140,n2141,n2150);
xor (n2141,n2142,n2146);
nand (n2142,n2143,n2144,n2145);
nand (n2143,n2072,n2076);
nand (n2144,n2080,n2076);
nand (n2145,n2072,n2080);
nand (n2146,n2147,n2148,n2149);
nand (n2147,n1991,n2004);
nand (n2148,n2008,n2004);
nand (n2149,n1991,n2008);
xor (n2150,n2151,n89);
xor (n2151,n2152,n2156);
nand (n2152,n2153,n2154,n2155);
nand (n2153,n2026,n2030);
nand (n2154,n2034,n2030);
nand (n2155,n2026,n2034);
xor (n2156,n2157,n2162);
not (n2157,n2158);
xor (n2158,n2159,n349);
or (n2159,n2160,n2161);
and (n2160,n49,n486);
and (n2161,n53,n490);
xor (n2162,n2163,n711);
or (n2163,n833,n2164);
and (n2164,n27,n838);
xor (n2165,n2166,n2202);
xor (n2166,n2167,n2171);
nand (n2167,n2168,n2169,n2170);
nand (n2168,n2024,n2038);
nand (n2169,n2045,n2038);
nand (n2170,n2024,n2045);
xor (n2171,n2172,n2191);
xor (n2172,n2173,n2177);
nand (n2173,n2174,n2175,n2176);
nand (n2174,n2047,n2051);
nand (n2175,n2055,n2051);
nand (n2176,n2047,n2055);
xor (n2177,n2178,n2187);
xor (n2178,n2179,n2183);
xor (n2179,n2180,n16);
or (n2180,n2181,n2182);
and (n2181,n86,n265);
and (n2182,n144,n269);
xor (n2183,n2184,n20);
or (n2184,n2185,n2186);
and (n2185,n176,n14);
and (n2186,n252,n18);
xor (n2187,n2188,n30);
or (n2188,n2189,n2190);
and (n2189,n339,n24);
and (n2190,n385,n28);
xor (n2191,n2192,n2198);
xor (n2192,n2193,n2197);
xor (n2193,n2194,n488);
or (n2194,n2195,n2196);
and (n2195,n35,n709);
and (n2196,n39,n713);
not (n2197,n2001);
xor (n2198,n2199,n267);
or (n2199,n2200,n2201);
and (n2200,n61,n347);
and (n2201,n65,n351);
nand (n2202,n2203,n2204,n2205);
nand (n2203,n2062,n2066);
nand (n2204,n2070,n2066);
nand (n2205,n2062,n2070);
nor (n2206,n2207,n2314);
nor (n2207,n2208,n2212);
nand (n2208,n2209,n2210,n2211);
nand (n2209,n2099,n2103);
nand (n2210,n2107,n2103);
nand (n2211,n2099,n2107);
xor (n2212,n2213,n2310);
xor (n2213,n2214,n2254);
xor (n2214,n2215,n2250);
xor (n2215,n2216,n2246);
xor (n2216,n2217,n2242);
xor (n2217,n2218,n2232);
xor (n2218,n2219,n2228);
xor (n2219,n2220,n2224);
xor (n2220,n2221,n16);
or (n2221,n2222,n2223);
and (n2222,n65,n265);
and (n2223,n86,n269);
xor (n2224,n2225,n20);
or (n2225,n2226,n2227);
and (n2226,n144,n14);
and (n2227,n176,n18);
xor (n2228,n2229,n42);
or (n2229,n2230,n2231);
and (n2230,n385,n36);
and (n2231,n457,n40);
xor (n2232,n2233,n2238);
xor (n2233,n2234,n831);
xor (n2234,n2235,n349);
or (n2235,n2236,n2237);
and (n2236,n39,n486);
and (n2237,n49,n490);
xor (n2238,n2239,n267);
or (n2239,n2240,n2241);
and (n2240,n53,n347);
and (n2241,n61,n351);
nand (n2242,n2243,n2244,n2245);
nand (n2243,n2117,n2121);
nand (n2244,n2122,n2121);
nand (n2245,n2117,n2122);
nand (n2246,n2247,n2248,n2249);
nand (n2247,n2111,n2115);
nand (n2248,n2126,n2115);
nand (n2249,n2111,n2126);
nand (n2250,n2251,n2252,n2253);
nand (n2251,n2142,n2146);
nand (n2252,n2150,n2146);
nand (n2253,n2142,n2150);
xor (n2254,n2255,n2306);
xor (n2255,n2256,n2277);
xor (n2256,n2257,n2273);
xor (n2257,n2258,n2269);
xor (n2258,n2259,n2265);
xor (n2259,n2260,n2261);
not (n2260,n872);
xor (n2261,n2262,n30);
or (n2262,n2263,n2264);
and (n2263,n252,n24);
and (n2264,n339,n28);
xor (n2265,n2266,n56);
or (n2266,n2267,n2268);
and (n2267,n678,n50);
and (n2268,n682,n54);
nand (n2269,n2270,n2271,n2272);
nand (n2270,n2128,n2132);
nand (n2271,n2136,n2132);
nand (n2272,n2128,n2136);
nand (n2273,n2274,n2275,n2276);
nand (n2274,n2152,n2156);
nand (n2275,n89,n2156);
nand (n2276,n2152,n89);
xor (n2277,n2278,n2302);
xor (n2278,n2279,n2292);
xor (n2279,n2280,n2289);
xor (n2280,n2281,n2285);
xor (n2281,n2282,n68);
or (n2282,n2283,n2284);
and (n2283,n684,n62);
and (n2284,n818,n66);
xor (n2285,n2286,n89);
or (n2286,n2287,n2288);
and (n2287,n1022,n83);
and (n2288,n1026,n87);
nand (n2289,n2157,n2290,n2291);
nand (n2290,n2162,n2158);
not (n2291,n2162);
xor (n2292,n2293,n2298);
xor (n2293,n89,n2294);
nand (n2294,n2295,n2296,n2297);
nand (n2295,n2193,n2197);
nand (n2296,n2198,n2197);
nand (n2297,n2193,n2198);
nand (n2298,n2299,n2300,n2301);
nand (n2299,n2179,n2183);
nand (n2300,n2187,n2183);
nand (n2301,n2179,n2187);
nand (n2302,n2303,n2304,n2305);
nand (n2303,n2173,n2177);
nand (n2304,n2191,n2177);
nand (n2305,n2173,n2191);
nand (n2306,n2307,n2308,n2309);
nand (n2307,n2167,n2171);
nand (n2308,n2202,n2171);
nand (n2309,n2167,n2202);
nand (n2310,n2311,n2312,n2313);
nand (n2311,n2109,n2140);
nand (n2312,n2165,n2140);
nand (n2313,n2109,n2165);
nor (n2314,n2315,n2319);
nand (n2315,n2316,n2317,n2318);
nand (n2316,n2214,n2254);
nand (n2317,n2310,n2254);
nand (n2318,n2214,n2310);
xor (n2319,n2320,n2329);
xor (n2320,n2321,n2325);
nand (n2321,n2322,n2323,n2324);
nand (n2322,n2216,n2246);
nand (n2323,n2250,n2246);
nand (n2324,n2216,n2250);
nand (n2325,n2326,n2327,n2328);
nand (n2326,n2256,n2277);
nand (n2327,n2306,n2277);
nand (n2328,n2256,n2306);
xor (n2329,n2330,n2361);
xor (n2330,n2331,n2335);
nand (n2331,n2332,n2333,n2334);
nand (n2332,n2279,n2292);
nand (n2333,n2302,n2292);
nand (n2334,n2279,n2302);
xor (n2335,n2336,n2349);
xor (n2336,n2337,n2341);
nand (n2337,n2338,n2339,n2340);
nand (n2338,n89,n2294);
nand (n2339,n2298,n2294);
nand (n2340,n89,n2298);
xor (n2341,n2342,n2345);
xor (n2342,n2343,n89);
xor (n2343,n2344,n830);
xor (n2344,n822,n825);
nand (n2345,n2346,n2347,n2348);
nand (n2346,n2234,n831);
nand (n2347,n2238,n831);
nand (n2348,n2234,n2238);
xor (n2349,n2350,n2357);
xor (n2350,n2351,n2353);
xor (n2351,n2352,n858);
xor (n2352,n849,n853);
nand (n2353,n2354,n2355,n2356);
nand (n2354,n2220,n2224);
nand (n2355,n2228,n2224);
nand (n2356,n2220,n2228);
nand (n2357,n2358,n2359,n2360);
nand (n2358,n2281,n2285);
nand (n2359,n2289,n2285);
nand (n2360,n2281,n2289);
xor (n2361,n2362,n2371);
xor (n2362,n2363,n2367);
nand (n2363,n2364,n2365,n2366);
nand (n2364,n2218,n2232);
nand (n2365,n2242,n2232);
nand (n2366,n2218,n2242);
nand (n2367,n2368,n2369,n2370);
nand (n2368,n2258,n2269);
nand (n2369,n2273,n2269);
nand (n2370,n2258,n2273);
xor (n2371,n2372,n2379);
xor (n2372,n2373,n2377);
nand (n2373,n2374,n2375,n2376);
nand (n2374,n2260,n2261);
nand (n2375,n2265,n2261);
nand (n2376,n2260,n2265);
xor (n2377,n2378,n877);
xor (n2378,n868,n872);
xor (n2379,n2380,n2389);
xor (n2380,n2381,n2385);
xor (n2381,n2382,n56);
or (n2382,n2383,n2384);
and (n2383,n457,n50);
and (n2384,n678,n54);
xor (n2385,n2386,n68);
or (n2386,n2387,n2388);
and (n2387,n682,n62);
and (n2388,n684,n66);
xor (n2389,n2390,n89);
or (n2390,n2391,n2392);
and (n2391,n818,n83);
and (n2392,n1022,n87);
nand (n2393,n2394,n2478);
nor (n2394,n2395,n2445);
nor (n2395,n2396,n2400);
nand (n2396,n2397,n2398,n2399);
nand (n2397,n2321,n2325);
nand (n2398,n2329,n2325);
nand (n2399,n2321,n2329);
xor (n2400,n2401,n2441);
xor (n2401,n2402,n2422);
xor (n2402,n2403,n2410);
xor (n2403,n2404,n2406);
xor (n2404,n2405,n866);
xor (n2405,n847,n863);
nand (n2406,n2407,n2408,n2409);
nand (n2407,n2373,n2377);
nand (n2408,n2379,n2377);
nand (n2409,n2373,n2379);
xor (n2410,n2411,n2418);
xor (n2411,n2412,n2416);
nand (n2412,n2413,n2414,n2415);
nand (n2413,n2381,n2385);
nand (n2414,n2389,n2385);
nand (n2415,n2381,n2389);
xor (n2416,n2417,n776);
xor (n2417,n770,n774);
nand (n2418,n2419,n2420,n2421);
nand (n2419,n2343,n89);
nand (n2420,n2345,n89);
nand (n2421,n2343,n2345);
xor (n2422,n2423,n2437);
xor (n2423,n2424,n2428);
nand (n2424,n2425,n2426,n2427);
nand (n2425,n2337,n2341);
nand (n2426,n2349,n2341);
nand (n2427,n2337,n2349);
xor (n2428,n2429,n2433);
xor (n2429,n2430,n2432);
xor (n2430,n2431,n792);
xor (n2431,n783,n787);
xor (n2432,n815,n820);
nand (n2433,n2434,n2435,n2436);
nand (n2434,n2351,n2353);
nand (n2435,n2357,n2353);
nand (n2436,n2351,n2357);
nand (n2437,n2438,n2439,n2440);
nand (n2438,n2363,n2367);
nand (n2439,n2371,n2367);
nand (n2440,n2363,n2371);
nand (n2441,n2442,n2443,n2444);
nand (n2442,n2331,n2335);
nand (n2443,n2361,n2335);
nand (n2444,n2331,n2361);
nor (n2445,n2446,n2450);
nand (n2446,n2447,n2448,n2449);
nand (n2447,n2402,n2422);
nand (n2448,n2441,n2422);
nand (n2449,n2402,n2441);
xor (n2450,n2451,n2474);
xor (n2451,n2452,n2462);
xor (n2452,n2453,n2460);
xor (n2453,n2454,n2456);
xor (n2454,n2455,n763);
xor (n2455,n748,n760);
nand (n2456,n2457,n2458,n2459);
nand (n2457,n2412,n2416);
nand (n2458,n2418,n2416);
nand (n2459,n2412,n2418);
xor (n2460,n2461,n798);
xor (n2461,n768,n781);
xor (n2462,n2463,n2470);
xor (n2463,n2464,n2466);
xor (n2464,n2465,n845);
xor (n2465,n812,n842);
nand (n2466,n2467,n2468,n2469);
nand (n2467,n2430,n2432);
nand (n2468,n2433,n2432);
nand (n2469,n2430,n2433);
nand (n2470,n2471,n2472,n2473);
nand (n2471,n2404,n2406);
nand (n2472,n2410,n2406);
nand (n2473,n2404,n2410);
nand (n2474,n2475,n2476,n2477);
nand (n2475,n2424,n2428);
nand (n2476,n2437,n2428);
nand (n2477,n2424,n2437);
nor (n2478,n2479,n2496);
nor (n2479,n2480,n2484);
nand (n2480,n2481,n2482,n2483);
nand (n2481,n2452,n2462);
nand (n2482,n2474,n2462);
nand (n2483,n2452,n2474);
xor (n2484,n2485,n2492);
xor (n2485,n2486,n2490);
nand (n2486,n2487,n2488,n2489);
nand (n2487,n2454,n2456);
nand (n2488,n2460,n2456);
nand (n2489,n2454,n2460);
xor (n2490,n2491,n885);
xor (n2491,n808,n810);
nand (n2492,n2493,n2494,n2495);
nand (n2493,n2464,n2466);
nand (n2494,n2470,n2466);
nand (n2495,n2464,n2470);
nor (n2496,n2497,n2501);
nand (n2497,n2498,n2499,n2500);
nand (n2498,n2486,n2490);
nand (n2499,n2492,n2490);
nand (n2500,n2486,n2492);
xor (n2501,n2502,n806);
xor (n2502,n584,n668);
not (n2503,n2504);
nor (n2504,n2505,n2520);
nor (n2505,n2393,n2506);
nor (n2506,n2507,n2514);
nor (n2507,n2508,n2513);
nor (n2508,n2509,n2511);
nor (n2509,n2510,n2092);
nand (n2510,n1981,n1985);
not (n2511,n2512);
nand (n2512,n2093,n2097);
not (n2513,n2206);
not (n2514,n2515);
nor (n2515,n2516,n2518);
nor (n2516,n2517,n2314);
nand (n2517,n2208,n2212);
not (n2518,n2519);
nand (n2519,n2315,n2319);
not (n2520,n2521);
nor (n2521,n2522,n2529);
nor (n2522,n2523,n2528);
nor (n2523,n2524,n2526);
nor (n2524,n2525,n2445);
nand (n2525,n2396,n2400);
not (n2526,n2527);
nand (n2527,n2446,n2450);
not (n2528,n2478);
not (n2529,n2530);
nor (n2530,n2531,n2533);
nor (n2531,n2532,n2496);
nand (n2532,n2480,n2484);
not (n2533,n2534);
nand (n2534,n2497,n2501);
nand (n2535,n2536,n2955);
nand (n2536,n2537,n2848);
nor (n2537,n2538,n2833);
nor (n2538,n2539,n2704);
nand (n2539,n2540,n2681);
nor (n2540,n2541,n2658);
nor (n2541,n2542,n2631);
nand (n2542,n2543,n2588,n2630);
nand (n2543,n2544,n2556);
xor (n2544,n2545,n2551);
xor (n2545,n2546,n2547);
xor (n2546,n1849,n1853);
xor (n2547,n2548,n16);
or (n2548,n2549,n2550);
and (n2549,n1051,n265);
and (n2550,n1065,n269);
and (n2551,n16,n2552);
xor (n2552,n2553,n711);
or (n2553,n2554,n2555);
and (n2554,n678,n834);
and (n2555,n682,n838);
nand (n2556,n2557,n2574,n2587);
nand (n2557,n2558,n2559);
xor (n2558,n16,n2552);
nand (n2559,n2560,n2569,n2573);
nand (n2560,n2561,n2565);
xor (n2561,n2562,n349);
or (n2562,n2563,n2564);
and (n2563,n1026,n486);
and (n2564,n1028,n490);
xor (n2565,n2566,n488);
or (n2566,n2567,n2568);
and (n2567,n818,n709);
and (n2568,n1022,n713);
nand (n2569,n2570,n2565);
and (n2570,n267,n2571);
xnor (n2571,n2572,n267);
nand (n2572,n1065,n347);
nand (n2573,n2561,n2570);
nand (n2574,n2575,n2559);
xor (n2575,n2576,n2583);
xor (n2576,n2577,n2581);
xnor (n2577,n2578,n836);
nor (n2578,n2579,n2580);
and (n2579,n457,n1037);
and (n2580,n385,n1039);
xnor (n2581,n2582,n16);
nand (n2582,n1065,n265);
xor (n2583,n2584,n349);
or (n2584,n2585,n2586);
and (n2585,n1022,n486);
and (n2586,n1026,n490);
nand (n2587,n2558,n2575);
nand (n2588,n2589,n2556);
xor (n2589,n2590,n2609);
xor (n2590,n2591,n2595);
nand (n2591,n2592,n2593,n2594);
nand (n2592,n2577,n2581);
nand (n2593,n2583,n2581);
nand (n2594,n2577,n2583);
xor (n2595,n2596,n2605);
xor (n2596,n2597,n2601);
xor (n2597,n2598,n349);
or (n2598,n2599,n2600);
and (n2599,n818,n486);
and (n2600,n1022,n490);
xor (n2601,n2602,n488);
or (n2602,n2603,n2604);
and (n2603,n682,n709);
and (n2604,n684,n713);
xor (n2605,n2606,n267);
or (n2606,n2607,n2608);
and (n2607,n1026,n347);
and (n2608,n1028,n351);
nand (n2609,n2610,n2624,n2629);
nand (n2610,n2611,n2615);
xor (n2611,n2612,n488);
or (n2612,n2613,n2614);
and (n2613,n684,n709);
and (n2614,n818,n713);
and (n2615,n2616,n2620);
xnor (n2616,n2617,n836);
nor (n2617,n2618,n2619);
and (n2618,n678,n1037);
and (n2619,n457,n1039);
xor (n2620,n2621,n711);
or (n2621,n2622,n2623);
and (n2622,n682,n834);
and (n2623,n684,n838);
nand (n2624,n2625,n2615);
xor (n2625,n2626,n267);
or (n2626,n2627,n2628);
and (n2627,n1028,n347);
and (n2628,n1051,n351);
nand (n2629,n2611,n2625);
nand (n2630,n2544,n2589);
xor (n2631,n2632,n2646);
xor (n2632,n2633,n2642);
xor (n2633,n2634,n2640);
xor (n2634,n2635,n2639);
xor (n2635,n2636,n16);
or (n2636,n2637,n2638);
and (n2637,n1028,n265);
and (n2638,n1051,n269);
xor (n2639,n1793,n20);
xor (n2640,n2641,n1836);
xor (n2641,n1829,n1833);
nand (n2642,n2643,n2644,n2645);
nand (n2643,n2591,n2595);
nand (n2644,n2609,n2595);
nand (n2645,n2591,n2609);
xor (n2646,n2647,n2656);
xor (n2647,n2648,n2652);
nand (n2648,n2649,n2650,n2651);
nand (n2649,n2546,n2547);
nand (n2650,n2551,n2547);
nand (n2651,n2546,n2551);
nand (n2652,n2653,n2654,n2655);
nand (n2653,n2597,n2601);
nand (n2654,n2605,n2601);
nand (n2655,n2597,n2605);
xor (n2656,n2657,n1858);
xor (n2657,n1844,n1848);
nor (n2658,n2659,n2663);
nand (n2659,n2660,n2661,n2662);
nand (n2660,n2633,n2642);
nand (n2661,n2646,n2642);
nand (n2662,n2633,n2646);
xor (n2663,n2664,n2671);
xor (n2664,n2665,n2667);
xor (n2665,n2666,n1842);
xor (n2666,n1823,n1827);
nand (n2667,n2668,n2669,n2670);
nand (n2668,n2648,n2652);
nand (n2669,n2656,n2652);
nand (n2670,n2648,n2656);
xor (n2671,n2672,n2677);
xor (n2672,n2673,n2675);
xor (n2673,n2674,n1792);
xor (n2674,n1783,n1787);
xor (n2675,n2676,n1807);
xor (n2676,n1801,n1805);
nand (n2677,n2678,n2679,n2680);
nand (n2678,n2635,n2639);
nand (n2679,n2640,n2639);
nand (n2680,n2635,n2640);
nor (n2681,n2682,n2697);
nor (n2682,n2683,n2687);
nand (n2683,n2684,n2685,n2686);
nand (n2684,n2665,n2667);
nand (n2685,n2671,n2667);
nand (n2686,n2665,n2671);
xor (n2687,n2688,n2695);
xor (n2688,n2689,n2691);
xor (n2689,n2690,n1799);
xor (n2690,n1779,n1781);
nand (n2691,n2692,n2693,n2694);
nand (n2692,n2673,n2675);
nand (n2693,n2677,n2675);
nand (n2694,n2673,n2677);
xor (n2695,n2696,n1821);
xor (n2696,n1816,n1818);
nor (n2697,n2698,n2702);
nand (n2698,n2699,n2700,n2701);
nand (n2699,n2689,n2691);
nand (n2700,n2695,n2691);
nand (n2701,n2689,n2695);
xor (n2702,n2703,n1814);
xor (n2703,n1689,n1740);
nor (n2704,n2705,n2827);
nor (n2705,n2706,n2803);
nor (n2706,n2707,n2800);
nor (n2707,n2708,n2776);
nand (n2708,n2709,n2748);
or (n2709,n2710,n2734,n2747);
and (n2710,n2711,n2720);
xor (n2711,n2712,n2716);
xnor (n2712,n2713,n836);
nor (n2713,n2714,n2715);
and (n2714,n684,n1037);
and (n2715,n682,n1039);
xnor (n2716,n2717,n711);
nor (n2717,n2718,n2719);
and (n2718,n1022,n838);
and (n2719,n818,n834);
or (n2720,n2721,n2728,n2733);
and (n2721,n2722,n2724);
not (n2722,n2723);
nand (n2723,n1065,n486);
xnor (n2724,n2725,n836);
nor (n2725,n2726,n2727);
and (n2726,n818,n1037);
and (n2727,n684,n1039);
and (n2728,n2724,n2729);
xnor (n2729,n2730,n711);
nor (n2730,n2731,n2732);
and (n2731,n1026,n838);
and (n2732,n1022,n834);
and (n2733,n2722,n2729);
and (n2734,n2720,n2735);
xor (n2735,n2736,n2743);
xor (n2736,n2737,n2739);
and (n2737,n349,n2738);
xnor (n2738,n2723,n349);
xnor (n2739,n2740,n488);
nor (n2740,n2741,n2742);
and (n2741,n1028,n713);
and (n2742,n1026,n709);
xnor (n2743,n2744,n349);
nor (n2744,n2745,n2746);
and (n2745,n1065,n490);
and (n2746,n1051,n486);
and (n2747,n2711,n2735);
xor (n2748,n2749,n2765);
xor (n2749,n2750,n2754);
or (n2750,n2751,n2752,n2753);
and (n2751,n2737,n2739);
and (n2752,n2739,n2743);
and (n2753,n2737,n2743);
xor (n2754,n2755,n2761);
xor (n2755,n2756,n2757);
and (n2756,n2712,n2716);
xnor (n2757,n2758,n488);
nor (n2758,n2759,n2760);
and (n2759,n1026,n713);
and (n2760,n1022,n709);
xnor (n2761,n2762,n349);
nor (n2762,n2763,n2764);
and (n2763,n1051,n490);
and (n2764,n1028,n486);
xor (n2765,n2766,n2772);
xor (n2766,n2767,n2768);
not (n2767,n2572);
xnor (n2768,n2769,n836);
nor (n2769,n2770,n2771);
and (n2770,n682,n1037);
and (n2771,n678,n1039);
xnor (n2772,n2773,n711);
nor (n2773,n2774,n2775);
and (n2774,n818,n838);
and (n2775,n684,n834);
nor (n2776,n2777,n2781);
or (n2777,n2778,n2779,n2780);
and (n2778,n2750,n2754);
and (n2779,n2754,n2765);
and (n2780,n2750,n2765);
xor (n2781,n2782,n2789);
xor (n2782,n2783,n2787);
or (n2783,n2784,n2785,n2786);
and (n2784,n2756,n2757);
and (n2785,n2757,n2761);
and (n2786,n2756,n2761);
xor (n2787,n2788,n2570);
xor (n2788,n2561,n2565);
xor (n2789,n2790,n2796);
xor (n2790,n2791,n2795);
xor (n2791,n2792,n267);
or (n2792,n2793,n2794);
and (n2793,n1051,n347);
and (n2794,n1065,n351);
xor (n2795,n2616,n2620);
or (n2796,n2797,n2798,n2799);
and (n2797,n2767,n2768);
and (n2798,n2768,n2772);
and (n2799,n2767,n2772);
not (n2800,n2801);
not (n2801,n2802);
and (n2802,n2777,n2781);
not (n2803,n2804);
nor (n2804,n2805,n2820);
nor (n2805,n2806,n2810);
nand (n2806,n2807,n2808,n2809);
nand (n2807,n2783,n2787);
nand (n2808,n2789,n2787);
nand (n2809,n2783,n2789);
xor (n2810,n2811,n2818);
xor (n2811,n2812,n2814);
xor (n2812,n2813,n2625);
xor (n2813,n2611,n2615);
nand (n2814,n2815,n2816,n2817);
nand (n2815,n2791,n2795);
nand (n2816,n2796,n2795);
nand (n2817,n2791,n2796);
xor (n2818,n2819,n2575);
xor (n2819,n2558,n2559);
nor (n2820,n2821,n2825);
nand (n2821,n2822,n2823,n2824);
nand (n2822,n2812,n2814);
nand (n2823,n2818,n2814);
nand (n2824,n2812,n2818);
xor (n2825,n2826,n2589);
xor (n2826,n2544,n2556);
not (n2827,n2828);
nor (n2828,n2829,n2831);
nor (n2829,n2830,n2820);
nand (n2830,n2806,n2810);
not (n2831,n2832);
nand (n2832,n2821,n2825);
not (n2833,n2834);
nor (n2834,n2835,n2842);
nor (n2835,n2836,n2841);
nor (n2836,n2837,n2839);
nor (n2837,n2838,n2658);
nand (n2838,n2542,n2631);
not (n2839,n2840);
nand (n2840,n2659,n2663);
not (n2841,n2681);
not (n2842,n2843);
nor (n2843,n2844,n2846);
nor (n2844,n2845,n2697);
nand (n2845,n2683,n2687);
not (n2846,n2847);
nand (n2847,n2698,n2702);
nand (n2848,n2849,n2853);
nor (n2849,n2850,n2539);
nand (n2850,n2851,n2804);
nor (n2851,n2852,n2776);
nor (n2852,n2709,n2748);
or (n2853,n2854,n2876);
and (n2854,n2855,n2857);
xor (n2855,n2856,n2735);
xor (n2856,n2711,n2720);
or (n2857,n2858,n2872,n2875);
and (n2858,n2859,n2868);
and (n2859,n2860,n2864);
xnor (n2860,n2861,n836);
nor (n2861,n2862,n2863);
and (n2862,n1022,n1037);
and (n2863,n818,n1039);
xnor (n2864,n2865,n711);
nor (n2865,n2866,n2867);
and (n2866,n1028,n838);
and (n2867,n1026,n834);
xnor (n2868,n2869,n488);
nor (n2869,n2870,n2871);
and (n2870,n1051,n713);
and (n2871,n1028,n709);
and (n2872,n2868,n2873);
xor (n2873,n2874,n2729);
xor (n2874,n2722,n2724);
and (n2875,n2859,n2873);
and (n2876,n2877,n2878);
xor (n2877,n2855,n2857);
or (n2878,n2879,n2894);
and (n2879,n2880,n2892);
or (n2880,n2881,n2886,n2891);
and (n2881,n2882,n2883);
xor (n2882,n2860,n2864);
and (n2883,n488,n2884);
xnor (n2884,n2885,n488);
nand (n2885,n1065,n709);
and (n2886,n2883,n2887);
xnor (n2887,n2888,n488);
nor (n2888,n2889,n2890);
and (n2889,n1065,n713);
and (n2890,n1051,n709);
and (n2891,n2882,n2887);
xor (n2892,n2893,n2873);
xor (n2893,n2859,n2868);
and (n2894,n2895,n2896);
xor (n2895,n2880,n2892);
or (n2896,n2897,n2913);
and (n2897,n2898,n2900);
xor (n2898,n2899,n2887);
xor (n2899,n2882,n2883);
or (n2900,n2901,n2907,n2912);
and (n2901,n2902,n2903);
not (n2902,n2885);
xnor (n2903,n2904,n836);
nor (n2904,n2905,n2906);
and (n2905,n1026,n1037);
and (n2906,n1022,n1039);
and (n2907,n2903,n2908);
xnor (n2908,n2909,n711);
nor (n2909,n2910,n2911);
and (n2910,n1051,n838);
and (n2911,n1028,n834);
and (n2912,n2902,n2908);
and (n2913,n2914,n2915);
xor (n2914,n2898,n2900);
or (n2915,n2916,n2927);
and (n2916,n2917,n2919);
xor (n2917,n2918,n2908);
xor (n2918,n2902,n2903);
and (n2919,n2920,n2923);
and (n2920,n711,n2921);
xnor (n2921,n2922,n711);
nand (n2922,n1065,n834);
xnor (n2923,n2924,n836);
nor (n2924,n2925,n2926);
and (n2925,n1028,n1037);
and (n2926,n1026,n1039);
and (n2927,n2928,n2929);
xor (n2928,n2917,n2919);
or (n2929,n2930,n2936);
and (n2930,n2931,n2935);
xnor (n2931,n2932,n711);
nor (n2932,n2933,n2934);
and (n2933,n1065,n838);
and (n2934,n1051,n834);
xor (n2935,n2920,n2923);
and (n2936,n2937,n2938);
xor (n2937,n2931,n2935);
or (n2938,n2939,n2945);
and (n2939,n2940,n2944);
xnor (n2940,n2941,n836);
nor (n2941,n2942,n2943);
and (n2942,n1051,n1037);
and (n2943,n1028,n1039);
not (n2944,n2922);
and (n2945,n2946,n2947);
xor (n2946,n2940,n2944);
and (n2947,n2948,n2952);
xnor (n2948,n2949,n836);
nor (n2949,n2950,n2951);
and (n2950,n1065,n1037);
and (n2951,n1051,n1039);
and (n2952,n2953,n836);
xnor (n2953,n2954,n836);
nand (n2954,n1065,n1039);
not (n2955,n2956);
nand (n2956,n2957,n1977);
nor (n2957,n2958,n1009);
nand (n2958,n2959,n1932);
nor (n2959,n2960,n1904);
nor (n2960,n1687,n1866);
not (n2961,n2962);
nor (n2962,n3,n187);
nand (n2963,n2964,n3002);
not (n2964,n2965);
nor (n2965,n2966,n2998);
xor (n2966,n2967,n2994);
xor (n2967,n2968,n2972);
nand (n2968,n2969,n2970,n2971);
nand (n2969,n215,n89);
nand (n2970,n219,n89);
nand (n2971,n215,n219);
xor (n2972,n2973,n2988);
xor (n2973,n2974,n2978);
nand (n2974,n2975,n2976,n2977);
nand (n2975,n197,n201);
nand (n2976,n205,n201);
nand (n2977,n197,n205);
xor (n2978,n2979,n2984);
xor (n2979,n215,n2980);
xor (n2980,n2981,n56);
or (n2981,n2982,n2983);
and (n2982,n13,n50);
and (n2983,n27,n54);
xor (n2984,n2985,n89);
or (n2985,n2986,n2987);
and (n2986,n49,n83);
and (n2987,n53,n87);
xor (n2988,n2989,n216);
xor (n2989,n2990,n89);
xor (n2990,n2991,n68);
or (n2991,n2992,n2993);
and (n2992,n35,n62);
and (n2993,n39,n66);
nand (n2994,n2995,n2996,n2997);
nand (n2995,n195,n209);
nand (n2996,n213,n209);
nand (n2997,n195,n213);
nand (n2998,n2999,n3000,n3001);
nand (n2999,n189,n193);
nand (n3000,n223,n193);
nand (n3001,n189,n223);
nand (n3002,n2966,n2998);
xor (n3003,n3004,n3262);
xor (n3004,n3005,n3059);
xor (n3005,n3006,n3031);
xor (n3006,n3007,n3016);
xor (n3007,n3008,n3013);
or (n3008,n3009,n3010,n3012);
and (n3009,n216,n195);
and (n3010,n195,n3011);
not (n3011,n210);
and (n3012,n216,n3011);
xor (n3013,n3014,n3015);
xor (n3014,n2984,n2974);
xor (n3015,n2979,n2990);
or (n3016,n3017,n3027,n3030);
and (n3017,n3018,n3022);
or (n3018,n3019,n3020,n3021);
and (n3019,n73,n125);
not (n3020,n221);
and (n3021,n73,n129);
or (n3022,n3023,n3024,n3026);
and (n3023,n124,n107);
and (n3024,n107,n3025);
not (n3025,n94);
and (n3026,n124,n3025);
and (n3027,n3022,n3028);
xor (n3028,n3029,n3011);
xor (n3029,n216,n195);
and (n3030,n3018,n3028);
or (n3031,n3032,n3044,n3058);
and (n3032,n3033,n3042);
or (n3033,n3034,n3039,n3041);
and (n3034,n3035,n100);
or (n3035,n3036,n3037,n3038);
and (n3036,n124,n76);
not (n3037,n120);
and (n3038,n124,n80);
and (n3039,n100,n3040);
not (n3040,n122);
and (n3041,n3035,n3040);
xor (n3042,n3043,n3028);
xor (n3043,n3018,n3022);
and (n3044,n3042,n3045);
or (n3045,n3046,n3054,n3057);
and (n3046,n3047,n3052);
or (n3047,n3048,n3050,n3051);
and (n3048,n3049,n137);
not (n3049,n71);
and (n3050,n137,n7);
and (n3051,n3049,n7);
xor (n3052,n3053,n3025);
xor (n3053,n124,n107);
and (n3054,n3052,n3055);
xor (n3055,n3056,n3040);
xor (n3056,n3035,n100);
and (n3057,n3047,n3055);
and (n3058,n3033,n3045);
or (n3059,n3060,n3148,n3261);
and (n3060,n3061,n3063);
xor (n3061,n3062,n3045);
xor (n3062,n3033,n3042);
or (n3063,n3064,n3085,n3147);
and (n3064,n3065,n3083);
or (n3065,n3066,n3079,n3082);
and (n3066,n3067,n3071);
or (n3067,n3068,n3069,n3070);
not (n3068,n69);
and (n3069,n58,n140);
and (n3070,n46,n140);
or (n3071,n3072,n3077,n3078);
and (n3072,n146,n3073);
or (n3073,n3074,n3075,n3076);
and (n3074,n10,n168);
not (n3075,n167);
and (n3076,n10,n172);
and (n3077,n3073,n179);
and (n3078,n146,n179);
and (n3079,n3071,n3080);
xor (n3080,n3081,n7);
xor (n3081,n3049,n137);
and (n3082,n3067,n3080);
xor (n3083,n3084,n3055);
xor (n3084,n3047,n3052);
and (n3085,n3083,n3086);
or (n3086,n3087,n3100,n3146);
and (n3087,n3088,n3098);
or (n3088,n3089,n3094,n3097);
and (n3089,n3090,n3092);
xor (n3090,n3091,n140);
xor (n3091,n46,n58);
and (n3092,n238,n3093);
not (n3093,n240);
and (n3094,n3092,n3095);
xor (n3095,n3096,n179);
xor (n3096,n146,n3073);
and (n3097,n3090,n3095);
xor (n3098,n3099,n3080);
xor (n3099,n3067,n3071);
and (n3100,n3098,n3101);
or (n3101,n3102,n3115,n3145);
and (n3102,n3103,n3113);
or (n3103,n3104,n3110,n3112);
and (n3104,n3105,n3106);
not (n3105,n243);
or (n3106,n3107,n3108,n3109);
not (n3107,n260);
and (n3108,n271,n282);
and (n3109,n261,n282);
and (n3110,n3106,n3111);
not (n3111,n237);
and (n3112,n3105,n3111);
xor (n3113,n3114,n3095);
xor (n3114,n3090,n3092);
and (n3115,n3113,n3116);
or (n3116,n3117,n3131,n3144);
and (n3117,n3118,n3122);
or (n3118,n3119,n3120,n3121);
and (n3119,n275,n287);
and (n3120,n287,n329);
and (n3121,n275,n329);
or (n3122,n3123,n3128,n3130);
and (n3123,n296,n3124);
or (n3124,n3125,n3126,n3127);
and (n3125,n262,n315);
not (n3126,n319);
and (n3127,n262,n320);
and (n3128,n3124,n3129);
xor (n3129,n295,n282);
and (n3130,n296,n3129);
and (n3131,n3122,n3132);
or (n3132,n3133,n3140,n3143);
and (n3133,n3134,n3135);
not (n3134,n367);
or (n3135,n3136,n3138,n3139);
and (n3136,n335,n3137);
not (n3137,n411);
and (n3138,n3137,n341);
not (n3139,n362);
and (n3140,n3135,n3141);
xor (n3141,n3142,n329);
xor (n3142,n275,n287);
and (n3143,n3134,n3141);
and (n3144,n3118,n3132);
and (n3145,n3103,n3116);
and (n3146,n3088,n3101);
and (n3147,n3065,n3086);
and (n3148,n3063,n3149);
or (n3149,n3150,n3152);
xor (n3150,n3151,n3086);
xor (n3151,n3065,n3083);
or (n3152,n3153,n3155);
xor (n3153,n3154,n3101);
xor (n3154,n3088,n3098);
or (n3155,n3156,n3188,n3260);
and (n3156,n3157,n3186);
or (n3157,n3158,n3182,n3185);
and (n3158,n3159,n3161);
xor (n3159,n3160,n3111);
xor (n3160,n3105,n3106);
or (n3161,n3162,n3178,n3181);
and (n3162,n3163,n3165);
xor (n3163,n3164,n3129);
xor (n3164,n296,n3124);
or (n3165,n3166,n3172,n3177);
and (n3166,n444,n3167);
and (n3167,n3168,n460);
or (n3168,n3169,n3170,n3171);
and (n3169,n344,n449);
not (n3170,n448);
and (n3171,n344,n453);
and (n3172,n3167,n3173);
or (n3173,n3174,n3175,n3176);
not (n3174,n394);
and (n3175,n395,n420);
and (n3176,n390,n420);
and (n3177,n444,n3173);
and (n3178,n3165,n3179);
xor (n3179,n3180,n3141);
xor (n3180,n3134,n3135);
and (n3181,n3163,n3179);
and (n3182,n3161,n3183);
xor (n3183,n3184,n3132);
xor (n3184,n3118,n3122);
and (n3185,n3159,n3183);
xor (n3186,n3187,n3116);
xor (n3187,n3103,n3113);
and (n3188,n3186,n3189);
or (n3189,n3190,n3192);
xor (n3190,n3191,n3183);
xor (n3191,n3159,n3161);
or (n3192,n3193,n3224,n3259);
and (n3193,n3194,n3222);
or (n3194,n3195,n3204,n3221);
and (n3195,n3196,n3198);
xor (n3196,n3197,n341);
xor (n3197,n335,n3137);
or (n3198,n3199,n3201,n3203);
and (n3199,n3200,n417);
not (n3200,n470);
and (n3201,n417,n3202);
xor (n3202,n3168,n460);
and (n3203,n3200,n3202);
and (n3204,n3198,n3205);
or (n3205,n3206,n3217,n3220);
and (n3206,n3207,n3212);
or (n3207,n3208,n3210,n3211);
and (n3208,n504,n3209);
not (n3209,n909);
and (n3210,n3209,n908);
and (n3211,n504,n908);
or (n3212,n3213,n3215,n3216);
and (n3213,n507,n3214);
not (n3214,n904);
and (n3215,n3214,n480);
and (n3216,n507,n480);
and (n3217,n3212,n3218);
xor (n3218,n3219,n420);
xor (n3219,n390,n395);
and (n3220,n3207,n3218);
and (n3221,n3196,n3205);
xor (n3222,n3223,n3179);
xor (n3223,n3163,n3165);
and (n3224,n3222,n3225);
or (n3225,n3226,n3255,n3258);
and (n3226,n3227,n3229);
xor (n3227,n3228,n3173);
xor (n3228,n444,n3167);
or (n3229,n3230,n3251,n3254);
and (n3230,n3231,n3249);
or (n3231,n3232,n3245,n3248);
and (n3232,n3233,n3237);
or (n3233,n3234,n3235,n3236);
and (n3234,n588,n662);
and (n3235,n662,n731);
and (n3236,n588,n731);
or (n3237,n3238,n3239,n3244);
and (n3238,n592,n664);
and (n3239,n664,n3240);
or (n3240,n3241,n3242,n3243);
and (n3241,n483,n693);
not (n3242,n729);
and (n3243,n483,n689);
and (n3244,n592,n3240);
and (n3245,n3237,n3246);
xor (n3246,n3247,n908);
xor (n3247,n504,n3209);
and (n3248,n3233,n3246);
xor (n3249,n3250,n3202);
xor (n3250,n3200,n417);
and (n3251,n3249,n3252);
xor (n3252,n3253,n3218);
xor (n3253,n3207,n3212);
and (n3254,n3231,n3252);
and (n3255,n3229,n3256);
xor (n3256,n3257,n3205);
xor (n3257,n3196,n3198);
and (n3258,n3227,n3256);
and (n3259,n3194,n3225);
and (n3260,n3157,n3189);
and (n3261,n3061,n3149);
and (n3262,n3263,n3265);
xor (n3263,n3264,n3149);
xor (n3264,n3061,n3063);
and (n3265,n3266,n3267);
xnor (n3266,n3150,n3152);
and (n3267,n3268,n3269);
xnor (n3268,n3153,n3155);
and (n3269,n3270,n3272);
xor (n3270,n3271,n3189);
xor (n3271,n3157,n3186);
and (n3272,n3273,n3274);
xnor (n3273,n3190,n3192);
or (n3274,n3275,n3355);
and (n3275,n3276,n3278);
xor (n3276,n3277,n3225);
xor (n3277,n3194,n3222);
or (n3278,n3279,n3281);
xor (n3279,n3280,n3256);
xor (n3280,n3227,n3229);
or (n3281,n3282,n3305,n3354);
and (n3282,n3283,n3303);
or (n3283,n3284,n3299,n3302);
and (n3284,n3285,n3287);
xor (n3285,n3286,n480);
xor (n3286,n507,n3214);
or (n3287,n3288,n3295,n3298);
and (n3288,n660,n3289);
or (n3289,n3290,n3292,n3294);
and (n3290,n721,n3291);
not (n3291,n687);
and (n3292,n3291,n3293);
not (n3293,n673);
and (n3294,n721,n3293);
and (n3295,n3289,n3296);
xor (n3296,n3297,n731);
xor (n3297,n588,n662);
and (n3298,n660,n3296);
and (n3299,n3287,n3300);
xor (n3300,n3301,n3246);
xor (n3301,n3233,n3237);
and (n3302,n3285,n3300);
xor (n3303,n3304,n3252);
xor (n3304,n3231,n3249);
and (n3305,n3303,n3306);
or (n3306,n3307,n3318,n3353);
and (n3307,n3308,n3316);
or (n3308,n3309,n3312,n3315);
and (n3309,n3310,n608);
xor (n3310,n3311,n3240);
xor (n3311,n592,n664);
and (n3312,n608,n3313);
xor (n3313,n3314,n3296);
xor (n3314,n660,n3289);
and (n3315,n3310,n3313);
xor (n3316,n3317,n3300);
xor (n3317,n3285,n3287);
and (n3318,n3316,n3319);
or (n3319,n3320,n3349,n3352);
and (n3320,n3321,n3334);
or (n3321,n3322,n3332,n3333);
and (n3322,n3323,n766);
or (n3323,n3324,n3329,n3331);
and (n3324,n3325,n760);
or (n3325,n3326,n3327,n3328);
and (n3326,n705,n750);
not (n3327,n754);
and (n3328,n705,n755);
and (n3329,n760,n3330);
not (n3330,n763);
and (n3331,n3325,n3330);
not (n3332,n801);
and (n3333,n3323,n802);
or (n3334,n3335,n3342,n3348);
and (n3335,n3336,n3340);
or (n3336,n3337,n3338,n3339);
and (n3337,n706,n702);
not (n3338,n720);
and (n3339,n706,n716);
xor (n3340,n3341,n3293);
xor (n3341,n721,n3291);
and (n3342,n3340,n3343);
or (n3343,n3344,n3345,n3347);
and (n3344,n705,n843);
and (n3345,n843,n3346);
not (n3346,n2457);
and (n3347,n705,n3346);
and (n3348,n3336,n3343);
and (n3349,n3334,n3350);
xor (n3350,n3351,n3313);
xor (n3351,n3310,n608);
and (n3352,n3321,n3350);
and (n3353,n3308,n3319);
and (n3354,n3283,n3306);
and (n3355,n3356,n3357);
xor (n3356,n3276,n3278);
and (n3357,n3358,n3359);
xnor (n3358,n3279,n3281);
or (n3359,n3360,n3445);
and (n3360,n3361,n3363);
xor (n3361,n3362,n3306);
xor (n3362,n3283,n3303);
or (n3363,n3364,n3366);
xor (n3364,n3365,n3319);
xor (n3365,n3308,n3316);
or (n3366,n3367,n3389,n3444);
and (n3367,n3368,n3387);
or (n3368,n3369,n3383,n3386);
and (n3369,n3370,n3372);
xor (n3370,n3371,n802);
xor (n3371,n3323,n766);
or (n3372,n3373,n3376,n3382);
and (n3373,n3374,n2460);
xor (n3374,n3375,n3330);
xor (n3375,n3325,n760);
and (n3376,n2460,n3377);
or (n3377,n3378,n3379,n3381);
not (n3378,n882);
and (n3379,n866,n3380);
not (n3380,n863);
and (n3381,n847,n3380);
and (n3382,n3374,n3377);
and (n3383,n3372,n3384);
xor (n3384,n3385,n3343);
xor (n3385,n3336,n3340);
and (n3386,n3370,n3384);
xor (n3387,n3388,n3350);
xor (n3388,n3321,n3334);
and (n3389,n3387,n3390);
or (n3390,n3391,n3406,n3443);
and (n3391,n3392,n3404);
or (n3392,n3393,n3400,n3403);
and (n3393,n3394,n3398);
or (n3394,n3395,n3396,n3397);
and (n3395,n814,n2430);
and (n3396,n2430,n2411);
and (n3397,n814,n2411);
xor (n3398,n3399,n3346);
xor (n3399,n705,n843);
and (n3400,n3398,n3401);
and (n3401,n2406,n3402);
not (n3402,n2404);
and (n3403,n3394,n3401);
xor (n3404,n3405,n3384);
xor (n3405,n3370,n3372);
and (n3406,n3404,n3407);
or (n3407,n3408,n3428,n3442);
and (n3408,n3409,n3426);
or (n3409,n3410,n3415,n3425);
and (n3410,n3411,n2433);
or (n3411,n3412,n3413,n3414);
and (n3412,n831,n822);
not (n3413,n821);
and (n3414,n831,n825);
and (n3415,n2433,n3416);
or (n3416,n3417,n3422,n3424);
and (n3417,n830,n3418);
or (n3418,n3419,n3420,n3421);
and (n3419,n830,n2234);
not (n3420,n2348);
and (n3421,n830,n2238);
and (n3422,n3418,n3423);
not (n3423,n2343);
and (n3424,n830,n3423);
and (n3425,n3411,n3416);
xor (n3426,n3427,n3377);
xor (n3427,n3374,n2460);
and (n3428,n3426,n3429);
or (n3429,n3430,n3434,n3441);
and (n3430,n3431,n3433);
xor (n3431,n3432,n2411);
xor (n3432,n814,n2430);
not (n3433,n2403);
and (n3434,n3433,n3435);
or (n3435,n3436,n3439,n3440);
and (n3436,n3437,n2349);
and (n3437,n2218,n3438);
not (n3438,n2232);
and (n3439,n2349,n2371);
and (n3440,n3437,n2371);
and (n3441,n3431,n3435);
and (n3442,n3409,n3429);
and (n3443,n3392,n3407);
and (n3444,n3368,n3390);
and (n3445,n3446,n3447);
xor (n3446,n3361,n3363);
and (n3447,n3448,n3449);
xnor (n3448,n3364,n3366);
or (n3449,n3450,n3654);
and (n3450,n3451,n3453);
xor (n3451,n3452,n3390);
xor (n3452,n3368,n3387);
or (n3453,n3454,n3529,n3653);
and (n3454,n3455,n3527);
or (n3455,n3456,n3523,n3526);
and (n3456,n3457,n3459);
xor (n3457,n3458,n3401);
xor (n3458,n3394,n3398);
or (n3459,n3460,n3494,n3522);
and (n3460,n3461,n3492);
or (n3461,n3462,n3480,n3491);
and (n3462,n3463,n3472);
and (n3463,n3464,n2258);
or (n3464,n3465,n3470,n3471);
and (n3465,n3466,n2128);
or (n3466,n3467,n3468,n3469);
and (n3467,n2197,n1993);
not (n3468,n2137);
and (n3469,n2197,n1997);
not (n3470,n2270);
and (n3471,n3466,n2132);
or (n3472,n3473,n3478,n3479);
and (n3473,n2298,n3474);
or (n3474,n3475,n3476,n3477);
and (n3475,n2197,n2117);
not (n3476,n2245);
and (n3477,n2197,n2122);
and (n3478,n3474,n2279);
and (n3479,n2298,n2279);
and (n3480,n3472,n3481);
or (n3481,n3482,n3488,n3490);
and (n3482,n3483,n3484);
not (n3483,n2217);
or (n3484,n3485,n3486,n3487);
and (n3485,n2001,n2193);
not (n3486,n2297);
and (n3487,n2001,n2198);
and (n3488,n3484,n3489);
not (n3489,n2274);
and (n3490,n3483,n3489);
and (n3491,n3463,n3481);
xor (n3492,n3493,n3416);
xor (n3493,n3411,n2433);
and (n3494,n3492,n3495);
or (n3495,n3496,n3518,n3521);
and (n3496,n3497,n3499);
xor (n3497,n3498,n3423);
xor (n3498,n830,n3418);
or (n3499,n3500,n3509,n3517);
and (n3500,n3501,n3508);
or (n3501,n3502,n3504,n3507);
and (n3502,n2177,n3503);
not (n3503,n2174);
and (n3504,n3503,n3505);
xor (n3505,n3506,n2122);
xor (n3506,n2197,n2117);
and (n3507,n2177,n3505);
xor (n3508,n3464,n2258);
and (n3509,n3508,n3510);
or (n3510,n3511,n3515,n3516);
and (n3511,n3512,n3513);
not (n3512,n2191);
xor (n3513,n3514,n2132);
xor (n3514,n3466,n2128);
and (n3515,n3513,n2151);
and (n3516,n3512,n2151);
and (n3517,n3501,n3510);
and (n3518,n3499,n3519);
xor (n3519,n3520,n2371);
xor (n3520,n3437,n2349);
and (n3521,n3497,n3519);
and (n3522,n3461,n3495);
and (n3523,n3459,n3524);
xor (n3524,n3525,n3429);
xor (n3525,n3409,n3426);
and (n3526,n3457,n3524);
xor (n3527,n3528,n3407);
xor (n3528,n3392,n3404);
and (n3529,n3527,n3530);
or (n3530,n3531,n3564,n3652);
and (n3531,n3532,n3562);
or (n3532,n3533,n3558,n3561);
and (n3533,n3534,n3536);
xor (n3534,n3535,n3435);
xor (n3535,n3431,n3433);
or (n3536,n3537,n3554,n3557);
and (n3537,n3538,n3540);
xor (n3538,n3539,n3481);
xor (n3539,n3463,n3472);
or (n3540,n3541,n3546,n3553);
and (n3541,n3542,n3544);
xor (n3542,n3543,n2279);
xor (n3543,n2298,n3474);
xor (n3544,n3545,n3489);
xor (n3545,n3483,n3484);
and (n3546,n3544,n3547);
and (n3547,n2142,n3548);
or (n3548,n3549,n3550,n3552);
not (n3549,n2148);
and (n3550,n2008,n3551);
not (n3551,n1991);
and (n3552,n2004,n3551);
and (n3553,n3542,n3547);
and (n3554,n3540,n3555);
xor (n3555,n3556,n3519);
xor (n3556,n3497,n3499);
and (n3557,n3538,n3555);
and (n3558,n3536,n3559);
xor (n3559,n3560,n3495);
xor (n3560,n3461,n3492);
and (n3561,n3534,n3559);
xor (n3562,n3563,n3524);
xor (n3563,n3457,n3459);
and (n3564,n3562,n3565);
or (n3565,n3566,n3623,n3651);
and (n3566,n3567,n3569);
xor (n3567,n3568,n3559);
xor (n3568,n3534,n3536);
or (n3569,n3570,n3602,n3622);
and (n3570,n3571,n3600);
or (n3571,n3572,n3585,n3599);
and (n3572,n3573,n3583);
or (n3573,n3574,n3581,n3582);
and (n3574,n3575,n3579);
or (n3575,n3576,n3577,n3578);
and (n3576,n2056,n2041);
and (n3577,n2041,n2024);
and (n3578,n2056,n2024);
xor (n3579,n3580,n3505);
xor (n3580,n2177,n3503);
and (n3581,n3579,n2202);
and (n3582,n3575,n2202);
xor (n3583,n3584,n3510);
xor (n3584,n3501,n3508);
and (n3585,n3583,n3586);
or (n3586,n3587,n3596,n3598);
and (n3587,n3588,n3594);
or (n3588,n3589,n3590,n3593);
and (n3589,n2046,n2040);
and (n3590,n2040,n3591);
xor (n3591,n3592,n2024);
xor (n3592,n2056,n2041);
and (n3593,n2046,n3591);
xor (n3594,n3595,n2151);
xor (n3595,n3512,n3513);
and (n3596,n3594,n3597);
xor (n3597,n2142,n3548);
and (n3598,n3588,n3597);
and (n3599,n3573,n3586);
xor (n3600,n3601,n3555);
xor (n3601,n3538,n3540);
and (n3602,n3600,n3603);
or (n3603,n3604,n3618,n3621);
and (n3604,n3605,n3607);
xor (n3605,n3606,n3547);
xor (n3606,n3542,n3544);
or (n3607,n3608,n3616,n3617);
and (n3608,n3609,n3611);
xor (n3609,n3610,n2202);
xor (n3610,n3575,n3579);
or (n3611,n3612,n3613,n3615);
not (n3612,n2101);
and (n3613,n2016,n3614);
not (n3614,n1989);
and (n3615,n2012,n3614);
and (n3616,n3611,n2103);
and (n3617,n3609,n2103);
and (n3618,n3607,n3619);
xor (n3619,n3620,n3586);
xor (n3620,n3573,n3583);
and (n3621,n3605,n3619);
and (n3622,n3571,n3603);
and (n3623,n3569,n3624);
or (n3624,n3625,n3627);
xor (n3625,n3626,n3603);
xor (n3626,n3571,n3600);
or (n3627,n3628,n3644,n3650);
and (n3628,n3629,n3642);
or (n3629,n3630,n3638,n3641);
and (n3630,n3631,n3633);
xor (n3631,n3632,n3597);
xor (n3632,n3588,n3594);
or (n3633,n3634,n3636,n3637);
and (n3634,n3635,n2088);
not (n3635,n1987);
not (n3636,n2095);
and (n3637,n3635,n2020);
and (n3638,n3633,n3639);
xor (n3639,n3640,n2103);
xor (n3640,n3609,n3611);
and (n3641,n3631,n3639);
xor (n3642,n3643,n3619);
xor (n3643,n3605,n3607);
and (n3644,n3642,n3645);
or (n3645,n3646,n3648);
or (n3646,n1981,n3647);
not (n3647,n1985);
xor (n3648,n3649,n3639);
xor (n3649,n3631,n3633);
and (n3650,n3629,n3645);
and (n3651,n3567,n3624);
and (n3652,n3532,n3565);
and (n3653,n3455,n3530);
and (n3654,n3655,n3656);
xor (n3655,n3451,n3453);
and (n3656,n3657,n3659);
xor (n3657,n3658,n3530);
xor (n3658,n3455,n3527);
or (n3659,n3660,n3662);
xor (n3660,n3661,n3565);
xor (n3661,n3532,n3562);
and (n3662,n3663,n3664);
not (n3663,n3660);
and (n3664,n3665,n3667);
xor (n3665,n3666,n3624);
xor (n3666,n3567,n3569);
and (n3667,n3668,n3669);
xnor (n3668,n3625,n3627);
and (n3669,n3670,n3672);
xor (n3670,n3671,n3645);
xor (n3671,n3629,n3642);
and (n3672,n3673,n3674);
xnor (n3673,n3646,n3648);
and (n3674,n3675,n3678);
not (n3675,n3676);
nand (n3676,n3677,n2510);
not (n3677,n1980);
nand (n3678,n1007,n3679);
nand (n3679,n2957,n2536);
endmodule
