module top (out,n16,n17,n22,n27,n35,n40,n45,n52,n63
        ,n65,n71,n77,n83,n92,n97,n102,n108,n115,n123
        ,n129,n163,n168,n173,n181,n189,n208,n273,n341,n421
        ,n468,n498);
output out;
input n16;
input n17;
input n22;
input n27;
input n35;
input n40;
input n45;
input n52;
input n63;
input n65;
input n71;
input n77;
input n83;
input n92;
input n97;
input n102;
input n108;
input n115;
input n123;
input n129;
input n163;
input n168;
input n173;
input n181;
input n189;
input n208;
input n273;
input n341;
input n421;
input n468;
input n498;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
xor (out,n0,n1064);
nand (n0,n1,n1063);
or (n1,n2,n392);
not (n2,n3);
nand (n3,n4,n390);
not (n4,n5);
nor (n5,n6,n321);
xor (n6,n7,n256);
xor (n7,n8,n154);
xor (n8,n9,n133);
xor (n9,n10,n55);
and (n10,n11,n29);
nand (n11,n12,n23);
or (n12,n13,n20);
nor (n13,n14,n18);
and (n14,n15,n17);
not (n15,n16);
and (n18,n16,n19);
not (n19,n17);
nand (n20,n16,n21);
not (n21,n22);
or (n23,n24,n21);
nor (n24,n25,n28);
and (n25,n26,n16);
not (n26,n27);
and (n28,n27,n15);
nand (n29,n30,n48);
or (n30,n31,n43);
not (n31,n32);
nor (n32,n33,n37);
nand (n33,n34,n36);
or (n34,n15,n35);
nand (n36,n15,n35);
nor (n37,n38,n41);
and (n38,n39,n35);
not (n39,n40);
and (n41,n40,n42);
not (n42,n35);
nor (n43,n44,n46);
and (n44,n39,n45);
and (n46,n40,n47);
not (n47,n45);
or (n48,n49,n50);
not (n49,n33);
nor (n50,n51,n53);
and (n51,n39,n52);
and (n53,n40,n54);
not (n54,n52);
or (n55,n56,n132);
and (n56,n57,n110);
xor (n57,n58,n85);
nand (n58,n59,n79);
or (n59,n60,n68);
not (n60,n61);
nand (n61,n62,n66);
or (n62,n63,n64);
not (n64,n65);
or (n66,n67,n65);
not (n67,n63);
nand (n68,n69,n73);
nand (n69,n70,n72);
or (n70,n71,n67);
nand (n72,n67,n71);
not (n73,n74);
nand (n74,n75,n78);
or (n75,n76,n71);
not (n76,n77);
nand (n78,n76,n71);
nand (n79,n74,n80);
nor (n80,n81,n84);
and (n81,n82,n67);
not (n82,n83);
and (n84,n63,n83);
nand (n85,n86,n104);
or (n86,n87,n99);
not (n87,n88);
and (n88,n89,n94);
not (n89,n90);
nand (n90,n91,n93);
or (n91,n92,n67);
nand (n93,n92,n67);
nand (n94,n95,n98);
or (n95,n92,n96);
not (n96,n97);
nand (n98,n96,n92);
nor (n99,n100,n103);
and (n100,n101,n97);
not (n101,n102);
and (n103,n102,n96);
or (n104,n89,n105);
nor (n105,n106,n109);
and (n106,n107,n97);
not (n107,n108);
and (n109,n108,n96);
nand (n110,n111,n126);
or (n111,n112,n121);
nand (n112,n113,n118);
nor (n113,n114,n116);
and (n114,n39,n115);
and (n116,n40,n117);
not (n117,n115);
nand (n118,n119,n120);
or (n119,n115,n76);
nand (n120,n76,n115);
nor (n121,n122,n124);
and (n122,n76,n123);
and (n124,n77,n125);
not (n125,n123);
or (n126,n113,n127);
nor (n127,n128,n130);
and (n128,n76,n129);
and (n130,n77,n131);
not (n131,n129);
and (n132,n58,n85);
xor (n133,n134,n148);
xor (n134,n135,n142);
nand (n135,n136,n138);
or (n136,n137,n68);
not (n137,n80);
nand (n138,n74,n139);
nor (n139,n140,n141);
and (n140,n125,n67);
and (n141,n63,n123);
nand (n142,n143,n144);
or (n143,n87,n105);
or (n144,n89,n145);
nor (n145,n146,n147);
and (n146,n65,n96);
and (n147,n64,n97);
nand (n148,n149,n150);
or (n149,n112,n127);
or (n150,n113,n151);
nor (n151,n152,n153);
and (n152,n76,n45);
and (n153,n77,n47);
xor (n154,n155,n211);
xor (n155,n156,n197);
xor (n156,n157,n182);
xor (n157,n158,n180);
nand (n158,n159,n176);
or (n159,n160,n170);
nand (n160,n161,n166);
nor (n161,n162,n164);
and (n162,n96,n163);
and (n164,n97,n165);
not (n165,n163);
nand (n166,n167,n169);
or (n167,n165,n168);
nand (n169,n165,n168);
nor (n170,n171,n174);
and (n171,n172,n173);
not (n172,n168);
and (n174,n168,n175);
not (n175,n173);
or (n176,n161,n177);
nor (n177,n178,n179);
and (n178,n172,n102);
and (n179,n168,n101);
and (n180,n168,n181);
xor (n182,n183,n191);
nand (n183,n184,n185);
or (n184,n20,n24);
or (n185,n186,n21);
nor (n186,n187,n190);
and (n187,n188,n16);
not (n188,n189);
and (n190,n189,n15);
nand (n191,n192,n193);
or (n192,n31,n50);
or (n193,n49,n194);
nor (n194,n195,n196);
and (n195,n39,n17);
and (n196,n40,n19);
or (n197,n198,n210);
and (n198,n199,n209);
xor (n199,n200,n207);
nand (n200,n201,n206);
or (n201,n160,n202);
nor (n202,n203,n204);
and (n203,n172,n181);
and (n204,n168,n205);
not (n205,n181);
or (n206,n161,n170);
and (n207,n168,n208);
xor (n209,n11,n29);
and (n210,n200,n207);
or (n211,n212,n255);
and (n212,n213,n254);
xor (n213,n214,n230);
and (n214,n215,n222);
nand (n215,n216,n221);
or (n216,n217,n20);
not (n217,n218);
nor (n218,n219,n220);
and (n219,n54,n15);
and (n220,n16,n52);
or (n221,n13,n21);
nand (n222,n223,n228);
or (n223,n224,n31);
not (n224,n225);
nor (n225,n226,n227);
and (n226,n40,n129);
and (n227,n131,n39);
nand (n228,n229,n33);
not (n229,n43);
or (n230,n231,n253);
and (n231,n232,n247);
xor (n232,n233,n240);
nand (n233,n234,n239);
or (n234,n235,n68);
not (n235,n236);
nor (n236,n237,n238);
and (n237,n63,n108);
and (n238,n107,n67);
nand (n239,n74,n61);
nand (n240,n241,n246);
or (n241,n242,n87);
not (n242,n243);
nand (n243,n244,n245);
or (n244,n97,n175);
or (n245,n96,n173);
or (n246,n89,n99);
nand (n247,n248,n252);
or (n248,n112,n249);
nor (n249,n250,n251);
and (n250,n76,n83);
and (n251,n77,n82);
or (n252,n113,n121);
and (n253,n233,n240);
xor (n254,n57,n110);
and (n255,n214,n230);
or (n256,n257,n320);
and (n257,n258,n276);
xor (n258,n259,n260);
xor (n259,n199,n209);
or (n260,n261,n275);
and (n261,n262,n274);
xor (n262,n263,n272);
nand (n263,n264,n269);
or (n264,n265,n160);
nor (n265,n266,n267);
and (n266,n208,n172);
and (n267,n268,n168);
not (n268,n208);
nand (n269,n270,n271);
not (n270,n202);
not (n271,n161);
and (n272,n168,n273);
xor (n274,n215,n222);
and (n275,n263,n272);
or (n276,n277,n319);
and (n277,n278,n318);
xor (n278,n279,n294);
and (n279,n280,n287);
nand (n280,n281,n282);
or (n281,n21,n217);
nand (n282,n283,n286);
nand (n283,n284,n285);
or (n284,n45,n15);
nand (n285,n15,n45);
not (n286,n20);
nand (n287,n288,n293);
or (n288,n289,n31);
not (n289,n290);
nand (n290,n291,n292);
or (n291,n40,n125);
or (n292,n39,n123);
nand (n293,n33,n225);
or (n294,n295,n317);
and (n295,n296,n311);
xor (n296,n297,n304);
nand (n297,n298,n303);
or (n298,n299,n68);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n101,n67);
and (n302,n63,n102);
nand (n303,n236,n74);
nand (n304,n305,n310);
or (n305,n306,n87);
not (n306,n307);
nand (n307,n308,n309);
or (n308,n97,n205);
or (n309,n96,n181);
nand (n310,n90,n243);
nand (n311,n312,n316);
or (n312,n112,n313);
nor (n313,n314,n315);
and (n314,n76,n65);
and (n315,n77,n64);
or (n316,n249,n113);
and (n317,n297,n304);
xor (n318,n232,n247);
and (n319,n279,n294);
and (n320,n259,n260);
or (n321,n322,n389);
and (n322,n323,n326);
xor (n323,n324,n325);
xor (n324,n213,n254);
xor (n325,n258,n276);
or (n326,n327,n388);
and (n327,n328,n344);
xor (n328,n329,n330);
xor (n329,n262,n274);
or (n330,n331,n343);
and (n331,n332,n342);
xor (n332,n333,n340);
nand (n333,n334,n339);
or (n334,n160,n335);
nor (n335,n336,n337);
and (n336,n273,n172);
and (n337,n338,n168);
not (n338,n273);
or (n339,n161,n265);
and (n340,n168,n341);
xor (n342,n280,n287);
and (n343,n333,n340);
or (n344,n345,n387);
and (n345,n346,n386);
xor (n346,n347,n362);
and (n347,n348,n355);
nand (n348,n349,n353);
or (n349,n350,n20);
nor (n350,n351,n352);
and (n351,n131,n16);
and (n352,n129,n15);
or (n353,n354,n21);
not (n354,n283);
nand (n355,n356,n361);
or (n356,n357,n31);
not (n357,n358);
nor (n358,n359,n360);
and (n359,n40,n83);
and (n360,n82,n39);
nand (n361,n33,n290);
or (n362,n363,n385);
and (n363,n364,n378);
xor (n364,n365,n372);
nand (n365,n366,n371);
or (n366,n367,n68);
not (n367,n368);
nor (n368,n369,n370);
and (n369,n175,n67);
and (n370,n63,n173);
nand (n371,n300,n74);
nand (n372,n373,n377);
or (n373,n87,n374);
nor (n374,n375,n376);
and (n375,n96,n208);
and (n376,n97,n268);
nand (n377,n90,n307);
nand (n378,n379,n384);
or (n379,n380,n112);
not (n380,n381);
nor (n381,n382,n383);
and (n382,n107,n76);
and (n383,n77,n108);
or (n384,n113,n313);
and (n385,n365,n372);
xor (n386,n296,n311);
and (n387,n347,n362);
and (n388,n329,n330);
and (n389,n324,n325);
not (n390,n391);
and (n391,n6,n321);
not (n392,n393);
nand (n393,n394,n1057);
or (n394,n395,n540);
not (n395,n396);
nor (n396,n397,n473);
not (n397,n398);
nand (n398,n399,n401);
not (n399,n400);
xor (n400,n323,n326);
not (n401,n402);
or (n402,n403,n472);
and (n403,n404,n471);
xor (n404,n405,n406);
xor (n405,n278,n318);
or (n406,n407,n470);
and (n407,n408,n424);
xor (n408,n409,n410);
xor (n409,n332,n342);
or (n410,n411,n423);
and (n411,n412,n422);
xor (n412,n413,n420);
nand (n413,n414,n419);
or (n414,n415,n160);
nor (n415,n416,n417);
and (n416,n172,n341);
and (n417,n168,n418);
not (n418,n341);
or (n419,n161,n335);
and (n420,n168,n421);
xor (n422,n348,n355);
and (n423,n413,n420);
and (n424,n425,n449);
or (n425,n426,n448);
and (n426,n427,n442);
xor (n427,n428,n435);
nand (n428,n429,n434);
or (n429,n430,n31);
not (n430,n431);
nor (n431,n432,n433);
and (n432,n64,n39);
and (n433,n40,n65);
nand (n434,n33,n358);
nand (n435,n436,n441);
or (n436,n437,n68);
not (n437,n438);
nor (n438,n439,n440);
and (n439,n205,n67);
and (n440,n63,n181);
nand (n441,n74,n368);
nand (n442,n443,n447);
or (n443,n87,n444);
nor (n444,n445,n446);
and (n445,n96,n273);
and (n446,n97,n338);
or (n447,n89,n374);
and (n448,n428,n435);
or (n449,n450,n469);
and (n450,n451,n467);
xor (n451,n452,n460);
nand (n452,n453,n458);
or (n453,n454,n112);
not (n454,n455);
nand (n455,n456,n457);
or (n456,n77,n101);
or (n457,n76,n102);
nand (n458,n381,n459);
not (n459,n113);
nand (n460,n461,n466);
or (n461,n160,n462);
nor (n462,n463,n464);
and (n463,n172,n421);
and (n464,n465,n168);
not (n465,n421);
or (n466,n161,n415);
and (n467,n168,n468);
and (n469,n452,n460);
and (n470,n409,n410);
xor (n471,n328,n344);
and (n472,n405,n406);
nor (n473,n474,n475);
xor (n474,n404,n471);
or (n475,n476,n539);
and (n476,n477,n480);
xor (n477,n478,n479);
xor (n478,n346,n386);
xor (n479,n408,n424);
or (n480,n481,n538);
and (n481,n482,n485);
xor (n482,n483,n484);
xor (n483,n364,n378);
xor (n484,n412,n422);
or (n485,n486,n537);
and (n486,n487,n513);
xor (n487,n488,n494);
nand (n488,n489,n493);
or (n489,n490,n20);
nor (n490,n491,n492);
and (n491,n125,n16);
and (n492,n123,n15);
or (n493,n350,n21);
or (n494,n495,n512);
and (n495,n496,n506);
xor (n496,n497,n499);
and (n497,n168,n498);
nand (n499,n500,n505);
or (n500,n501,n31);
not (n501,n502);
nand (n502,n503,n504);
or (n503,n40,n107);
or (n504,n39,n108);
nand (n505,n431,n33);
nand (n506,n507,n508);
or (n507,n437,n73);
or (n508,n68,n509);
nor (n509,n510,n511);
and (n510,n67,n208);
and (n511,n63,n268);
and (n512,n497,n499);
or (n513,n514,n536);
and (n514,n515,n528);
xor (n515,n516,n522);
nand (n516,n517,n521);
or (n517,n87,n518);
nor (n518,n519,n520);
and (n519,n96,n341);
and (n520,n97,n418);
or (n521,n89,n444);
nand (n522,n523,n527);
or (n523,n524,n20);
nor (n524,n525,n526);
and (n525,n82,n16);
and (n526,n83,n15);
or (n527,n490,n21);
nand (n528,n529,n534);
or (n529,n530,n160);
nor (n530,n531,n532);
and (n531,n468,n172);
and (n532,n533,n168);
not (n533,n468);
nand (n534,n535,n271);
not (n535,n462);
and (n536,n516,n522);
and (n537,n488,n494);
and (n538,n483,n484);
and (n539,n478,n479);
not (n540,n541);
nand (n541,n542,n767);
nor (n542,n543,n762);
and (n543,n544,n650);
and (n544,n545,n614);
nand (n545,n546,n548);
not (n546,n547);
xor (n547,n477,n480);
not (n548,n549);
or (n549,n550,n613);
and (n550,n551,n557);
xor (n551,n552,n556);
nand (n552,n553,n555);
or (n553,n449,n554);
not (n554,n425);
nand (n555,n554,n449);
xor (n556,n482,n485);
or (n557,n558,n612);
and (n558,n559,n562);
xor (n559,n560,n561);
xor (n560,n451,n467);
xor (n561,n427,n442);
or (n562,n563,n611);
and (n563,n564,n586);
xor (n564,n565,n571);
nand (n565,n566,n570);
or (n566,n112,n567);
nor (n567,n568,n569);
and (n568,n76,n173);
and (n569,n77,n175);
or (n570,n113,n454);
nor (n571,n572,n580);
not (n572,n573);
nand (n573,n574,n579);
or (n574,n575,n31);
not (n575,n576);
nor (n576,n577,n578);
and (n577,n101,n39);
and (n578,n40,n102);
nand (n579,n33,n502);
nand (n580,n581,n168);
nand (n581,n582,n583);
or (n582,n97,n163);
nand (n583,n584,n585);
or (n584,n165,n96);
not (n585,n498);
or (n586,n587,n610);
and (n587,n588,n604);
xor (n588,n589,n597);
nand (n589,n590,n595);
or (n590,n591,n68);
not (n591,n592);
nand (n592,n593,n594);
or (n593,n63,n338);
or (n594,n67,n273);
nand (n595,n596,n74);
not (n596,n509);
nand (n597,n598,n603);
or (n598,n599,n87);
not (n599,n600);
nand (n600,n601,n602);
or (n601,n97,n465);
or (n602,n96,n421);
or (n603,n89,n518);
nand (n604,n605,n609);
or (n605,n606,n20);
nor (n606,n607,n608);
and (n607,n15,n65);
and (n608,n16,n64);
or (n609,n524,n21);
and (n610,n589,n597);
and (n611,n565,n571);
and (n612,n560,n561);
and (n613,n552,n556);
nand (n614,n615,n617);
not (n615,n616);
xor (n616,n551,n557);
not (n617,n618);
or (n618,n619,n649);
and (n619,n620,n648);
xor (n620,n621,n622);
xor (n621,n487,n513);
or (n622,n623,n647);
and (n623,n624,n627);
xor (n624,n625,n626);
xor (n625,n515,n528);
xor (n626,n496,n506);
or (n627,n628,n646);
and (n628,n629,n642);
xor (n629,n630,n636);
nand (n630,n631,n635);
or (n631,n160,n632);
nor (n632,n633,n634);
and (n633,n172,n498);
and (n634,n585,n168);
or (n635,n161,n530);
nand (n636,n637,n641);
or (n637,n112,n638);
nor (n638,n639,n640);
and (n639,n76,n181);
and (n640,n77,n205);
or (n641,n113,n567);
nand (n642,n643,n645);
or (n643,n644,n572);
not (n644,n580);
or (n645,n573,n580);
and (n646,n630,n636);
and (n647,n625,n626);
xor (n648,n559,n562);
and (n649,n621,n622);
not (n650,n651);
nand (n651,n652,n759);
or (n652,n653,n753);
not (n653,n654);
nand (n654,n655,n706);
xor (n655,n656,n705);
xor (n656,n657,n658);
xor (n657,n564,n586);
or (n658,n659,n704);
and (n659,n660,n703);
xor (n660,n661,n680);
or (n661,n662,n679);
and (n662,n663,n672);
xor (n663,n664,n665);
and (n664,n271,n498);
nand (n665,n666,n671);
or (n666,n667,n31);
not (n667,n668);
nand (n668,n669,n670);
or (n669,n40,n175);
or (n670,n39,n173);
nand (n671,n33,n576);
nand (n672,n673,n678);
or (n673,n674,n68);
not (n674,n675);
nor (n675,n676,n677);
and (n676,n418,n67);
and (n677,n63,n341);
nand (n678,n74,n592);
and (n679,n664,n665);
or (n680,n681,n702);
and (n681,n682,n696);
xor (n682,n683,n690);
nand (n683,n684,n689);
or (n684,n685,n87);
not (n685,n686);
nand (n686,n687,n688);
or (n687,n97,n533);
or (n688,n96,n468);
nand (n689,n90,n600);
nand (n690,n691,n695);
or (n691,n692,n20);
nor (n692,n693,n694);
and (n693,n15,n108);
and (n694,n16,n107);
or (n695,n606,n21);
nand (n696,n697,n701);
or (n697,n112,n698);
nor (n698,n699,n700);
and (n699,n76,n208);
and (n700,n77,n268);
or (n701,n638,n113);
and (n702,n683,n690);
xor (n703,n588,n604);
and (n704,n661,n680);
xor (n705,n624,n627);
or (n706,n707,n752);
and (n707,n708,n711);
xor (n708,n709,n710);
xor (n709,n629,n642);
xor (n710,n660,n703);
or (n711,n712,n751);
and (n712,n713,n750);
xor (n713,n714,n728);
and (n714,n715,n721);
and (n715,n716,n97);
nand (n716,n717,n718);
or (n717,n63,n92);
nand (n718,n719,n585);
or (n719,n720,n67);
not (n720,n92);
nand (n721,n722,n723);
or (n722,n49,n667);
nand (n723,n724,n32);
not (n724,n725);
nor (n725,n726,n727);
and (n726,n39,n181);
and (n727,n40,n205);
or (n728,n729,n749);
and (n729,n730,n743);
xor (n730,n731,n737);
nand (n731,n732,n736);
or (n732,n68,n733);
nor (n733,n734,n735);
and (n734,n465,n63);
and (n735,n421,n67);
nand (n736,n675,n74);
nand (n737,n738,n739);
or (n738,n89,n685);
nand (n739,n88,n740);
nand (n740,n741,n742);
or (n741,n97,n585);
or (n742,n96,n498);
nand (n743,n744,n748);
or (n744,n20,n745);
nor (n745,n746,n747);
and (n746,n15,n102);
and (n747,n16,n101);
or (n748,n692,n21);
and (n749,n731,n737);
xor (n750,n663,n672);
and (n751,n714,n728);
and (n752,n709,n710);
not (n753,n754);
nand (n754,n755,n756);
xor (n755,n620,n648);
or (n756,n757,n758);
and (n757,n656,n705);
and (n758,n657,n658);
nand (n759,n760,n761);
not (n760,n755);
not (n761,n756);
nand (n762,n763,n766);
or (n763,n764,n765);
not (n764,n545);
nand (n765,n616,n618);
nand (n766,n547,n549);
nand (n767,n768,n1055,n544);
nand (n768,n769,n1045,n1054);
nand (n769,n770,n905,n912);
nor (n770,n771,n844);
not (n771,n772);
nand (n772,n773,n807);
not (n773,n774);
xor (n774,n775,n806);
xor (n775,n776,n777);
xor (n776,n682,n696);
or (n777,n778,n805);
and (n778,n779,n787);
xor (n779,n780,n786);
nand (n780,n781,n785);
or (n781,n112,n782);
nor (n782,n783,n784);
and (n783,n273,n76);
and (n784,n77,n338);
or (n785,n698,n113);
xor (n786,n715,n721);
or (n787,n788,n804);
and (n788,n789,n797);
xor (n789,n790,n791);
and (n790,n90,n498);
nand (n791,n792,n796);
or (n792,n793,n20);
nor (n793,n794,n795);
and (n794,n175,n16);
and (n795,n173,n15);
or (n796,n745,n21);
nand (n797,n798,n803);
or (n798,n68,n799);
not (n799,n800);
nor (n800,n801,n802);
and (n801,n533,n67);
and (n802,n63,n468);
or (n803,n73,n733);
and (n804,n790,n791);
and (n805,n780,n786);
xor (n806,n713,n750);
not (n807,n808);
or (n808,n809,n843);
and (n809,n810,n842);
xor (n810,n811,n812);
xor (n811,n730,n743);
or (n812,n813,n841);
and (n813,n814,n827);
xor (n814,n815,n821);
nand (n815,n816,n820);
or (n816,n31,n817);
nor (n817,n818,n819);
and (n818,n268,n40);
and (n819,n208,n39);
or (n820,n49,n725);
nand (n821,n822,n826);
or (n822,n112,n823);
nor (n823,n824,n825);
and (n824,n341,n76);
and (n825,n77,n418);
or (n826,n113,n782);
and (n827,n828,n834);
nor (n828,n829,n67);
nor (n829,n830,n832);
and (n830,n831,n585);
nand (n831,n77,n71);
and (n832,n76,n833);
not (n833,n71);
nand (n834,n835,n840);
or (n835,n20,n836);
not (n836,n837);
nor (n837,n838,n839);
and (n838,n16,n181);
and (n839,n205,n15);
or (n840,n793,n21);
and (n841,n815,n821);
xor (n842,n779,n787);
and (n843,n811,n812);
nand (n844,n845,n879);
not (n845,n846);
nor (n846,n847,n848);
xor (n847,n810,n842);
or (n848,n849,n878);
and (n849,n850,n877);
xor (n850,n851,n876);
or (n851,n852,n875);
and (n852,n853,n869);
xor (n853,n854,n861);
nand (n854,n855,n860);
or (n855,n856,n68);
not (n856,n857);
nand (n857,n858,n859);
or (n858,n63,n585);
or (n859,n67,n498);
nand (n860,n800,n74);
nand (n861,n862,n867);
or (n862,n863,n31);
not (n863,n864);
nand (n864,n865,n866);
or (n865,n40,n338);
or (n866,n39,n273);
nand (n867,n868,n33);
not (n868,n817);
nand (n869,n870,n874);
or (n870,n112,n871);
nor (n871,n872,n873);
and (n872,n76,n421);
and (n873,n77,n465);
or (n874,n113,n823);
and (n875,n854,n861);
xor (n876,n789,n797);
xor (n877,n814,n827);
and (n878,n851,n876);
or (n879,n880,n881);
xor (n880,n850,n877);
or (n881,n882,n904);
and (n882,n883,n903);
xor (n883,n884,n885);
xor (n884,n828,n834);
or (n885,n886,n902);
and (n886,n887,n895);
xor (n887,n888,n889);
and (n888,n74,n498);
nand (n889,n890,n891);
or (n890,n21,n836);
or (n891,n20,n892);
nor (n892,n893,n894);
and (n893,n15,n208);
and (n894,n16,n268);
nand (n895,n896,n901);
or (n896,n897,n31);
not (n897,n898);
nor (n898,n899,n900);
and (n899,n40,n341);
and (n900,n418,n39);
nand (n901,n33,n864);
and (n902,n888,n889);
xor (n903,n853,n869);
and (n904,n884,n885);
nand (n905,n906,n908);
not (n906,n907);
xor (n907,n708,n711);
not (n908,n909);
or (n909,n910,n911);
and (n910,n775,n806);
and (n911,n776,n777);
or (n912,n913,n1044);
and (n913,n914,n939);
xor (n914,n915,n938);
or (n915,n916,n937);
and (n916,n917,n936);
xor (n917,n918,n924);
nand (n918,n919,n923);
or (n919,n112,n920);
nor (n920,n921,n922);
and (n921,n76,n468);
and (n922,n77,n533);
or (n923,n113,n871);
and (n924,n925,n930);
and (n925,n926,n77);
nand (n926,n927,n928);
or (n927,n40,n115);
nand (n928,n929,n585);
or (n929,n117,n39);
nand (n930,n931,n935);
or (n931,n932,n20);
nor (n932,n933,n934);
and (n933,n15,n273);
and (n934,n16,n338);
or (n935,n892,n21);
xor (n936,n887,n895);
and (n937,n918,n924);
xor (n938,n883,n903);
or (n939,n940,n1043);
and (n940,n941,n962);
xor (n941,n942,n961);
or (n942,n943,n960);
and (n943,n944,n959);
xor (n944,n945,n952);
nand (n945,n946,n951);
or (n946,n947,n31);
not (n947,n948);
nor (n948,n949,n950);
and (n949,n465,n39);
and (n950,n40,n421);
nand (n951,n33,n898);
nand (n952,n953,n958);
or (n953,n954,n112);
not (n954,n955);
nand (n955,n956,n957);
or (n956,n585,n77);
or (n957,n76,n498);
or (n958,n113,n920);
xor (n959,n925,n930);
and (n960,n945,n952);
xor (n961,n917,n936);
or (n962,n963,n1042);
and (n963,n964,n984);
xor (n964,n965,n983);
or (n965,n966,n982);
and (n966,n967,n975);
xor (n967,n968,n969);
nor (n968,n113,n585);
nand (n969,n970,n974);
or (n970,n971,n31);
nor (n971,n972,n973);
and (n972,n468,n39);
and (n973,n533,n40);
nand (n974,n948,n33);
nand (n975,n976,n981);
or (n976,n20,n977);
not (n977,n978);
nand (n978,n979,n980);
or (n979,n341,n15);
nand (n980,n15,n341);
or (n981,n932,n21);
and (n982,n968,n969);
xor (n983,n944,n959);
or (n984,n985,n1041);
and (n985,n986,n1040);
xor (n986,n987,n1002);
nor (n987,n988,n996);
not (n988,n989);
nand (n989,n990,n995);
or (n990,n20,n991);
not (n991,n992);
nand (n992,n993,n994);
or (n993,n421,n15);
nand (n994,n15,n421);
nand (n995,n978,n22);
nand (n996,n997,n40);
nand (n997,n998,n1001);
nand (n998,n999,n585);
not (n999,n1000);
and (n1000,n16,n35);
or (n1001,n35,n16);
nand (n1002,n1003,n1039);
nand (n1003,n1004,n1017);
or (n1004,n1005,n1012);
not (n1005,n1006);
nor (n1006,n1007,n1011);
and (n1007,n32,n1008);
nand (n1008,n1009,n1010);
or (n1009,n40,n585);
or (n1010,n39,n498);
nor (n1011,n49,n971);
not (n1012,n1013);
nor (n1013,n1014,n1015);
and (n1014,n996,n989);
and (n1015,n1016,n988);
not (n1016,n996);
nand (n1017,n1018,n1038);
or (n1018,n1019,n1028);
nor (n1019,n1020,n1022);
not (n1020,n1021);
nand (n1021,n33,n498);
nand (n1022,n1023,n1024);
or (n1023,n21,n991);
nand (n1024,n1025,n286);
nand (n1025,n1026,n1027);
or (n1026,n533,n16);
nand (n1027,n16,n533);
nand (n1028,n1029,n1036);
nand (n1029,n1030,n1034);
or (n1030,n1031,n20);
nor (n1031,n1032,n1033);
and (n1032,n585,n16);
and (n1033,n498,n15);
or (n1034,n1035,n21);
not (n1035,n1025);
nor (n1036,n1037,n15);
and (n1037,n498,n22);
nand (n1038,n1020,n1022);
or (n1039,n1013,n1006);
xor (n1040,n967,n975);
and (n1041,n987,n1002);
and (n1042,n965,n983);
and (n1043,n942,n961);
and (n1044,n915,n938);
nand (n1045,n1046,n905);
nand (n1046,n1047,n1053);
or (n1047,n1048,n771);
not (n1048,n1049);
nand (n1049,n1050,n1052);
or (n1050,n846,n1051);
nand (n1051,n880,n881);
nand (n1052,n847,n848);
nand (n1053,n774,n808);
nand (n1054,n907,n909);
and (n1055,n759,n1056);
or (n1056,n655,n706);
nand (n1057,n1058,n398);
or (n1058,n1059,n1061);
not (n1059,n1060);
nand (n1060,n474,n475);
not (n1061,n1062);
nand (n1062,n400,n402);
or (n1063,n393,n3);
xor (n1064,n1065,n1843);
xor (n1065,n1066,n1840);
xor (n1066,n1067,n1839);
xor (n1067,n1068,n1830);
xor (n1068,n1069,n1829);
xor (n1069,n1070,n1815);
xor (n1070,n1071,n1814);
xor (n1071,n1072,n1793);
xor (n1072,n1073,n1792);
xor (n1073,n1074,n1766);
xor (n1074,n1075,n1765);
xor (n1075,n1076,n1732);
xor (n1076,n1077,n1731);
xor (n1077,n1078,n1693);
xor (n1078,n1079,n84);
xor (n1079,n1080,n1649);
xor (n1080,n1081,n1648);
xor (n1081,n1082,n1599);
xor (n1082,n1083,n1598);
xor (n1083,n1084,n1543);
xor (n1084,n1085,n1542);
xor (n1085,n1086,n1480);
xor (n1086,n1087,n1479);
or (n1087,n1088,n1416);
and (n1088,n1089,n180);
or (n1089,n1090,n1351);
and (n1090,n1091,n207);
or (n1091,n1092,n1286);
and (n1092,n1093,n272);
or (n1093,n1094,n1223);
and (n1094,n1095,n340);
or (n1095,n1096,n1159);
and (n1096,n1097,n420);
and (n1097,n467,n1098);
or (n1098,n1099,n1101);
and (n1099,n497,n1100);
and (n1100,n163,n468);
and (n1101,n1102,n1103);
xor (n1102,n497,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n163,n498);
and (n1106,n97,n468);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n97,n498);
and (n1112,n92,n468);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1118);
and (n1116,n1117,n802);
and (n1117,n92,n498);
and (n1118,n1119,n1120);
xor (n1119,n1117,n802);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
and (n1122,n63,n498);
and (n1123,n71,n468);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
and (n1128,n71,n498);
and (n1129,n77,n468);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
and (n1134,n77,n498);
and (n1135,n115,n468);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n115,n498);
and (n1141,n40,n468);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
and (n1146,n40,n498);
and (n1147,n35,n468);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
and (n1152,n35,n498);
and (n1153,n16,n468);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
and (n1156,n1157,n1158);
and (n1157,n16,n498);
and (n1158,n22,n468);
and (n1159,n1160,n1161);
xor (n1160,n1097,n420);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n467,n1098);
and (n1164,n163,n421);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1102,n1103);
and (n1170,n97,n421);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1108,n1109);
and (n1176,n92,n421);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1114,n1115);
and (n1182,n63,n421);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1119,n1120);
and (n1188,n71,n421);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1125,n1126);
and (n1194,n77,n421);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1131,n1132);
and (n1200,n115,n421);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1206);
and (n1204,n1205,n950);
xor (n1205,n1137,n1138);
and (n1206,n1207,n1208);
xor (n1207,n1205,n950);
or (n1208,n1209,n1212);
and (n1209,n1210,n1211);
xor (n1210,n1143,n1144);
and (n1211,n35,n421);
and (n1212,n1213,n1214);
xor (n1213,n1210,n1211);
or (n1214,n1215,n1218);
and (n1215,n1216,n1217);
xor (n1216,n1149,n1150);
and (n1217,n16,n421);
and (n1218,n1219,n1220);
xor (n1219,n1216,n1217);
and (n1220,n1221,n1222);
xor (n1221,n1155,n1156);
and (n1222,n22,n421);
and (n1223,n1224,n1225);
xor (n1224,n1095,n340);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1160,n1161);
and (n1228,n163,n341);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1166,n1167);
and (n1234,n97,n341);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1172,n1173);
and (n1240,n92,n341);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1246);
and (n1244,n1245,n677);
xor (n1245,n1178,n1179);
and (n1246,n1247,n1248);
xor (n1247,n1245,n677);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1184,n1185);
and (n1251,n71,n341);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1190,n1191);
and (n1257,n77,n341);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1196,n1197);
and (n1263,n115,n341);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
or (n1266,n1267,n1269);
and (n1267,n1268,n899);
xor (n1268,n1202,n1203);
and (n1269,n1270,n1271);
xor (n1270,n1268,n899);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1207,n1208);
and (n1274,n35,n341);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1213,n1214);
and (n1280,n16,n341);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
and (n1283,n1284,n1285);
xor (n1284,n1219,n1220);
and (n1285,n22,n341);
and (n1286,n1287,n1288);
xor (n1287,n1093,n272);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1224,n1225);
and (n1291,n163,n273);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1230,n1231);
and (n1297,n97,n273);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1236,n1237);
and (n1303,n92,n273);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1242,n1243);
and (n1309,n63,n273);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1247,n1248);
and (n1315,n71,n273);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1322);
and (n1319,n1320,n1321);
xor (n1320,n1253,n1254);
and (n1321,n77,n273);
and (n1322,n1323,n1324);
xor (n1323,n1320,n1321);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1259,n1260);
and (n1327,n115,n273);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1334);
and (n1331,n1332,n1333);
xor (n1332,n1265,n1266);
and (n1333,n40,n273);
and (n1334,n1335,n1336);
xor (n1335,n1332,n1333);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1270,n1271);
and (n1339,n35,n273);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1276,n1277);
and (n1345,n16,n273);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
and (n1348,n1349,n1350);
xor (n1349,n1282,n1283);
and (n1350,n22,n273);
and (n1351,n1352,n1353);
xor (n1352,n1091,n207);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1287,n1288);
and (n1356,n163,n208);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
or (n1359,n1360,n1363);
and (n1360,n1361,n1362);
xor (n1361,n1293,n1294);
and (n1362,n97,n208);
and (n1363,n1364,n1365);
xor (n1364,n1361,n1362);
or (n1365,n1366,n1369);
and (n1366,n1367,n1368);
xor (n1367,n1299,n1300);
and (n1368,n92,n208);
and (n1369,n1370,n1371);
xor (n1370,n1367,n1368);
or (n1371,n1372,n1375);
and (n1372,n1373,n1374);
xor (n1373,n1305,n1306);
and (n1374,n63,n208);
and (n1375,n1376,n1377);
xor (n1376,n1373,n1374);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1311,n1312);
and (n1380,n71,n208);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1317,n1318);
and (n1386,n77,n208);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1323,n1324);
and (n1392,n115,n208);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1329,n1330);
and (n1398,n40,n208);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
or (n1401,n1402,n1405);
and (n1402,n1403,n1404);
xor (n1403,n1335,n1336);
and (n1404,n35,n208);
and (n1405,n1406,n1407);
xor (n1406,n1403,n1404);
or (n1407,n1408,n1411);
and (n1408,n1409,n1410);
xor (n1409,n1341,n1342);
and (n1410,n16,n208);
and (n1411,n1412,n1413);
xor (n1412,n1409,n1410);
and (n1413,n1414,n1415);
xor (n1414,n1347,n1348);
and (n1415,n22,n208);
and (n1416,n1417,n1418);
xor (n1417,n1089,n180);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1352,n1353);
and (n1421,n163,n181);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1358,n1359);
and (n1427,n97,n181);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1364,n1365);
and (n1433,n92,n181);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1439);
and (n1437,n1438,n440);
xor (n1438,n1370,n1371);
and (n1439,n1440,n1441);
xor (n1440,n1438,n440);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1376,n1377);
and (n1444,n71,n181);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1382,n1383);
and (n1450,n77,n181);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1388,n1389);
and (n1456,n115,n181);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
or (n1459,n1460,n1463);
and (n1460,n1461,n1462);
xor (n1461,n1394,n1395);
and (n1462,n40,n181);
and (n1463,n1464,n1465);
xor (n1464,n1461,n1462);
or (n1465,n1466,n1469);
and (n1466,n1467,n1468);
xor (n1467,n1400,n1401);
and (n1468,n35,n181);
and (n1469,n1470,n1471);
xor (n1470,n1467,n1468);
or (n1471,n1472,n1474);
and (n1472,n1473,n838);
xor (n1473,n1406,n1407);
and (n1474,n1475,n1476);
xor (n1475,n1473,n838);
and (n1476,n1477,n1478);
xor (n1477,n1412,n1413);
and (n1478,n22,n181);
and (n1479,n168,n173);
or (n1480,n1481,n1484);
and (n1481,n1482,n1483);
xor (n1482,n1417,n1418);
and (n1483,n163,n173);
and (n1484,n1485,n1486);
xor (n1485,n1482,n1483);
or (n1486,n1487,n1490);
and (n1487,n1488,n1489);
xor (n1488,n1423,n1424);
and (n1489,n97,n173);
and (n1490,n1491,n1492);
xor (n1491,n1488,n1489);
or (n1492,n1493,n1496);
and (n1493,n1494,n1495);
xor (n1494,n1429,n1430);
and (n1495,n92,n173);
and (n1496,n1497,n1498);
xor (n1497,n1494,n1495);
or (n1498,n1499,n1501);
and (n1499,n1500,n370);
xor (n1500,n1435,n1436);
and (n1501,n1502,n1503);
xor (n1502,n1500,n370);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1440,n1441);
and (n1506,n71,n173);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1446,n1447);
and (n1512,n77,n173);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1452,n1453);
and (n1518,n115,n173);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1458,n1459);
and (n1524,n40,n173);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1464,n1465);
and (n1530,n35,n173);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1470,n1471);
and (n1536,n16,n173);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
and (n1539,n1540,n1541);
xor (n1540,n1475,n1476);
and (n1541,n22,n173);
and (n1542,n163,n102);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1485,n1486);
and (n1546,n97,n102);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1491,n1492);
and (n1552,n92,n102);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1558);
and (n1556,n1557,n302);
xor (n1557,n1497,n1498);
and (n1558,n1559,n1560);
xor (n1559,n1557,n302);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1502,n1503);
and (n1563,n71,n102);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
or (n1566,n1567,n1570);
and (n1567,n1568,n1569);
xor (n1568,n1508,n1509);
and (n1569,n77,n102);
and (n1570,n1571,n1572);
xor (n1571,n1568,n1569);
or (n1572,n1573,n1576);
and (n1573,n1574,n1575);
xor (n1574,n1514,n1515);
and (n1575,n115,n102);
and (n1576,n1577,n1578);
xor (n1577,n1574,n1575);
or (n1578,n1579,n1581);
and (n1579,n1580,n578);
xor (n1580,n1520,n1521);
and (n1581,n1582,n1583);
xor (n1582,n1580,n578);
or (n1583,n1584,n1587);
and (n1584,n1585,n1586);
xor (n1585,n1526,n1527);
and (n1586,n35,n102);
and (n1587,n1588,n1589);
xor (n1588,n1585,n1586);
or (n1589,n1590,n1593);
and (n1590,n1591,n1592);
xor (n1591,n1532,n1533);
and (n1592,n16,n102);
and (n1593,n1594,n1595);
xor (n1594,n1591,n1592);
and (n1595,n1596,n1597);
xor (n1596,n1538,n1539);
and (n1597,n22,n102);
and (n1598,n97,n108);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
xor (n1601,n1548,n1549);
and (n1602,n92,n108);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1608);
and (n1606,n1607,n237);
xor (n1607,n1554,n1555);
and (n1608,n1609,n1610);
xor (n1609,n1607,n237);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1559,n1560);
and (n1613,n71,n108);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1619);
and (n1617,n1618,n383);
xor (n1618,n1565,n1566);
and (n1619,n1620,n1621);
xor (n1620,n1618,n383);
or (n1621,n1622,n1625);
and (n1622,n1623,n1624);
xor (n1623,n1571,n1572);
and (n1624,n115,n108);
and (n1625,n1626,n1627);
xor (n1626,n1623,n1624);
or (n1627,n1628,n1631);
and (n1628,n1629,n1630);
xor (n1629,n1577,n1578);
and (n1630,n40,n108);
and (n1631,n1632,n1633);
xor (n1632,n1629,n1630);
or (n1633,n1634,n1637);
and (n1634,n1635,n1636);
xor (n1635,n1582,n1583);
and (n1636,n35,n108);
and (n1637,n1638,n1639);
xor (n1638,n1635,n1636);
or (n1639,n1640,n1643);
and (n1640,n1641,n1642);
xor (n1641,n1588,n1589);
and (n1642,n16,n108);
and (n1643,n1644,n1645);
xor (n1644,n1641,n1642);
and (n1645,n1646,n1647);
xor (n1646,n1594,n1595);
and (n1647,n22,n108);
and (n1648,n92,n65);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1604,n1605);
and (n1652,n63,n65);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1609,n1610);
and (n1658,n71,n65);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1615,n1616);
and (n1664,n77,n65);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
or (n1667,n1668,n1671);
and (n1668,n1669,n1670);
xor (n1669,n1620,n1621);
and (n1670,n115,n65);
and (n1671,n1672,n1673);
xor (n1672,n1669,n1670);
or (n1673,n1674,n1676);
and (n1674,n1675,n433);
xor (n1675,n1626,n1627);
and (n1676,n1677,n1678);
xor (n1677,n1675,n433);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1632,n1633);
and (n1681,n35,n65);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1638,n1639);
and (n1687,n16,n65);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
and (n1690,n1691,n1692);
xor (n1691,n1644,n1645);
and (n1692,n22,n65);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1654,n1655);
and (n1696,n71,n83);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1660,n1661);
and (n1702,n77,n83);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
or (n1705,n1706,n1709);
and (n1706,n1707,n1708);
xor (n1707,n1666,n1667);
and (n1708,n115,n83);
and (n1709,n1710,n1711);
xor (n1710,n1707,n1708);
or (n1711,n1712,n1714);
and (n1712,n1713,n359);
xor (n1713,n1672,n1673);
and (n1714,n1715,n1716);
xor (n1715,n1713,n359);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
xor (n1718,n1677,n1678);
and (n1719,n35,n83);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
xor (n1724,n1683,n1684);
and (n1725,n16,n83);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
and (n1728,n1729,n1730);
xor (n1729,n1689,n1690);
and (n1730,n22,n83);
and (n1731,n71,n123);
or (n1732,n1733,n1736);
and (n1733,n1734,n1735);
xor (n1734,n1698,n1699);
and (n1735,n77,n123);
and (n1736,n1737,n1738);
xor (n1737,n1734,n1735);
or (n1738,n1739,n1742);
and (n1739,n1740,n1741);
xor (n1740,n1704,n1705);
and (n1741,n115,n123);
and (n1742,n1743,n1744);
xor (n1743,n1740,n1741);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1710,n1711);
and (n1747,n40,n123);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
or (n1750,n1751,n1754);
and (n1751,n1752,n1753);
xor (n1752,n1715,n1716);
and (n1753,n35,n123);
and (n1754,n1755,n1756);
xor (n1755,n1752,n1753);
or (n1756,n1757,n1760);
and (n1757,n1758,n1759);
xor (n1758,n1721,n1722);
and (n1759,n16,n123);
and (n1760,n1761,n1762);
xor (n1761,n1758,n1759);
and (n1762,n1763,n1764);
xor (n1763,n1727,n1728);
and (n1764,n22,n123);
and (n1765,n77,n129);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1737,n1738);
and (n1769,n115,n129);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
or (n1772,n1773,n1775);
and (n1773,n1774,n226);
xor (n1774,n1743,n1744);
and (n1775,n1776,n1777);
xor (n1776,n1774,n226);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1749,n1750);
and (n1780,n35,n129);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1755,n1756);
and (n1786,n16,n129);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
and (n1789,n1790,n1791);
xor (n1790,n1761,n1762);
and (n1791,n22,n129);
and (n1792,n115,n45);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1771,n1772);
and (n1796,n40,n45);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1776,n1777);
and (n1802,n35,n45);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1782,n1783);
and (n1808,n16,n45);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
and (n1811,n1812,n1813);
xor (n1812,n1788,n1789);
and (n1813,n22,n45);
and (n1814,n40,n52);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1798,n1799);
and (n1818,n35,n52);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1824);
and (n1822,n1823,n220);
xor (n1823,n1804,n1805);
and (n1824,n1825,n1826);
xor (n1825,n1823,n220);
and (n1826,n1827,n1828);
xor (n1827,n1810,n1811);
and (n1828,n22,n52);
and (n1829,n35,n17);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1820,n1821);
and (n1833,n16,n17);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
and (n1836,n1837,n1838);
xor (n1837,n1825,n1826);
and (n1838,n22,n17);
and (n1839,n16,n27);
and (n1840,n1841,n1842);
xor (n1841,n1835,n1836);
and (n1842,n22,n27);
and (n1843,n22,n189);
endmodule
