module top (out,n14,n15,n22,n24,n33,n42,n44,n49,n51
        ,n62,n70,n77,n87,n97,n103,n106,n112,n130,n173
        ,n189);
output out;
input n14;
input n15;
input n22;
input n24;
input n33;
input n42;
input n44;
input n49;
input n51;
input n62;
input n70;
input n77;
input n87;
input n97;
input n103;
input n106;
input n112;
input n130;
input n173;
input n189;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
xor (out,n0,n398);
xor (n0,n1,n220);
xor (n1,n2,n156);
or (n2,n3,n155);
and (n3,n4,n123);
xor (n4,n5,n90);
or (n5,n6,n89);
and (n6,n7,n65);
xor (n7,n8,n36);
nand (n8,n9,n30);
or (n9,n10,n18);
not (n10,n11);
nand (n11,n12,n16);
or (n12,n13,n15);
not (n13,n14);
or (n16,n17,n14);
not (n17,n15);
not (n18,n19);
nor (n19,n20,n26);
nand (n20,n21,n25);
or (n21,n22,n23);
not (n23,n24);
nand (n25,n22,n23);
nor (n26,n27,n28);
and (n27,n13,n22);
and (n28,n14,n29);
not (n29,n22);
nand (n30,n20,n31);
nor (n31,n32,n34);
and (n32,n33,n14);
and (n34,n35,n13);
not (n35,n33);
nand (n36,n37,n57);
or (n37,n38,n46);
not (n38,n39);
nor (n39,n40,n45);
and (n40,n41,n43);
not (n41,n42);
not (n43,n44);
and (n45,n42,n44);
nand (n46,n47,n54);
nor (n47,n48,n52);
and (n48,n49,n50);
not (n50,n51);
and (n52,n53,n51);
not (n53,n49);
nand (n54,n55,n56);
or (n55,n51,n43);
nand (n56,n43,n51);
nand (n57,n58,n64);
not (n58,n59);
nor (n59,n60,n63);
and (n60,n61,n44);
not (n61,n62);
and (n63,n62,n43);
not (n64,n47);
nand (n65,n66,n83);
or (n66,n67,n73);
not (n67,n68);
nor (n68,n69,n71);
and (n69,n70,n24);
and (n71,n72,n23);
not (n72,n70);
not (n73,n74);
nor (n74,n75,n80);
nand (n75,n76,n78);
or (n76,n77,n43);
or (n78,n44,n79);
not (n79,n77);
nor (n80,n81,n82);
and (n81,n23,n77);
and (n82,n24,n79);
nand (n83,n75,n84);
nand (n84,n85,n88);
or (n85,n24,n86);
not (n86,n87);
or (n88,n23,n87);
and (n89,n8,n36);
xor (n90,n91,n115);
xor (n91,n92,n99);
and (n92,n93,n15);
not (n93,n94);
and (n94,n95,n98);
nand (n95,n14,n96);
not (n96,n97);
nand (n98,n97,n13);
nand (n99,n100,n109);
or (n100,n101,n104);
nand (n101,n102,n49);
not (n102,n103);
nor (n104,n105,n107);
and (n105,n53,n106);
and (n107,n49,n108);
not (n108,n106);
or (n109,n110,n102);
nor (n110,n111,n113);
and (n111,n53,n112);
and (n113,n49,n114);
not (n114,n112);
nand (n115,n116,n118);
or (n116,n117,n18);
not (n117,n31);
nand (n118,n119,n20);
not (n119,n120);
nor (n120,n121,n122);
and (n121,n13,n70);
and (n122,n14,n72);
xor (n123,n124,n141);
xor (n124,n125,n133);
nand (n125,n126,n127);
or (n126,n46,n59);
or (n127,n47,n128);
nor (n128,n129,n131);
and (n129,n43,n130);
and (n131,n44,n132);
not (n132,n130);
nand (n133,n134,n136);
or (n134,n135,n73);
not (n135,n84);
nand (n136,n137,n75);
not (n137,n138);
nor (n138,n139,n140);
and (n139,n23,n42);
and (n140,n24,n41);
and (n141,n142,n148);
nor (n142,n143,n13);
nor (n143,n144,n147);
and (n144,n145,n23);
not (n145,n146);
and (n146,n15,n22);
and (n147,n17,n29);
nand (n148,n149,n154);
or (n149,n101,n150);
not (n150,n151);
nor (n151,n152,n153);
and (n152,n132,n53);
and (n153,n130,n49);
or (n154,n104,n102);
and (n155,n5,n90);
xor (n156,n157,n195);
xor (n157,n158,n192);
xor (n158,n159,n184);
xor (n159,n160,n167);
nand (n160,n161,n162);
or (n161,n18,n120);
or (n162,n163,n164);
not (n163,n20);
nor (n164,n165,n166);
and (n165,n13,n87);
and (n166,n14,n86);
nand (n167,n168,n179);
or (n168,n169,n175);
not (n169,n170);
nand (n170,n171,n174);
or (n171,n172,n15);
not (n172,n173);
or (n174,n17,n173);
nand (n175,n94,n176);
nand (n176,n177,n178);
or (n177,n97,n172);
nand (n178,n172,n97);
nand (n179,n180,n93);
not (n180,n181);
nor (n181,n182,n183);
and (n182,n172,n33);
and (n183,n173,n35);
nand (n184,n185,n186);
or (n185,n101,n110);
or (n186,n187,n102);
nor (n187,n188,n190);
and (n188,n53,n189);
and (n190,n49,n191);
not (n191,n189);
or (n192,n193,n194);
and (n193,n124,n141);
and (n194,n125,n133);
xor (n195,n196,n217);
xor (n196,n197,n204);
nand (n197,n198,n199);
or (n198,n73,n138);
or (n199,n200,n201);
not (n200,n75);
nor (n201,n202,n203);
and (n202,n23,n62);
and (n203,n24,n61);
xor (n204,n205,n211);
and (n205,n206,n173);
nand (n206,n207,n208);
or (n207,n15,n97);
nand (n208,n209,n13);
not (n209,n210);
and (n210,n15,n97);
nand (n211,n212,n213);
or (n212,n46,n128);
or (n213,n47,n214);
nor (n214,n215,n216);
and (n215,n43,n106);
and (n216,n44,n108);
or (n217,n218,n219);
and (n218,n91,n115);
and (n219,n92,n99);
nand (n220,n221,n397);
or (n221,n222,n252);
not (n222,n223);
nand (n223,n224,n226);
not (n224,n225);
xor (n225,n4,n123);
not (n226,n227);
or (n227,n228,n251);
and (n228,n229,n250);
xor (n229,n230,n231);
xor (n230,n142,n148);
or (n231,n232,n249);
and (n232,n233,n242);
xor (n233,n234,n235);
and (n234,n20,n15);
nand (n235,n236,n241);
or (n236,n101,n237);
not (n237,n238);
nor (n238,n239,n240);
and (n239,n62,n49);
and (n240,n61,n53);
nand (n241,n151,n103);
nand (n242,n243,n248);
or (n243,n244,n46);
not (n244,n245);
nor (n245,n246,n247);
and (n246,n86,n43);
and (n247,n87,n44);
nand (n248,n64,n39);
and (n249,n234,n235);
xor (n250,n7,n65);
and (n251,n230,n231);
not (n252,n253);
nand (n253,n254,n396);
or (n254,n255,n286);
not (n255,n256);
nand (n256,n257,n259);
not (n257,n258);
xor (n258,n229,n250);
not (n259,n260);
or (n260,n261,n285);
and (n261,n262,n284);
xor (n262,n263,n270);
nand (n263,n264,n269);
or (n264,n265,n73);
not (n265,n266);
nor (n266,n267,n268);
and (n267,n33,n24);
and (n268,n35,n23);
nand (n269,n75,n68);
and (n270,n271,n276);
and (n271,n272,n24);
nand (n272,n273,n275);
or (n273,n274,n44);
and (n274,n15,n77);
or (n275,n15,n77);
nand (n276,n277,n278);
or (n277,n102,n237);
nand (n278,n279,n283);
not (n279,n280);
nor (n280,n281,n282);
and (n281,n42,n53);
and (n282,n41,n49);
not (n283,n101);
xor (n284,n233,n242);
and (n285,n263,n270);
not (n286,n287);
nand (n287,n288,n395);
or (n288,n289,n313);
not (n289,n290);
nand (n290,n291,n293);
not (n291,n292);
xor (n292,n262,n284);
not (n293,n294);
or (n294,n295,n312);
and (n295,n296,n311);
xor (n296,n297,n304);
nand (n297,n298,n303);
or (n298,n299,n46);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n72,n43);
and (n302,n70,n44);
nand (n303,n64,n245);
nand (n304,n305,n310);
or (n305,n306,n73);
not (n306,n307);
nand (n307,n308,n309);
or (n308,n23,n15);
or (n309,n24,n17);
nand (n310,n75,n266);
xor (n311,n271,n276);
and (n312,n297,n304);
not (n313,n314);
nand (n314,n315,n394);
or (n315,n316,n340);
not (n316,n317);
nand (n317,n318,n320);
not (n318,n319);
xor (n319,n296,n311);
not (n320,n321);
or (n321,n322,n339);
and (n322,n323,n332);
xor (n323,n324,n325);
and (n324,n75,n15);
nand (n325,n326,n331);
or (n326,n327,n46);
not (n327,n328);
nor (n328,n329,n330);
and (n329,n33,n44);
and (n330,n35,n43);
nand (n331,n64,n300);
nand (n332,n333,n338);
or (n333,n101,n334);
not (n334,n335);
nor (n335,n336,n337);
and (n336,n86,n53);
and (n337,n87,n49);
or (n338,n280,n102);
and (n339,n324,n325);
not (n340,n341);
nand (n341,n342,n393);
or (n342,n343,n359);
nor (n343,n344,n345);
xor (n344,n323,n332);
and (n345,n346,n352);
nor (n346,n347,n43);
nor (n347,n348,n349);
and (n348,n50,n17);
and (n349,n350,n53);
not (n350,n351);
and (n351,n15,n51);
nand (n352,n353,n354);
or (n353,n102,n334);
nand (n354,n355,n283);
not (n355,n356);
nor (n356,n357,n358);
and (n357,n53,n70);
and (n358,n49,n72);
not (n359,n360);
or (n360,n361,n392);
and (n361,n362,n371);
xor (n362,n363,n370);
nand (n363,n364,n369);
or (n364,n365,n46);
not (n365,n366);
nand (n366,n367,n368);
or (n367,n43,n15);
or (n368,n44,n17);
nand (n369,n64,n328);
xor (n370,n346,n352);
or (n371,n372,n391);
and (n372,n373,n381);
xor (n373,n374,n375);
nor (n374,n47,n17);
nand (n375,n376,n380);
or (n376,n377,n101);
nor (n377,n378,n379);
and (n378,n53,n33);
and (n379,n49,n35);
or (n380,n356,n102);
nor (n381,n382,n389);
nor (n382,n383,n385);
and (n383,n384,n103);
not (n384,n377);
nor (n385,n386,n101);
nor (n386,n387,n388);
and (n387,n15,n53);
and (n388,n17,n49);
or (n389,n390,n53);
and (n390,n15,n103);
and (n391,n374,n375);
and (n392,n363,n370);
nand (n393,n344,n345);
nand (n394,n319,n321);
nand (n395,n292,n294);
nand (n396,n258,n260);
nand (n397,n225,n227);
xor (n398,n399,n602);
xor (n399,n400,n600);
xor (n400,n401,n599);
xor (n401,n402,n591);
xor (n402,n403,n590);
xor (n403,n404,n576);
xor (n404,n405,n575);
xor (n405,n406,n556);
xor (n406,n407,n555);
xor (n407,n408,n529);
xor (n408,n409,n528);
xor (n409,n410,n499);
xor (n410,n411,n498);
xor (n411,n412,n460);
xor (n412,n413,n459);
xor (n413,n414,n417);
xor (n414,n415,n416);
and (n415,n189,n103);
and (n416,n112,n49);
or (n417,n418,n421);
and (n418,n419,n420);
and (n419,n112,n103);
and (n420,n106,n49);
and (n421,n422,n423);
xor (n422,n419,n420);
or (n423,n424,n426);
and (n424,n425,n153);
and (n425,n106,n103);
and (n426,n427,n428);
xor (n427,n425,n153);
or (n428,n429,n431);
and (n429,n430,n239);
and (n430,n130,n103);
and (n431,n432,n433);
xor (n432,n430,n239);
or (n433,n434,n437);
and (n434,n435,n436);
and (n435,n62,n103);
and (n436,n42,n49);
and (n437,n438,n439);
xor (n438,n435,n436);
or (n439,n440,n442);
and (n440,n441,n337);
and (n441,n42,n103);
and (n442,n443,n444);
xor (n443,n441,n337);
or (n444,n445,n448);
and (n445,n446,n447);
and (n446,n87,n103);
and (n447,n70,n49);
and (n448,n449,n450);
xor (n449,n446,n447);
or (n450,n451,n454);
and (n451,n452,n453);
and (n452,n70,n103);
and (n453,n33,n49);
and (n454,n455,n456);
xor (n455,n452,n453);
and (n456,n457,n458);
and (n457,n33,n103);
and (n458,n15,n49);
and (n459,n106,n51);
or (n460,n461,n464);
and (n461,n462,n463);
xor (n462,n422,n423);
and (n463,n130,n51);
and (n464,n465,n466);
xor (n465,n462,n463);
or (n466,n467,n470);
and (n467,n468,n469);
xor (n468,n427,n428);
and (n469,n62,n51);
and (n470,n471,n472);
xor (n471,n468,n469);
or (n472,n473,n476);
and (n473,n474,n475);
xor (n474,n432,n433);
and (n475,n42,n51);
and (n476,n477,n478);
xor (n477,n474,n475);
or (n478,n479,n482);
and (n479,n480,n481);
xor (n480,n438,n439);
and (n481,n87,n51);
and (n482,n483,n484);
xor (n483,n480,n481);
or (n484,n485,n488);
and (n485,n486,n487);
xor (n486,n443,n444);
and (n487,n70,n51);
and (n488,n489,n490);
xor (n489,n486,n487);
or (n490,n491,n494);
and (n491,n492,n493);
xor (n492,n449,n450);
and (n493,n33,n51);
and (n494,n495,n496);
xor (n495,n492,n493);
and (n496,n497,n351);
xor (n497,n455,n456);
and (n498,n130,n44);
or (n499,n500,n503);
and (n500,n501,n502);
xor (n501,n465,n466);
and (n502,n62,n44);
and (n503,n504,n505);
xor (n504,n501,n502);
or (n505,n506,n508);
and (n506,n507,n45);
xor (n507,n471,n472);
and (n508,n509,n510);
xor (n509,n507,n45);
or (n510,n511,n513);
and (n511,n512,n247);
xor (n512,n477,n478);
and (n513,n514,n515);
xor (n514,n512,n247);
or (n515,n516,n518);
and (n516,n517,n302);
xor (n517,n483,n484);
and (n518,n519,n520);
xor (n519,n517,n302);
or (n520,n521,n523);
and (n521,n522,n329);
xor (n522,n489,n490);
and (n523,n524,n525);
xor (n524,n522,n329);
and (n525,n526,n527);
xor (n526,n495,n496);
and (n527,n15,n44);
and (n528,n62,n77);
or (n529,n530,n533);
and (n530,n531,n532);
xor (n531,n504,n505);
and (n532,n42,n77);
and (n533,n534,n535);
xor (n534,n531,n532);
or (n535,n536,n539);
and (n536,n537,n538);
xor (n537,n509,n510);
and (n538,n87,n77);
and (n539,n540,n541);
xor (n540,n537,n538);
or (n541,n542,n545);
and (n542,n543,n544);
xor (n543,n514,n515);
and (n544,n70,n77);
and (n545,n546,n547);
xor (n546,n543,n544);
or (n547,n548,n551);
and (n548,n549,n550);
xor (n549,n519,n520);
and (n550,n33,n77);
and (n551,n552,n553);
xor (n552,n549,n550);
and (n553,n554,n274);
xor (n554,n524,n525);
and (n555,n42,n24);
or (n556,n557,n560);
and (n557,n558,n559);
xor (n558,n534,n535);
and (n559,n87,n24);
and (n560,n561,n562);
xor (n561,n558,n559);
or (n562,n563,n565);
and (n563,n564,n69);
xor (n564,n540,n541);
and (n565,n566,n567);
xor (n566,n564,n69);
or (n567,n568,n570);
and (n568,n569,n267);
xor (n569,n546,n547);
and (n570,n571,n572);
xor (n571,n569,n267);
and (n572,n573,n574);
xor (n573,n552,n553);
and (n574,n15,n24);
and (n575,n87,n22);
or (n576,n577,n580);
and (n577,n578,n579);
xor (n578,n561,n562);
and (n579,n70,n22);
and (n580,n581,n582);
xor (n581,n578,n579);
or (n582,n583,n586);
and (n583,n584,n585);
xor (n584,n566,n567);
and (n585,n33,n22);
and (n586,n587,n588);
xor (n587,n584,n585);
and (n588,n589,n146);
xor (n589,n571,n572);
and (n590,n70,n14);
or (n591,n592,n594);
and (n592,n593,n32);
xor (n593,n581,n582);
and (n594,n595,n596);
xor (n595,n593,n32);
and (n596,n597,n598);
xor (n597,n587,n588);
and (n598,n15,n14);
and (n599,n33,n97);
and (n600,n601,n210);
xor (n601,n595,n596);
and (n602,n15,n173);
endmodule
