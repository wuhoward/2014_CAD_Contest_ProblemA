module top (out,n3,n20,n22,n23,n32,n33,n35,n36,n46
        ,n56,n60,n70,n71,n73,n74,n81,n87,n99,n100
        ,n102,n103,n106,n112,n124,n125,n134,n140,n170,n210
        ,n241,n272,n596,n602,n612);
output out;
input n3;
input n20;
input n22;
input n23;
input n32;
input n33;
input n35;
input n36;
input n46;
input n56;
input n60;
input n70;
input n71;
input n73;
input n74;
input n81;
input n87;
input n99;
input n100;
input n102;
input n103;
input n106;
input n112;
input n124;
input n125;
input n134;
input n140;
input n170;
input n210;
input n241;
input n272;
input n596;
input n602;
input n612;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n101;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
xor (out,n0,n949);
nand (n0,n1,n553);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nand (n5,n6,n552);
or (n6,n7,n252);
not (n7,n8);
nand (n8,n9,n251);
nand (n9,n10,n220);
not (n10,n11);
xor (n11,n12,n179);
xor (n12,n13,n90);
xor (n13,n14,n62);
xor (n14,n15,n50);
nand (n15,n16,n42);
or (n16,n17,n27);
not (n17,n18);
nor (n18,n19,n24);
and (n19,n20,n21);
wire s0n21,s1n21,notn21;
or (n21,s0n21,s1n21);
not(notn21,n3);
and (s0n21,notn21,n22);
and (s1n21,n3,n23);
and (n24,n25,n26);
not (n25,n20);
not (n26,n21);
nand (n27,n28,n39);
nor (n28,n29,n37);
and (n29,n30,n34);
not (n30,n31);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n3);
and (s0n31,notn31,n32);
and (s1n31,n3,n33);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n3);
and (s0n34,notn34,n35);
and (s1n34,n3,n36);
and (n37,n31,n38);
not (n38,n34);
nand (n39,n40,n41);
or (n40,n30,n21);
nand (n41,n21,n30);
nand (n42,n43,n49);
not (n43,n44);
nor (n44,n45,n47);
and (n45,n26,n46);
and (n47,n21,n48);
not (n48,n46);
not (n49,n28);
nor (n50,n51,n57);
nand (n51,n21,n52);
not (n52,n53);
wire s0n53,s1n53,notn53;
or (n53,s0n53,s1n53);
not(notn53,n3);
and (s0n53,notn53,1'b0);
and (s1n53,n3,n55);
and (n55,n56,n23);
nor (n57,n58,n61);
and (n58,n53,n59);
not (n59,n60);
and (n61,n52,n60);
nand (n62,n63,n84);
or (n63,n64,n79);
nand (n64,n65,n76);
not (n65,n66);
nand (n66,n67,n75);
or (n67,n68,n72);
not (n68,n69);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n3);
and (s0n69,notn69,n70);
and (s1n69,n3,n71);
wire s0n72,s1n72,notn72;
or (n72,s0n72,s1n72);
not(notn72,n3);
and (s0n72,notn72,n73);
and (s1n72,n3,n74);
nand (n75,n72,n68);
nand (n76,n77,n78);
or (n77,n68,n34);
nand (n78,n34,n68);
nor (n79,n80,n82);
and (n80,n38,n81);
and (n82,n34,n83);
not (n83,n81);
or (n84,n65,n85);
nor (n85,n86,n88);
and (n86,n38,n87);
and (n88,n34,n89);
not (n89,n87);
xor (n90,n91,n156);
xor (n91,n92,n143);
xor (n92,n93,n116);
nand (n93,n94,n109);
or (n94,n95,n104);
not (n95,n96);
nor (n96,n97,n101);
not (n97,n98);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n3);
and (s0n98,notn98,n99);
and (s1n98,n3,n100);
wire s0n101,s1n101,notn101;
or (n101,s0n101,s1n101);
not(notn101,n3);
and (s0n101,notn101,n102);
and (s1n101,n3,n103);
nor (n104,n105,n107);
and (n105,n97,n106);
and (n107,n98,n108);
not (n108,n106);
or (n109,n110,n115);
nor (n110,n111,n113);
and (n111,n97,n112);
and (n113,n98,n114);
not (n114,n112);
not (n115,n101);
nand (n116,n117,n137);
or (n117,n118,n131);
not (n118,n119);
and (n119,n120,n127);
nand (n120,n121,n126);
or (n121,n122,n72);
not (n122,n123);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n3);
and (s0n123,notn123,n124);
and (s1n123,n3,n125);
nand (n126,n72,n122);
not (n127,n128);
nand (n128,n129,n130);
or (n129,n122,n98);
nand (n130,n98,n122);
nor (n131,n132,n135);
and (n132,n133,n134);
not (n133,n72);
and (n135,n72,n136);
not (n136,n134);
or (n137,n138,n127);
nor (n138,n139,n141);
and (n139,n133,n140);
and (n141,n72,n142);
not (n142,n140);
and (n143,n144,n150);
nand (n144,n145,n149);
or (n145,n95,n146);
nor (n146,n147,n148);
and (n147,n97,n140);
and (n148,n98,n142);
or (n149,n104,n115);
nand (n150,n151,n155);
or (n151,n118,n152);
nor (n152,n153,n154);
and (n153,n133,n87);
and (n154,n72,n89);
or (n155,n127,n131);
or (n156,n157,n178);
and (n157,n158,n172);
xor (n158,n159,n166);
nand (n159,n160,n165);
or (n160,n161,n27);
not (n161,n162);
nor (n162,n163,n164);
and (n163,n60,n21);
and (n164,n59,n26);
nand (n165,n49,n18);
nor (n166,n51,n167);
nor (n167,n168,n171);
and (n168,n53,n169);
not (n169,n170);
and (n171,n52,n170);
nand (n172,n173,n177);
or (n173,n64,n174);
nor (n174,n175,n176);
and (n175,n38,n46);
and (n176,n34,n48);
or (n177,n65,n79);
and (n178,n159,n166);
or (n179,n180,n219);
and (n180,n181,n196);
xor (n181,n182,n183);
xor (n182,n144,n150);
and (n183,n184,n190);
nand (n184,n185,n189);
or (n185,n95,n186);
nor (n186,n187,n188);
and (n187,n97,n134);
and (n188,n98,n136);
or (n189,n146,n115);
nand (n190,n191,n195);
or (n191,n118,n192);
nor (n192,n193,n194);
and (n193,n133,n81);
and (n194,n72,n83);
or (n195,n152,n127);
or (n196,n197,n218);
and (n197,n198,n212);
xor (n198,n199,n206);
nand (n199,n200,n205);
or (n200,n201,n27);
not (n201,n202);
nor (n202,n203,n204);
and (n203,n170,n21);
and (n204,n169,n26);
nand (n205,n49,n162);
nor (n206,n51,n207);
nor (n207,n208,n211);
and (n208,n53,n209);
not (n209,n210);
and (n211,n52,n210);
nand (n212,n213,n217);
or (n213,n64,n214);
nor (n214,n215,n216);
and (n215,n38,n20);
and (n216,n34,n25);
or (n217,n65,n174);
and (n218,n199,n206);
and (n219,n182,n183);
not (n220,n221);
or (n221,n222,n250);
and (n222,n223,n226);
xor (n223,n224,n225);
xor (n224,n158,n172);
xor (n225,n181,n196);
and (n226,n227,n228);
xor (n227,n184,n190);
or (n228,n229,n249);
and (n229,n230,n243);
xor (n230,n231,n237);
nand (n231,n232,n236);
or (n232,n233,n27);
nor (n233,n234,n235);
and (n234,n210,n26);
and (n235,n209,n21);
nand (n236,n202,n49);
nor (n237,n51,n238);
nor (n238,n239,n242);
and (n239,n53,n240);
not (n240,n241);
and (n242,n52,n241);
nand (n243,n244,n248);
or (n244,n95,n245);
nor (n245,n246,n247);
and (n246,n97,n87);
and (n247,n98,n89);
or (n248,n186,n115);
and (n249,n231,n237);
and (n250,n224,n225);
nand (n251,n11,n221);
not (n252,n253);
nand (n253,n254,n407,n551);
nand (n254,n255,n400);
nand (n255,n256,n399);
or (n256,n257,n388);
nor (n257,n258,n387);
and (n258,n259,n359);
not (n259,n260);
nor (n260,n261,n342);
or (n261,n262,n341);
and (n262,n263,n312);
xor (n263,n264,n299);
or (n264,n265,n298);
and (n265,n266,n289);
xor (n266,n267,n279);
nand (n267,n268,n275);
or (n268,n269,n27);
not (n269,n270);
nand (n270,n271,n273);
or (n271,n26,n272);
or (n273,n21,n274);
not (n274,n272);
or (n275,n28,n276);
nor (n276,n277,n278);
and (n277,n241,n26);
and (n278,n240,n21);
nand (n279,n280,n285);
or (n280,n281,n118);
not (n281,n282);
nand (n282,n283,n284);
or (n283,n72,n59);
or (n284,n133,n60);
nand (n285,n128,n286);
nor (n286,n287,n288);
and (n287,n20,n72);
and (n288,n25,n133);
nand (n289,n290,n294);
or (n290,n64,n291);
nor (n291,n292,n293);
and (n292,n38,n210);
and (n293,n34,n209);
or (n294,n65,n295);
nor (n295,n296,n297);
and (n296,n38,n170);
and (n297,n34,n169);
and (n298,n267,n279);
xor (n299,n300,n309);
xor (n300,n301,n303);
and (n301,n302,n272);
not (n302,n51);
nand (n303,n304,n308);
or (n304,n95,n305);
nor (n305,n306,n307);
and (n306,n83,n98);
and (n307,n81,n97);
or (n308,n245,n115);
nand (n309,n310,n311);
or (n310,n27,n276);
or (n311,n28,n233);
xor (n312,n313,n327);
xor (n313,n314,n321);
nand (n314,n315,n317);
or (n315,n118,n316);
not (n316,n286);
or (n317,n127,n318);
nor (n318,n319,n320);
and (n319,n133,n46);
and (n320,n72,n48);
nand (n321,n322,n323);
or (n322,n64,n295);
or (n323,n65,n324);
nor (n324,n325,n326);
and (n325,n38,n60);
and (n326,n34,n59);
and (n327,n328,n333);
nor (n328,n329,n26);
nor (n329,n330,n332);
and (n330,n38,n331);
nand (n331,n31,n272);
and (n332,n30,n274);
nand (n333,n334,n339);
or (n334,n335,n95);
not (n335,n336);
nor (n336,n337,n338);
and (n337,n46,n98);
and (n338,n48,n97);
nand (n339,n340,n101);
not (n340,n305);
and (n341,n264,n299);
xor (n342,n343,n348);
xor (n343,n344,n345);
xor (n344,n230,n243);
or (n345,n346,n347);
and (n346,n313,n327);
and (n347,n314,n321);
xor (n348,n349,n356);
xor (n349,n350,n353);
nand (n350,n351,n352);
or (n351,n64,n324);
or (n352,n65,n214);
nand (n353,n354,n355);
or (n354,n118,n318);
or (n355,n192,n127);
or (n356,n357,n358);
and (n357,n300,n309);
and (n358,n301,n303);
not (n359,n360);
nand (n360,n361,n362);
xor (n361,n263,n312);
or (n362,n363,n386);
and (n363,n364,n385);
xor (n364,n365,n366);
xor (n365,n328,n333);
or (n366,n367,n384);
and (n367,n368,n377);
xor (n368,n369,n370);
and (n369,n49,n272);
nand (n370,n371,n372);
or (n371,n115,n335);
nand (n372,n373,n96);
not (n373,n374);
nor (n374,n375,n376);
and (n375,n20,n97);
and (n376,n25,n98);
nand (n377,n378,n383);
or (n378,n379,n118);
not (n379,n380);
nor (n380,n381,n382);
and (n381,n170,n72);
and (n382,n133,n169);
nand (n383,n128,n282);
and (n384,n369,n370);
xor (n385,n266,n289);
and (n386,n365,n366);
and (n387,n261,n342);
nor (n388,n389,n396);
xor (n389,n390,n393);
xor (n390,n391,n392);
xor (n391,n198,n212);
xor (n392,n227,n228);
or (n393,n394,n395);
and (n394,n349,n356);
and (n395,n350,n353);
or (n396,n397,n398);
and (n397,n343,n348);
and (n398,n344,n345);
nand (n399,n389,n396);
nand (n400,n401,n403);
not (n401,n402);
xor (n402,n223,n226);
not (n403,n404);
or (n404,n405,n406);
and (n405,n390,n393);
and (n406,n391,n392);
nand (n407,n400,n408,n550);
nor (n408,n409,n547);
nor (n409,n410,n545);
and (n410,n411,n540);
or (n411,n412,n539);
and (n412,n413,n455);
xor (n413,n414,n448);
or (n414,n415,n447);
and (n415,n416,n435);
xor (n416,n417,n424);
nand (n417,n418,n423);
or (n418,n419,n118);
not (n419,n420);
nor (n420,n421,n422);
and (n421,n209,n133);
and (n422,n210,n72);
nand (n423,n128,n380);
nand (n424,n425,n430);
or (n425,n426,n65);
not (n426,n427);
nor (n427,n428,n429);
and (n428,n241,n34);
and (n429,n240,n38);
nand (n430,n431,n432);
not (n431,n64);
nand (n432,n433,n434);
or (n433,n38,n272);
or (n434,n34,n274);
xor (n435,n436,n441);
and (n436,n437,n34);
nand (n437,n438,n440);
or (n438,n72,n439);
and (n439,n272,n69);
or (n440,n69,n272);
nand (n441,n442,n446);
or (n442,n95,n443);
nor (n443,n444,n445);
and (n444,n97,n60);
and (n445,n98,n59);
or (n446,n374,n115);
and (n447,n417,n424);
xor (n448,n449,n454);
xor (n449,n450,n453);
nand (n450,n451,n452);
or (n451,n426,n64);
or (n452,n65,n291);
and (n453,n436,n441);
xor (n454,n368,n377);
or (n455,n456,n538);
and (n456,n457,n478);
xor (n457,n458,n477);
or (n458,n459,n476);
and (n459,n460,n469);
xor (n460,n461,n462);
and (n461,n66,n272);
nand (n462,n463,n468);
or (n463,n464,n118);
not (n464,n465);
nor (n465,n466,n467);
and (n466,n241,n72);
and (n467,n240,n133);
nand (n468,n420,n128);
nand (n469,n470,n475);
or (n470,n95,n471);
not (n471,n472);
nor (n472,n473,n474);
and (n473,n169,n97);
and (n474,n170,n98);
or (n475,n443,n115);
and (n476,n461,n462);
xor (n477,n416,n435);
or (n478,n479,n537);
and (n479,n480,n536);
xor (n480,n481,n495);
nor (n481,n482,n490);
not (n482,n483);
nand (n483,n484,n489);
or (n484,n485,n95);
not (n485,n486);
nand (n486,n487,n488);
or (n487,n209,n98);
nand (n488,n98,n209);
nand (n489,n472,n101);
nand (n490,n491,n72);
nand (n491,n492,n494);
or (n492,n98,n493);
and (n493,n272,n123);
or (n494,n123,n272);
nand (n495,n496,n534);
or (n496,n497,n520);
not (n497,n498);
nand (n498,n499,n519);
or (n499,n500,n509);
nor (n500,n501,n508);
nand (n501,n502,n507);
or (n502,n503,n95);
not (n503,n504);
nand (n504,n505,n506);
or (n505,n240,n98);
nand (n506,n98,n240);
nand (n507,n486,n101);
nor (n508,n127,n274);
nand (n509,n510,n517);
nand (n510,n511,n516);
or (n511,n512,n95);
not (n512,n513);
nand (n513,n514,n515);
or (n514,n97,n272);
or (n515,n98,n274);
nand (n516,n504,n101);
nor (n517,n518,n97);
and (n518,n272,n101);
nand (n519,n501,n508);
not (n520,n521);
nand (n521,n522,n530);
not (n522,n523);
nand (n523,n524,n529);
or (n524,n525,n118);
not (n525,n526);
nand (n526,n527,n528);
or (n527,n133,n272);
or (n528,n72,n274);
nand (n529,n128,n465);
nor (n530,n531,n533);
and (n531,n482,n532);
not (n532,n490);
and (n533,n483,n490);
nand (n534,n535,n523);
not (n535,n530);
xor (n536,n460,n469);
and (n537,n481,n495);
and (n538,n458,n477);
and (n539,n414,n448);
or (n540,n541,n542);
xor (n541,n364,n385);
or (n542,n543,n544);
and (n543,n449,n454);
and (n544,n450,n453);
not (n545,n546);
nand (n546,n541,n542);
nand (n547,n548,n259);
not (n548,n549);
nor (n549,n361,n362);
not (n550,n388);
nand (n551,n402,n404);
or (n552,n253,n8);
nand (n553,n554,n2);
xnor (n554,n555,n915);
nand (n555,n556,n902);
or (n556,n557,n848);
not (n557,n558);
and (n558,n559,n770,n842);
nor (n559,n560,n719);
nor (n560,n561,n674);
or (n561,n562,n673);
and (n562,n563,n647);
xor (n563,n564,n589);
xor (n564,n565,n580);
xor (n565,n566,n576);
nand (n566,n567,n572);
or (n567,n568,n27);
not (n568,n569);
nor (n569,n570,n571);
and (n570,n87,n21);
and (n571,n89,n26);
nand (n572,n49,n573);
nor (n573,n574,n575);
and (n574,n134,n21);
and (n575,n136,n26);
nor (n576,n51,n577);
nor (n577,n578,n579);
and (n578,n53,n83);
and (n579,n52,n81);
nand (n580,n581,n585);
or (n581,n64,n582);
nor (n582,n583,n584);
and (n583,n38,n140);
and (n584,n34,n142);
or (n585,n65,n586);
nor (n586,n587,n588);
and (n587,n38,n106);
and (n588,n34,n108);
xor (n589,n590,n627);
xor (n590,n591,n613);
xor (n591,n592,n605);
nand (n592,n593,n599);
or (n593,n95,n594);
nor (n594,n595,n597);
and (n595,n97,n596);
and (n597,n98,n598);
not (n598,n596);
or (n599,n600,n115);
nor (n600,n601,n603);
and (n601,n97,n602);
and (n603,n98,n604);
not (n604,n602);
nand (n605,n606,n610);
or (n606,n118,n607);
nor (n607,n608,n609);
and (n608,n133,n112);
and (n609,n72,n114);
or (n610,n611,n127);
xor (n611,n612,n133);
and (n613,n614,n621);
nand (n614,n615,n620);
or (n615,n95,n616);
nor (n616,n617,n618);
and (n617,n97,n612);
and (n618,n98,n619);
not (n619,n612);
or (n620,n594,n115);
nand (n621,n622,n626);
or (n622,n118,n623);
nor (n623,n624,n625);
and (n624,n133,n106);
and (n625,n72,n108);
or (n626,n127,n607);
or (n627,n628,n646);
and (n628,n629,n640);
xor (n629,n630,n636);
nand (n630,n631,n635);
or (n631,n632,n27);
nor (n632,n633,n634);
and (n633,n81,n26);
and (n634,n83,n21);
nand (n635,n49,n569);
nor (n636,n51,n637);
nor (n637,n638,n639);
and (n638,n53,n48);
and (n639,n52,n46);
nand (n640,n641,n645);
or (n641,n64,n642);
nor (n642,n643,n644);
and (n643,n38,n134);
and (n644,n34,n136);
or (n645,n65,n582);
and (n646,n630,n636);
or (n647,n648,n672);
and (n648,n649,n658);
xor (n649,n650,n651);
xor (n650,n614,n621);
and (n651,n652,n655);
nand (n652,n653,n654);
or (n653,n95,n110);
or (n654,n616,n115);
nand (n655,n656,n657);
or (n656,n118,n138);
or (n657,n623,n127);
or (n658,n659,n671);
and (n659,n660,n668);
xor (n660,n661,n664);
nand (n661,n662,n663);
or (n662,n27,n44);
or (n663,n28,n632);
nor (n664,n51,n665);
nor (n665,n666,n667);
and (n666,n53,n25);
and (n667,n52,n20);
nand (n668,n669,n670);
or (n669,n642,n65);
or (n670,n64,n85);
and (n671,n661,n664);
and (n672,n650,n651);
and (n673,n564,n589);
xor (n674,n675,n716);
xor (n675,n676,n695);
xor (n676,n677,n689);
xor (n677,n678,n685);
nand (n678,n679,n681);
or (n679,n680,n27);
not (n680,n573);
or (n681,n28,n682);
nor (n682,n683,n684);
and (n683,n26,n140);
and (n684,n21,n142);
nor (n685,n51,n686);
nor (n686,n687,n688);
and (n687,n53,n89);
and (n688,n52,n87);
nand (n689,n690,n691);
or (n690,n64,n586);
or (n691,n65,n692);
nor (n692,n693,n694);
and (n693,n38,n112);
and (n694,n34,n114);
xor (n695,n696,n713);
xor (n696,n697,n712);
xor (n697,n698,n706);
nand (n698,n699,n700);
or (n699,n95,n600);
or (n700,n701,n115);
nor (n701,n702,n704);
and (n702,n97,n703);
and (n703,n56,n602);
and (n704,n98,n705);
not (n705,n703);
nand (n706,n707,n708);
or (n707,n611,n118);
nand (n708,n128,n709);
nand (n709,n710,n711);
or (n710,n72,n598);
or (n711,n133,n596);
and (n712,n592,n605);
or (n713,n714,n715);
and (n714,n565,n580);
and (n715,n566,n576);
or (n716,n717,n718);
and (n717,n590,n627);
and (n718,n591,n613);
not (n719,n720);
nand (n720,n721,n766);
not (n721,n722);
xor (n722,n723,n742);
xor (n723,n724,n739);
xor (n724,n725,n733);
xor (n725,n726,n730);
nor (n726,n51,n727);
nor (n727,n728,n729);
and (n728,n53,n136);
and (n729,n52,n134);
nand (n730,n731,n732);
or (n731,n101,n96);
not (n732,n701);
nand (n733,n734,n738);
or (n734,n735,n65);
nor (n735,n736,n737);
and (n736,n612,n38);
and (n737,n619,n34);
or (n738,n64,n692);
or (n739,n740,n741);
and (n740,n696,n713);
and (n741,n697,n712);
xor (n742,n743,n748);
xor (n743,n744,n745);
and (n744,n698,n706);
or (n745,n746,n747);
and (n746,n677,n689);
and (n747,n678,n685);
nand (n748,n749,n765);
or (n749,n750,n758);
not (n750,n751);
nand (n751,n752,n754);
or (n752,n118,n753);
not (n753,n709);
or (n754,n127,n755);
nor (n755,n756,n757);
and (n756,n133,n602);
and (n757,n72,n604);
not (n758,n759);
nand (n759,n760,n761);
or (n760,n27,n682);
or (n761,n28,n762);
nor (n762,n763,n764);
and (n763,n26,n106);
and (n764,n21,n108);
or (n765,n759,n751);
not (n766,n767);
or (n767,n768,n769);
and (n768,n675,n716);
and (n769,n676,n695);
nand (n770,n771,n832);
not (n771,n772);
xor (n772,n773,n824);
xor (n773,n774,n794);
xor (n774,n775,n790);
xor (n775,n776,n781);
nand (n776,n777,n778);
or (n777,n119,n128);
nand (n778,n779,n780);
or (n779,n72,n705);
or (n780,n133,n703);
nand (n781,n782,n786);
or (n782,n64,n783);
nor (n783,n784,n785);
and (n784,n38,n596);
and (n785,n34,n598);
or (n786,n65,n787);
nor (n787,n788,n789);
and (n788,n38,n602);
and (n789,n34,n604);
nor (n790,n51,n791);
nor (n791,n792,n793);
and (n792,n53,n108);
and (n793,n52,n106);
xor (n794,n795,n810);
xor (n795,n796,n805);
nand (n796,n797,n801);
or (n797,n27,n798);
nor (n798,n799,n800);
and (n799,n26,n112);
and (n800,n21,n114);
or (n801,n28,n802);
nor (n802,n803,n804);
and (n803,n26,n612);
and (n804,n21,n619);
nand (n805,n806,n808);
or (n806,n807,n127);
not (n807,n778);
nand (n808,n809,n119);
not (n809,n755);
or (n810,n811,n823);
and (n811,n812,n820);
xor (n812,n813,n817);
nor (n813,n51,n814);
nor (n814,n815,n816);
and (n815,n53,n142);
and (n816,n52,n140);
nand (n817,n818,n819);
or (n818,n64,n735);
or (n819,n65,n783);
nand (n820,n821,n822);
or (n821,n27,n762);
or (n822,n28,n798);
and (n823,n813,n817);
or (n824,n825,n831);
and (n825,n826,n828);
xor (n826,n827,n765);
not (n827,n805);
or (n828,n829,n830);
and (n829,n725,n733);
and (n830,n726,n730);
and (n831,n827,n765);
not (n832,n833);
or (n833,n834,n841);
and (n834,n835,n838);
xor (n835,n836,n837);
xor (n836,n812,n820);
xor (n837,n826,n828);
or (n838,n839,n840);
and (n839,n743,n748);
and (n840,n744,n745);
and (n841,n836,n837);
not (n842,n843);
nor (n843,n844,n845);
xor (n844,n835,n838);
or (n845,n846,n847);
and (n846,n723,n742);
and (n847,n724,n739);
not (n848,n849);
nand (n849,n850,n892,n901);
nand (n850,n253,n851);
nor (n851,n852,n871);
nand (n852,n853,n9);
not (n853,n854);
nor (n854,n855,n868);
xor (n855,n856,n865);
xor (n856,n857,n858);
xor (n857,n660,n668);
xor (n858,n859,n862);
xor (n859,n860,n861);
xor (n860,n652,n655);
and (n861,n93,n116);
or (n862,n863,n864);
and (n863,n14,n62);
and (n864,n15,n50);
or (n865,n866,n867);
and (n866,n91,n156);
and (n867,n92,n143);
or (n868,n869,n870);
and (n869,n12,n179);
and (n870,n13,n90);
nand (n871,n872,n885);
nand (n872,n873,n881);
not (n873,n874);
xor (n874,n875,n878);
xor (n875,n876,n877);
xor (n876,n629,n640);
xor (n877,n649,n658);
or (n878,n879,n880);
and (n879,n859,n862);
and (n880,n860,n861);
not (n881,n882);
or (n882,n883,n884);
and (n883,n856,n865);
and (n884,n857,n858);
nand (n885,n886,n888);
not (n886,n887);
xor (n887,n563,n647);
not (n888,n889);
or (n889,n890,n891);
and (n890,n875,n878);
and (n891,n876,n877);
nand (n892,n893,n885);
nand (n893,n894,n900);
or (n894,n895,n896);
not (n895,n872);
not (n896,n897);
nand (n897,n898,n899);
or (n898,n854,n251);
nand (n899,n855,n868);
nand (n900,n874,n882);
nand (n901,n889,n887);
not (n902,n903);
nand (n903,n904,n914);
or (n904,n905,n906);
not (n905,n770);
not (n906,n907);
nand (n907,n908,n913);
or (n908,n909,n843);
nor (n909,n910,n912);
and (n910,n911,n720);
and (n911,n561,n674);
nor (n912,n721,n766);
nand (n913,n844,n845);
or (n914,n771,n832);
nand (n915,n916,n948);
not (n916,n917);
nor (n917,n918,n921);
or (n918,n919,n920);
and (n919,n773,n824);
and (n920,n774,n794);
xor (n921,n922,n945);
xor (n922,n923,n926);
or (n923,n924,n925);
and (n924,n775,n790);
and (n925,n776,n781);
xor (n926,n927,n938);
xor (n927,n928,n934);
nand (n928,n929,n930);
or (n929,n27,n802);
or (n930,n28,n931);
nor (n931,n932,n933);
and (n932,n26,n596);
and (n933,n21,n598);
nor (n934,n51,n935);
nor (n935,n936,n937);
and (n936,n53,n114);
and (n937,n52,n112);
nor (n938,n939,n941);
and (n939,n431,n940);
not (n940,n787);
and (n941,n66,n942);
nand (n942,n943,n944);
or (n943,n34,n705);
or (n944,n38,n703);
or (n945,n946,n947);
and (n946,n795,n810);
and (n947,n796,n805);
nand (n948,n918,n921);
wire s0n949,s1n949,notn949;
or (n949,s0n949,s1n949);
not(notn949,n3);
and (s0n949,notn949,n950);
and (s1n949,n3,n1968);
xor (n950,n951,n1670);
xor (n951,n952,n1966);
xor (n952,n953,n1665);
xor (n953,n954,n1959);
xor (n954,n955,n1659);
xor (n955,n956,n1947);
xor (n956,n957,n1653);
xor (n957,n958,n1930);
xor (n958,n959,n1647);
xor (n959,n960,n1908);
xor (n960,n961,n1641);
xor (n961,n962,n1881);
xor (n962,n963,n1635);
xor (n963,n964,n1849);
xor (n964,n965,n1629);
xor (n965,n966,n1812);
xor (n966,n967,n1623);
xor (n967,n968,n1770);
xor (n968,n969,n1617);
xor (n969,n970,n1723);
xor (n970,n971,n1611);
xor (n971,n972,n1671);
xor (n972,n973,n1605);
xor (n973,n974,n1602);
xor (n974,n975,n1601);
xor (n975,n976,n1531);
xor (n976,n977,n1530);
xor (n977,n978,n1449);
xor (n978,n979,n1448);
xor (n979,n980,n1362);
xor (n980,n981,n1361);
xor (n981,n982,n1269);
xor (n982,n983,n1268);
xor (n983,n984,n995);
xor (n984,n985,n994);
xor (n985,n986,n993);
xor (n986,n987,n992);
xor (n987,n988,n991);
xor (n988,n989,n990);
and (n989,n703,n101);
and (n990,n703,n98);
and (n991,n989,n990);
and (n992,n703,n123);
and (n993,n987,n992);
and (n994,n703,n72);
or (n995,n996,n997);
and (n996,n985,n994);
and (n997,n984,n998);
or (n998,n999,n1183);
and (n999,n1000,n1182);
xor (n1000,n986,n1001);
or (n1001,n1002,n1094);
and (n1002,n1003,n1093);
xor (n1003,n988,n1004);
or (n1004,n991,n1005);
and (n1005,n1006,n1008);
xor (n1006,n989,n1007);
and (n1007,n602,n98);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
and (n1010,n602,n101);
and (n1011,n596,n98);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
and (n1016,n596,n101);
and (n1017,n612,n98);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1024);
and (n1021,n1022,n1023);
and (n1022,n612,n101);
and (n1023,n112,n98);
and (n1024,n1025,n1026);
xor (n1025,n1022,n1023);
or (n1026,n1027,n1030);
and (n1027,n1028,n1029);
and (n1028,n112,n101);
and (n1029,n106,n98);
and (n1030,n1031,n1032);
xor (n1031,n1028,n1029);
or (n1032,n1033,n1036);
and (n1033,n1034,n1035);
and (n1034,n106,n101);
and (n1035,n140,n98);
and (n1036,n1037,n1038);
xor (n1037,n1034,n1035);
or (n1038,n1039,n1042);
and (n1039,n1040,n1041);
and (n1040,n140,n101);
and (n1041,n134,n98);
and (n1042,n1043,n1044);
xor (n1043,n1040,n1041);
or (n1044,n1045,n1048);
and (n1045,n1046,n1047);
and (n1046,n134,n101);
and (n1047,n87,n98);
and (n1048,n1049,n1050);
xor (n1049,n1046,n1047);
or (n1050,n1051,n1054);
and (n1051,n1052,n1053);
and (n1052,n87,n101);
and (n1053,n81,n98);
and (n1054,n1055,n1056);
xor (n1055,n1052,n1053);
or (n1056,n1057,n1059);
and (n1057,n1058,n337);
and (n1058,n81,n101);
and (n1059,n1060,n1061);
xor (n1060,n1058,n337);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
and (n1063,n46,n101);
and (n1064,n20,n98);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
and (n1069,n20,n101);
and (n1070,n60,n98);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1076);
and (n1074,n1075,n474);
and (n1075,n60,n101);
and (n1076,n1077,n1078);
xor (n1077,n1075,n474);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
and (n1080,n170,n101);
and (n1081,n210,n98);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
and (n1086,n210,n101);
and (n1087,n241,n98);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
and (n1090,n1091,n1092);
and (n1091,n241,n101);
and (n1092,n272,n98);
and (n1093,n602,n123);
and (n1094,n1095,n1096);
xor (n1095,n1003,n1093);
or (n1096,n1097,n1100);
and (n1097,n1098,n1099);
xor (n1098,n1006,n1008);
and (n1099,n596,n123);
and (n1100,n1101,n1102);
xor (n1101,n1098,n1099);
or (n1102,n1103,n1106);
and (n1103,n1104,n1105);
xor (n1104,n1013,n1014);
and (n1105,n612,n123);
and (n1106,n1107,n1108);
xor (n1107,n1104,n1105);
or (n1108,n1109,n1112);
and (n1109,n1110,n1111);
xor (n1110,n1019,n1020);
and (n1111,n112,n123);
and (n1112,n1113,n1114);
xor (n1113,n1110,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
xor (n1116,n1025,n1026);
and (n1117,n106,n123);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1031,n1032);
and (n1123,n140,n123);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1037,n1038);
and (n1129,n134,n123);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
xor (n1134,n1043,n1044);
and (n1135,n87,n123);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
xor (n1140,n1049,n1050);
and (n1141,n81,n123);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1055,n1056);
and (n1147,n46,n123);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1060,n1061);
and (n1153,n20,n123);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1066,n1067);
and (n1159,n60,n123);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1072,n1073);
and (n1165,n170,n123);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1077,n1078);
and (n1171,n210,n123);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1083,n1084);
and (n1177,n241,n123);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
and (n1180,n1181,n493);
xor (n1181,n1089,n1090);
and (n1182,n602,n72);
and (n1183,n1184,n1185);
xor (n1184,n1000,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1095,n1096);
and (n1188,n596,n72);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1101,n1102);
and (n1194,n612,n72);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1107,n1108);
and (n1200,n112,n72);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1113,n1114);
and (n1206,n106,n72);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1119,n1120);
and (n1212,n140,n72);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1125,n1126);
and (n1218,n134,n72);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1131,n1132);
and (n1224,n87,n72);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1137,n1138);
and (n1230,n81,n72);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1143,n1144);
and (n1236,n46,n72);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1242);
and (n1240,n1241,n287);
xor (n1241,n1149,n1150);
and (n1242,n1243,n1244);
xor (n1243,n1241,n287);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1155,n1156);
and (n1247,n60,n72);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1253);
and (n1251,n1252,n381);
xor (n1252,n1161,n1162);
and (n1253,n1254,n1255);
xor (n1254,n1252,n381);
or (n1255,n1256,n1258);
and (n1256,n1257,n422);
xor (n1257,n1167,n1168);
and (n1258,n1259,n1260);
xor (n1259,n1257,n422);
or (n1260,n1261,n1263);
and (n1261,n1262,n466);
xor (n1262,n1173,n1174);
and (n1263,n1264,n1265);
xor (n1264,n1262,n466);
and (n1265,n1266,n1267);
xor (n1266,n1179,n1180);
and (n1267,n272,n72);
and (n1268,n703,n69);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n984,n998);
and (n1272,n602,n69);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1184,n1185);
and (n1278,n596,n69);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1190,n1191);
and (n1284,n612,n69);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1196,n1197);
and (n1290,n112,n69);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1202,n1203);
and (n1296,n106,n69);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1208,n1209);
and (n1302,n140,n69);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1214,n1215);
and (n1308,n134,n69);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1220,n1221);
and (n1314,n87,n69);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1226,n1227);
and (n1320,n81,n69);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1232,n1233);
and (n1326,n46,n69);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1238,n1239);
and (n1332,n20,n69);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
or (n1335,n1336,n1339);
and (n1336,n1337,n1338);
xor (n1337,n1243,n1244);
and (n1338,n60,n69);
and (n1339,n1340,n1341);
xor (n1340,n1337,n1338);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1249,n1250);
and (n1344,n170,n69);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1351);
and (n1348,n1349,n1350);
xor (n1349,n1254,n1255);
and (n1350,n210,n69);
and (n1351,n1352,n1353);
xor (n1352,n1349,n1350);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1259,n1260);
and (n1356,n241,n69);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
and (n1359,n1360,n439);
xor (n1360,n1264,n1265);
and (n1361,n602,n34);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1274,n1275);
and (n1365,n596,n34);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1280,n1281);
and (n1371,n612,n34);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1286,n1287);
and (n1377,n112,n34);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1292,n1293);
and (n1383,n106,n34);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1298,n1299);
and (n1389,n140,n34);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
or (n1392,n1393,n1396);
and (n1393,n1394,n1395);
xor (n1394,n1304,n1305);
and (n1395,n134,n34);
and (n1396,n1397,n1398);
xor (n1397,n1394,n1395);
or (n1398,n1399,n1402);
and (n1399,n1400,n1401);
xor (n1400,n1310,n1311);
and (n1401,n87,n34);
and (n1402,n1403,n1404);
xor (n1403,n1400,n1401);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1316,n1317);
and (n1407,n81,n34);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1414);
and (n1411,n1412,n1413);
xor (n1412,n1322,n1323);
and (n1413,n46,n34);
and (n1414,n1415,n1416);
xor (n1415,n1412,n1413);
or (n1416,n1417,n1420);
and (n1417,n1418,n1419);
xor (n1418,n1328,n1329);
and (n1419,n20,n34);
and (n1420,n1421,n1422);
xor (n1421,n1418,n1419);
or (n1422,n1423,n1426);
and (n1423,n1424,n1425);
xor (n1424,n1334,n1335);
and (n1425,n60,n34);
and (n1426,n1427,n1428);
xor (n1427,n1424,n1425);
or (n1428,n1429,n1432);
and (n1429,n1430,n1431);
xor (n1430,n1340,n1341);
and (n1431,n170,n34);
and (n1432,n1433,n1434);
xor (n1433,n1430,n1431);
or (n1434,n1435,n1438);
and (n1435,n1436,n1437);
xor (n1436,n1346,n1347);
and (n1437,n210,n34);
and (n1438,n1439,n1440);
xor (n1439,n1436,n1437);
or (n1440,n1441,n1443);
and (n1441,n1442,n428);
xor (n1442,n1352,n1353);
and (n1443,n1444,n1445);
xor (n1444,n1442,n428);
and (n1445,n1446,n1447);
xor (n1446,n1358,n1359);
and (n1447,n272,n34);
and (n1448,n596,n31);
or (n1449,n1450,n1453);
and (n1450,n1451,n1452);
xor (n1451,n1367,n1368);
and (n1452,n612,n31);
and (n1453,n1454,n1455);
xor (n1454,n1451,n1452);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1373,n1374);
and (n1458,n112,n31);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1379,n1380);
and (n1464,n106,n31);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1385,n1386);
and (n1470,n140,n31);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1391,n1392);
and (n1476,n134,n31);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1397,n1398);
and (n1482,n87,n31);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1403,n1404);
and (n1488,n81,n31);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1409,n1410);
and (n1494,n46,n31);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1415,n1416);
and (n1500,n20,n31);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1421,n1422);
and (n1506,n60,n31);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1427,n1428);
and (n1512,n170,n31);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1433,n1434);
and (n1518,n210,n31);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1439,n1440);
and (n1524,n241,n31);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
and (n1527,n1528,n1529);
xor (n1528,n1444,n1445);
not (n1529,n331);
and (n1530,n612,n21);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1454,n1455);
and (n1534,n112,n21);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1460,n1461);
and (n1540,n106,n21);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1466,n1467);
and (n1546,n140,n21);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1552);
and (n1550,n1551,n574);
xor (n1551,n1472,n1473);
and (n1552,n1553,n1554);
xor (n1553,n1551,n574);
or (n1554,n1555,n1557);
and (n1555,n1556,n570);
xor (n1556,n1478,n1479);
and (n1557,n1558,n1559);
xor (n1558,n1556,n570);
or (n1559,n1560,n1563);
and (n1560,n1561,n1562);
xor (n1561,n1484,n1485);
and (n1562,n81,n21);
and (n1563,n1564,n1565);
xor (n1564,n1561,n1562);
or (n1565,n1566,n1569);
and (n1566,n1567,n1568);
xor (n1567,n1490,n1491);
and (n1568,n46,n21);
and (n1569,n1570,n1571);
xor (n1570,n1567,n1568);
or (n1571,n1572,n1574);
and (n1572,n1573,n19);
xor (n1573,n1496,n1497);
and (n1574,n1575,n1576);
xor (n1575,n1573,n19);
or (n1576,n1577,n1579);
and (n1577,n1578,n163);
xor (n1578,n1502,n1503);
and (n1579,n1580,n1581);
xor (n1580,n1578,n163);
or (n1581,n1582,n1584);
and (n1582,n1583,n203);
xor (n1583,n1508,n1509);
and (n1584,n1585,n1586);
xor (n1585,n1583,n203);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
xor (n1588,n1514,n1515);
and (n1589,n210,n21);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1520,n1521);
and (n1595,n241,n21);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
and (n1598,n1599,n1600);
xor (n1599,n1526,n1527);
and (n1600,n272,n21);
and (n1601,n112,n53);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1536,n1537);
and (n1605,n106,n53);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1542,n1543);
and (n1611,n140,n53);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1548,n1549);
and (n1617,n134,n53);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
or (n1620,n1621,n1624);
and (n1621,n1622,n1623);
xor (n1622,n1553,n1554);
and (n1623,n87,n53);
and (n1624,n1625,n1626);
xor (n1625,n1622,n1623);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1558,n1559);
and (n1629,n81,n53);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1564,n1565);
and (n1635,n46,n53);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1570,n1571);
and (n1641,n20,n53);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
xor (n1646,n1575,n1576);
and (n1647,n60,n53);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
or (n1650,n1651,n1654);
and (n1651,n1652,n1653);
xor (n1652,n1580,n1581);
and (n1653,n170,n53);
and (n1654,n1655,n1656);
xor (n1655,n1652,n1653);
or (n1656,n1657,n1660);
and (n1657,n1658,n1659);
xor (n1658,n1585,n1586);
and (n1659,n210,n53);
and (n1660,n1661,n1662);
xor (n1661,n1658,n1659);
or (n1662,n1663,n1666);
and (n1663,n1664,n1665);
xor (n1664,n1591,n1592);
and (n1665,n241,n53);
and (n1666,n1667,n1668);
xor (n1667,n1664,n1665);
and (n1668,n1669,n1670);
xor (n1669,n1597,n1598);
and (n1670,n272,n53);
or (n1671,n1672,n1674);
and (n1672,n1673,n1611);
xor (n1673,n1607,n1608);
and (n1674,n1675,n1676);
xor (n1675,n1673,n1611);
or (n1676,n1677,n1679);
and (n1677,n1678,n1617);
xor (n1678,n1613,n1614);
and (n1679,n1680,n1681);
xor (n1680,n1678,n1617);
or (n1681,n1682,n1684);
and (n1682,n1683,n1623);
xor (n1683,n1619,n1620);
and (n1684,n1685,n1686);
xor (n1685,n1683,n1623);
or (n1686,n1687,n1689);
and (n1687,n1688,n1629);
xor (n1688,n1625,n1626);
and (n1689,n1690,n1691);
xor (n1690,n1688,n1629);
or (n1691,n1692,n1694);
and (n1692,n1693,n1635);
xor (n1693,n1631,n1632);
and (n1694,n1695,n1696);
xor (n1695,n1693,n1635);
or (n1696,n1697,n1699);
and (n1697,n1698,n1641);
xor (n1698,n1637,n1638);
and (n1699,n1700,n1701);
xor (n1700,n1698,n1641);
or (n1701,n1702,n1704);
and (n1702,n1703,n1647);
xor (n1703,n1643,n1644);
and (n1704,n1705,n1706);
xor (n1705,n1703,n1647);
or (n1706,n1707,n1709);
and (n1707,n1708,n1653);
xor (n1708,n1649,n1650);
and (n1709,n1710,n1711);
xor (n1710,n1708,n1653);
or (n1711,n1712,n1714);
and (n1712,n1713,n1659);
xor (n1713,n1655,n1656);
and (n1714,n1715,n1716);
xor (n1715,n1713,n1659);
or (n1716,n1717,n1719);
and (n1717,n1718,n1665);
xor (n1718,n1661,n1662);
and (n1719,n1720,n1721);
xor (n1720,n1718,n1665);
and (n1721,n1722,n1670);
xor (n1722,n1667,n1668);
or (n1723,n1724,n1726);
and (n1724,n1725,n1617);
xor (n1725,n1675,n1676);
and (n1726,n1727,n1728);
xor (n1727,n1725,n1617);
or (n1728,n1729,n1731);
and (n1729,n1730,n1623);
xor (n1730,n1680,n1681);
and (n1731,n1732,n1733);
xor (n1732,n1730,n1623);
or (n1733,n1734,n1736);
and (n1734,n1735,n1629);
xor (n1735,n1685,n1686);
and (n1736,n1737,n1738);
xor (n1737,n1735,n1629);
or (n1738,n1739,n1741);
and (n1739,n1740,n1635);
xor (n1740,n1690,n1691);
and (n1741,n1742,n1743);
xor (n1742,n1740,n1635);
or (n1743,n1744,n1746);
and (n1744,n1745,n1641);
xor (n1745,n1695,n1696);
and (n1746,n1747,n1748);
xor (n1747,n1745,n1641);
or (n1748,n1749,n1751);
and (n1749,n1750,n1647);
xor (n1750,n1700,n1701);
and (n1751,n1752,n1753);
xor (n1752,n1750,n1647);
or (n1753,n1754,n1756);
and (n1754,n1755,n1653);
xor (n1755,n1705,n1706);
and (n1756,n1757,n1758);
xor (n1757,n1755,n1653);
or (n1758,n1759,n1761);
and (n1759,n1760,n1659);
xor (n1760,n1710,n1711);
and (n1761,n1762,n1763);
xor (n1762,n1760,n1659);
or (n1763,n1764,n1766);
and (n1764,n1765,n1665);
xor (n1765,n1715,n1716);
and (n1766,n1767,n1768);
xor (n1767,n1765,n1665);
and (n1768,n1769,n1670);
xor (n1769,n1720,n1721);
or (n1770,n1771,n1773);
and (n1771,n1772,n1623);
xor (n1772,n1727,n1728);
and (n1773,n1774,n1775);
xor (n1774,n1772,n1623);
or (n1775,n1776,n1778);
and (n1776,n1777,n1629);
xor (n1777,n1732,n1733);
and (n1778,n1779,n1780);
xor (n1779,n1777,n1629);
or (n1780,n1781,n1783);
and (n1781,n1782,n1635);
xor (n1782,n1737,n1738);
and (n1783,n1784,n1785);
xor (n1784,n1782,n1635);
or (n1785,n1786,n1788);
and (n1786,n1787,n1641);
xor (n1787,n1742,n1743);
and (n1788,n1789,n1790);
xor (n1789,n1787,n1641);
or (n1790,n1791,n1793);
and (n1791,n1792,n1647);
xor (n1792,n1747,n1748);
and (n1793,n1794,n1795);
xor (n1794,n1792,n1647);
or (n1795,n1796,n1798);
and (n1796,n1797,n1653);
xor (n1797,n1752,n1753);
and (n1798,n1799,n1800);
xor (n1799,n1797,n1653);
or (n1800,n1801,n1803);
and (n1801,n1802,n1659);
xor (n1802,n1757,n1758);
and (n1803,n1804,n1805);
xor (n1804,n1802,n1659);
or (n1805,n1806,n1808);
and (n1806,n1807,n1665);
xor (n1807,n1762,n1763);
and (n1808,n1809,n1810);
xor (n1809,n1807,n1665);
and (n1810,n1811,n1670);
xor (n1811,n1767,n1768);
or (n1812,n1813,n1815);
and (n1813,n1814,n1629);
xor (n1814,n1774,n1775);
and (n1815,n1816,n1817);
xor (n1816,n1814,n1629);
or (n1817,n1818,n1820);
and (n1818,n1819,n1635);
xor (n1819,n1779,n1780);
and (n1820,n1821,n1822);
xor (n1821,n1819,n1635);
or (n1822,n1823,n1825);
and (n1823,n1824,n1641);
xor (n1824,n1784,n1785);
and (n1825,n1826,n1827);
xor (n1826,n1824,n1641);
or (n1827,n1828,n1830);
and (n1828,n1829,n1647);
xor (n1829,n1789,n1790);
and (n1830,n1831,n1832);
xor (n1831,n1829,n1647);
or (n1832,n1833,n1835);
and (n1833,n1834,n1653);
xor (n1834,n1794,n1795);
and (n1835,n1836,n1837);
xor (n1836,n1834,n1653);
or (n1837,n1838,n1840);
and (n1838,n1839,n1659);
xor (n1839,n1799,n1800);
and (n1840,n1841,n1842);
xor (n1841,n1839,n1659);
or (n1842,n1843,n1845);
and (n1843,n1844,n1665);
xor (n1844,n1804,n1805);
and (n1845,n1846,n1847);
xor (n1846,n1844,n1665);
and (n1847,n1848,n1670);
xor (n1848,n1809,n1810);
or (n1849,n1850,n1852);
and (n1850,n1851,n1635);
xor (n1851,n1816,n1817);
and (n1852,n1853,n1854);
xor (n1853,n1851,n1635);
or (n1854,n1855,n1857);
and (n1855,n1856,n1641);
xor (n1856,n1821,n1822);
and (n1857,n1858,n1859);
xor (n1858,n1856,n1641);
or (n1859,n1860,n1862);
and (n1860,n1861,n1647);
xor (n1861,n1826,n1827);
and (n1862,n1863,n1864);
xor (n1863,n1861,n1647);
or (n1864,n1865,n1867);
and (n1865,n1866,n1653);
xor (n1866,n1831,n1832);
and (n1867,n1868,n1869);
xor (n1868,n1866,n1653);
or (n1869,n1870,n1872);
and (n1870,n1871,n1659);
xor (n1871,n1836,n1837);
and (n1872,n1873,n1874);
xor (n1873,n1871,n1659);
or (n1874,n1875,n1877);
and (n1875,n1876,n1665);
xor (n1876,n1841,n1842);
and (n1877,n1878,n1879);
xor (n1878,n1876,n1665);
and (n1879,n1880,n1670);
xor (n1880,n1846,n1847);
or (n1881,n1882,n1884);
and (n1882,n1883,n1641);
xor (n1883,n1853,n1854);
and (n1884,n1885,n1886);
xor (n1885,n1883,n1641);
or (n1886,n1887,n1889);
and (n1887,n1888,n1647);
xor (n1888,n1858,n1859);
and (n1889,n1890,n1891);
xor (n1890,n1888,n1647);
or (n1891,n1892,n1894);
and (n1892,n1893,n1653);
xor (n1893,n1863,n1864);
and (n1894,n1895,n1896);
xor (n1895,n1893,n1653);
or (n1896,n1897,n1899);
and (n1897,n1898,n1659);
xor (n1898,n1868,n1869);
and (n1899,n1900,n1901);
xor (n1900,n1898,n1659);
or (n1901,n1902,n1904);
and (n1902,n1903,n1665);
xor (n1903,n1873,n1874);
and (n1904,n1905,n1906);
xor (n1905,n1903,n1665);
and (n1906,n1907,n1670);
xor (n1907,n1878,n1879);
or (n1908,n1909,n1911);
and (n1909,n1910,n1647);
xor (n1910,n1885,n1886);
and (n1911,n1912,n1913);
xor (n1912,n1910,n1647);
or (n1913,n1914,n1916);
and (n1914,n1915,n1653);
xor (n1915,n1890,n1891);
and (n1916,n1917,n1918);
xor (n1917,n1915,n1653);
or (n1918,n1919,n1921);
and (n1919,n1920,n1659);
xor (n1920,n1895,n1896);
and (n1921,n1922,n1923);
xor (n1922,n1920,n1659);
or (n1923,n1924,n1926);
and (n1924,n1925,n1665);
xor (n1925,n1900,n1901);
and (n1926,n1927,n1928);
xor (n1927,n1925,n1665);
and (n1928,n1929,n1670);
xor (n1929,n1905,n1906);
or (n1930,n1931,n1933);
and (n1931,n1932,n1653);
xor (n1932,n1912,n1913);
and (n1933,n1934,n1935);
xor (n1934,n1932,n1653);
or (n1935,n1936,n1938);
and (n1936,n1937,n1659);
xor (n1937,n1917,n1918);
and (n1938,n1939,n1940);
xor (n1939,n1937,n1659);
or (n1940,n1941,n1943);
and (n1941,n1942,n1665);
xor (n1942,n1922,n1923);
and (n1943,n1944,n1945);
xor (n1944,n1942,n1665);
and (n1945,n1946,n1670);
xor (n1946,n1927,n1928);
or (n1947,n1948,n1950);
and (n1948,n1949,n1659);
xor (n1949,n1934,n1935);
and (n1950,n1951,n1952);
xor (n1951,n1949,n1659);
or (n1952,n1953,n1955);
and (n1953,n1954,n1665);
xor (n1954,n1939,n1940);
and (n1955,n1956,n1957);
xor (n1956,n1954,n1665);
and (n1957,n1958,n1670);
xor (n1958,n1944,n1945);
or (n1959,n1960,n1962);
and (n1960,n1961,n1665);
xor (n1961,n1951,n1952);
and (n1962,n1963,n1964);
xor (n1963,n1961,n1665);
and (n1964,n1965,n1670);
xor (n1965,n1956,n1957);
and (n1966,n1967,n1670);
xor (n1967,n1963,n1964);
xor (n1968,n1848,n1670);
endmodule
