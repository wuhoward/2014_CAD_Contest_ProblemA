module top (out,n4,n22,n23,n25,n26,n32,n33,n39,n40
        ,n51,n52,n57,n58,n63,n74,n75,n83,n94,n95
        ,n103,n109,n127,n168,n173,n174,n225,n281,n332,n371
        ,n419,n425,n434,n444,n450,n1031);
output out;
input n4;
input n22;
input n23;
input n25;
input n26;
input n32;
input n33;
input n39;
input n40;
input n51;
input n52;
input n57;
input n58;
input n63;
input n74;
input n75;
input n83;
input n94;
input n95;
input n103;
input n109;
input n127;
input n168;
input n173;
input n174;
input n225;
input n281;
input n332;
input n371;
input n419;
input n425;
input n434;
input n444;
input n450;
input n1031;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n53;
wire n54;
wire n55;
wire n56;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
xnor (out,n0,n1032);
nand (n0,n1,n1031);
nand (n1,n2,n906);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
nand (n6,n7,n905);
or (n7,n8,n241);
nand (n8,n9,n240);
nand (n9,n10,n189);
not (n10,n11);
xor (n11,n12,n142);
xor (n12,n13,n85);
xor (n13,n14,n71);
xor (n14,n15,n43);
nand (n15,n16,n35);
or (n16,n17,n29);
and (n17,n18,n28);
nand (n18,n19,n27);
or (n19,n20,n24);
not (n20,n21);
wire s0n21,s1n21,notn21;
or (n21,s0n21,s1n21);
not(notn21,n4);
and (s0n21,notn21,n22);
and (s1n21,n4,n23);
wire s0n24,s1n24,notn24;
or (n24,s0n24,s1n24);
not(notn24,n4);
and (s0n24,notn24,n25);
and (s1n24,n4,n26);
nand (n27,n24,n20);
not (n28,n29);
nand (n29,n30,n34);
or (n30,n20,n31);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n4);
and (s0n31,notn31,n32);
and (s1n31,n4,n33);
nand (n34,n31,n20);
nand (n35,n36,n41);
or (n36,n24,n37);
not (n37,n38);
and (n38,n39,n40);
or (n41,n42,n38);
not (n42,n24);
nand (n43,n44,n66);
or (n44,n45,n60);
nand (n45,n46,n54);
not (n46,n47);
nand (n47,n48,n53);
or (n48,n49,n24);
not (n49,n50);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n4);
and (s0n50,notn50,n51);
and (s1n50,n4,n52);
nand (n53,n24,n49);
nand (n54,n55,n59);
or (n55,n49,n56);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n4);
and (s0n56,notn56,n57);
and (s1n56,n4,n58);
nand (n59,n56,n49);
nor (n60,n61,n64);
and (n61,n62,n63);
not (n62,n56);
and (n64,n56,n65);
not (n65,n63);
or (n66,n46,n67);
nor (n67,n68,n69);
and (n68,n62,n40);
and (n69,n56,n70);
not (n70,n40);
nor (n71,n72,n80);
nand (n72,n73,n76);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n4);
and (s0n73,notn73,n74);
and (s1n73,n4,n75);
not (n76,n77);
wire s0n77,s1n77,notn77;
or (n77,s0n77,s1n77);
not(notn77,n4);
and (s0n77,notn77,1'b0);
and (s1n77,n4,n79);
and (n79,n39,n75);
nor (n80,n81,n84);
and (n81,n77,n82);
not (n82,n83);
and (n84,n76,n83);
xor (n85,n86,n120);
xor (n86,n87,n112);
nand (n87,n88,n106);
or (n88,n89,n100);
nand (n89,n90,n97);
nor (n90,n91,n96);
and (n91,n92,n56);
not (n92,n93);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n4);
and (s0n93,notn93,n94);
and (s1n93,n4,n95);
and (n96,n93,n62);
nand (n97,n98,n99);
or (n98,n92,n73);
nand (n99,n73,n92);
nor (n100,n101,n104);
and (n101,n102,n103);
not (n102,n73);
and (n104,n73,n105);
not (n105,n103);
or (n106,n90,n107);
nor (n107,n108,n110);
and (n108,n102,n109);
and (n110,n73,n111);
not (n111,n109);
nand (n112,n113,n115);
or (n113,n114,n28);
not (n114,n35);
nand (n115,n116,n17);
not (n116,n117);
nor (n117,n118,n119);
and (n118,n42,n40);
and (n119,n24,n70);
or (n120,n121,n141);
and (n121,n122,n135);
xor (n122,n123,n129);
nor (n123,n72,n124);
nor (n124,n125,n128);
and (n125,n77,n126);
not (n126,n127);
and (n128,n76,n127);
nand (n129,n130,n134);
or (n130,n45,n131);
nor (n131,n132,n133);
and (n132,n109,n62);
and (n133,n111,n56);
or (n134,n46,n60);
nand (n135,n136,n140);
or (n136,n89,n137);
nor (n137,n138,n139);
and (n138,n102,n83);
and (n139,n73,n82);
or (n140,n90,n100);
and (n141,n123,n129);
or (n142,n143,n188);
and (n143,n144,n161);
xor (n144,n145,n146);
not (n145,n112);
or (n146,n147,n153);
nand (n147,n148,n152);
or (n148,n89,n149);
nor (n149,n150,n151);
and (n150,n102,n127);
and (n151,n73,n126);
or (n152,n90,n137);
nand (n153,n154,n160);
or (n154,n155,n156);
not (n155,n17);
not (n156,n157);
nand (n157,n158,n159);
or (n158,n24,n65);
or (n159,n42,n63);
or (n160,n28,n117);
or (n161,n162,n187);
and (n162,n163,n181);
xor (n163,n164,n170);
nor (n164,n72,n165);
nor (n165,n166,n169);
and (n166,n77,n167);
not (n167,n168);
and (n169,n76,n168);
nand (n170,n171,n177);
or (n171,n172,n175);
wire s0n172,s1n172,notn172;
or (n172,s0n172,s1n172);
not(notn172,n4);
and (s0n172,notn172,n173);
and (s1n172,n4,n174);
nor (n175,n176,n172);
not (n176,n31);
not (n177,n178);
nor (n178,n179,n180);
and (n179,n176,n38);
and (n180,n31,n37);
nand (n181,n182,n183);
or (n182,n131,n46);
or (n183,n45,n184);
nor (n184,n185,n186);
and (n185,n62,n103);
and (n186,n56,n105);
and (n187,n164,n170);
and (n188,n145,n146);
not (n189,n190);
or (n190,n191,n239);
and (n191,n192,n195);
xor (n192,n193,n194);
xor (n193,n122,n135);
xor (n194,n144,n161);
or (n195,n196,n238);
and (n196,n197,n234);
xor (n197,n198,n211);
and (n198,n199,n207);
nand (n199,n200,n205);
or (n200,n201,n202);
not (n201,n175);
nor (n202,n203,n204);
and (n203,n176,n40);
and (n204,n31,n70);
or (n205,n178,n206);
not (n206,n172);
nand (n207,n208,n210);
or (n208,n209,n155);
xor (n209,n109,n42);
nand (n210,n29,n157);
or (n211,n212,n233);
and (n212,n213,n227);
xor (n213,n214,n221);
nand (n214,n215,n220);
or (n215,n216,n89);
not (n216,n217);
nor (n217,n218,n219);
and (n218,n168,n73);
and (n219,n167,n102);
or (n220,n90,n149);
nor (n221,n72,n222);
nor (n222,n223,n226);
and (n223,n77,n224);
not (n224,n225);
and (n226,n76,n225);
nand (n227,n228,n232);
or (n228,n45,n229);
nor (n229,n230,n231);
and (n230,n62,n83);
and (n231,n56,n82);
or (n232,n46,n184);
and (n233,n214,n221);
nand (n234,n235,n146);
or (n235,n236,n237);
not (n236,n153);
not (n237,n147);
and (n238,n198,n211);
and (n239,n193,n194);
or (n240,n10,n189);
nand (n241,n242,n904);
or (n242,n243,n293);
nor (n243,n244,n245);
xor (n244,n192,n195);
or (n245,n246,n292);
and (n246,n247,n291);
xor (n247,n248,n249);
xor (n248,n163,n181);
or (n249,n250,n290);
and (n250,n251,n266);
xor (n251,n252,n253);
xor (n252,n199,n207);
and (n253,n254,n260);
nand (n254,n255,n259);
or (n255,n201,n256);
nor (n256,n257,n258);
and (n257,n176,n63);
and (n258,n31,n65);
or (n259,n202,n206);
nand (n260,n261,n265);
or (n261,n155,n262);
nor (n262,n263,n264);
and (n263,n42,n103);
and (n264,n24,n105);
or (n265,n209,n28);
or (n266,n267,n289);
and (n267,n268,n283);
xor (n268,n269,n277);
nand (n269,n270,n275);
or (n270,n271,n89);
not (n271,n272);
nor (n272,n273,n274);
and (n273,n225,n73);
and (n274,n224,n102);
nand (n275,n276,n217);
not (n276,n90);
nor (n277,n72,n278);
nor (n278,n279,n282);
and (n279,n77,n280);
not (n280,n281);
and (n282,n76,n281);
nand (n283,n284,n288);
or (n284,n45,n285);
nor (n285,n286,n287);
and (n286,n62,n127);
and (n287,n56,n126);
or (n288,n46,n229);
and (n289,n269,n277);
and (n290,n252,n253);
xor (n291,n197,n234);
and (n292,n248,n249);
not (n293,n294);
nand (n294,n295,n900);
or (n295,n296,n397);
not (n296,n297);
nor (n297,n298,n389);
nor (n298,n299,n382);
or (n299,n300,n381);
and (n300,n301,n341);
xor (n301,n302,n303);
xor (n302,n268,n283);
xor (n303,n304,n319);
xor (n304,n305,n306);
xor (n305,n254,n260);
and (n306,n307,n313);
nand (n307,n308,n312);
or (n308,n201,n309);
nor (n309,n310,n311);
and (n310,n176,n109);
and (n311,n31,n111);
or (n312,n256,n206);
nand (n313,n314,n318);
or (n314,n155,n315);
nor (n315,n316,n317);
and (n316,n42,n83);
and (n317,n24,n82);
or (n318,n28,n262);
or (n319,n320,n340);
and (n320,n321,n334);
xor (n321,n322,n328);
nand (n322,n323,n327);
or (n323,n324,n89);
nor (n324,n325,n326);
and (n325,n281,n102);
and (n326,n280,n73);
nand (n327,n276,n272);
nor (n328,n72,n329);
nor (n329,n330,n333);
and (n330,n77,n331);
not (n331,n332);
and (n333,n76,n332);
nand (n334,n335,n339);
or (n335,n45,n336);
nor (n336,n337,n338);
and (n337,n62,n168);
and (n338,n56,n167);
or (n339,n46,n285);
and (n340,n322,n328);
or (n341,n342,n380);
and (n342,n343,n358);
xor (n343,n344,n345);
xor (n344,n307,n313);
and (n345,n346,n352);
nand (n346,n347,n351);
or (n347,n201,n348);
nor (n348,n349,n350);
and (n349,n176,n103);
and (n350,n31,n105);
or (n351,n309,n206);
nand (n352,n353,n357);
or (n353,n155,n354);
nor (n354,n355,n356);
and (n355,n42,n127);
and (n356,n24,n126);
or (n357,n315,n28);
or (n358,n359,n379);
and (n359,n360,n373);
xor (n360,n361,n367);
nand (n361,n362,n366);
or (n362,n89,n363);
nor (n363,n364,n365);
and (n364,n102,n332);
and (n365,n73,n331);
or (n366,n90,n324);
nor (n367,n72,n368);
nor (n368,n369,n372);
and (n369,n77,n370);
not (n370,n371);
and (n372,n76,n371);
nand (n373,n374,n375);
or (n374,n336,n46);
or (n375,n45,n376);
nor (n376,n377,n378);
and (n377,n62,n225);
and (n378,n56,n224);
and (n379,n361,n367);
and (n380,n344,n345);
and (n381,n302,n303);
xor (n382,n383,n386);
xor (n383,n384,n385);
xor (n384,n213,n227);
xor (n385,n251,n266);
or (n386,n387,n388);
and (n387,n304,n319);
and (n388,n305,n306);
not (n389,n390);
nand (n390,n391,n393);
not (n391,n392);
xor (n392,n247,n291);
not (n393,n394);
or (n394,n395,n396);
and (n395,n383,n386);
and (n396,n384,n385);
not (n397,n398);
nand (n398,n399,n889,n899);
nand (n399,n400,n810);
nand (n400,n401,n665,n809);
nand (n401,n402,n618);
nand (n402,n403,n617);
or (n403,n404,n572);
nor (n404,n405,n571);
and (n405,n406,n543);
not (n406,n407);
nor (n407,n408,n503);
or (n408,n409,n502);
and (n409,n410,n473);
xor (n410,n411,n454);
or (n411,n412,n453);
and (n412,n413,n440);
xor (n413,n414,n428);
nand (n414,n415,n422);
or (n415,n416,n89);
not (n416,n417);
nand (n417,n418,n420);
or (n418,n102,n419);
or (n420,n73,n421);
not (n421,n419);
or (n422,n90,n423);
nor (n423,n424,n426);
and (n424,n425,n102);
and (n426,n427,n73);
not (n427,n425);
nand (n428,n429,n436);
or (n429,n430,n155);
not (n430,n431);
nand (n431,n432,n435);
or (n432,n24,n433);
not (n433,n434);
or (n435,n42,n434);
nand (n436,n29,n437);
nor (n437,n438,n439);
and (n438,n371,n24);
and (n439,n370,n42);
nand (n440,n441,n447);
or (n441,n45,n442);
nor (n442,n443,n445);
and (n443,n62,n444);
and (n445,n56,n446);
not (n446,n444);
or (n447,n46,n448);
nor (n448,n449,n451);
and (n449,n62,n450);
and (n451,n56,n452);
not (n452,n450);
and (n453,n414,n428);
xor (n454,n455,n467);
xor (n455,n456,n458);
and (n456,n457,n419);
not (n457,n72);
nand (n458,n459,n463);
or (n459,n201,n460);
nor (n460,n461,n462);
and (n461,n280,n31);
and (n462,n281,n176);
or (n463,n464,n206);
nor (n464,n465,n466);
and (n465,n176,n225);
and (n466,n31,n224);
nand (n467,n468,n469);
or (n468,n89,n423);
or (n469,n90,n470);
nor (n470,n471,n472);
and (n471,n444,n102);
and (n472,n446,n73);
xor (n473,n474,n488);
xor (n474,n475,n482);
nand (n475,n476,n478);
or (n476,n155,n477);
not (n477,n437);
or (n478,n28,n479);
nor (n479,n480,n481);
and (n480,n42,n332);
and (n481,n24,n331);
nand (n482,n483,n484);
or (n483,n45,n448);
or (n484,n46,n485);
nor (n485,n486,n487);
and (n486,n62,n434);
and (n487,n56,n433);
and (n488,n489,n494);
nor (n489,n490,n102);
nor (n490,n491,n493);
and (n491,n62,n492);
nand (n492,n93,n419);
and (n493,n92,n421);
nand (n494,n495,n500);
or (n495,n496,n201);
not (n496,n497);
nor (n497,n498,n499);
and (n498,n332,n31);
and (n499,n331,n176);
nand (n500,n501,n172);
not (n501,n460);
and (n502,n411,n454);
xor (n503,n504,n526);
xor (n504,n505,n523);
xor (n505,n506,n517);
xor (n506,n507,n513);
nand (n507,n508,n509);
or (n508,n470,n89);
nand (n509,n510,n276);
nor (n510,n511,n512);
and (n511,n450,n73);
and (n512,n452,n102);
nor (n513,n72,n514);
nor (n514,n515,n516);
and (n515,n77,n427);
and (n516,n76,n425);
nand (n517,n518,n519);
or (n518,n201,n464);
or (n519,n520,n206);
nor (n520,n521,n522);
and (n521,n176,n168);
and (n522,n31,n167);
or (n523,n524,n525);
and (n524,n474,n488);
and (n525,n475,n482);
xor (n526,n527,n540);
xor (n527,n528,n534);
nand (n528,n529,n530);
or (n529,n45,n485);
or (n530,n46,n531);
nor (n531,n532,n533);
and (n532,n62,n371);
and (n533,n56,n370);
nand (n534,n535,n536);
or (n535,n155,n479);
or (n536,n537,n28);
nor (n537,n538,n539);
and (n538,n42,n281);
and (n539,n24,n280);
or (n540,n541,n542);
and (n541,n455,n467);
and (n542,n456,n458);
not (n543,n544);
nand (n544,n545,n546);
xor (n545,n410,n473);
or (n546,n547,n570);
and (n547,n548,n569);
xor (n548,n549,n550);
xor (n549,n489,n494);
or (n550,n551,n568);
and (n551,n552,n561);
xor (n552,n553,n554);
and (n553,n276,n419);
nand (n554,n555,n556);
or (n555,n206,n496);
nand (n556,n557,n175);
not (n557,n558);
nor (n558,n559,n560);
and (n559,n371,n176);
and (n560,n370,n31);
nand (n561,n562,n567);
or (n562,n563,n155);
not (n563,n564);
nor (n564,n565,n566);
and (n565,n450,n24);
and (n566,n42,n452);
nand (n567,n29,n431);
and (n568,n553,n554);
xor (n569,n413,n440);
and (n570,n549,n550);
and (n571,n408,n503);
nor (n572,n573,n614);
xor (n573,n574,n611);
xor (n574,n575,n594);
xor (n575,n576,n588);
xor (n576,n577,n584);
nand (n577,n578,n580);
or (n578,n579,n89);
not (n579,n510);
nand (n580,n276,n581);
nor (n581,n582,n583);
and (n582,n434,n73);
and (n583,n433,n102);
nor (n584,n72,n585);
nor (n585,n586,n587);
and (n586,n77,n446);
and (n587,n76,n444);
nand (n588,n589,n590);
or (n589,n45,n531);
or (n590,n46,n591);
nor (n591,n592,n593);
and (n592,n62,n332);
and (n593,n56,n331);
xor (n594,n595,n608);
xor (n595,n596,n602);
nand (n596,n597,n598);
or (n597,n201,n520);
or (n598,n599,n206);
nor (n599,n600,n601);
and (n600,n176,n127);
and (n601,n31,n126);
nand (n602,n603,n604);
or (n603,n155,n537);
or (n604,n605,n28);
nor (n605,n606,n607);
and (n606,n42,n225);
and (n607,n24,n224);
or (n608,n609,n610);
and (n609,n506,n517);
and (n610,n507,n513);
or (n611,n612,n613);
and (n612,n527,n540);
and (n613,n528,n534);
or (n614,n615,n616);
and (n615,n504,n526);
and (n616,n505,n523);
nand (n617,n573,n614);
nand (n618,n619,n661);
not (n619,n620);
xor (n620,n621,n660);
xor (n621,n622,n641);
xor (n622,n623,n635);
xor (n623,n624,n631);
nand (n624,n625,n627);
or (n625,n626,n89);
not (n626,n581);
nand (n627,n276,n628);
nor (n628,n629,n630);
and (n629,n371,n73);
and (n630,n370,n102);
nor (n631,n72,n632);
nor (n632,n633,n634);
and (n633,n77,n452);
and (n634,n76,n450);
nand (n635,n636,n637);
or (n636,n45,n591);
or (n637,n46,n638);
nor (n638,n639,n640);
and (n639,n62,n281);
and (n640,n56,n280);
xor (n641,n642,n657);
xor (n642,n643,n656);
xor (n643,n644,n650);
nand (n644,n645,n646);
or (n645,n201,n599);
or (n646,n647,n206);
nor (n647,n648,n649);
and (n648,n176,n83);
and (n649,n31,n82);
nand (n650,n651,n652);
or (n651,n155,n605);
or (n652,n28,n653);
nor (n653,n654,n655);
and (n654,n42,n168);
and (n655,n24,n167);
and (n656,n596,n602);
or (n657,n658,n659);
and (n658,n576,n588);
and (n659,n577,n584);
and (n660,n595,n608);
not (n661,n662);
or (n662,n663,n664);
and (n663,n574,n611);
and (n664,n575,n594);
nand (n665,n618,n666,n808);
nor (n666,n667,n805);
nor (n667,n668,n803);
and (n668,n669,n798);
or (n669,n670,n797);
and (n670,n671,n713);
xor (n671,n672,n706);
or (n672,n673,n705);
and (n673,n674,n693);
xor (n674,n675,n682);
nand (n675,n676,n681);
or (n676,n677,n155);
not (n677,n678);
nor (n678,n679,n680);
and (n679,n446,n42);
and (n680,n444,n24);
nand (n681,n29,n564);
nand (n682,n683,n688);
or (n683,n684,n46);
not (n684,n685);
nor (n685,n686,n687);
and (n686,n425,n56);
and (n687,n427,n62);
nand (n688,n689,n690);
not (n689,n45);
nand (n690,n691,n692);
or (n691,n62,n419);
or (n692,n56,n421);
xor (n693,n694,n699);
and (n694,n695,n56);
nand (n695,n696,n698);
or (n696,n24,n697);
and (n697,n419,n50);
or (n698,n50,n419);
nand (n699,n700,n704);
or (n700,n201,n701);
nor (n701,n702,n703);
and (n702,n176,n434);
and (n703,n31,n433);
or (n704,n558,n206);
and (n705,n675,n682);
xor (n706,n707,n712);
xor (n707,n708,n711);
nand (n708,n709,n710);
or (n709,n684,n45);
or (n710,n46,n442);
and (n711,n694,n699);
xor (n712,n552,n561);
or (n713,n714,n796);
and (n714,n715,n736);
xor (n715,n716,n735);
or (n716,n717,n734);
and (n717,n718,n727);
xor (n718,n719,n720);
and (n719,n47,n419);
nand (n720,n721,n726);
or (n721,n722,n155);
not (n722,n723);
nor (n723,n724,n725);
and (n724,n425,n24);
and (n725,n427,n42);
nand (n726,n678,n29);
nand (n727,n728,n733);
or (n728,n201,n729);
not (n729,n730);
nor (n730,n731,n732);
and (n731,n452,n176);
and (n732,n450,n31);
or (n733,n701,n206);
and (n734,n719,n720);
xor (n735,n674,n693);
or (n736,n737,n795);
and (n737,n738,n794);
xor (n738,n739,n753);
nor (n739,n740,n748);
not (n740,n741);
nand (n741,n742,n747);
or (n742,n743,n201);
not (n743,n744);
nand (n744,n745,n746);
or (n745,n446,n31);
nand (n746,n31,n446);
nand (n747,n730,n172);
nand (n748,n749,n24);
nand (n749,n750,n752);
or (n750,n31,n751);
and (n751,n419,n21);
or (n752,n21,n419);
nand (n753,n754,n792);
or (n754,n755,n778);
not (n755,n756);
nand (n756,n757,n777);
or (n757,n758,n767);
nor (n758,n759,n766);
nand (n759,n760,n765);
or (n760,n761,n201);
not (n761,n762);
nand (n762,n763,n764);
or (n763,n427,n31);
nand (n764,n31,n427);
nand (n765,n744,n172);
nor (n766,n28,n421);
nand (n767,n768,n775);
nand (n768,n769,n774);
or (n769,n770,n201);
not (n770,n771);
nand (n771,n772,n773);
or (n772,n176,n419);
or (n773,n31,n421);
nand (n774,n762,n172);
nor (n775,n776,n176);
and (n776,n419,n172);
nand (n777,n759,n766);
not (n778,n779);
nand (n779,n780,n788);
not (n780,n781);
nand (n781,n782,n787);
or (n782,n783,n155);
not (n783,n784);
nand (n784,n785,n786);
or (n785,n42,n419);
or (n786,n24,n421);
nand (n787,n29,n723);
nor (n788,n789,n791);
and (n789,n740,n790);
not (n790,n748);
and (n791,n741,n748);
nand (n792,n793,n781);
not (n793,n788);
xor (n794,n718,n727);
and (n795,n739,n753);
and (n796,n716,n735);
and (n797,n672,n706);
or (n798,n799,n800);
xor (n799,n548,n569);
or (n800,n801,n802);
and (n801,n707,n712);
and (n802,n708,n711);
not (n803,n804);
nand (n804,n799,n800);
nand (n805,n806,n406);
not (n806,n807);
nor (n807,n545,n546);
not (n808,n572);
nand (n809,n620,n662);
nor (n810,n811,n868);
nand (n811,n812,n861);
not (n812,n813);
nor (n813,n814,n852);
xor (n814,n815,n843);
xor (n815,n816,n817);
xor (n816,n360,n373);
xor (n817,n818,n827);
xor (n818,n819,n820);
xor (n819,n346,n352);
and (n820,n821,n824);
nand (n821,n822,n823);
or (n822,n201,n647);
or (n823,n348,n206);
nand (n824,n825,n826);
or (n825,n155,n653);
or (n826,n354,n28);
or (n827,n828,n842);
and (n828,n829,n839);
xor (n829,n830,n835);
nand (n830,n831,n833);
or (n831,n832,n89);
not (n832,n628);
nand (n833,n834,n276);
not (n834,n363);
nor (n835,n72,n836);
nor (n836,n837,n838);
and (n837,n77,n433);
and (n838,n76,n434);
nand (n839,n840,n841);
or (n840,n45,n638);
or (n841,n46,n376);
and (n842,n830,n835);
or (n843,n844,n851);
and (n844,n845,n848);
xor (n845,n846,n847);
xor (n846,n821,n824);
and (n847,n644,n650);
or (n848,n849,n850);
and (n849,n623,n635);
and (n850,n624,n631);
and (n851,n846,n847);
or (n852,n853,n860);
and (n853,n854,n857);
xor (n854,n855,n856);
xor (n855,n829,n839);
xor (n856,n845,n848);
or (n857,n858,n859);
and (n858,n642,n657);
and (n859,n643,n656);
and (n860,n855,n856);
nand (n861,n862,n864);
not (n862,n863);
xor (n863,n854,n857);
not (n864,n865);
or (n865,n866,n867);
and (n866,n621,n660);
and (n867,n622,n641);
nand (n868,n869,n882);
nand (n869,n870,n878);
not (n870,n871);
xor (n871,n872,n875);
xor (n872,n873,n874);
xor (n873,n321,n334);
xor (n874,n343,n358);
or (n875,n876,n877);
and (n876,n818,n827);
and (n877,n819,n820);
not (n878,n879);
or (n879,n880,n881);
and (n880,n815,n843);
and (n881,n816,n817);
nand (n882,n883,n885);
not (n883,n884);
xor (n884,n301,n341);
not (n885,n886);
or (n886,n887,n888);
and (n887,n872,n875);
and (n888,n873,n874);
nand (n889,n890,n882);
nand (n890,n891,n898);
or (n891,n892,n893);
not (n892,n869);
not (n893,n894);
nand (n894,n895,n897);
or (n895,n813,n896);
nand (n896,n863,n865);
nand (n897,n814,n852);
nand (n898,n871,n879);
nand (n899,n886,n884);
nor (n900,n901,n903);
and (n901,n902,n390);
and (n902,n299,n382);
nor (n903,n391,n393);
nand (n904,n244,n245);
nand (n905,n241,n8);
not (n906,n907);
and (n907,n908,n3,n39);
nand (n908,n909,n1030);
or (n909,n910,n963);
not (n910,n911);
nor (n911,n912,n962);
and (n912,n913,n951);
not (n913,n914);
or (n914,n915,n950);
and (n915,n916,n931);
xor (n916,n917,n927);
nand (n917,n918,n923);
or (n918,n919,n90);
not (n919,n920);
nand (n920,n921,n922);
or (n921,n73,n37);
or (n922,n102,n38);
or (n923,n89,n924);
nor (n924,n925,n926);
and (n925,n102,n40);
and (n926,n73,n70);
nand (n927,n928,n929,n457);
or (n928,n77,n63);
not (n929,n930);
and (n930,n63,n77);
or (n931,n932,n949);
and (n932,n933,n945);
xor (n933,n934,n939);
nand (n934,n935,n936);
or (n935,n689,n47);
nand (n936,n937,n938);
or (n937,n56,n37);
or (n938,n62,n38);
nand (n939,n940,n944);
or (n940,n89,n941);
nor (n941,n942,n943);
and (n942,n102,n63);
and (n943,n73,n65);
or (n944,n90,n924);
nor (n945,n72,n946);
nor (n946,n947,n948);
and (n947,n77,n111);
and (n948,n76,n109);
and (n949,n934,n939);
and (n950,n917,n927);
not (n951,n952);
xor (n952,n953,n961);
xor (n953,n954,n957);
nand (n954,n955,n920);
or (n955,n956,n276);
not (n956,n89);
nor (n957,n72,n958);
nor (n958,n959,n960);
and (n959,n77,n70);
and (n960,n76,n40);
not (n961,n927);
and (n962,n914,n952);
nand (n963,n964,n1012,n1029);
nand (n964,n398,n965);
and (n965,n966,n968,n1007);
and (n966,n297,n9,n967);
not (n967,n243);
nor (n968,n969,n994);
nor (n969,n970,n973);
or (n970,n971,n972);
and (n971,n12,n142);
and (n972,n13,n85);
xor (n973,n974,n991);
xor (n974,n975,n978);
or (n975,n976,n977);
and (n976,n14,n71);
and (n977,n15,n43);
xor (n978,n979,n987);
xor (n979,n980,n983);
nand (n980,n981,n982);
or (n981,n89,n107);
or (n982,n90,n941);
nor (n983,n72,n984);
nor (n984,n985,n986);
and (n985,n77,n105);
and (n986,n76,n103);
nor (n987,n988,n990);
and (n988,n689,n989);
not (n989,n67);
and (n990,n47,n936);
or (n991,n992,n993);
and (n992,n86,n120);
and (n993,n87,n112);
and (n994,n995,n999);
not (n995,n996);
or (n996,n997,n998);
and (n997,n974,n991);
and (n998,n975,n978);
not (n999,n1000);
xor (n1000,n1001,n1004);
xor (n1001,n1002,n1003);
not (n1002,n987);
xor (n1003,n933,n945);
or (n1004,n1005,n1006);
and (n1005,n979,n987);
and (n1006,n980,n983);
or (n1007,n1008,n1011);
or (n1008,n1009,n1010);
and (n1009,n1001,n1004);
and (n1010,n1002,n1003);
xor (n1011,n916,n931);
nand (n1012,n1013,n1007);
nand (n1013,n1014,n1023);
or (n1014,n1015,n1016);
not (n1015,n968);
not (n1016,n1017);
nand (n1017,n1018,n240);
or (n1018,n1019,n1020);
not (n1019,n9);
not (n1020,n1021);
nand (n1021,n1022,n904);
or (n1022,n900,n243);
nor (n1023,n1024,n1028);
and (n1024,n1025,n1027);
not (n1025,n1026);
nand (n1026,n970,n973);
not (n1027,n994);
nor (n1028,n995,n999);
nand (n1029,n1008,n1011);
nand (n1030,n910,n963);
and (n1032,n1031,n1033);
wire s0n1033,s1n1033,notn1033;
or (n1033,s0n1033,s1n1033);
not(notn1033,n4);
and (s0n1033,notn1033,n1034);
and (s1n1033,n4,n2334);
and (n1034,n39,n1035);
xor (n1035,n1036,n1850);
xor (n1036,n1037,n2332);
xor (n1037,n1038,n1845);
xor (n1038,n1039,n2325);
xor (n1039,n1040,n1839);
xor (n1040,n1041,n2313);
xor (n1041,n1042,n1833);
xor (n1042,n1043,n2296);
xor (n1043,n1044,n1827);
xor (n1044,n1045,n2274);
xor (n1045,n1046,n1821);
xor (n1046,n1047,n2247);
xor (n1047,n1048,n1815);
xor (n1048,n1049,n2215);
xor (n1049,n1050,n1809);
xor (n1050,n1051,n2178);
xor (n1051,n1052,n1803);
xor (n1052,n1053,n2136);
xor (n1053,n1054,n1797);
xor (n1054,n1055,n2089);
xor (n1055,n1056,n1791);
xor (n1056,n1057,n2037);
xor (n1057,n1058,n1785);
xor (n1058,n1059,n1980);
xor (n1059,n1060,n1779);
xor (n1060,n1061,n1918);
xor (n1061,n1062,n1773);
xor (n1062,n1063,n1851);
xor (n1063,n1064,n930);
xor (n1064,n1065,n1765);
xor (n1065,n1066,n1764);
xor (n1066,n1067,n1676);
xor (n1067,n1068,n1675);
xor (n1068,n1069,n1577);
xor (n1069,n1070,n1576);
xor (n1070,n1071,n1474);
xor (n1071,n1072,n1473);
xor (n1072,n1073,n1366);
xor (n1073,n1074,n1365);
xor (n1074,n1075,n1086);
xor (n1075,n1076,n1085);
xor (n1076,n1077,n1084);
xor (n1077,n1078,n1083);
xor (n1078,n1079,n1082);
xor (n1079,n1080,n1081);
and (n1080,n38,n172);
and (n1081,n38,n31);
and (n1082,n1080,n1081);
and (n1083,n38,n21);
and (n1084,n1078,n1083);
and (n1085,n38,n24);
or (n1086,n1087,n1088);
and (n1087,n1076,n1085);
and (n1088,n1075,n1089);
or (n1089,n1087,n1090);
and (n1090,n1075,n1091);
or (n1091,n1087,n1092);
and (n1092,n1075,n1093);
or (n1093,n1087,n1094);
and (n1094,n1075,n1095);
or (n1095,n1096,n1280);
and (n1096,n1097,n1279);
xor (n1097,n1077,n1098);
or (n1098,n1099,n1191);
and (n1099,n1100,n1190);
xor (n1100,n1079,n1101);
or (n1101,n1082,n1102);
and (n1102,n1103,n1105);
xor (n1103,n1080,n1104);
and (n1104,n40,n31);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
and (n1107,n40,n172);
and (n1108,n63,n31);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
and (n1113,n63,n172);
and (n1114,n109,n31);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
and (n1119,n109,n172);
and (n1120,n103,n31);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
and (n1125,n103,n172);
and (n1126,n83,n31);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
and (n1131,n83,n172);
and (n1132,n127,n31);
and (n1133,n1134,n1135);
xor (n1134,n1131,n1132);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
and (n1137,n127,n172);
and (n1138,n168,n31);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
and (n1143,n168,n172);
and (n1144,n225,n31);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
and (n1149,n225,n172);
and (n1150,n281,n31);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1156);
and (n1154,n1155,n498);
and (n1155,n281,n172);
and (n1156,n1157,n1158);
xor (n1157,n1155,n498);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
and (n1160,n332,n172);
and (n1161,n371,n31);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
and (n1166,n371,n172);
and (n1167,n434,n31);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1173);
and (n1171,n1172,n732);
and (n1172,n434,n172);
and (n1173,n1174,n1175);
xor (n1174,n1172,n732);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
and (n1177,n450,n172);
and (n1178,n444,n31);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
and (n1183,n444,n172);
and (n1184,n425,n31);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
and (n1187,n1188,n1189);
and (n1188,n425,n172);
and (n1189,n419,n31);
and (n1190,n40,n21);
and (n1191,n1192,n1193);
xor (n1192,n1100,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1103,n1105);
and (n1196,n63,n21);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1203);
and (n1200,n1201,n1202);
xor (n1201,n1110,n1111);
and (n1202,n109,n21);
and (n1203,n1204,n1205);
xor (n1204,n1201,n1202);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1116,n1117);
and (n1208,n103,n21);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1122,n1123);
and (n1214,n83,n21);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1128,n1129);
and (n1220,n127,n21);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
or (n1223,n1224,n1227);
and (n1224,n1225,n1226);
xor (n1225,n1134,n1135);
and (n1226,n168,n21);
and (n1227,n1228,n1229);
xor (n1228,n1225,n1226);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1140,n1141);
and (n1232,n225,n21);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1146,n1147);
and (n1238,n281,n21);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1152,n1153);
and (n1244,n332,n21);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1157,n1158);
and (n1250,n371,n21);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1163,n1164);
and (n1256,n434,n21);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1169,n1170);
and (n1262,n450,n21);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1174,n1175);
and (n1268,n444,n21);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1180,n1181);
and (n1274,n425,n21);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
and (n1277,n1278,n751);
xor (n1278,n1186,n1187);
and (n1279,n40,n24);
and (n1280,n1281,n1282);
xor (n1281,n1097,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1192,n1193);
and (n1285,n63,n24);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1198,n1199);
and (n1291,n109,n24);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1204,n1205);
and (n1297,n103,n24);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1210,n1211);
and (n1303,n83,n24);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1216,n1217);
and (n1309,n127,n24);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1222,n1223);
and (n1315,n168,n24);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1322);
and (n1319,n1320,n1321);
xor (n1320,n1228,n1229);
and (n1321,n225,n24);
and (n1322,n1323,n1324);
xor (n1323,n1320,n1321);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1234,n1235);
and (n1327,n281,n24);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1334);
and (n1331,n1332,n1333);
xor (n1332,n1240,n1241);
and (n1333,n332,n24);
and (n1334,n1335,n1336);
xor (n1335,n1332,n1333);
or (n1336,n1337,n1339);
and (n1337,n1338,n438);
xor (n1338,n1246,n1247);
and (n1339,n1340,n1341);
xor (n1340,n1338,n438);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1252,n1253);
and (n1344,n434,n24);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1350);
and (n1348,n1349,n565);
xor (n1349,n1258,n1259);
and (n1350,n1351,n1352);
xor (n1351,n1349,n565);
or (n1352,n1353,n1355);
and (n1353,n1354,n680);
xor (n1354,n1264,n1265);
and (n1355,n1356,n1357);
xor (n1356,n1354,n680);
or (n1357,n1358,n1360);
and (n1358,n1359,n724);
xor (n1359,n1270,n1271);
and (n1360,n1361,n1362);
xor (n1361,n1359,n724);
and (n1362,n1363,n1364);
xor (n1363,n1276,n1277);
and (n1364,n419,n24);
and (n1365,n38,n50);
or (n1366,n1367,n1369);
and (n1367,n1368,n1365);
xor (n1368,n1075,n1089);
and (n1369,n1370,n1371);
xor (n1370,n1368,n1365);
or (n1371,n1372,n1374);
and (n1372,n1373,n1365);
xor (n1373,n1075,n1091);
and (n1374,n1375,n1376);
xor (n1375,n1373,n1365);
or (n1376,n1377,n1379);
and (n1377,n1378,n1365);
xor (n1378,n1075,n1093);
and (n1379,n1380,n1381);
xor (n1380,n1378,n1365);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1075,n1095);
and (n1384,n40,n50);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1281,n1282);
and (n1390,n63,n50);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1287,n1288);
and (n1396,n109,n50);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1293,n1294);
and (n1402,n103,n50);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1299,n1300);
and (n1408,n83,n50);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1305,n1306);
and (n1414,n127,n50);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1311,n1312);
and (n1420,n168,n50);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1317,n1318);
and (n1426,n225,n50);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1323,n1324);
and (n1432,n281,n50);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1329,n1330);
and (n1438,n332,n50);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1335,n1336);
and (n1444,n371,n50);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1340,n1341);
and (n1450,n434,n50);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1346,n1347);
and (n1456,n450,n50);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
or (n1459,n1460,n1463);
and (n1460,n1461,n1462);
xor (n1461,n1351,n1352);
and (n1462,n444,n50);
and (n1463,n1464,n1465);
xor (n1464,n1461,n1462);
or (n1465,n1466,n1469);
and (n1466,n1467,n1468);
xor (n1467,n1356,n1357);
and (n1468,n425,n50);
and (n1469,n1470,n1471);
xor (n1470,n1467,n1468);
and (n1471,n1472,n697);
xor (n1472,n1361,n1362);
and (n1473,n38,n56);
or (n1474,n1475,n1477);
and (n1475,n1476,n1473);
xor (n1476,n1370,n1371);
and (n1477,n1478,n1479);
xor (n1478,n1476,n1473);
or (n1479,n1480,n1482);
and (n1480,n1481,n1473);
xor (n1481,n1375,n1376);
and (n1482,n1483,n1484);
xor (n1483,n1481,n1473);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1380,n1381);
and (n1487,n40,n56);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1386,n1387);
and (n1493,n63,n56);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1392,n1393);
and (n1499,n109,n56);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1398,n1399);
and (n1505,n103,n56);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1404,n1405);
and (n1511,n83,n56);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1410,n1411);
and (n1517,n127,n56);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
or (n1520,n1521,n1524);
and (n1521,n1522,n1523);
xor (n1522,n1416,n1417);
and (n1523,n168,n56);
and (n1524,n1525,n1526);
xor (n1525,n1522,n1523);
or (n1526,n1527,n1530);
and (n1527,n1528,n1529);
xor (n1528,n1422,n1423);
and (n1529,n225,n56);
and (n1530,n1531,n1532);
xor (n1531,n1528,n1529);
or (n1532,n1533,n1536);
and (n1533,n1534,n1535);
xor (n1534,n1428,n1429);
and (n1535,n281,n56);
and (n1536,n1537,n1538);
xor (n1537,n1534,n1535);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1434,n1435);
and (n1541,n332,n56);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
or (n1544,n1545,n1548);
and (n1545,n1546,n1547);
xor (n1546,n1440,n1441);
and (n1547,n371,n56);
and (n1548,n1549,n1550);
xor (n1549,n1546,n1547);
or (n1550,n1551,n1554);
and (n1551,n1552,n1553);
xor (n1552,n1446,n1447);
and (n1553,n434,n56);
and (n1554,n1555,n1556);
xor (n1555,n1552,n1553);
or (n1556,n1557,n1560);
and (n1557,n1558,n1559);
xor (n1558,n1452,n1453);
and (n1559,n450,n56);
and (n1560,n1561,n1562);
xor (n1561,n1558,n1559);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
xor (n1564,n1458,n1459);
and (n1565,n444,n56);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
or (n1568,n1569,n1571);
and (n1569,n1570,n686);
xor (n1570,n1464,n1465);
and (n1571,n1572,n1573);
xor (n1572,n1570,n686);
and (n1573,n1574,n1575);
xor (n1574,n1470,n1471);
and (n1575,n419,n56);
and (n1576,n38,n93);
or (n1577,n1578,n1580);
and (n1578,n1579,n1576);
xor (n1579,n1478,n1479);
and (n1580,n1581,n1582);
xor (n1581,n1579,n1576);
or (n1582,n1583,n1586);
and (n1583,n1584,n1585);
xor (n1584,n1483,n1484);
and (n1585,n40,n93);
and (n1586,n1587,n1588);
xor (n1587,n1584,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n1489,n1490);
and (n1591,n63,n93);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1495,n1496);
and (n1597,n109,n93);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1501,n1502);
and (n1603,n103,n93);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1507,n1508);
and (n1609,n83,n93);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1513,n1514);
and (n1615,n127,n93);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1519,n1520);
and (n1621,n168,n93);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1525,n1526);
and (n1627,n225,n93);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1531,n1532);
and (n1633,n281,n93);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1537,n1538);
and (n1639,n332,n93);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1543,n1544);
and (n1645,n371,n93);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1549,n1550);
and (n1651,n434,n93);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1555,n1556);
and (n1657,n450,n93);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1561,n1562);
and (n1663,n444,n93);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1567,n1568);
and (n1669,n425,n93);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
and (n1672,n1673,n1674);
xor (n1673,n1572,n1573);
not (n1674,n492);
and (n1675,n38,n73);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1581,n1582);
and (n1679,n40,n73);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1587,n1588);
and (n1685,n63,n73);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1593,n1594);
and (n1691,n109,n73);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1599,n1600);
and (n1697,n103,n73);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1605,n1606);
and (n1703,n83,n73);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1611,n1612);
and (n1709,n127,n73);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1715);
and (n1713,n1714,n218);
xor (n1714,n1617,n1618);
and (n1715,n1716,n1717);
xor (n1716,n1714,n218);
or (n1717,n1718,n1720);
and (n1718,n1719,n273);
xor (n1719,n1623,n1624);
and (n1720,n1721,n1722);
xor (n1721,n1719,n273);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
xor (n1724,n1629,n1630);
and (n1725,n281,n73);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
or (n1728,n1729,n1732);
and (n1729,n1730,n1731);
xor (n1730,n1635,n1636);
and (n1731,n332,n73);
and (n1732,n1733,n1734);
xor (n1733,n1730,n1731);
or (n1734,n1735,n1737);
and (n1735,n1736,n629);
xor (n1736,n1641,n1642);
and (n1737,n1738,n1739);
xor (n1738,n1736,n629);
or (n1739,n1740,n1742);
and (n1740,n1741,n582);
xor (n1741,n1647,n1648);
and (n1742,n1743,n1744);
xor (n1743,n1741,n582);
or (n1744,n1745,n1747);
and (n1745,n1746,n511);
xor (n1746,n1653,n1654);
and (n1747,n1748,n1749);
xor (n1748,n1746,n511);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
xor (n1751,n1659,n1660);
and (n1752,n444,n73);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
or (n1755,n1756,n1759);
and (n1756,n1757,n1758);
xor (n1757,n1665,n1666);
and (n1758,n425,n73);
and (n1759,n1760,n1761);
xor (n1760,n1757,n1758);
and (n1761,n1762,n1763);
xor (n1762,n1671,n1672);
and (n1763,n419,n73);
and (n1764,n40,n77);
or (n1765,n1766,n1768);
and (n1766,n1767,n930);
xor (n1767,n1681,n1682);
and (n1768,n1769,n1770);
xor (n1769,n1767,n930);
or (n1770,n1771,n1774);
and (n1771,n1772,n1773);
xor (n1772,n1687,n1688);
and (n1773,n109,n77);
and (n1774,n1775,n1776);
xor (n1775,n1772,n1773);
or (n1776,n1777,n1780);
and (n1777,n1778,n1779);
xor (n1778,n1693,n1694);
and (n1779,n103,n77);
and (n1780,n1781,n1782);
xor (n1781,n1778,n1779);
or (n1782,n1783,n1786);
and (n1783,n1784,n1785);
xor (n1784,n1699,n1700);
and (n1785,n83,n77);
and (n1786,n1787,n1788);
xor (n1787,n1784,n1785);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1705,n1706);
and (n1791,n127,n77);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1711,n1712);
and (n1797,n168,n77);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
xor (n1802,n1716,n1717);
and (n1803,n225,n77);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
xor (n1808,n1721,n1722);
and (n1809,n281,n77);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
xor (n1814,n1727,n1728);
and (n1815,n332,n77);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
xor (n1820,n1733,n1734);
and (n1821,n371,n77);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
xor (n1826,n1738,n1739);
and (n1827,n434,n77);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1743,n1744);
and (n1833,n450,n77);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1748,n1749);
and (n1839,n444,n77);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1754,n1755);
and (n1845,n425,n77);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
and (n1848,n1849,n1850);
xor (n1849,n1760,n1761);
and (n1850,n419,n77);
or (n1851,n1852,n1854);
and (n1852,n1853,n1773);
xor (n1853,n1769,n1770);
and (n1854,n1855,n1856);
xor (n1855,n1853,n1773);
or (n1856,n1857,n1859);
and (n1857,n1858,n1779);
xor (n1858,n1775,n1776);
and (n1859,n1860,n1861);
xor (n1860,n1858,n1779);
or (n1861,n1862,n1864);
and (n1862,n1863,n1785);
xor (n1863,n1781,n1782);
and (n1864,n1865,n1866);
xor (n1865,n1863,n1785);
or (n1866,n1867,n1869);
and (n1867,n1868,n1791);
xor (n1868,n1787,n1788);
and (n1869,n1870,n1871);
xor (n1870,n1868,n1791);
or (n1871,n1872,n1874);
and (n1872,n1873,n1797);
xor (n1873,n1793,n1794);
and (n1874,n1875,n1876);
xor (n1875,n1873,n1797);
or (n1876,n1877,n1879);
and (n1877,n1878,n1803);
xor (n1878,n1799,n1800);
and (n1879,n1880,n1881);
xor (n1880,n1878,n1803);
or (n1881,n1882,n1884);
and (n1882,n1883,n1809);
xor (n1883,n1805,n1806);
and (n1884,n1885,n1886);
xor (n1885,n1883,n1809);
or (n1886,n1887,n1889);
and (n1887,n1888,n1815);
xor (n1888,n1811,n1812);
and (n1889,n1890,n1891);
xor (n1890,n1888,n1815);
or (n1891,n1892,n1894);
and (n1892,n1893,n1821);
xor (n1893,n1817,n1818);
and (n1894,n1895,n1896);
xor (n1895,n1893,n1821);
or (n1896,n1897,n1899);
and (n1897,n1898,n1827);
xor (n1898,n1823,n1824);
and (n1899,n1900,n1901);
xor (n1900,n1898,n1827);
or (n1901,n1902,n1904);
and (n1902,n1903,n1833);
xor (n1903,n1829,n1830);
and (n1904,n1905,n1906);
xor (n1905,n1903,n1833);
or (n1906,n1907,n1909);
and (n1907,n1908,n1839);
xor (n1908,n1835,n1836);
and (n1909,n1910,n1911);
xor (n1910,n1908,n1839);
or (n1911,n1912,n1914);
and (n1912,n1913,n1845);
xor (n1913,n1841,n1842);
and (n1914,n1915,n1916);
xor (n1915,n1913,n1845);
and (n1916,n1917,n1850);
xor (n1917,n1847,n1848);
or (n1918,n1919,n1921);
and (n1919,n1920,n1779);
xor (n1920,n1855,n1856);
and (n1921,n1922,n1923);
xor (n1922,n1920,n1779);
or (n1923,n1924,n1926);
and (n1924,n1925,n1785);
xor (n1925,n1860,n1861);
and (n1926,n1927,n1928);
xor (n1927,n1925,n1785);
or (n1928,n1929,n1931);
and (n1929,n1930,n1791);
xor (n1930,n1865,n1866);
and (n1931,n1932,n1933);
xor (n1932,n1930,n1791);
or (n1933,n1934,n1936);
and (n1934,n1935,n1797);
xor (n1935,n1870,n1871);
and (n1936,n1937,n1938);
xor (n1937,n1935,n1797);
or (n1938,n1939,n1941);
and (n1939,n1940,n1803);
xor (n1940,n1875,n1876);
and (n1941,n1942,n1943);
xor (n1942,n1940,n1803);
or (n1943,n1944,n1946);
and (n1944,n1945,n1809);
xor (n1945,n1880,n1881);
and (n1946,n1947,n1948);
xor (n1947,n1945,n1809);
or (n1948,n1949,n1951);
and (n1949,n1950,n1815);
xor (n1950,n1885,n1886);
and (n1951,n1952,n1953);
xor (n1952,n1950,n1815);
or (n1953,n1954,n1956);
and (n1954,n1955,n1821);
xor (n1955,n1890,n1891);
and (n1956,n1957,n1958);
xor (n1957,n1955,n1821);
or (n1958,n1959,n1961);
and (n1959,n1960,n1827);
xor (n1960,n1895,n1896);
and (n1961,n1962,n1963);
xor (n1962,n1960,n1827);
or (n1963,n1964,n1966);
and (n1964,n1965,n1833);
xor (n1965,n1900,n1901);
and (n1966,n1967,n1968);
xor (n1967,n1965,n1833);
or (n1968,n1969,n1971);
and (n1969,n1970,n1839);
xor (n1970,n1905,n1906);
and (n1971,n1972,n1973);
xor (n1972,n1970,n1839);
or (n1973,n1974,n1976);
and (n1974,n1975,n1845);
xor (n1975,n1910,n1911);
and (n1976,n1977,n1978);
xor (n1977,n1975,n1845);
and (n1978,n1979,n1850);
xor (n1979,n1915,n1916);
or (n1980,n1981,n1983);
and (n1981,n1982,n1785);
xor (n1982,n1922,n1923);
and (n1983,n1984,n1985);
xor (n1984,n1982,n1785);
or (n1985,n1986,n1988);
and (n1986,n1987,n1791);
xor (n1987,n1927,n1928);
and (n1988,n1989,n1990);
xor (n1989,n1987,n1791);
or (n1990,n1991,n1993);
and (n1991,n1992,n1797);
xor (n1992,n1932,n1933);
and (n1993,n1994,n1995);
xor (n1994,n1992,n1797);
or (n1995,n1996,n1998);
and (n1996,n1997,n1803);
xor (n1997,n1937,n1938);
and (n1998,n1999,n2000);
xor (n1999,n1997,n1803);
or (n2000,n2001,n2003);
and (n2001,n2002,n1809);
xor (n2002,n1942,n1943);
and (n2003,n2004,n2005);
xor (n2004,n2002,n1809);
or (n2005,n2006,n2008);
and (n2006,n2007,n1815);
xor (n2007,n1947,n1948);
and (n2008,n2009,n2010);
xor (n2009,n2007,n1815);
or (n2010,n2011,n2013);
and (n2011,n2012,n1821);
xor (n2012,n1952,n1953);
and (n2013,n2014,n2015);
xor (n2014,n2012,n1821);
or (n2015,n2016,n2018);
and (n2016,n2017,n1827);
xor (n2017,n1957,n1958);
and (n2018,n2019,n2020);
xor (n2019,n2017,n1827);
or (n2020,n2021,n2023);
and (n2021,n2022,n1833);
xor (n2022,n1962,n1963);
and (n2023,n2024,n2025);
xor (n2024,n2022,n1833);
or (n2025,n2026,n2028);
and (n2026,n2027,n1839);
xor (n2027,n1967,n1968);
and (n2028,n2029,n2030);
xor (n2029,n2027,n1839);
or (n2030,n2031,n2033);
and (n2031,n2032,n1845);
xor (n2032,n1972,n1973);
and (n2033,n2034,n2035);
xor (n2034,n2032,n1845);
and (n2035,n2036,n1850);
xor (n2036,n1977,n1978);
or (n2037,n2038,n2040);
and (n2038,n2039,n1791);
xor (n2039,n1984,n1985);
and (n2040,n2041,n2042);
xor (n2041,n2039,n1791);
or (n2042,n2043,n2045);
and (n2043,n2044,n1797);
xor (n2044,n1989,n1990);
and (n2045,n2046,n2047);
xor (n2046,n2044,n1797);
or (n2047,n2048,n2050);
and (n2048,n2049,n1803);
xor (n2049,n1994,n1995);
and (n2050,n2051,n2052);
xor (n2051,n2049,n1803);
or (n2052,n2053,n2055);
and (n2053,n2054,n1809);
xor (n2054,n1999,n2000);
and (n2055,n2056,n2057);
xor (n2056,n2054,n1809);
or (n2057,n2058,n2060);
and (n2058,n2059,n1815);
xor (n2059,n2004,n2005);
and (n2060,n2061,n2062);
xor (n2061,n2059,n1815);
or (n2062,n2063,n2065);
and (n2063,n2064,n1821);
xor (n2064,n2009,n2010);
and (n2065,n2066,n2067);
xor (n2066,n2064,n1821);
or (n2067,n2068,n2070);
and (n2068,n2069,n1827);
xor (n2069,n2014,n2015);
and (n2070,n2071,n2072);
xor (n2071,n2069,n1827);
or (n2072,n2073,n2075);
and (n2073,n2074,n1833);
xor (n2074,n2019,n2020);
and (n2075,n2076,n2077);
xor (n2076,n2074,n1833);
or (n2077,n2078,n2080);
and (n2078,n2079,n1839);
xor (n2079,n2024,n2025);
and (n2080,n2081,n2082);
xor (n2081,n2079,n1839);
or (n2082,n2083,n2085);
and (n2083,n2084,n1845);
xor (n2084,n2029,n2030);
and (n2085,n2086,n2087);
xor (n2086,n2084,n1845);
and (n2087,n2088,n1850);
xor (n2088,n2034,n2035);
or (n2089,n2090,n2092);
and (n2090,n2091,n1797);
xor (n2091,n2041,n2042);
and (n2092,n2093,n2094);
xor (n2093,n2091,n1797);
or (n2094,n2095,n2097);
and (n2095,n2096,n1803);
xor (n2096,n2046,n2047);
and (n2097,n2098,n2099);
xor (n2098,n2096,n1803);
or (n2099,n2100,n2102);
and (n2100,n2101,n1809);
xor (n2101,n2051,n2052);
and (n2102,n2103,n2104);
xor (n2103,n2101,n1809);
or (n2104,n2105,n2107);
and (n2105,n2106,n1815);
xor (n2106,n2056,n2057);
and (n2107,n2108,n2109);
xor (n2108,n2106,n1815);
or (n2109,n2110,n2112);
and (n2110,n2111,n1821);
xor (n2111,n2061,n2062);
and (n2112,n2113,n2114);
xor (n2113,n2111,n1821);
or (n2114,n2115,n2117);
and (n2115,n2116,n1827);
xor (n2116,n2066,n2067);
and (n2117,n2118,n2119);
xor (n2118,n2116,n1827);
or (n2119,n2120,n2122);
and (n2120,n2121,n1833);
xor (n2121,n2071,n2072);
and (n2122,n2123,n2124);
xor (n2123,n2121,n1833);
or (n2124,n2125,n2127);
and (n2125,n2126,n1839);
xor (n2126,n2076,n2077);
and (n2127,n2128,n2129);
xor (n2128,n2126,n1839);
or (n2129,n2130,n2132);
and (n2130,n2131,n1845);
xor (n2131,n2081,n2082);
and (n2132,n2133,n2134);
xor (n2133,n2131,n1845);
and (n2134,n2135,n1850);
xor (n2135,n2086,n2087);
or (n2136,n2137,n2139);
and (n2137,n2138,n1803);
xor (n2138,n2093,n2094);
and (n2139,n2140,n2141);
xor (n2140,n2138,n1803);
or (n2141,n2142,n2144);
and (n2142,n2143,n1809);
xor (n2143,n2098,n2099);
and (n2144,n2145,n2146);
xor (n2145,n2143,n1809);
or (n2146,n2147,n2149);
and (n2147,n2148,n1815);
xor (n2148,n2103,n2104);
and (n2149,n2150,n2151);
xor (n2150,n2148,n1815);
or (n2151,n2152,n2154);
and (n2152,n2153,n1821);
xor (n2153,n2108,n2109);
and (n2154,n2155,n2156);
xor (n2155,n2153,n1821);
or (n2156,n2157,n2159);
and (n2157,n2158,n1827);
xor (n2158,n2113,n2114);
and (n2159,n2160,n2161);
xor (n2160,n2158,n1827);
or (n2161,n2162,n2164);
and (n2162,n2163,n1833);
xor (n2163,n2118,n2119);
and (n2164,n2165,n2166);
xor (n2165,n2163,n1833);
or (n2166,n2167,n2169);
and (n2167,n2168,n1839);
xor (n2168,n2123,n2124);
and (n2169,n2170,n2171);
xor (n2170,n2168,n1839);
or (n2171,n2172,n2174);
and (n2172,n2173,n1845);
xor (n2173,n2128,n2129);
and (n2174,n2175,n2176);
xor (n2175,n2173,n1845);
and (n2176,n2177,n1850);
xor (n2177,n2133,n2134);
or (n2178,n2179,n2181);
and (n2179,n2180,n1809);
xor (n2180,n2140,n2141);
and (n2181,n2182,n2183);
xor (n2182,n2180,n1809);
or (n2183,n2184,n2186);
and (n2184,n2185,n1815);
xor (n2185,n2145,n2146);
and (n2186,n2187,n2188);
xor (n2187,n2185,n1815);
or (n2188,n2189,n2191);
and (n2189,n2190,n1821);
xor (n2190,n2150,n2151);
and (n2191,n2192,n2193);
xor (n2192,n2190,n1821);
or (n2193,n2194,n2196);
and (n2194,n2195,n1827);
xor (n2195,n2155,n2156);
and (n2196,n2197,n2198);
xor (n2197,n2195,n1827);
or (n2198,n2199,n2201);
and (n2199,n2200,n1833);
xor (n2200,n2160,n2161);
and (n2201,n2202,n2203);
xor (n2202,n2200,n1833);
or (n2203,n2204,n2206);
and (n2204,n2205,n1839);
xor (n2205,n2165,n2166);
and (n2206,n2207,n2208);
xor (n2207,n2205,n1839);
or (n2208,n2209,n2211);
and (n2209,n2210,n1845);
xor (n2210,n2170,n2171);
and (n2211,n2212,n2213);
xor (n2212,n2210,n1845);
and (n2213,n2214,n1850);
xor (n2214,n2175,n2176);
or (n2215,n2216,n2218);
and (n2216,n2217,n1815);
xor (n2217,n2182,n2183);
and (n2218,n2219,n2220);
xor (n2219,n2217,n1815);
or (n2220,n2221,n2223);
and (n2221,n2222,n1821);
xor (n2222,n2187,n2188);
and (n2223,n2224,n2225);
xor (n2224,n2222,n1821);
or (n2225,n2226,n2228);
and (n2226,n2227,n1827);
xor (n2227,n2192,n2193);
and (n2228,n2229,n2230);
xor (n2229,n2227,n1827);
or (n2230,n2231,n2233);
and (n2231,n2232,n1833);
xor (n2232,n2197,n2198);
and (n2233,n2234,n2235);
xor (n2234,n2232,n1833);
or (n2235,n2236,n2238);
and (n2236,n2237,n1839);
xor (n2237,n2202,n2203);
and (n2238,n2239,n2240);
xor (n2239,n2237,n1839);
or (n2240,n2241,n2243);
and (n2241,n2242,n1845);
xor (n2242,n2207,n2208);
and (n2243,n2244,n2245);
xor (n2244,n2242,n1845);
and (n2245,n2246,n1850);
xor (n2246,n2212,n2213);
or (n2247,n2248,n2250);
and (n2248,n2249,n1821);
xor (n2249,n2219,n2220);
and (n2250,n2251,n2252);
xor (n2251,n2249,n1821);
or (n2252,n2253,n2255);
and (n2253,n2254,n1827);
xor (n2254,n2224,n2225);
and (n2255,n2256,n2257);
xor (n2256,n2254,n1827);
or (n2257,n2258,n2260);
and (n2258,n2259,n1833);
xor (n2259,n2229,n2230);
and (n2260,n2261,n2262);
xor (n2261,n2259,n1833);
or (n2262,n2263,n2265);
and (n2263,n2264,n1839);
xor (n2264,n2234,n2235);
and (n2265,n2266,n2267);
xor (n2266,n2264,n1839);
or (n2267,n2268,n2270);
and (n2268,n2269,n1845);
xor (n2269,n2239,n2240);
and (n2270,n2271,n2272);
xor (n2271,n2269,n1845);
and (n2272,n2273,n1850);
xor (n2273,n2244,n2245);
or (n2274,n2275,n2277);
and (n2275,n2276,n1827);
xor (n2276,n2251,n2252);
and (n2277,n2278,n2279);
xor (n2278,n2276,n1827);
or (n2279,n2280,n2282);
and (n2280,n2281,n1833);
xor (n2281,n2256,n2257);
and (n2282,n2283,n2284);
xor (n2283,n2281,n1833);
or (n2284,n2285,n2287);
and (n2285,n2286,n1839);
xor (n2286,n2261,n2262);
and (n2287,n2288,n2289);
xor (n2288,n2286,n1839);
or (n2289,n2290,n2292);
and (n2290,n2291,n1845);
xor (n2291,n2266,n2267);
and (n2292,n2293,n2294);
xor (n2293,n2291,n1845);
and (n2294,n2295,n1850);
xor (n2295,n2271,n2272);
or (n2296,n2297,n2299);
and (n2297,n2298,n1833);
xor (n2298,n2278,n2279);
and (n2299,n2300,n2301);
xor (n2300,n2298,n1833);
or (n2301,n2302,n2304);
and (n2302,n2303,n1839);
xor (n2303,n2283,n2284);
and (n2304,n2305,n2306);
xor (n2305,n2303,n1839);
or (n2306,n2307,n2309);
and (n2307,n2308,n1845);
xor (n2308,n2288,n2289);
and (n2309,n2310,n2311);
xor (n2310,n2308,n1845);
and (n2311,n2312,n1850);
xor (n2312,n2293,n2294);
or (n2313,n2314,n2316);
and (n2314,n2315,n1839);
xor (n2315,n2300,n2301);
and (n2316,n2317,n2318);
xor (n2317,n2315,n1839);
or (n2318,n2319,n2321);
and (n2319,n2320,n1845);
xor (n2320,n2305,n2306);
and (n2321,n2322,n2323);
xor (n2322,n2320,n1845);
and (n2323,n2324,n1850);
xor (n2324,n2310,n2311);
or (n2325,n2326,n2328);
and (n2326,n2327,n1845);
xor (n2327,n2317,n2318);
and (n2328,n2329,n2330);
xor (n2329,n2327,n1845);
and (n2330,n2331,n1850);
xor (n2331,n2322,n2323);
and (n2332,n2333,n1850);
xor (n2333,n2329,n2330);
xor (n2334,n2312,n1850);
endmodule
