module top (out,n17,n19,n26,n27,n37,n45,n46,n52,n53
        ,n61,n73,n78,n82,n88,n97,n98,n100,n105,n106
        ,n110,n117,n125,n131,n140,n151,n157,n166,n174,n176
        ,n181,n187,n201,n212,n219,n1078);
output out;
input n17;
input n19;
input n26;
input n27;
input n37;
input n45;
input n46;
input n52;
input n53;
input n61;
input n73;
input n78;
input n82;
input n88;
input n97;
input n98;
input n100;
input n105;
input n106;
input n110;
input n117;
input n125;
input n131;
input n140;
input n151;
input n157;
input n166;
input n174;
input n176;
input n181;
input n187;
input n201;
input n212;
input n219;
input n1078;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
xor (out,n0,n1108);
nand (n0,n1,n1107);
or (n1,n2,n1008);
nand (n2,n3,n1007);
or (n3,n4,n494);
nor (n4,n5,n433);
xor (n5,n6,n363);
xor (n6,n7,n221);
xor (n7,n8,n143);
xor (n8,n9,n91);
xor (n9,n10,n67);
xor (n10,n11,n39);
nand (n11,n12,n33);
or (n12,n13,n21);
not (n13,n14);
nor (n14,n15,n20);
and (n15,n16,n18);
not (n16,n17);
not (n18,n19);
and (n20,n17,n19);
not (n21,n22);
nor (n22,n23,n29);
nand (n23,n24,n28);
or (n24,n25,n27);
not (n25,n26);
nand (n28,n27,n25);
nor (n29,n30,n32);
and (n30,n31,n19);
not (n31,n27);
and (n32,n27,n18);
nand (n33,n23,n34);
nand (n34,n35,n38);
or (n35,n36,n19);
not (n36,n37);
or (n38,n18,n37);
nand (n39,n40,n56);
or (n40,n41,n48);
not (n41,n42);
nand (n42,n43,n47);
or (n43,n44,n46);
not (n44,n45);
nand (n47,n46,n44);
not (n48,n49);
nand (n49,n50,n54);
or (n50,n51,n53);
not (n51,n52);
or (n54,n55,n52);
not (n55,n53);
nand (n56,n57,n63);
not (n57,n58);
nor (n58,n59,n62);
and (n59,n53,n60);
not (n60,n61);
and (n62,n55,n61);
and (n63,n41,n64);
nand (n64,n65,n66);
nand (n65,n53,n44);
nand (n66,n45,n55);
nand (n67,n68,n85);
or (n68,n69,n80);
nand (n69,n70,n75);
nor (n70,n71,n74);
and (n71,n72,n53);
not (n72,n73);
and (n74,n73,n55);
nor (n75,n76,n79);
and (n76,n72,n77);
not (n77,n78);
and (n79,n73,n78);
nor (n80,n81,n83);
and (n81,n82,n77);
and (n83,n78,n84);
not (n84,n82);
or (n85,n86,n70);
nor (n86,n87,n89);
and (n87,n88,n77);
and (n89,n78,n90);
not (n90,n88);
xor (n91,n92,n119);
xor (n92,n93,n101);
and (n93,n94,n100);
nand (n94,n95,n99);
or (n95,n96,n98);
not (n96,n97);
nand (n99,n98,n96);
nand (n101,n102,n113);
or (n102,n103,n107);
nand (n103,n104,n106);
not (n104,n105);
nor (n107,n108,n111);
and (n108,n109,n110);
not (n109,n106);
and (n111,n106,n112);
not (n112,n110);
nand (n113,n114,n105);
nor (n114,n115,n118);
and (n115,n116,n109);
not (n116,n117);
and (n118,n117,n106);
nand (n119,n120,n133);
or (n120,n121,n127);
not (n121,n122);
nor (n122,n123,n126);
and (n123,n124,n25);
not (n124,n125);
and (n126,n125,n26);
not (n127,n128);
nand (n128,n129,n132);
or (n129,n130,n106);
not (n130,n131);
nand (n132,n106,n130);
or (n133,n134,n138);
nand (n134,n127,n135);
nand (n135,n136,n137);
or (n136,n130,n26);
nand (n137,n130,n26);
nor (n138,n139,n141);
and (n139,n25,n140);
and (n141,n26,n142);
not (n142,n140);
xor (n143,n144,n195);
xor (n144,n145,n168);
nand (n145,n146,n162);
or (n146,n147,n153);
not (n147,n148);
nor (n148,n149,n152);
and (n149,n150,n96);
not (n150,n151);
and (n152,n151,n97);
nand (n153,n154,n159);
not (n154,n155);
nand (n155,n156,n158);
or (n156,n77,n157);
nand (n158,n77,n157);
nand (n159,n160,n161);
or (n160,n157,n96);
nand (n161,n96,n157);
nand (n162,n155,n163);
nor (n163,n164,n167);
and (n164,n165,n96);
not (n165,n166);
and (n167,n166,n97);
nand (n168,n169,n183);
or (n169,n170,n178);
not (n170,n171);
nor (n171,n172,n177);
and (n172,n173,n175);
not (n173,n174);
not (n175,n176);
and (n177,n174,n176);
not (n178,n179);
nand (n179,n180,n182);
or (n180,n18,n181);
nand (n182,n181,n18);
nand (n183,n184,n190);
not (n184,n185);
nor (n185,n186,n188);
and (n186,n175,n187);
and (n188,n176,n189);
not (n189,n187);
not (n190,n191);
nand (n191,n178,n192);
nand (n192,n193,n194);
or (n193,n181,n175);
nand (n194,n175,n181);
nand (n195,n196,n214);
or (n196,n197,n208);
not (n197,n198);
nor (n198,n199,n203);
nand (n199,n200,n202);
or (n200,n175,n201);
nand (n202,n201,n175);
nor (n203,n204,n206);
and (n204,n205,n201);
not (n205,n46);
and (n206,n46,n207);
not (n207,n201);
not (n208,n209);
nor (n209,n210,n213);
and (n210,n211,n205);
not (n211,n212);
and (n213,n212,n46);
or (n214,n215,n216);
not (n215,n199);
nor (n216,n217,n220);
and (n217,n218,n46);
not (n218,n219);
and (n220,n219,n205);
or (n221,n222,n362);
and (n222,n223,n301);
xor (n223,n224,n264);
or (n224,n225,n263);
and (n225,n226,n246);
xor (n226,n227,n237);
nand (n227,n228,n233);
or (n228,n229,n230);
not (n229,n63);
nor (n230,n231,n232);
and (n231,n55,n82);
and (n232,n53,n84);
or (n233,n41,n234);
nor (n234,n235,n236);
and (n235,n55,n88);
and (n236,n53,n90);
nand (n237,n238,n242);
or (n238,n69,n239);
nor (n239,n240,n241);
and (n240,n77,n151);
and (n241,n78,n150);
or (n242,n70,n243);
nor (n243,n244,n245);
and (n244,n77,n166);
and (n245,n78,n165);
and (n246,n247,n253);
nor (n247,n248,n77);
nor (n248,n249,n251);
and (n249,n250,n55);
nand (n250,n100,n73);
and (n251,n252,n72);
not (n252,n100);
nand (n253,n254,n259);
or (n254,n103,n255);
not (n255,n256);
nor (n256,n257,n258);
and (n257,n36,n109);
and (n258,n37,n106);
or (n259,n260,n104);
nor (n260,n261,n262);
and (n261,n109,n140);
and (n262,n106,n142);
and (n263,n227,n237);
xor (n264,n265,n283);
xor (n265,n266,n269);
nand (n266,n267,n268);
or (n267,n69,n243);
or (n268,n70,n80);
xor (n269,n270,n276);
nor (n270,n271,n96);
nor (n271,n272,n274);
and (n272,n273,n77);
nand (n273,n100,n157);
and (n274,n252,n275);
not (n275,n157);
nand (n276,n277,n282);
or (n277,n103,n278);
not (n278,n279);
nor (n279,n280,n281);
and (n280,n125,n106);
and (n281,n124,n109);
or (n282,n107,n104);
or (n283,n284,n300);
and (n284,n285,n290);
xor (n285,n286,n287);
nor (n286,n154,n252);
nand (n287,n288,n289);
or (n288,n104,n278);
or (n289,n260,n103);
nand (n290,n291,n295);
or (n291,n134,n292);
nor (n292,n293,n294);
and (n293,n17,n25);
and (n294,n16,n26);
or (n295,n127,n296);
not (n296,n297);
nor (n297,n298,n299);
and (n298,n37,n26);
and (n299,n36,n25);
and (n300,n286,n287);
or (n301,n302,n361);
and (n302,n303,n360);
xor (n303,n304,n334);
or (n304,n305,n333);
and (n305,n306,n324);
xor (n306,n307,n314);
nand (n307,n308,n312);
or (n308,n134,n309);
nor (n309,n310,n311);
and (n310,n174,n25);
and (n311,n173,n26);
nand (n312,n313,n128);
not (n313,n292);
nand (n314,n315,n320);
or (n315,n316,n178);
not (n316,n317);
nor (n317,n318,n319);
and (n318,n212,n176);
and (n319,n211,n175);
or (n320,n191,n321);
nor (n321,n322,n323);
and (n322,n51,n176);
and (n323,n52,n175);
nand (n324,n325,n329);
or (n325,n197,n326);
nor (n326,n327,n328);
and (n327,n205,n88);
and (n328,n90,n46);
or (n329,n215,n330);
nor (n330,n331,n332);
and (n331,n205,n61);
and (n332,n46,n60);
and (n333,n307,n314);
or (n334,n335,n359);
and (n335,n336,n353);
xor (n336,n337,n347);
nand (n337,n338,n342);
or (n338,n339,n21);
nor (n339,n340,n341);
and (n340,n18,n219);
and (n341,n19,n218);
nand (n342,n343,n23);
not (n343,n344);
nor (n344,n345,n346);
and (n345,n18,n187);
and (n346,n19,n189);
nand (n347,n348,n352);
or (n348,n229,n349);
nor (n349,n350,n351);
and (n350,n55,n166);
and (n351,n53,n165);
or (n352,n41,n230);
nand (n353,n354,n358);
or (n354,n69,n355);
nor (n355,n356,n357);
and (n356,n252,n78);
and (n357,n100,n77);
or (n358,n239,n70);
and (n359,n337,n347);
xor (n360,n285,n290);
and (n361,n304,n334);
and (n362,n224,n264);
xor (n363,n364,n414);
xor (n364,n365,n368);
or (n365,n366,n367);
and (n366,n265,n283);
and (n367,n266,n269);
xor (n368,n369,n393);
xor (n369,n370,n371);
and (n370,n270,n276);
or (n371,n372,n392);
and (n372,n373,n385);
xor (n373,n374,n378);
nand (n374,n375,n376);
or (n375,n296,n134);
nand (n376,n377,n128);
not (n377,n138);
nand (n378,n379,n384);
or (n379,n380,n153);
not (n380,n381);
nand (n381,n382,n383);
or (n382,n96,n100);
or (n383,n252,n97);
nand (n384,n155,n148);
nand (n385,n386,n391);
or (n386,n191,n387);
not (n387,n388);
nor (n388,n389,n390);
and (n389,n219,n176);
and (n390,n218,n175);
or (n391,n178,n185);
and (n392,n374,n378);
or (n393,n394,n413);
and (n394,n395,n410);
xor (n395,n396,n403);
nand (n396,n397,n402);
or (n397,n398,n197);
not (n398,n399);
nor (n399,n400,n401);
and (n400,n51,n205);
and (n401,n52,n46);
nand (n402,n199,n209);
nand (n403,n404,n406);
or (n404,n13,n405);
not (n405,n23);
or (n406,n21,n407);
nor (n407,n408,n409);
and (n408,n18,n174);
and (n409,n19,n173);
nand (n410,n411,n412);
or (n411,n229,n234);
or (n412,n41,n58);
and (n413,n396,n403);
or (n414,n415,n432);
and (n415,n416,n431);
xor (n416,n417,n430);
or (n417,n418,n429);
and (n418,n419,n426);
xor (n419,n420,n423);
nand (n420,n421,n422);
or (n421,n316,n191);
nand (n422,n179,n388);
nand (n423,n424,n425);
or (n424,n197,n330);
nand (n425,n199,n399);
nand (n426,n427,n428);
or (n427,n21,n344);
or (n428,n405,n407);
and (n429,n420,n423);
xor (n430,n395,n410);
xor (n431,n373,n385);
and (n432,n417,n430);
or (n433,n434,n493);
and (n434,n435,n492);
xor (n435,n436,n437);
xor (n436,n416,n431);
or (n437,n438,n491);
and (n438,n439,n442);
xor (n439,n440,n441);
xor (n440,n419,n426);
xor (n441,n226,n246);
or (n442,n443,n490);
and (n443,n444,n465);
xor (n444,n445,n446);
xor (n445,n247,n253);
or (n446,n447,n464);
and (n447,n448,n457);
xor (n448,n449,n450);
nor (n449,n70,n252);
nand (n450,n451,n455);
or (n451,n134,n452);
nor (n452,n453,n454);
and (n453,n187,n25);
and (n454,n189,n26);
nand (n455,n456,n128);
not (n456,n309);
nand (n457,n458,n463);
or (n458,n191,n459);
not (n459,n460);
nor (n460,n461,n462);
and (n461,n60,n175);
and (n462,n61,n176);
or (n463,n178,n321);
and (n464,n449,n450);
or (n465,n466,n489);
and (n466,n467,n483);
xor (n467,n468,n476);
nand (n468,n469,n474);
or (n469,n470,n197);
not (n470,n471);
nand (n471,n472,n473);
or (n472,n46,n84);
or (n473,n82,n205);
nand (n474,n475,n199);
not (n475,n326);
nand (n476,n477,n482);
or (n477,n103,n478);
not (n478,n479);
nor (n479,n480,n481);
and (n480,n16,n109);
and (n481,n17,n106);
nand (n482,n256,n105);
nand (n483,n484,n488);
or (n484,n229,n485);
nor (n485,n486,n487);
and (n486,n55,n151);
and (n487,n53,n150);
or (n488,n41,n349);
and (n489,n468,n476);
and (n490,n445,n446);
and (n491,n440,n441);
xor (n492,n223,n301);
and (n493,n436,n437);
not (n494,n495);
nand (n495,n496,n711);
nor (n496,n497,n710);
and (n497,n498,n562);
nand (n498,n499,n501);
not (n499,n500);
xor (n500,n435,n492);
not (n501,n502);
or (n502,n503,n561);
and (n503,n504,n507);
xor (n504,n505,n506);
xor (n505,n303,n360);
xor (n506,n439,n442);
or (n507,n508,n560);
and (n508,n509,n512);
xor (n509,n510,n511);
xor (n510,n336,n353);
xor (n511,n306,n324);
or (n512,n513,n559);
and (n513,n514,n535);
xor (n514,n515,n521);
nand (n515,n516,n520);
or (n516,n21,n517);
nor (n517,n518,n519);
and (n518,n18,n212);
and (n519,n19,n211);
or (n520,n405,n339);
nor (n521,n522,n529);
not (n522,n523);
nand (n523,n524,n525);
or (n524,n452,n127);
or (n525,n134,n526);
nor (n526,n527,n528);
and (n527,n219,n25);
and (n528,n218,n26);
nand (n529,n530,n53);
nand (n530,n531,n532);
or (n531,n100,n45);
nand (n532,n533,n205);
not (n533,n534);
and (n534,n100,n45);
or (n535,n536,n558);
and (n536,n537,n552);
xor (n537,n538,n545);
nand (n538,n539,n544);
or (n539,n540,n191);
not (n540,n541);
nand (n541,n542,n543);
or (n542,n176,n90);
or (n543,n175,n88);
nand (n544,n179,n460);
nand (n545,n546,n551);
or (n546,n547,n197);
not (n547,n548);
nand (n548,n549,n550);
or (n549,n46,n165);
or (n550,n205,n166);
nand (n551,n199,n471);
nand (n552,n553,n554);
or (n553,n104,n478);
or (n554,n555,n103);
nor (n555,n556,n557);
and (n556,n109,n174);
and (n557,n106,n173);
and (n558,n538,n545);
and (n559,n515,n521);
and (n560,n510,n511);
and (n561,n505,n506);
nand (n562,n563,n709);
or (n563,n564,n701);
not (n564,n565);
nand (n565,n566,n700);
or (n566,n567,n650);
nor (n567,n568,n598);
xor (n568,n569,n597);
xor (n569,n570,n571);
xor (n570,n444,n465);
or (n571,n572,n596);
and (n572,n573,n576);
xor (n573,n574,n575);
xor (n574,n467,n483);
xor (n575,n448,n457);
or (n576,n577,n595);
and (n577,n578,n591);
xor (n578,n579,n585);
nand (n579,n580,n584);
or (n580,n229,n581);
nor (n581,n582,n583);
and (n582,n252,n53);
and (n583,n100,n55);
or (n584,n41,n485);
nand (n585,n586,n590);
or (n586,n21,n587);
nor (n587,n588,n589);
and (n588,n18,n52);
and (n589,n19,n51);
or (n590,n405,n517);
nand (n591,n592,n594);
or (n592,n593,n522);
not (n593,n529);
or (n594,n523,n529);
and (n595,n579,n585);
and (n596,n574,n575);
xor (n597,n509,n512);
or (n598,n599,n649);
and (n599,n600,n648);
xor (n600,n601,n602);
xor (n601,n514,n535);
or (n602,n603,n647);
and (n603,n604,n646);
xor (n604,n605,n623);
or (n605,n606,n622);
and (n606,n607,n616);
xor (n607,n608,n609);
nor (n608,n41,n252);
nand (n609,n610,n614);
or (n610,n611,n134);
nor (n611,n612,n613);
and (n612,n25,n212);
and (n613,n26,n211);
nand (n614,n615,n128);
not (n615,n526);
nand (n616,n617,n618);
or (n617,n540,n178);
or (n618,n191,n619);
nor (n619,n620,n621);
and (n620,n175,n82);
and (n621,n176,n84);
and (n622,n608,n609);
or (n623,n624,n645);
and (n624,n625,n639);
xor (n625,n626,n633);
nand (n626,n627,n632);
or (n627,n628,n197);
not (n628,n629);
nand (n629,n630,n631);
or (n630,n46,n150);
or (n631,n205,n151);
nand (n632,n199,n548);
nand (n633,n634,n638);
or (n634,n635,n103);
nor (n635,n636,n637);
and (n636,n109,n187);
and (n637,n106,n189);
or (n638,n555,n104);
nand (n639,n640,n644);
or (n640,n21,n641);
nor (n641,n642,n643);
and (n642,n18,n61);
and (n643,n19,n60);
or (n644,n405,n587);
and (n645,n626,n633);
xor (n646,n537,n552);
and (n647,n605,n623);
xor (n648,n573,n576);
and (n649,n601,n602);
nand (n650,n651,n699);
or (n651,n652,n698);
and (n652,n653,n656);
xor (n653,n654,n655);
xor (n654,n578,n591);
xor (n655,n604,n646);
or (n656,n657,n697);
and (n657,n658,n696);
xor (n658,n659,n672);
and (n659,n660,n666);
and (n660,n661,n46);
nand (n661,n662,n663);
or (n662,n100,n201);
nand (n663,n664,n175);
not (n664,n665);
and (n665,n100,n201);
nand (n666,n667,n671);
or (n667,n134,n668);
nor (n668,n669,n670);
and (n669,n25,n52);
and (n670,n26,n51);
or (n671,n127,n611);
or (n672,n673,n695);
and (n673,n674,n689);
xor (n674,n675,n682);
nand (n675,n676,n680);
or (n676,n677,n191);
nor (n677,n678,n679);
and (n678,n175,n166);
and (n679,n176,n165);
nand (n680,n681,n179);
not (n681,n619);
nand (n682,n683,n684);
or (n683,n628,n215);
nand (n684,n685,n198);
not (n685,n686);
nor (n686,n687,n688);
and (n687,n252,n46);
and (n688,n205,n100);
nand (n689,n690,n694);
or (n690,n103,n691);
nor (n691,n692,n693);
and (n692,n109,n219);
and (n693,n106,n218);
or (n694,n635,n104);
and (n695,n675,n682);
xor (n696,n607,n616);
and (n697,n659,n672);
and (n698,n654,n655);
xor (n699,n600,n648);
nand (n700,n568,n598);
not (n701,n702);
nand (n702,n703,n705);
not (n703,n704);
xor (n704,n504,n507);
not (n705,n706);
or (n706,n707,n708);
and (n707,n569,n597);
and (n708,n570,n571);
nand (n709,n704,n706);
nor (n710,n499,n501);
nand (n711,n498,n712,n1003);
nand (n712,n713,n1002);
or (n713,n714,n751);
not (n714,n715);
or (n715,n716,n717);
xor (n716,n653,n656);
or (n717,n718,n750);
and (n718,n719,n749);
xor (n719,n720,n721);
xor (n720,n625,n639);
or (n721,n722,n748);
and (n722,n723,n731);
xor (n723,n724,n730);
nand (n724,n725,n729);
or (n725,n21,n726);
nor (n726,n727,n728);
and (n727,n18,n88);
and (n728,n19,n90);
or (n729,n405,n641);
xor (n730,n660,n666);
or (n731,n732,n747);
and (n732,n733,n741);
xor (n733,n734,n735);
nor (n734,n215,n252);
nand (n735,n736,n740);
or (n736,n737,n103);
nor (n737,n738,n739);
and (n738,n211,n106);
and (n739,n212,n109);
or (n740,n691,n104);
nand (n741,n742,n746);
or (n742,n191,n743);
nor (n743,n744,n745);
and (n744,n175,n151);
and (n745,n176,n150);
or (n746,n178,n677);
and (n747,n734,n735);
and (n748,n724,n730);
xor (n749,n658,n696);
and (n750,n720,n721);
not (n751,n752);
or (n752,n753,n1001);
and (n753,n754,n794);
xor (n754,n755,n793);
or (n755,n756,n792);
and (n756,n757,n791);
xor (n757,n758,n759);
xor (n758,n674,n689);
or (n759,n760,n790);
and (n760,n761,n776);
xor (n761,n762,n770);
nand (n762,n763,n768);
or (n763,n764,n134);
not (n764,n765);
nand (n765,n766,n767);
or (n766,n26,n60);
or (n767,n25,n61);
nand (n768,n769,n128);
not (n769,n668);
nand (n770,n771,n775);
or (n771,n21,n772);
nor (n772,n773,n774);
and (n773,n18,n82);
and (n774,n19,n84);
or (n775,n405,n726);
and (n776,n777,n783);
nor (n777,n778,n175);
nor (n778,n779,n781);
and (n779,n252,n780);
not (n780,n181);
nor (n781,n782,n19);
and (n782,n100,n181);
nand (n783,n784,n789);
or (n784,n103,n785);
not (n785,n786);
nor (n786,n787,n788);
and (n787,n51,n109);
and (n788,n52,n106);
or (n789,n737,n104);
and (n790,n762,n770);
xor (n791,n723,n731);
and (n792,n758,n759);
xor (n793,n719,n749);
nand (n794,n795,n998,n1000);
nand (n795,n796,n831,n991);
nand (n796,n797,n799);
not (n797,n798);
xor (n798,n757,n791);
not (n799,n800);
or (n800,n801,n830);
and (n801,n802,n829);
xor (n802,n803,n828);
or (n803,n804,n827);
and (n804,n805,n821);
xor (n805,n806,n814);
nand (n806,n807,n812);
or (n807,n808,n191);
not (n808,n809);
nand (n809,n810,n811);
or (n810,n175,n100);
or (n811,n252,n176);
nand (n812,n813,n179);
not (n813,n743);
nand (n814,n815,n820);
or (n815,n816,n134);
not (n816,n817);
nand (n817,n818,n819);
or (n818,n26,n90);
or (n819,n25,n88);
nand (n820,n128,n765);
nand (n821,n822,n826);
or (n822,n21,n823);
nor (n823,n824,n825);
and (n824,n18,n166);
and (n825,n19,n165);
or (n826,n405,n772);
and (n827,n806,n814);
xor (n828,n733,n741);
xor (n829,n761,n776);
and (n830,n803,n828);
nand (n831,n832,n990);
or (n832,n833,n883);
not (n833,n834);
nand (n834,n835,n859);
not (n835,n836);
xor (n836,n837,n858);
xor (n837,n838,n839);
xor (n838,n777,n783);
or (n839,n840,n857);
and (n840,n841,n850);
xor (n841,n842,n843);
and (n842,n179,n100);
nand (n843,n844,n849);
or (n844,n103,n845);
not (n845,n846);
nor (n846,n847,n848);
and (n847,n60,n109);
and (n848,n61,n106);
nand (n849,n786,n105);
nand (n850,n851,n856);
or (n851,n852,n134);
not (n852,n853);
nor (n853,n854,n855);
and (n854,n84,n25);
and (n855,n82,n26);
nand (n856,n128,n817);
and (n857,n842,n843);
xor (n858,n805,n821);
not (n859,n860);
or (n860,n861,n882);
and (n861,n862,n881);
xor (n862,n863,n869);
nand (n863,n864,n868);
or (n864,n21,n865);
nor (n865,n866,n867);
and (n866,n150,n19);
and (n867,n151,n18);
or (n868,n405,n823);
and (n869,n870,n875);
and (n870,n871,n19);
nand (n871,n872,n874);
or (n872,n873,n26);
and (n873,n100,n27);
or (n874,n100,n27);
nand (n875,n876,n877);
or (n876,n104,n845);
or (n877,n878,n103);
nor (n878,n879,n880);
and (n879,n109,n88);
and (n880,n106,n90);
xor (n881,n841,n850);
and (n882,n863,n869);
not (n883,n884);
nand (n884,n885,n989);
or (n885,n886,n909);
not (n886,n887);
nand (n887,n888,n890);
not (n888,n889);
xor (n889,n862,n881);
not (n890,n891);
or (n891,n892,n908);
and (n892,n893,n907);
xor (n893,n894,n901);
nand (n894,n895,n900);
or (n895,n896,n134);
not (n896,n897);
nor (n897,n898,n899);
and (n898,n165,n25);
and (n899,n166,n26);
nand (n900,n853,n128);
nand (n901,n902,n903);
or (n902,n405,n865);
nand (n903,n22,n904);
nand (n904,n905,n906);
or (n905,n100,n18);
or (n906,n252,n19);
xor (n907,n870,n875);
and (n908,n894,n901);
not (n909,n910);
or (n910,n911,n988);
and (n911,n912,n933);
xor (n912,n913,n932);
or (n913,n914,n931);
and (n914,n915,n924);
xor (n915,n916,n917);
and (n916,n23,n100);
nand (n917,n918,n923);
or (n918,n919,n134);
not (n919,n920);
nor (n920,n921,n922);
and (n921,n150,n25);
and (n922,n151,n26);
nand (n923,n897,n128);
nand (n924,n925,n930);
or (n925,n103,n926);
not (n926,n927);
nor (n927,n928,n929);
and (n928,n84,n109);
and (n929,n82,n106);
or (n930,n878,n104);
and (n931,n916,n917);
xor (n932,n893,n907);
nand (n933,n934,n987);
or (n934,n935,n951);
nor (n935,n936,n937);
xor (n936,n915,n924);
nor (n937,n938,n946);
not (n938,n939);
nand (n939,n940,n941);
or (n940,n104,n926);
nand (n941,n942,n945);
nand (n942,n943,n944);
or (n943,n166,n109);
nand (n944,n109,n166);
not (n945,n103);
nand (n946,n947,n26);
nand (n947,n948,n950);
or (n948,n949,n106);
and (n949,n100,n131);
or (n950,n100,n131);
nor (n951,n952,n986);
and (n952,n953,n965);
nand (n953,n954,n961);
not (n954,n955);
nand (n955,n956,n960);
or (n956,n134,n957);
nor (n957,n958,n959);
and (n958,n26,n252);
and (n959,n100,n25);
or (n960,n127,n919);
nor (n961,n962,n963);
and (n962,n946,n939);
and (n963,n964,n938);
not (n964,n946);
or (n965,n966,n985);
and (n966,n967,n976);
xor (n967,n968,n969);
nor (n968,n127,n252);
nand (n969,n970,n975);
or (n970,n103,n971);
not (n971,n972);
nand (n972,n973,n974);
or (n973,n150,n106);
nand (n974,n106,n150);
nand (n975,n942,n105);
nor (n976,n977,n983);
nor (n977,n978,n979);
and (n978,n972,n105);
nor (n979,n980,n103);
nor (n980,n981,n982);
and (n981,n252,n106);
and (n982,n100,n109);
or (n983,n984,n109);
and (n984,n100,n105);
and (n985,n968,n969);
nor (n986,n954,n961);
nand (n987,n936,n937);
and (n988,n913,n932);
nand (n989,n889,n891);
nand (n990,n836,n860);
nand (n991,n992,n996);
not (n992,n993);
or (n993,n994,n995);
and (n994,n837,n858);
and (n995,n838,n839);
not (n996,n997);
xor (n997,n802,n829);
nand (n998,n796,n999);
and (n999,n997,n993);
nand (n1000,n800,n798);
and (n1001,n755,n793);
nand (n1002,n716,n717);
nor (n1003,n701,n1004);
nand (n1004,n1005,n1006);
not (n1005,n567);
or (n1006,n651,n699);
nand (n1007,n5,n433);
nand (n1008,n1009,n1106);
not (n1009,n1010);
nor (n1010,n1011,n1103);
xor (n1011,n1012,n1084);
xor (n1012,n1013,n1081);
xor (n1013,n1014,n1058);
xor (n1014,n1015,n1037);
xor (n1015,n1016,n1030);
xor (n1016,n1017,n1023);
nand (n1017,n1018,n1019);
or (n1018,n170,n191);
nand (n1019,n179,n1020);
nand (n1020,n1021,n1022);
or (n1021,n17,n175);
nand (n1022,n175,n17);
nand (n1023,n1024,n1026);
or (n1024,n1025,n153);
not (n1025,n163);
nand (n1026,n155,n1027);
nor (n1027,n1028,n1029);
and (n1028,n84,n96);
and (n1029,n82,n97);
nand (n1030,n1031,n1035);
or (n1031,n1032,n252);
not (n1032,n1033);
nor (n1033,n1034,n94);
not (n1034,n98);
or (n1035,n1036,n150);
not (n1036,n94);
xor (n1037,n1038,n1051);
xor (n1038,n1039,n1045);
nand (n1039,n1040,n1041);
or (n1040,n121,n134);
nand (n1041,n128,n1042);
nand (n1042,n1043,n1044);
or (n1043,n110,n25);
nand (n1044,n25,n110);
nand (n1045,n1046,n1047);
or (n1046,n197,n216);
nand (n1047,n199,n1048);
nor (n1048,n1049,n1050);
and (n1049,n187,n46);
and (n1050,n189,n205);
nand (n1051,n1052,n1054);
or (n1052,n21,n1053);
not (n1053,n34);
or (n1054,n405,n1055);
nor (n1055,n1056,n1057);
and (n1056,n142,n19);
and (n1057,n140,n18);
xor (n1058,n1059,n1072);
xor (n1059,n1060,n1066);
nand (n1060,n1061,n1062);
or (n1061,n48,n229);
or (n1062,n1063,n41);
nor (n1063,n1064,n1065);
and (n1064,n55,n212);
and (n1065,n53,n211);
nand (n1066,n1067,n1068);
or (n1067,n69,n86);
or (n1068,n1069,n70);
nor (n1069,n1070,n1071);
and (n1070,n77,n61);
and (n1071,n78,n60);
nand (n1072,n1073,n1075);
or (n1073,n103,n1074);
not (n1074,n114);
or (n1075,n1076,n104);
nor (n1076,n1077,n1079);
and (n1077,n1078,n109);
and (n1079,n1080,n106);
not (n1080,n1078);
or (n1081,n1082,n1083);
and (n1082,n364,n414);
and (n1083,n365,n368);
xor (n1084,n1085,n1100);
xor (n1085,n1086,n1089);
or (n1086,n1087,n1088);
and (n1087,n369,n393);
and (n1088,n370,n371);
xor (n1089,n1090,n1097);
xor (n1090,n1091,n1094);
or (n1091,n1092,n1093);
and (n1092,n92,n119);
and (n1093,n93,n101);
or (n1094,n1095,n1096);
and (n1095,n10,n67);
and (n1096,n11,n39);
or (n1097,n1098,n1099);
and (n1098,n144,n195);
and (n1099,n145,n168);
or (n1100,n1101,n1102);
and (n1101,n8,n143);
and (n1102,n9,n91);
or (n1103,n1104,n1105);
and (n1104,n6,n363);
and (n1105,n7,n221);
nand (n1106,n1011,n1103);
nand (n1107,n2,n1008);
xor (n1108,n1109,n1896);
xor (n1109,n1110,n1895);
xor (n1110,n1111,n1887);
xor (n1111,n1112,n167);
xor (n1112,n1113,n1872);
xor (n1113,n1114,n1871);
xor (n1114,n1115,n1850);
xor (n1115,n1116,n1849);
xor (n1116,n1117,n1822);
xor (n1117,n1118,n1821);
xor (n1118,n1119,n1788);
xor (n1119,n1120,n1787);
xor (n1120,n1121,n1749);
xor (n1121,n1122,n1748);
xor (n1122,n1123,n1705);
xor (n1123,n1124,n1704);
xor (n1124,n1125,n1654);
xor (n1125,n1126,n1653);
xor (n1126,n1127,n1599);
xor (n1127,n1128,n177);
xor (n1128,n1129,n1537);
xor (n1129,n1130,n1536);
xor (n1130,n1131,n1468);
xor (n1131,n1132,n1467);
xor (n1132,n1133,n1393);
xor (n1133,n1134,n1392);
xor (n1134,n1135,n1315);
xor (n1135,n1136,n126);
xor (n1136,n1137,n1229);
xor (n1137,n1138,n1228);
xor (n1138,n1139,n1141);
xor (n1139,n1140,n118);
and (n1140,n1078,n105);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
and (n1143,n117,n105);
and (n1144,n110,n106);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1150);
and (n1148,n1149,n280);
and (n1149,n110,n105);
and (n1150,n1151,n1152);
xor (n1151,n1149,n280);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
and (n1154,n125,n105);
and (n1155,n140,n106);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1161);
and (n1159,n1160,n258);
and (n1160,n140,n105);
and (n1161,n1162,n1163);
xor (n1162,n1160,n258);
or (n1163,n1164,n1166);
and (n1164,n1165,n481);
and (n1165,n37,n105);
and (n1166,n1167,n1168);
xor (n1167,n1165,n481);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
and (n1170,n17,n105);
and (n1171,n174,n106);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
and (n1176,n174,n105);
and (n1177,n187,n106);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
and (n1182,n187,n105);
and (n1183,n219,n106);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
and (n1188,n219,n105);
and (n1189,n212,n106);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1195);
and (n1193,n1194,n788);
and (n1194,n212,n105);
and (n1195,n1196,n1197);
xor (n1196,n1194,n788);
or (n1197,n1198,n1200);
and (n1198,n1199,n848);
and (n1199,n52,n105);
and (n1200,n1201,n1202);
xor (n1201,n1199,n848);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
and (n1204,n61,n105);
and (n1205,n88,n106);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
or (n1208,n1209,n1211);
and (n1209,n1210,n929);
and (n1210,n88,n105);
and (n1211,n1212,n1213);
xor (n1212,n1210,n929);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
and (n1215,n82,n105);
and (n1216,n166,n106);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
and (n1221,n166,n105);
and (n1222,n151,n106);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
and (n1225,n1226,n1227);
and (n1226,n151,n105);
and (n1227,n100,n106);
and (n1228,n110,n131);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1146,n1147);
and (n1232,n125,n131);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1151,n1152);
and (n1238,n140,n131);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1157,n1158);
and (n1244,n37,n131);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1162,n1163);
and (n1250,n17,n131);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1167,n1168);
and (n1256,n174,n131);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1173,n1174);
and (n1262,n187,n131);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1179,n1180);
and (n1268,n219,n131);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1185,n1186);
and (n1274,n212,n131);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1191,n1192);
and (n1280,n52,n131);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1196,n1197);
and (n1286,n61,n131);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1201,n1202);
and (n1292,n88,n131);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1207,n1208);
and (n1298,n82,n131);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1212,n1213);
and (n1304,n166,n131);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1218,n1219);
and (n1310,n151,n131);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
and (n1313,n1314,n949);
xor (n1314,n1224,n1225);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1234,n1235);
and (n1318,n140,n26);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
or (n1321,n1322,n1324);
and (n1322,n1323,n298);
xor (n1323,n1240,n1241);
and (n1324,n1325,n1326);
xor (n1325,n1323,n298);
or (n1326,n1327,n1330);
and (n1327,n1328,n1329);
xor (n1328,n1246,n1247);
and (n1329,n17,n26);
and (n1330,n1331,n1332);
xor (n1331,n1328,n1329);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1252,n1253);
and (n1335,n174,n26);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1258,n1259);
and (n1341,n187,n26);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1264,n1265);
and (n1347,n219,n26);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1270,n1271);
and (n1353,n212,n26);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1276,n1277);
and (n1359,n52,n26);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1282,n1283);
and (n1365,n61,n26);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1288,n1289);
and (n1371,n88,n26);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1377);
and (n1375,n1376,n855);
xor (n1376,n1294,n1295);
and (n1377,n1378,n1379);
xor (n1378,n1376,n855);
or (n1379,n1380,n1382);
and (n1380,n1381,n899);
xor (n1381,n1300,n1301);
and (n1382,n1383,n1384);
xor (n1383,n1381,n899);
or (n1384,n1385,n1387);
and (n1385,n1386,n922);
xor (n1386,n1306,n1307);
and (n1387,n1388,n1389);
xor (n1388,n1386,n922);
and (n1389,n1390,n1391);
xor (n1390,n1312,n1313);
and (n1391,n100,n26);
and (n1392,n140,n27);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1320,n1321);
and (n1396,n37,n27);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1325,n1326);
and (n1402,n17,n27);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1331,n1332);
and (n1408,n174,n27);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1337,n1338);
and (n1414,n187,n27);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1343,n1344);
and (n1420,n219,n27);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1349,n1350);
and (n1426,n212,n27);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1355,n1356);
and (n1432,n52,n27);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1361,n1362);
and (n1438,n61,n27);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1367,n1368);
and (n1444,n88,n27);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1373,n1374);
and (n1450,n82,n27);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1378,n1379);
and (n1456,n166,n27);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
or (n1459,n1460,n1463);
and (n1460,n1461,n1462);
xor (n1461,n1383,n1384);
and (n1462,n151,n27);
and (n1463,n1464,n1465);
xor (n1464,n1461,n1462);
and (n1465,n1466,n873);
xor (n1466,n1388,n1389);
and (n1467,n37,n19);
or (n1468,n1469,n1471);
and (n1469,n1470,n20);
xor (n1470,n1398,n1399);
and (n1471,n1472,n1473);
xor (n1472,n1470,n20);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1404,n1405);
and (n1476,n174,n19);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1410,n1411);
and (n1482,n187,n19);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1416,n1417);
and (n1488,n219,n19);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1422,n1423);
and (n1494,n212,n19);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1428,n1429);
and (n1500,n52,n19);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1434,n1435);
and (n1506,n61,n19);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1440,n1441);
and (n1512,n88,n19);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1446,n1447);
and (n1518,n82,n19);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1452,n1453);
and (n1524,n166,n19);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1458,n1459);
and (n1530,n151,n19);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
and (n1533,n1534,n1535);
xor (n1534,n1464,n1465);
and (n1535,n100,n19);
and (n1536,n17,n181);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1472,n1473);
and (n1540,n174,n181);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1478,n1479);
and (n1546,n187,n181);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1484,n1485);
and (n1552,n219,n181);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1490,n1491);
and (n1558,n212,n181);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1496,n1497);
and (n1564,n52,n181);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1502,n1503);
and (n1570,n61,n181);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1508,n1509);
and (n1576,n88,n181);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1514,n1515);
and (n1582,n82,n181);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1520,n1521);
and (n1588,n166,n181);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1526,n1527);
and (n1594,n151,n181);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
and (n1597,n1598,n782);
xor (n1598,n1532,n1533);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
xor (n1601,n1542,n1543);
and (n1602,n187,n176);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1608);
and (n1606,n1607,n389);
xor (n1607,n1548,n1549);
and (n1608,n1609,n1610);
xor (n1609,n1607,n389);
or (n1610,n1611,n1613);
and (n1611,n1612,n318);
xor (n1612,n1554,n1555);
and (n1613,n1614,n1615);
xor (n1614,n1612,n318);
or (n1615,n1616,n1619);
and (n1616,n1617,n1618);
xor (n1617,n1560,n1561);
and (n1618,n52,n176);
and (n1619,n1620,n1621);
xor (n1620,n1617,n1618);
or (n1621,n1622,n1624);
and (n1622,n1623,n462);
xor (n1623,n1566,n1567);
and (n1624,n1625,n1626);
xor (n1625,n1623,n462);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1572,n1573);
and (n1629,n88,n176);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1578,n1579);
and (n1635,n82,n176);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1584,n1585);
and (n1641,n166,n176);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
xor (n1646,n1590,n1591);
and (n1647,n151,n176);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
and (n1650,n1651,n1652);
xor (n1651,n1596,n1597);
and (n1652,n100,n176);
and (n1653,n187,n201);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1604,n1605);
and (n1657,n219,n201);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1609,n1610);
and (n1663,n212,n201);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1614,n1615);
and (n1669,n52,n201);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1620,n1621);
and (n1675,n61,n201);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1625,n1626);
and (n1681,n88,n201);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1631,n1632);
and (n1687,n82,n201);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
or (n1690,n1691,n1694);
and (n1691,n1692,n1693);
xor (n1692,n1637,n1638);
and (n1693,n166,n201);
and (n1694,n1695,n1696);
xor (n1695,n1692,n1693);
or (n1696,n1697,n1700);
and (n1697,n1698,n1699);
xor (n1698,n1643,n1644);
and (n1699,n151,n201);
and (n1700,n1701,n1702);
xor (n1701,n1698,n1699);
and (n1702,n1703,n665);
xor (n1703,n1649,n1650);
and (n1704,n219,n46);
or (n1705,n1706,n1708);
and (n1706,n1707,n213);
xor (n1707,n1659,n1660);
and (n1708,n1709,n1710);
xor (n1709,n1707,n213);
or (n1710,n1711,n1713);
and (n1711,n1712,n401);
xor (n1712,n1665,n1666);
and (n1713,n1714,n1715);
xor (n1714,n1712,n401);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1671,n1672);
and (n1718,n61,n46);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1677,n1678);
and (n1724,n88,n46);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1683,n1684);
and (n1730,n82,n46);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1689,n1690);
and (n1736,n166,n46);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1695,n1696);
and (n1742,n151,n46);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
and (n1745,n1746,n1747);
xor (n1746,n1701,n1702);
and (n1747,n100,n46);
and (n1748,n212,n45);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
xor (n1751,n1709,n1710);
and (n1752,n52,n45);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
or (n1755,n1756,n1759);
and (n1756,n1757,n1758);
xor (n1757,n1714,n1715);
and (n1758,n61,n45);
and (n1759,n1760,n1761);
xor (n1760,n1757,n1758);
or (n1761,n1762,n1765);
and (n1762,n1763,n1764);
xor (n1763,n1720,n1721);
and (n1764,n88,n45);
and (n1765,n1766,n1767);
xor (n1766,n1763,n1764);
or (n1767,n1768,n1771);
and (n1768,n1769,n1770);
xor (n1769,n1726,n1727);
and (n1770,n82,n45);
and (n1771,n1772,n1773);
xor (n1772,n1769,n1770);
or (n1773,n1774,n1777);
and (n1774,n1775,n1776);
xor (n1775,n1732,n1733);
and (n1776,n166,n45);
and (n1777,n1778,n1779);
xor (n1778,n1775,n1776);
or (n1779,n1780,n1783);
and (n1780,n1781,n1782);
xor (n1781,n1738,n1739);
and (n1782,n151,n45);
and (n1783,n1784,n1785);
xor (n1784,n1781,n1782);
and (n1785,n1786,n534);
xor (n1786,n1744,n1745);
and (n1787,n52,n53);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1754,n1755);
and (n1791,n61,n53);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1760,n1761);
and (n1797,n88,n53);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
xor (n1802,n1766,n1767);
and (n1803,n82,n53);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
xor (n1808,n1772,n1773);
and (n1809,n166,n53);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
xor (n1814,n1778,n1779);
and (n1815,n151,n53);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
and (n1818,n1819,n1820);
xor (n1819,n1784,n1785);
and (n1820,n100,n53);
and (n1821,n61,n73);
or (n1822,n1823,n1826);
and (n1823,n1824,n1825);
xor (n1824,n1793,n1794);
and (n1825,n88,n73);
and (n1826,n1827,n1828);
xor (n1827,n1824,n1825);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1799,n1800);
and (n1831,n82,n73);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1838);
and (n1835,n1836,n1837);
xor (n1836,n1805,n1806);
and (n1837,n166,n73);
and (n1838,n1839,n1840);
xor (n1839,n1836,n1837);
or (n1840,n1841,n1844);
and (n1841,n1842,n1843);
xor (n1842,n1811,n1812);
and (n1843,n151,n73);
and (n1844,n1845,n1846);
xor (n1845,n1842,n1843);
and (n1846,n1847,n1848);
xor (n1847,n1817,n1818);
not (n1848,n250);
and (n1849,n88,n78);
or (n1850,n1851,n1854);
and (n1851,n1852,n1853);
xor (n1852,n1827,n1828);
and (n1853,n82,n78);
and (n1854,n1855,n1856);
xor (n1855,n1852,n1853);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n1833,n1834);
and (n1859,n166,n78);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1839,n1840);
and (n1865,n151,n78);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
and (n1868,n1869,n1870);
xor (n1869,n1845,n1846);
and (n1870,n100,n78);
and (n1871,n82,n157);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1855,n1856);
and (n1875,n166,n157);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1861,n1862);
and (n1881,n151,n157);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
and (n1884,n1885,n1886);
xor (n1885,n1867,n1868);
not (n1886,n273);
or (n1887,n1888,n1890);
and (n1888,n1889,n152);
xor (n1889,n1877,n1878);
and (n1890,n1891,n1892);
xor (n1891,n1889,n152);
and (n1892,n1893,n1894);
xor (n1893,n1883,n1884);
and (n1894,n100,n97);
and (n1895,n151,n98);
and (n1896,n1897,n1898);
xor (n1897,n1891,n1892);
and (n1898,n100,n98);
endmodule
