module top (out,n3,n4,n5,n26,n28,n35,n36,n45,n52
        ,n54,n60,n66,n71,n80,n85,n92,n99,n111,n119
        ,n125,n137,n141,n148,n154,n162,n167,n172,n177,n186
        ,n192,n197,n204,n214);
output out;
input n3;
input n4;
input n5;
input n26;
input n28;
input n35;
input n36;
input n45;
input n52;
input n54;
input n60;
input n66;
input n71;
input n80;
input n85;
input n92;
input n99;
input n111;
input n119;
input n125;
input n137;
input n141;
input n148;
input n154;
input n162;
input n167;
input n172;
input n177;
input n186;
input n192;
input n197;
input n204;
input n214;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
xnor (out,n0,n819);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n816);
nand (n7,n8,n815);
or (n8,n9,n408);
not (n9,n10);
nand (n10,n11,n407);
nand (n11,n12,n373);
not (n12,n13);
xor (n13,n14,n319);
xor (n14,n15,n216);
xor (n15,n16,n181);
xor (n16,n17,n102);
or (n17,n18,n101);
and (n18,n19,n74);
xor (n19,n20,n47);
nand (n20,n21,n41);
or (n21,n22,n30);
not (n22,n23);
nor (n23,n24,n29);
and (n24,n25,n27);
not (n25,n26);
not (n27,n28);
and (n29,n26,n28);
nand (n30,n31,n38);
not (n31,n32);
nand (n32,n33,n37);
or (n33,n34,n36);
not (n34,n35);
nand (n37,n36,n34);
nand (n38,n39,n40);
or (n39,n34,n28);
nand (n40,n34,n28);
nand (n41,n42,n32);
nor (n42,n43,n46);
and (n43,n27,n44);
not (n44,n45);
and (n46,n45,n28);
nand (n47,n48,n68);
or (n48,n49,n57);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n53);
not (n53,n54);
or (n55,n56,n54);
not (n56,n52);
nand (n57,n58,n62);
nand (n58,n59,n61);
or (n59,n60,n56);
nand (n61,n56,n60);
not (n62,n63);
nand (n63,n64,n67);
or (n64,n65,n60);
not (n65,n66);
nand (n67,n60,n65);
nand (n68,n63,n69);
nor (n69,n70,n72);
and (n70,n71,n52);
and (n72,n73,n56);
not (n73,n71);
nand (n74,n75,n94);
or (n75,n76,n88);
not (n76,n77);
nor (n77,n78,n82);
nand (n78,n79,n81);
or (n79,n56,n80);
nand (n81,n56,n80);
nor (n82,n83,n86);
and (n83,n84,n80);
not (n84,n85);
and (n86,n85,n87);
not (n87,n80);
not (n88,n89);
nor (n89,n90,n93);
and (n90,n91,n84);
not (n91,n92);
and (n93,n92,n85);
or (n94,n95,n96);
not (n95,n78);
nor (n96,n97,n100);
and (n97,n98,n85);
not (n98,n99);
and (n100,n99,n84);
and (n101,n20,n47);
or (n102,n103,n180);
and (n103,n104,n156);
xor (n104,n105,n129);
nand (n105,n106,n122);
or (n106,n107,n117);
not (n107,n108);
nor (n108,n109,n113);
nand (n109,n110,n112);
or (n110,n111,n27);
nand (n112,n111,n27);
nor (n113,n114,n116);
and (n114,n115,n66);
not (n115,n111);
and (n116,n111,n65);
nor (n117,n118,n120);
and (n118,n119,n65);
and (n120,n121,n66);
not (n121,n119);
or (n122,n123,n128);
nor (n123,n124,n126);
and (n124,n65,n125);
and (n126,n66,n127);
not (n127,n125);
not (n128,n109);
nand (n129,n130,n150);
or (n130,n131,n144);
not (n131,n132);
and (n132,n133,n139);
not (n133,n134);
nand (n134,n135,n138);
or (n135,n136,n85);
not (n136,n137);
nand (n138,n85,n136);
nand (n139,n140,n142);
nand (n140,n141,n136);
nand (n142,n137,n143);
not (n143,n141);
not (n144,n145);
nor (n145,n146,n149);
and (n146,n147,n143);
not (n147,n148);
and (n149,n148,n141);
or (n150,n151,n133);
nor (n151,n152,n155);
and (n152,n153,n141);
not (n153,n154);
and (n155,n154,n143);
nand (n156,n157,n174);
or (n157,n158,n169);
nand (n158,n159,n164);
nor (n159,n160,n163);
and (n160,n161,n141);
not (n161,n162);
and (n163,n162,n143);
nor (n164,n165,n168);
and (n165,n161,n166);
not (n166,n167);
and (n168,n162,n167);
nor (n169,n170,n173);
and (n170,n171,n167);
not (n171,n172);
and (n173,n172,n166);
or (n174,n175,n159);
nor (n175,n176,n178);
and (n176,n166,n177);
and (n178,n167,n179);
not (n179,n177);
and (n180,n105,n129);
xor (n181,n182,n206);
xor (n182,n183,n188);
and (n183,n184,n172);
nand (n184,n185,n187);
or (n185,n166,n186);
nand (n187,n186,n166);
nand (n188,n189,n200);
or (n189,n190,n193);
nand (n190,n191,n36);
not (n191,n192);
not (n193,n194);
nor (n194,n195,n199);
and (n195,n196,n198);
not (n196,n197);
not (n198,n36);
and (n199,n197,n36);
nand (n200,n201,n192);
nor (n201,n202,n205);
and (n202,n203,n198);
not (n203,n204);
and (n205,n204,n36);
nand (n206,n207,n209);
or (n207,n30,n208);
not (n208,n42);
or (n209,n31,n210);
not (n210,n211);
nor (n211,n212,n215);
and (n212,n213,n27);
not (n213,n214);
and (n215,n214,n28);
xor (n216,n217,n271);
xor (n217,n218,n241);
xor (n218,n219,n233);
xor (n219,n220,n227);
nand (n220,n221,n223);
or (n221,n222,n57);
not (n222,n69);
nand (n223,n63,n224);
nor (n224,n225,n226);
and (n225,n121,n56);
and (n226,n119,n52);
nand (n227,n228,n229);
or (n228,n76,n96);
nand (n229,n78,n230);
nor (n230,n231,n232);
and (n231,n53,n84);
and (n232,n54,n85);
nand (n233,n234,n239);
or (n234,n128,n235);
not (n235,n236);
nand (n236,n237,n238);
or (n237,n66,n25);
or (n238,n65,n26);
nand (n239,n240,n108);
not (n240,n123);
xor (n241,n242,n258);
xor (n242,n243,n250);
nand (n243,n244,n245);
or (n244,n151,n131);
nand (n245,n246,n134);
not (n246,n247);
nor (n247,n248,n249);
and (n248,n143,n92);
and (n249,n141,n91);
nand (n250,n251,n252);
or (n251,n158,n175);
nand (n252,n253,n257);
not (n253,n254);
nor (n254,n255,n256);
and (n255,n166,n148);
and (n256,n167,n147);
not (n257,n159);
and (n258,n259,n264);
nor (n259,n260,n166);
nor (n260,n261,n263);
and (n261,n262,n143);
nand (n262,n172,n162);
and (n263,n171,n161);
nand (n264,n265,n270);
or (n265,n190,n266);
not (n266,n267);
nor (n267,n268,n269);
and (n268,n213,n198);
and (n269,n214,n36);
nand (n270,n194,n192);
or (n271,n272,n318);
and (n272,n273,n293);
xor (n273,n274,n275);
xor (n274,n259,n264);
or (n275,n276,n292);
and (n276,n277,n286);
xor (n277,n278,n279);
and (n278,n257,n172);
nand (n279,n280,n285);
or (n280,n281,n30);
not (n281,n282);
nor (n282,n283,n284);
and (n283,n127,n27);
and (n284,n125,n28);
nand (n285,n32,n23);
nand (n286,n287,n288);
or (n287,n49,n62);
or (n288,n57,n289);
nor (n289,n290,n291);
and (n290,n56,n99);
and (n291,n52,n98);
and (n292,n278,n279);
or (n293,n294,n317);
and (n294,n295,n310);
xor (n295,n296,n303);
nand (n296,n297,n302);
or (n297,n298,n76);
not (n298,n299);
nand (n299,n300,n301);
or (n300,n153,n85);
or (n301,n84,n154);
nand (n302,n89,n78);
nand (n303,n304,n305);
or (n304,n191,n266);
nand (n305,n306,n309);
nor (n306,n307,n308);
and (n307,n44,n198);
and (n308,n45,n36);
not (n309,n190);
nand (n310,n311,n316);
or (n311,n312,n131);
not (n312,n313);
nand (n313,n314,n315);
or (n314,n141,n179);
or (n315,n143,n177);
nand (n316,n145,n134);
and (n317,n296,n303);
and (n318,n274,n275);
or (n319,n320,n372);
and (n320,n321,n324);
xor (n321,n322,n323);
xor (n322,n104,n156);
xor (n323,n19,n74);
or (n324,n325,n371);
and (n325,n326,n348);
xor (n326,n327,n333);
nand (n327,n328,n332);
or (n328,n107,n329);
nor (n329,n330,n331);
and (n330,n65,n71);
and (n331,n66,n73);
or (n332,n117,n128);
nor (n333,n334,n342);
not (n334,n335);
nand (n335,n336,n341);
or (n336,n337,n30);
not (n337,n338);
nand (n338,n339,n340);
or (n339,n28,n121);
or (n340,n27,n119);
nand (n341,n32,n282);
nand (n342,n343,n141);
nand (n343,n344,n345);
or (n344,n172,n137);
nand (n345,n346,n84);
not (n346,n347);
and (n347,n172,n137);
or (n348,n349,n370);
and (n349,n350,n363);
xor (n350,n351,n357);
nand (n351,n352,n356);
or (n352,n57,n353);
nor (n353,n354,n355);
and (n354,n56,n92);
and (n355,n52,n91);
or (n356,n289,n62);
nand (n357,n358,n359);
or (n358,n298,n95);
nand (n359,n77,n360);
nand (n360,n361,n362);
or (n361,n85,n147);
or (n362,n84,n148);
nand (n363,n364,n368);
or (n364,n365,n190);
nor (n365,n366,n367);
and (n366,n198,n26);
and (n367,n36,n25);
or (n368,n369,n191);
not (n369,n306);
and (n370,n351,n357);
and (n371,n327,n333);
and (n372,n322,n323);
not (n373,n374);
or (n374,n375,n406);
and (n375,n376,n405);
xor (n376,n377,n378);
xor (n377,n273,n293);
or (n378,n379,n404);
and (n379,n380,n383);
xor (n380,n381,n382);
xor (n381,n295,n310);
xor (n382,n277,n286);
or (n383,n384,n403);
and (n384,n385,n399);
xor (n385,n386,n393);
nand (n386,n387,n388);
or (n387,n312,n133);
nand (n388,n389,n132);
not (n389,n390);
nor (n390,n391,n392);
and (n391,n171,n141);
and (n392,n143,n172);
nand (n393,n394,n398);
or (n394,n107,n395);
nor (n395,n396,n397);
and (n396,n65,n54);
and (n397,n66,n53);
or (n398,n128,n329);
nand (n399,n400,n402);
or (n400,n401,n334);
not (n401,n342);
or (n402,n335,n342);
and (n403,n386,n393);
and (n404,n381,n382);
xor (n405,n321,n324);
and (n406,n377,n378);
nand (n407,n13,n374);
not (n408,n409);
nand (n409,n410,n810);
or (n410,n411,n522);
not (n411,n412);
nor (n412,n413,n469);
nor (n413,n414,n415);
xor (n414,n376,n405);
or (n415,n416,n468);
and (n416,n417,n467);
xor (n417,n418,n419);
xor (n418,n326,n348);
or (n419,n420,n466);
and (n420,n421,n465);
xor (n421,n422,n442);
or (n422,n423,n441);
and (n423,n424,n433);
xor (n424,n425,n426);
and (n425,n134,n172);
nand (n426,n427,n432);
or (n427,n428,n30);
not (n428,n429);
nand (n429,n430,n431);
or (n430,n28,n73);
or (n431,n27,n71);
nand (n432,n32,n338);
nand (n433,n434,n439);
or (n434,n435,n57);
not (n435,n436);
nor (n436,n437,n438);
and (n437,n153,n56);
and (n438,n154,n52);
nand (n439,n440,n63);
not (n440,n353);
and (n441,n425,n426);
or (n442,n443,n464);
and (n443,n444,n458);
xor (n444,n445,n452);
nand (n445,n446,n451);
or (n446,n447,n76);
not (n447,n448);
nor (n448,n449,n450);
and (n449,n179,n84);
and (n450,n177,n85);
nand (n451,n78,n360);
nand (n452,n453,n457);
or (n453,n454,n190);
nor (n454,n455,n456);
and (n455,n198,n125);
and (n456,n36,n127);
or (n457,n365,n191);
nand (n458,n459,n463);
or (n459,n107,n460);
nor (n460,n461,n462);
and (n461,n65,n99);
and (n462,n66,n98);
or (n463,n395,n128);
and (n464,n445,n452);
xor (n465,n350,n363);
and (n466,n422,n442);
xor (n467,n380,n383);
and (n468,n418,n419);
nor (n469,n470,n521);
or (n470,n471,n520);
and (n471,n472,n475);
xor (n472,n473,n474);
xor (n473,n385,n399);
xor (n474,n421,n465);
or (n475,n476,n519);
and (n476,n477,n518);
xor (n477,n478,n493);
and (n478,n479,n485);
and (n479,n480,n85);
nand (n480,n481,n482);
or (n481,n172,n80);
nand (n482,n483,n56);
not (n483,n484);
and (n484,n172,n80);
nand (n485,n486,n487);
or (n486,n428,n31);
nand (n487,n488,n492);
not (n488,n489);
nor (n489,n490,n491);
and (n490,n27,n54);
and (n491,n28,n53);
not (n492,n30);
or (n493,n494,n517);
and (n494,n495,n510);
xor (n495,n496,n503);
nand (n496,n497,n502);
or (n497,n498,n57);
not (n498,n499);
nor (n499,n500,n501);
and (n500,n148,n52);
and (n501,n147,n56);
nand (n502,n63,n436);
nand (n503,n504,n509);
or (n504,n505,n76);
not (n505,n506);
nand (n506,n507,n508);
or (n507,n84,n172);
or (n508,n171,n85);
nand (n509,n78,n448);
nand (n510,n511,n516);
or (n511,n190,n512);
not (n512,n513);
nor (n513,n514,n515);
and (n514,n121,n198);
and (n515,n119,n36);
or (n516,n454,n191);
and (n517,n496,n503);
xor (n518,n424,n433);
and (n519,n478,n493);
and (n520,n473,n474);
xor (n521,n417,n467);
not (n522,n523);
nand (n523,n524,n799,n809);
nand (n524,n525,n659,n666);
nor (n525,n526,n597);
not (n526,n527);
or (n527,n528,n560);
xor (n528,n529,n559);
xor (n529,n530,n531);
xor (n530,n444,n458);
or (n531,n532,n558);
and (n532,n533,n541);
xor (n533,n534,n540);
nand (n534,n535,n539);
or (n535,n107,n536);
nor (n536,n537,n538);
and (n537,n65,n92);
and (n538,n66,n91);
or (n539,n128,n460);
xor (n540,n479,n485);
or (n541,n542,n557);
and (n542,n543,n551);
xor (n543,n544,n545);
and (n544,n78,n172);
nand (n545,n546,n547);
or (n546,n191,n512);
or (n547,n548,n190);
nor (n548,n549,n550);
and (n549,n198,n71);
and (n550,n36,n73);
nand (n551,n552,n556);
or (n552,n57,n553);
nor (n553,n554,n555);
and (n554,n56,n177);
and (n555,n52,n179);
or (n556,n62,n498);
and (n557,n544,n545);
and (n558,n534,n540);
xor (n559,n477,n518);
or (n560,n561,n596);
and (n561,n562,n595);
xor (n562,n563,n564);
xor (n563,n495,n510);
or (n564,n565,n594);
and (n565,n566,n579);
xor (n566,n567,n573);
nand (n567,n568,n572);
or (n568,n30,n569);
nor (n569,n570,n571);
and (n570,n27,n99);
and (n571,n28,n98);
or (n572,n31,n489);
nand (n573,n574,n578);
or (n574,n107,n575);
nor (n575,n576,n577);
and (n576,n65,n154);
and (n577,n66,n153);
or (n578,n536,n128);
and (n579,n580,n587);
nor (n580,n581,n56);
nor (n581,n582,n585);
and (n582,n583,n65);
not (n583,n584);
and (n584,n172,n60);
and (n585,n171,n586);
not (n586,n60);
nand (n587,n588,n593);
or (n588,n589,n190);
not (n589,n590);
nor (n590,n591,n592);
and (n591,n53,n198);
and (n592,n54,n36);
or (n593,n548,n191);
and (n594,n567,n573);
xor (n595,n533,n541);
and (n596,n563,n564);
nand (n597,n598,n653);
not (n598,n599);
nor (n599,n600,n628);
xor (n600,n601,n627);
xor (n601,n602,n626);
or (n602,n603,n625);
and (n603,n604,n619);
xor (n604,n605,n613);
nand (n605,n606,n611);
or (n606,n607,n57);
not (n607,n608);
nand (n608,n609,n610);
or (n609,n56,n172);
or (n610,n52,n171);
nand (n611,n612,n63);
not (n612,n553);
nand (n613,n614,n618);
or (n614,n30,n615);
nor (n615,n616,n617);
and (n616,n27,n92);
and (n617,n28,n91);
or (n618,n569,n31);
nand (n619,n620,n624);
or (n620,n107,n621);
nor (n621,n622,n623);
and (n622,n65,n148);
and (n623,n66,n147);
or (n624,n575,n128);
and (n625,n605,n613);
xor (n626,n543,n551);
xor (n627,n566,n579);
or (n628,n629,n652);
and (n629,n630,n651);
xor (n630,n631,n632);
xor (n631,n580,n587);
or (n632,n633,n650);
and (n633,n634,n643);
xor (n634,n635,n636);
and (n635,n63,n172);
nand (n636,n637,n642);
or (n637,n190,n638);
not (n638,n639);
nor (n639,n640,n641);
and (n640,n99,n36);
and (n641,n98,n198);
nand (n642,n590,n192);
nand (n643,n644,n649);
or (n644,n30,n645);
not (n645,n646);
nor (n646,n647,n648);
and (n647,n153,n27);
and (n648,n154,n28);
or (n649,n31,n615);
and (n650,n635,n636);
xor (n651,n604,n619);
and (n652,n631,n632);
not (n653,n654);
nor (n654,n655,n656);
xor (n655,n562,n595);
or (n656,n657,n658);
and (n657,n601,n627);
and (n658,n602,n626);
nand (n659,n660,n662);
not (n660,n661);
xor (n661,n472,n475);
not (n662,n663);
or (n663,n664,n665);
and (n664,n529,n559);
and (n665,n530,n531);
or (n666,n667,n798);
and (n667,n668,n695);
xor (n668,n669,n694);
or (n669,n670,n693);
and (n670,n671,n692);
xor (n671,n672,n679);
nand (n672,n673,n678);
or (n673,n107,n674);
not (n674,n675);
nor (n675,n676,n677);
and (n676,n177,n66);
and (n677,n179,n65);
or (n678,n621,n128);
and (n679,n680,n686);
nor (n680,n681,n65);
nor (n681,n682,n685);
and (n682,n683,n27);
not (n683,n684);
and (n684,n172,n111);
and (n685,n171,n115);
nand (n686,n687,n688);
or (n687,n191,n638);
nand (n688,n689,n309);
nand (n689,n690,n691);
or (n690,n92,n198);
nand (n691,n198,n92);
xor (n692,n634,n643);
and (n693,n672,n679);
xor (n694,n630,n651);
or (n695,n696,n797);
and (n696,n697,n716);
xor (n697,n698,n715);
or (n698,n699,n714);
and (n699,n700,n713);
xor (n700,n701,n706);
nand (n701,n702,n705);
or (n702,n703,n30);
not (n703,n704);
xor (n704,n147,n27);
nand (n705,n32,n646);
nand (n706,n707,n712);
or (n707,n708,n107);
not (n708,n709);
nand (n709,n710,n711);
or (n710,n65,n172);
or (n711,n171,n66);
nand (n712,n675,n109);
xor (n713,n680,n686);
and (n714,n701,n706);
xor (n715,n671,n692);
or (n716,n717,n796);
and (n717,n718,n740);
xor (n718,n719,n739);
or (n719,n720,n738);
and (n720,n721,n730);
xor (n721,n722,n723);
and (n722,n109,n172);
nand (n723,n724,n729);
or (n724,n725,n30);
not (n725,n726);
nor (n726,n727,n728);
and (n727,n179,n27);
and (n728,n177,n28);
nand (n729,n32,n704);
nand (n730,n731,n736);
or (n731,n190,n732);
not (n732,n733);
nand (n733,n734,n735);
or (n734,n154,n198);
nand (n735,n198,n154);
or (n736,n737,n191);
not (n737,n689);
and (n738,n722,n723);
xor (n739,n700,n713);
nand (n740,n741,n795);
or (n741,n742,n757);
nor (n742,n743,n744);
xor (n743,n721,n730);
nor (n744,n745,n752);
not (n745,n746);
nand (n746,n747,n751);
or (n747,n190,n748);
nor (n748,n749,n750);
and (n749,n147,n36);
and (n750,n148,n198);
nand (n751,n733,n192);
nand (n752,n753,n28);
nand (n753,n754,n756);
or (n754,n755,n36);
and (n755,n172,n35);
or (n756,n172,n35);
nor (n757,n758,n794);
and (n758,n759,n770);
nand (n759,n760,n764);
nor (n760,n761,n762);
and (n761,n752,n746);
and (n762,n763,n745);
not (n763,n752);
nor (n764,n765,n769);
and (n765,n492,n766);
nand (n766,n767,n768);
or (n767,n27,n172);
or (n768,n171,n28);
and (n769,n32,n726);
nand (n770,n771,n793);
or (n771,n772,n787);
not (n772,n773);
nor (n773,n774,n785);
not (n774,n775);
nand (n775,n776,n781);
or (n776,n191,n777);
not (n777,n778);
nor (n778,n779,n780);
and (n779,n179,n198);
and (n780,n177,n36);
nand (n781,n782,n309);
nor (n782,n783,n784);
and (n783,n171,n198);
and (n784,n172,n36);
nand (n785,n786,n36);
nand (n786,n172,n192);
not (n787,n788);
nand (n788,n789,n792);
nor (n789,n790,n791);
nor (n790,n777,n190);
nor (n791,n748,n191);
nand (n792,n172,n32);
or (n793,n789,n792);
nor (n794,n764,n760);
nand (n795,n743,n744);
and (n796,n719,n739);
and (n797,n698,n715);
and (n798,n669,n694);
nand (n799,n800,n659);
or (n800,n801,n803);
not (n801,n802);
nand (n802,n528,n560);
not (n803,n804);
nand (n804,n527,n805);
nand (n805,n806,n808);
or (n806,n654,n807);
nand (n807,n600,n628);
nand (n808,n655,n656);
nand (n809,n661,n663);
not (n810,n811);
nand (n811,n812,n814);
or (n812,n413,n813);
nand (n813,n470,n521);
nand (n814,n414,n415);
or (n815,n409,n10);
not (n816,n817);
nand (n817,n818,n3);
not (n818,n4);
wire s0n819,s1n819,notn819;
or (n819,s0n819,s1n819);
not(notn819,n4);
and (s0n819,notn819,n820);
and (s1n819,n4,1'b0);
wire s0n820,s1n820,notn820;
or (n820,s0n820,s1n820);
not(notn820,n3);
and (s0n820,notn820,n5);
and (s1n820,n3,n821);
xor (n821,n822,n1344);
xor (n822,n823,n1341);
xor (n823,n824,n1340);
xor (n824,n825,n1331);
xor (n825,n826,n1330);
xor (n826,n827,n1316);
xor (n827,n828,n1315);
xor (n828,n829,n1295);
xor (n829,n830,n1294);
xor (n830,n831,n1269);
xor (n831,n832,n1268);
xor (n832,n833,n1236);
xor (n833,n834,n1235);
xor (n834,n835,n1198);
xor (n835,n836,n70);
xor (n836,n837,n1154);
xor (n837,n838,n1153);
xor (n838,n839,n1103);
xor (n839,n840,n1102);
xor (n840,n841,n1046);
xor (n841,n842,n1045);
xor (n842,n843,n986);
xor (n843,n844,n46);
xor (n844,n845,n918);
xor (n845,n846,n917);
xor (n846,n847,n849);
xor (n847,n848,n199);
and (n848,n204,n192);
or (n849,n850,n852);
and (n850,n851,n269);
and (n851,n197,n192);
and (n852,n853,n854);
xor (n853,n851,n269);
or (n854,n855,n857);
and (n855,n856,n308);
and (n856,n214,n192);
and (n857,n858,n859);
xor (n858,n856,n308);
or (n859,n860,n863);
and (n860,n861,n862);
and (n861,n45,n192);
and (n862,n26,n36);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n869);
and (n866,n867,n868);
and (n867,n26,n192);
and (n868,n125,n36);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n874);
and (n872,n873,n515);
and (n873,n125,n192);
and (n874,n875,n876);
xor (n875,n873,n515);
or (n876,n877,n880);
and (n877,n878,n879);
and (n878,n119,n192);
and (n879,n71,n36);
and (n880,n881,n882);
xor (n881,n878,n879);
or (n882,n883,n885);
and (n883,n884,n592);
and (n884,n71,n192);
and (n885,n886,n887);
xor (n886,n884,n592);
or (n887,n888,n890);
and (n888,n889,n640);
and (n889,n54,n192);
and (n890,n891,n892);
xor (n891,n889,n640);
or (n892,n893,n896);
and (n893,n894,n895);
and (n894,n99,n192);
and (n895,n92,n36);
and (n896,n897,n898);
xor (n897,n894,n895);
or (n898,n899,n902);
and (n899,n900,n901);
and (n900,n92,n192);
and (n901,n154,n36);
and (n902,n903,n904);
xor (n903,n900,n901);
or (n904,n905,n908);
and (n905,n906,n907);
and (n906,n154,n192);
and (n907,n148,n36);
and (n908,n909,n910);
xor (n909,n906,n907);
or (n910,n911,n913);
and (n911,n912,n780);
and (n912,n148,n192);
and (n913,n914,n915);
xor (n914,n912,n780);
and (n915,n916,n784);
and (n916,n177,n192);
and (n917,n214,n35);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n853,n854);
and (n921,n45,n35);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n858,n859);
and (n927,n26,n35);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n864,n865);
and (n933,n125,n35);
and (n934,n935,n936);
xor (n935,n932,n933);
or (n936,n937,n940);
and (n937,n938,n939);
xor (n938,n870,n871);
and (n939,n119,n35);
and (n940,n941,n942);
xor (n941,n938,n939);
or (n942,n943,n946);
and (n943,n944,n945);
xor (n944,n875,n876);
and (n945,n71,n35);
and (n946,n947,n948);
xor (n947,n944,n945);
or (n948,n949,n952);
and (n949,n950,n951);
xor (n950,n881,n882);
and (n951,n54,n35);
and (n952,n953,n954);
xor (n953,n950,n951);
or (n954,n955,n958);
and (n955,n956,n957);
xor (n956,n886,n887);
and (n957,n99,n35);
and (n958,n959,n960);
xor (n959,n956,n957);
or (n960,n961,n964);
and (n961,n962,n963);
xor (n962,n891,n892);
and (n963,n92,n35);
and (n964,n965,n966);
xor (n965,n962,n963);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n897,n898);
and (n969,n154,n35);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n903,n904);
and (n975,n148,n35);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n909,n910);
and (n981,n177,n35);
and (n982,n983,n984);
xor (n983,n980,n981);
and (n984,n985,n755);
xor (n985,n914,n915);
or (n986,n987,n989);
and (n987,n988,n29);
xor (n988,n923,n924);
and (n989,n990,n991);
xor (n990,n988,n29);
or (n991,n992,n994);
and (n992,n993,n284);
xor (n993,n929,n930);
and (n994,n995,n996);
xor (n995,n993,n284);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n935,n936);
and (n999,n119,n28);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n941,n942);
and (n1005,n71,n28);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n947,n948);
and (n1011,n54,n28);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
xor (n1016,n953,n954);
and (n1017,n99,n28);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1024);
and (n1021,n1022,n1023);
xor (n1022,n959,n960);
and (n1023,n92,n28);
and (n1024,n1025,n1026);
xor (n1025,n1022,n1023);
or (n1026,n1027,n1029);
and (n1027,n1028,n648);
xor (n1028,n965,n966);
and (n1029,n1030,n1031);
xor (n1030,n1028,n648);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
xor (n1033,n971,n972);
and (n1034,n148,n28);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1040);
and (n1038,n1039,n728);
xor (n1039,n977,n978);
and (n1040,n1041,n1042);
xor (n1041,n1039,n728);
and (n1042,n1043,n1044);
xor (n1043,n983,n984);
and (n1044,n172,n28);
and (n1045,n26,n111);
or (n1046,n1047,n1050);
and (n1047,n1048,n1049);
xor (n1048,n990,n991);
and (n1049,n125,n111);
and (n1050,n1051,n1052);
xor (n1051,n1048,n1049);
or (n1052,n1053,n1056);
and (n1053,n1054,n1055);
xor (n1054,n995,n996);
and (n1055,n119,n111);
and (n1056,n1057,n1058);
xor (n1057,n1054,n1055);
or (n1058,n1059,n1062);
and (n1059,n1060,n1061);
xor (n1060,n1001,n1002);
and (n1061,n71,n111);
and (n1062,n1063,n1064);
xor (n1063,n1060,n1061);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
xor (n1066,n1007,n1008);
and (n1067,n54,n111);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1074);
and (n1071,n1072,n1073);
xor (n1072,n1013,n1014);
and (n1073,n99,n111);
and (n1074,n1075,n1076);
xor (n1075,n1072,n1073);
or (n1076,n1077,n1080);
and (n1077,n1078,n1079);
xor (n1078,n1019,n1020);
and (n1079,n92,n111);
and (n1080,n1081,n1082);
xor (n1081,n1078,n1079);
or (n1082,n1083,n1086);
and (n1083,n1084,n1085);
xor (n1084,n1025,n1026);
and (n1085,n154,n111);
and (n1086,n1087,n1088);
xor (n1087,n1084,n1085);
or (n1088,n1089,n1092);
and (n1089,n1090,n1091);
xor (n1090,n1030,n1031);
and (n1091,n148,n111);
and (n1092,n1093,n1094);
xor (n1093,n1090,n1091);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
xor (n1096,n1036,n1037);
and (n1097,n177,n111);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
and (n1100,n1101,n684);
xor (n1101,n1041,n1042);
and (n1102,n125,n66);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1051,n1052);
and (n1106,n119,n66);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1057,n1058);
and (n1112,n71,n66);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1063,n1064);
and (n1118,n54,n66);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1069,n1070);
and (n1124,n99,n66);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1075,n1076);
and (n1130,n92,n66);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1081,n1082);
and (n1136,n154,n66);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1087,n1088);
and (n1142,n148,n66);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1148);
and (n1146,n1147,n676);
xor (n1147,n1093,n1094);
and (n1148,n1149,n1150);
xor (n1149,n1147,n676);
and (n1150,n1151,n1152);
xor (n1151,n1099,n1100);
and (n1152,n172,n66);
and (n1153,n119,n60);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1108,n1109);
and (n1157,n71,n60);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1114,n1115);
and (n1163,n54,n60);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1120,n1121);
and (n1169,n99,n60);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
or (n1172,n1173,n1176);
and (n1173,n1174,n1175);
xor (n1174,n1126,n1127);
and (n1175,n92,n60);
and (n1176,n1177,n1178);
xor (n1177,n1174,n1175);
or (n1178,n1179,n1182);
and (n1179,n1180,n1181);
xor (n1180,n1132,n1133);
and (n1181,n154,n60);
and (n1182,n1183,n1184);
xor (n1183,n1180,n1181);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1138,n1139);
and (n1187,n148,n60);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1144,n1145);
and (n1193,n177,n60);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
and (n1196,n1197,n584);
xor (n1197,n1149,n1150);
or (n1198,n1199,n1202);
and (n1199,n1200,n1201);
xor (n1200,n1159,n1160);
and (n1201,n54,n52);
and (n1202,n1203,n1204);
xor (n1203,n1200,n1201);
or (n1204,n1205,n1208);
and (n1205,n1206,n1207);
xor (n1206,n1165,n1166);
and (n1207,n99,n52);
and (n1208,n1209,n1210);
xor (n1209,n1206,n1207);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1171,n1172);
and (n1213,n92,n52);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1219);
and (n1217,n1218,n438);
xor (n1218,n1177,n1178);
and (n1219,n1220,n1221);
xor (n1220,n1218,n438);
or (n1221,n1222,n1224);
and (n1222,n1223,n500);
xor (n1223,n1183,n1184);
and (n1224,n1225,n1226);
xor (n1225,n1223,n500);
or (n1226,n1227,n1230);
and (n1227,n1228,n1229);
xor (n1228,n1189,n1190);
and (n1229,n177,n52);
and (n1230,n1231,n1232);
xor (n1231,n1228,n1229);
and (n1232,n1233,n1234);
xor (n1233,n1195,n1196);
and (n1234,n172,n52);
and (n1235,n54,n80);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1203,n1204);
and (n1239,n99,n80);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1246);
and (n1243,n1244,n1245);
xor (n1244,n1209,n1210);
and (n1245,n92,n80);
and (n1246,n1247,n1248);
xor (n1247,n1244,n1245);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1215,n1216);
and (n1251,n154,n80);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1220,n1221);
and (n1257,n148,n80);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1225,n1226);
and (n1263,n177,n80);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
and (n1266,n1267,n484);
xor (n1267,n1231,n1232);
and (n1268,n99,n85);
or (n1269,n1270,n1272);
and (n1270,n1271,n93);
xor (n1271,n1241,n1242);
and (n1272,n1273,n1274);
xor (n1273,n1271,n93);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1247,n1248);
and (n1277,n154,n85);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1253,n1254);
and (n1283,n148,n85);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1289);
and (n1287,n1288,n450);
xor (n1288,n1259,n1260);
and (n1289,n1290,n1291);
xor (n1290,n1288,n450);
and (n1291,n1292,n1293);
xor (n1292,n1265,n1266);
and (n1293,n172,n85);
and (n1294,n92,n137);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1273,n1274);
and (n1298,n154,n137);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1279,n1280);
and (n1304,n148,n137);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1285,n1286);
and (n1310,n177,n137);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
and (n1313,n1314,n347);
xor (n1314,n1290,n1291);
and (n1315,n154,n141);
or (n1316,n1317,n1319);
and (n1317,n1318,n149);
xor (n1318,n1300,n1301);
and (n1319,n1320,n1321);
xor (n1320,n1318,n149);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1306,n1307);
and (n1324,n177,n141);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
and (n1327,n1328,n1329);
xor (n1328,n1312,n1313);
and (n1329,n172,n141);
and (n1330,n148,n162);
or (n1331,n1332,n1335);
and (n1332,n1333,n1334);
xor (n1333,n1320,n1321);
and (n1334,n177,n162);
and (n1335,n1336,n1337);
xor (n1336,n1333,n1334);
and (n1337,n1338,n1339);
xor (n1338,n1326,n1327);
not (n1339,n262);
and (n1340,n177,n167);
and (n1341,n1342,n1343);
xor (n1342,n1336,n1337);
and (n1343,n172,n167);
not (n1344,n1345);
nand (n1345,n172,n186);
endmodule
