module top (out,n5,n6,n15,n19,n20,n23,n24,n53,n59
        ,n68,n105,n109,n157,n187,n240,n342,n351,n354,n357
        ,n385,n436,n511,n563);
output out;
input n5;
input n6;
input n15;
input n19;
input n20;
input n23;
input n24;
input n53;
input n59;
input n68;
input n105;
input n109;
input n157;
input n187;
input n240;
input n342;
input n351;
input n354;
input n357;
input n385;
input n436;
input n511;
input n563;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n352;
wire n353;
wire n355;
wire n356;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
xor (out,n0,n741);
xor (n0,n1,n662);
xor (n1,n2,n339);
xor (n2,n3,n41);
xor (n3,n4,n7);
and (n4,n5,n6);
or (n7,n8,n35,n40);
and (n8,n9,n32);
or (n9,n10,n29,n31);
and (n10,n11,n26);
or (n11,n12,n21,n25);
and (n12,n13,n18);
nor (n13,n14,n16);
not (n14,n15);
and (n16,n17,n15);
not (n17,n6);
and (n18,n19,n20);
and (n21,n18,n22);
and (n22,n23,n24);
and (n25,n13,n22);
nor (n26,n27,n28);
not (n27,n19);
and (n28,n17,n19);
and (n29,n26,n30);
and (n30,n23,n20);
and (n31,n11,n30);
nor (n32,n33,n34);
not (n33,n23);
and (n34,n17,n23);
and (n35,n32,n36);
nor (n36,n37,n39);
and (n37,n38,n20);
not (n38,n5);
not (n39,n20);
and (n40,n9,n36);
or (n41,n42,n87);
and (n42,n43,n45);
xor (n43,n44,n36);
xor (n44,n9,n32);
or (n45,n46,n83,n86);
and (n46,n47,n80);
or (n47,n48,n76,n79);
and (n48,n49,n62);
or (n49,n50,n56,n61);
and (n50,n51,n55);
nor (n51,n52,n54);
not (n52,n53);
and (n54,n17,n53);
and (n55,n15,n20);
and (n56,n55,n57);
nor (n57,n58,n60);
and (n58,n38,n59);
not (n60,n59);
and (n61,n51,n57);
or (n62,n63,n73,n75);
and (n63,n64,n72);
or (n64,n65,n69,n71);
and (n65,n66,n67);
and (n66,n15,n24);
and (n67,n19,n68);
and (n69,n67,n70);
and (n70,n23,n59);
and (n71,n66,n70);
and (n72,n19,n24);
and (n73,n72,n74);
and (n74,n23,n68);
and (n75,n64,n74);
and (n76,n62,n77);
xor (n77,n78,n22);
xor (n78,n13,n18);
and (n79,n49,n77);
nor (n80,n81,n82);
and (n81,n38,n24);
not (n82,n24);
and (n83,n80,n84);
xor (n84,n85,n30);
xor (n85,n11,n26);
and (n86,n47,n84);
and (n87,n88,n89);
xor (n88,n43,n45);
or (n89,n90,n128);
and (n90,n91,n93);
xor (n91,n92,n84);
xor (n92,n47,n80);
or (n93,n94,n124,n127);
and (n94,n95,n121);
or (n95,n96,n117,n120);
and (n96,n97,n115);
or (n97,n98,n111,n114);
and (n98,n99,n107);
or (n99,n100,n103,n106);
and (n100,n101,n102);
and (n101,n15,n68);
and (n102,n19,n59);
and (n103,n102,n104);
and (n104,n23,n105);
and (n106,n101,n104);
and (n107,n108,n110);
and (n108,n109,n20);
and (n110,n53,n24);
and (n111,n107,n112);
xor (n112,n113,n70);
xor (n113,n66,n67);
and (n114,n99,n112);
xor (n115,n116,n57);
xor (n116,n51,n55);
and (n117,n115,n118);
xor (n118,n119,n74);
xor (n119,n64,n72);
and (n120,n97,n118);
nor (n121,n122,n123);
and (n122,n38,n68);
not (n123,n68);
and (n124,n121,n125);
xor (n125,n126,n77);
xor (n126,n49,n62);
and (n127,n95,n125);
and (n128,n129,n130);
xor (n129,n91,n93);
or (n130,n131,n174);
and (n131,n132,n134);
xor (n132,n133,n125);
xor (n133,n95,n121);
or (n134,n135,n170,n173);
and (n135,n136,n147);
or (n136,n137,n142,n146);
and (n137,n138,n141);
nor (n138,n139,n140);
not (n139,n109);
and (n140,n17,n109);
and (n141,n53,n20);
and (n142,n141,n143);
nor (n143,n144,n145);
and (n144,n38,n105);
not (n145,n105);
and (n146,n138,n143);
or (n147,n148,n166,n169);
and (n148,n149,n164);
or (n149,n150,n161,n163);
and (n150,n151,n159);
or (n151,n152,n155,n158);
and (n152,n153,n154);
and (n153,n15,n59);
and (n154,n19,n105);
and (n155,n154,n156);
and (n156,n23,n157);
and (n158,n153,n156);
xor (n159,n160,n104);
xor (n160,n101,n102);
and (n161,n159,n162);
xor (n162,n108,n110);
and (n163,n151,n162);
xor (n164,n165,n143);
xor (n165,n138,n141);
and (n166,n164,n167);
xor (n167,n168,n112);
xor (n168,n99,n107);
and (n169,n149,n167);
and (n170,n147,n171);
xor (n171,n172,n118);
xor (n172,n97,n115);
and (n173,n136,n171);
and (n174,n175,n176);
xor (n175,n132,n134);
or (n176,n177,n223);
and (n177,n178,n180);
xor (n178,n179,n171);
xor (n179,n136,n147);
or (n180,n181,n219,n222);
and (n181,n182,n200);
or (n182,n183,n195,n199);
and (n183,n184,n192);
or (n184,n185,n189,n191);
and (n185,n186,n188);
and (n186,n187,n20);
and (n188,n109,n24);
and (n189,n188,n190);
and (n190,n53,n68);
and (n191,n186,n190);
nor (n192,n193,n194);
not (n193,n187);
and (n194,n17,n187);
and (n195,n192,n196);
nor (n196,n197,n198);
and (n197,n38,n157);
not (n198,n157);
and (n199,n184,n196);
or (n200,n201,n215,n218);
and (n201,n202,n213);
or (n202,n203,n209,n212);
and (n203,n204,n207);
and (n204,n205,n206);
and (n205,n15,n105);
and (n206,n19,n157);
xor (n207,n208,n190);
xor (n208,n186,n188);
and (n209,n207,n210);
xor (n210,n211,n156);
xor (n211,n153,n154);
and (n212,n204,n210);
xor (n213,n214,n196);
xor (n214,n184,n192);
and (n215,n213,n216);
xor (n216,n217,n162);
xor (n217,n151,n159);
and (n218,n202,n216);
and (n219,n200,n220);
xor (n220,n221,n167);
xor (n221,n149,n164);
and (n222,n182,n220);
and (n223,n224,n225);
xor (n224,n178,n180);
or (n225,n226,n245);
and (n226,n227,n229);
xor (n227,n228,n220);
xor (n228,n182,n200);
and (n229,n230,n243);
or (n230,n231,n237,n242);
and (n231,n232,n235);
and (n232,n233,n234);
and (n233,n53,n59);
xor (n234,n205,n206);
xor (n235,n236,n210);
xor (n236,n204,n207);
and (n237,n235,n238);
nor (n238,n239,n241);
not (n239,n240);
and (n241,n17,n240);
and (n242,n232,n238);
xor (n243,n244,n216);
xor (n244,n202,n213);
and (n245,n246,n247);
xor (n246,n227,n229);
or (n247,n248,n278);
and (n248,n249,n250);
xor (n249,n230,n243);
or (n250,n251,n274,n277);
and (n251,n252,n259);
or (n252,n253,n256,n258);
and (n253,n254,n255);
and (n254,n240,n20);
and (n255,n187,n24);
and (n256,n255,n257);
and (n257,n109,n68);
and (n258,n254,n257);
or (n259,n260,n271,n273);
and (n260,n261,n269);
or (n261,n262,n265,n268);
and (n262,n263,n264);
and (n263,n109,n105);
and (n264,n53,n157);
and (n265,n266,n267);
and (n266,n53,n105);
and (n267,n15,n157);
and (n268,n262,n267);
xor (n269,n270,n257);
xor (n270,n254,n255);
and (n271,n269,n272);
xor (n272,n233,n234);
and (n273,n261,n272);
and (n274,n259,n275);
xor (n275,n276,n238);
xor (n276,n232,n235);
and (n277,n252,n275);
and (n278,n279,n280);
xor (n279,n249,n250);
or (n280,n281,n309);
and (n281,n282,n284);
xor (n282,n283,n275);
xor (n283,n252,n259);
or (n284,n285,n305,n308);
and (n285,n286,n289);
and (n286,n287,n288);
and (n287,n187,n68);
and (n288,n109,n59);
or (n289,n290,n301,n304);
and (n290,n291,n300);
or (n291,n292,n297,n299);
and (n292,n293,n296);
and (n293,n294,n295);
and (n294,n187,n105);
and (n295,n109,n157);
and (n296,n187,n59);
and (n297,n296,n298);
xor (n298,n263,n264);
and (n299,n293,n298);
xor (n300,n287,n288);
and (n301,n300,n302);
xor (n302,n303,n267);
xor (n303,n262,n266);
and (n304,n291,n302);
and (n305,n289,n306);
xor (n306,n307,n272);
xor (n307,n261,n269);
and (n308,n286,n306);
and (n309,n310,n311);
xor (n310,n282,n284);
or (n311,n312,n334);
and (n312,n313,n315);
xor (n313,n314,n306);
xor (n314,n286,n289);
and (n315,n316,n332);
or (n316,n317,n328,n331);
and (n317,n318,n327);
or (n318,n319,n324,n326);
and (n319,n320,n323);
and (n320,n321,n322);
and (n321,n240,n105);
and (n322,n187,n157);
and (n323,n240,n59);
and (n324,n323,n325);
xor (n325,n294,n295);
and (n326,n320,n325);
and (n327,n240,n68);
and (n328,n327,n329);
xor (n329,n330,n298);
xor (n330,n293,n296);
and (n331,n318,n329);
xor (n332,n333,n302);
xor (n333,n291,n300);
and (n334,n335,n336);
xor (n335,n313,n315);
and (n336,n337,n338);
and (n337,n240,n24);
xor (n338,n316,n332);
xor (n339,n340,n373);
xor (n340,n341,n343);
and (n341,n342,n6);
or (n343,n344,n368,n372);
and (n344,n345,n365);
or (n345,n346,n362,n364);
and (n346,n347,n359);
or (n347,n348,n355,n358);
and (n348,n349,n353);
nor (n349,n350,n352);
not (n350,n351);
and (n352,n17,n351);
and (n353,n354,n20);
and (n355,n353,n356);
and (n356,n357,n24);
and (n358,n349,n356);
nor (n359,n360,n361);
not (n360,n354);
and (n361,n17,n354);
and (n362,n359,n363);
and (n363,n357,n20);
and (n364,n347,n363);
nor (n365,n366,n367);
not (n366,n357);
and (n367,n17,n357);
and (n368,n365,n369);
nor (n369,n370,n39);
and (n370,n371,n20);
not (n371,n342);
and (n372,n345,n369);
or (n373,n374,n415);
and (n374,n375,n377);
xor (n375,n376,n369);
xor (n376,n345,n365);
or (n377,n378,n411,n414);
and (n378,n379,n409);
or (n379,n380,n405,n408);
and (n380,n381,n392);
or (n381,n382,n388,n391);
and (n382,n383,n387);
nor (n383,n384,n386);
not (n384,n385);
and (n386,n17,n385);
and (n387,n351,n20);
and (n388,n387,n389);
nor (n389,n390,n60);
and (n390,n371,n59);
and (n391,n383,n389);
or (n392,n393,n402,n404);
and (n393,n394,n401);
or (n394,n395,n398,n400);
and (n395,n396,n397);
and (n396,n351,n24);
and (n397,n354,n68);
and (n398,n397,n399);
and (n399,n357,n59);
and (n400,n396,n399);
and (n401,n354,n24);
and (n402,n401,n403);
and (n403,n357,n68);
and (n404,n394,n403);
and (n405,n392,n406);
xor (n406,n407,n356);
xor (n407,n349,n353);
and (n408,n381,n406);
nor (n409,n410,n82);
and (n410,n371,n24);
and (n411,n409,n412);
xor (n412,n413,n363);
xor (n413,n347,n359);
and (n414,n379,n412);
and (n415,n416,n417);
xor (n416,n375,n377);
or (n417,n418,n454);
and (n418,n419,n421);
xor (n419,n420,n412);
xor (n420,n379,n409);
or (n421,n422,n450,n453);
and (n422,n423,n448);
or (n423,n424,n444,n447);
and (n424,n425,n442);
or (n425,n426,n438,n441);
and (n426,n427,n434);
or (n427,n428,n431,n433);
and (n428,n429,n430);
and (n429,n351,n68);
and (n430,n354,n59);
and (n431,n430,n432);
and (n432,n357,n105);
and (n433,n429,n432);
and (n434,n435,n437);
and (n435,n436,n20);
and (n437,n385,n24);
and (n438,n434,n439);
xor (n439,n440,n399);
xor (n440,n396,n397);
and (n441,n427,n439);
xor (n442,n443,n389);
xor (n443,n383,n387);
and (n444,n442,n445);
xor (n445,n446,n403);
xor (n446,n394,n401);
and (n447,n425,n445);
nor (n448,n449,n123);
and (n449,n371,n68);
and (n450,n448,n451);
xor (n451,n452,n406);
xor (n452,n381,n392);
and (n453,n423,n451);
and (n454,n455,n456);
xor (n455,n419,n421);
or (n456,n457,n498);
and (n457,n458,n460);
xor (n458,n459,n451);
xor (n459,n423,n448);
or (n460,n461,n494,n497);
and (n461,n462,n472);
or (n462,n463,n468,n471);
and (n463,n464,n467);
nor (n464,n465,n466);
not (n465,n436);
and (n466,n17,n436);
and (n467,n385,n20);
and (n468,n467,n469);
nor (n469,n470,n145);
and (n470,n371,n105);
and (n471,n464,n469);
or (n472,n473,n490,n493);
and (n473,n474,n488);
or (n474,n475,n485,n487);
and (n475,n476,n483);
or (n476,n477,n480,n482);
and (n477,n478,n479);
and (n478,n351,n59);
and (n479,n354,n105);
and (n480,n479,n481);
and (n481,n357,n157);
and (n482,n478,n481);
xor (n483,n484,n432);
xor (n484,n429,n430);
and (n485,n483,n486);
xor (n486,n435,n437);
and (n487,n476,n486);
xor (n488,n489,n469);
xor (n489,n464,n467);
and (n490,n488,n491);
xor (n491,n492,n439);
xor (n492,n427,n434);
and (n493,n474,n491);
and (n494,n472,n495);
xor (n495,n496,n445);
xor (n496,n425,n442);
and (n497,n462,n495);
and (n498,n499,n500);
xor (n499,n458,n460);
or (n500,n501,n546);
and (n501,n502,n504);
xor (n502,n503,n495);
xor (n503,n462,n472);
or (n504,n505,n542,n545);
and (n505,n506,n523);
or (n506,n507,n519,n522);
and (n507,n508,n516);
or (n508,n509,n513,n515);
and (n509,n510,n512);
and (n510,n511,n20);
and (n512,n436,n24);
and (n513,n512,n514);
and (n514,n385,n68);
and (n515,n510,n514);
nor (n516,n517,n518);
not (n517,n511);
and (n518,n17,n511);
and (n519,n516,n520);
nor (n520,n521,n198);
and (n521,n371,n157);
and (n522,n508,n520);
or (n523,n524,n538,n541);
and (n524,n525,n536);
or (n525,n526,n532,n535);
and (n526,n527,n530);
and (n527,n528,n529);
and (n528,n351,n105);
and (n529,n354,n157);
xor (n530,n531,n514);
xor (n531,n510,n512);
and (n532,n530,n533);
xor (n533,n534,n481);
xor (n534,n478,n479);
and (n535,n527,n533);
xor (n536,n537,n520);
xor (n537,n508,n516);
and (n538,n536,n539);
xor (n539,n540,n486);
xor (n540,n476,n483);
and (n541,n525,n539);
and (n542,n523,n543);
xor (n543,n544,n491);
xor (n544,n474,n488);
and (n545,n506,n543);
and (n546,n547,n548);
xor (n547,n502,n504);
or (n548,n549,n568);
and (n549,n550,n552);
xor (n550,n551,n543);
xor (n551,n506,n523);
and (n552,n553,n566);
or (n553,n554,n560,n565);
and (n554,n555,n558);
and (n555,n556,n557);
and (n556,n385,n59);
xor (n557,n528,n529);
xor (n558,n559,n533);
xor (n559,n527,n530);
and (n560,n558,n561);
nor (n561,n562,n564);
not (n562,n563);
and (n564,n17,n563);
and (n565,n555,n561);
xor (n566,n567,n539);
xor (n567,n525,n536);
and (n568,n569,n570);
xor (n569,n550,n552);
or (n570,n571,n601);
and (n571,n572,n573);
xor (n572,n553,n566);
or (n573,n574,n597,n600);
and (n574,n575,n582);
or (n575,n576,n579,n581);
and (n576,n577,n578);
and (n577,n563,n20);
and (n578,n511,n24);
and (n579,n578,n580);
and (n580,n436,n68);
and (n581,n577,n580);
or (n582,n583,n594,n596);
and (n583,n584,n592);
or (n584,n585,n588,n591);
and (n585,n586,n587);
and (n586,n436,n105);
and (n587,n385,n157);
and (n588,n589,n590);
and (n589,n385,n105);
and (n590,n351,n157);
and (n591,n585,n590);
xor (n592,n593,n580);
xor (n593,n577,n578);
and (n594,n592,n595);
xor (n595,n556,n557);
and (n596,n584,n595);
and (n597,n582,n598);
xor (n598,n599,n561);
xor (n599,n555,n558);
and (n600,n575,n598);
and (n601,n602,n603);
xor (n602,n572,n573);
or (n603,n604,n632);
and (n604,n605,n607);
xor (n605,n606,n598);
xor (n606,n575,n582);
or (n607,n608,n628,n631);
and (n608,n609,n612);
and (n609,n610,n611);
and (n610,n511,n68);
and (n611,n436,n59);
or (n612,n613,n624,n627);
and (n613,n614,n623);
or (n614,n615,n620,n622);
and (n615,n616,n619);
and (n616,n617,n618);
and (n617,n511,n105);
and (n618,n436,n157);
and (n619,n511,n59);
and (n620,n619,n621);
xor (n621,n586,n587);
and (n622,n616,n621);
xor (n623,n610,n611);
and (n624,n623,n625);
xor (n625,n626,n590);
xor (n626,n585,n589);
and (n627,n614,n625);
and (n628,n612,n629);
xor (n629,n630,n595);
xor (n630,n584,n592);
and (n631,n609,n629);
and (n632,n633,n634);
xor (n633,n605,n607);
or (n634,n635,n657);
and (n635,n636,n638);
xor (n636,n637,n629);
xor (n637,n609,n612);
and (n638,n639,n655);
or (n639,n640,n651,n654);
and (n640,n641,n650);
or (n641,n642,n647,n649);
and (n642,n643,n646);
and (n643,n644,n645);
and (n644,n563,n105);
and (n645,n511,n157);
and (n646,n563,n59);
and (n647,n646,n648);
xor (n648,n617,n618);
and (n649,n643,n648);
and (n650,n563,n68);
and (n651,n650,n652);
xor (n652,n653,n621);
xor (n653,n616,n619);
and (n654,n641,n652);
xor (n655,n656,n625);
xor (n656,n614,n623);
and (n657,n658,n659);
xor (n658,n636,n638);
and (n659,n660,n661);
and (n660,n563,n24);
xor (n661,n639,n655);
or (n662,n663,n666,n740);
and (n663,n664,n665);
xor (n664,n88,n89);
xor (n665,n416,n417);
and (n666,n665,n667);
or (n667,n668,n671,n739);
and (n668,n669,n670);
xor (n669,n129,n130);
xor (n670,n455,n456);
and (n671,n670,n672);
or (n672,n673,n676,n738);
and (n673,n674,n675);
xor (n674,n175,n176);
xor (n675,n499,n500);
and (n676,n675,n677);
or (n677,n678,n681,n737);
and (n678,n679,n680);
xor (n679,n224,n225);
xor (n680,n547,n548);
and (n681,n680,n682);
or (n682,n683,n686,n736);
and (n683,n684,n685);
xor (n684,n246,n247);
xor (n685,n569,n570);
and (n686,n685,n687);
or (n687,n688,n691,n735);
and (n688,n689,n690);
xor (n689,n279,n280);
xor (n690,n602,n603);
and (n691,n690,n692);
or (n692,n693,n696,n734);
and (n693,n694,n695);
xor (n694,n310,n311);
xor (n695,n633,n634);
and (n696,n695,n697);
or (n697,n698,n701,n733);
and (n698,n699,n700);
xor (n699,n335,n336);
xor (n700,n658,n659);
and (n701,n700,n702);
or (n702,n703,n706,n732);
and (n703,n704,n705);
xor (n704,n337,n338);
xor (n705,n660,n661);
and (n706,n705,n707);
or (n707,n708,n713,n731);
and (n708,n709,n711);
xor (n709,n710,n329);
xor (n710,n318,n327);
xor (n711,n712,n652);
xor (n712,n641,n650);
and (n713,n711,n714);
or (n714,n715,n720,n730);
and (n715,n716,n718);
xor (n716,n717,n325);
xor (n717,n320,n323);
xor (n718,n719,n648);
xor (n719,n643,n646);
and (n720,n718,n721);
or (n721,n722,n725,n729);
and (n722,n723,n724);
xor (n723,n321,n322);
xor (n724,n644,n645);
and (n725,n724,n726);
and (n726,n727,n728);
and (n727,n240,n157);
and (n728,n563,n157);
and (n729,n723,n726);
and (n730,n716,n721);
and (n731,n709,n714);
and (n732,n704,n707);
and (n733,n699,n702);
and (n734,n694,n697);
and (n735,n689,n692);
and (n736,n684,n687);
and (n737,n679,n682);
and (n738,n674,n677);
and (n739,n669,n672);
and (n740,n664,n667);
xor (n741,n742,n842);
xor (n742,n743,n803);
xor (n743,n744,n796);
xor (n744,n745,n793);
or (n745,n746,n790,n792);
and (n746,n747,n787);
or (n747,n748,n778,n786);
and (n748,n749,n771);
nor (n749,n750,n770);
not (n750,n751);
xor (n751,n752,n753);
xor (n752,n19,n354);
or (n753,n754,n755,n769);
and (n754,n15,n351);
and (n755,n351,n756);
or (n756,n757,n758,n768);
and (n757,n53,n385);
and (n758,n385,n759);
or (n759,n760,n761,n767);
and (n760,n109,n436);
and (n761,n436,n762);
or (n762,n763,n764,n766);
and (n763,n187,n511);
and (n764,n511,n765);
and (n765,n240,n563);
and (n766,n187,n765);
and (n767,n109,n762);
and (n768,n53,n759);
and (n769,n15,n756);
and (n770,n17,n751);
and (n771,n772,n20);
xor (n772,n773,n774);
xor (n773,n23,n357);
or (n774,n775,n776,n777);
and (n775,n19,n354);
and (n776,n354,n753);
and (n777,n19,n753);
and (n778,n771,n779);
and (n779,n780,n24);
xor (n780,n781,n782);
xor (n781,n5,n342);
or (n782,n783,n784,n785);
and (n783,n23,n357);
and (n784,n357,n774);
and (n785,n23,n774);
and (n786,n749,n779);
nor (n787,n788,n789);
not (n788,n772);
and (n789,n17,n772);
and (n790,n787,n791);
and (n791,n780,n20);
and (n792,n747,n791);
nor (n793,n794,n795);
not (n794,n780);
and (n795,n17,n780);
nor (n796,n797,n39);
and (n797,n798,n20);
not (n798,n799);
or (n799,n800,n801,n802);
and (n800,n5,n342);
and (n801,n342,n782);
and (n802,n5,n782);
or (n803,n804,n838,n841);
and (n804,n805,n836);
or (n805,n806,n832,n835);
and (n806,n807,n819);
or (n807,n808,n815,n818);
and (n808,n809,n814);
nor (n809,n810,n813);
not (n810,n811);
xor (n811,n812,n756);
xor (n812,n15,n351);
and (n813,n17,n811);
and (n814,n751,n20);
and (n815,n814,n816);
nor (n816,n817,n60);
and (n817,n798,n59);
and (n818,n809,n816);
or (n819,n820,n829,n831);
and (n820,n821,n828);
or (n821,n822,n825,n827);
and (n822,n823,n824);
and (n823,n751,n24);
and (n824,n772,n68);
and (n825,n824,n826);
and (n826,n780,n59);
and (n827,n823,n826);
and (n828,n772,n24);
and (n829,n828,n830);
and (n830,n780,n68);
and (n831,n821,n830);
and (n832,n819,n833);
xor (n833,n834,n779);
xor (n834,n749,n771);
and (n835,n807,n833);
nor (n836,n837,n82);
and (n837,n798,n24);
and (n838,n836,n839);
xor (n839,n840,n791);
xor (n840,n747,n787);
and (n841,n805,n839);
or (n842,n843,n888);
and (n843,n844,n846);
xor (n844,n845,n839);
xor (n845,n805,n836);
or (n846,n847,n884,n887);
and (n847,n848,n882);
or (n848,n849,n878,n881);
and (n849,n850,n876);
or (n850,n851,n872,n875);
and (n851,n852,n859);
or (n852,n853,n856,n858);
and (n853,n854,n855);
and (n854,n751,n68);
and (n855,n772,n59);
and (n856,n855,n857);
and (n857,n780,n105);
and (n858,n854,n857);
or (n859,n860,n869,n871);
and (n860,n861,n866);
nor (n861,n862,n865);
not (n862,n863);
xor (n863,n864,n762);
xor (n864,n109,n436);
and (n865,n17,n863);
and (n866,n867,n20);
xor (n867,n868,n759);
xor (n868,n53,n385);
and (n869,n866,n870);
and (n870,n811,n24);
and (n871,n861,n870);
and (n872,n859,n873);
xor (n873,n874,n826);
xor (n874,n823,n824);
and (n875,n852,n873);
xor (n876,n877,n816);
xor (n877,n809,n814);
and (n878,n876,n879);
xor (n879,n880,n830);
xor (n880,n821,n828);
and (n881,n850,n879);
nor (n882,n883,n123);
and (n883,n798,n68);
and (n884,n882,n885);
xor (n885,n886,n833);
xor (n886,n807,n819);
and (n887,n848,n885);
and (n888,n889,n890);
xor (n889,n844,n846);
or (n890,n891,n933);
and (n891,n892,n894);
xor (n892,n893,n885);
xor (n893,n848,n882);
or (n894,n895,n929,n932);
and (n895,n896,n906);
or (n896,n897,n902,n905);
and (n897,n898,n901);
nor (n898,n899,n900);
not (n899,n867);
and (n900,n17,n867);
and (n901,n811,n20);
and (n902,n901,n903);
nor (n903,n904,n145);
and (n904,n798,n105);
and (n905,n898,n903);
or (n906,n907,n925,n928);
and (n907,n908,n923);
or (n908,n909,n919,n922);
and (n909,n910,n917);
or (n910,n911,n914,n916);
and (n911,n912,n913);
and (n912,n751,n59);
and (n913,n772,n105);
and (n914,n913,n915);
and (n915,n780,n157);
and (n916,n912,n915);
xor (n917,n918,n857);
xor (n918,n854,n855);
and (n919,n917,n920);
xor (n920,n921,n870);
xor (n921,n861,n866);
and (n922,n910,n920);
xor (n923,n924,n903);
xor (n924,n898,n901);
and (n925,n923,n926);
xor (n926,n927,n873);
xor (n927,n852,n859);
and (n928,n908,n926);
and (n929,n906,n930);
xor (n930,n931,n879);
xor (n931,n850,n876);
and (n932,n896,n930);
and (n933,n934,n935);
xor (n934,n892,n894);
or (n935,n936,n975);
and (n936,n937,n939);
xor (n937,n938,n930);
xor (n938,n896,n906);
or (n939,n940,n971,n974);
and (n940,n941,n951);
and (n941,n942,n949);
or (n942,n943,n946,n948);
and (n943,n944,n945);
and (n944,n863,n20);
and (n945,n867,n24);
and (n946,n945,n947);
and (n947,n811,n68);
and (n948,n944,n947);
nor (n949,n950,n198);
and (n950,n798,n157);
or (n951,n952,n968,n970);
and (n952,n953,n966);
or (n953,n954,n962,n965);
and (n954,n955,n960);
nor (n955,n956,n959);
not (n956,n957);
xor (n957,n958,n765);
xor (n958,n187,n511);
and (n959,n17,n957);
xor (n960,n961,n915);
xor (n961,n912,n913);
and (n962,n960,n963);
xor (n963,n964,n947);
xor (n964,n944,n945);
and (n965,n955,n963);
xor (n966,n967,n920);
xor (n967,n910,n917);
and (n968,n966,n969);
xor (n969,n942,n949);
and (n970,n953,n969);
and (n971,n951,n972);
xor (n972,n973,n926);
xor (n973,n908,n923);
and (n974,n941,n972);
and (n975,n976,n977);
xor (n976,n937,n939);
or (n977,n978,n1015);
and (n978,n979,n981);
xor (n979,n980,n972);
xor (n980,n941,n951);
or (n981,n982,n1011,n1014);
and (n982,n983,n994);
and (n983,n984,n991);
or (n984,n985,n988,n990);
and (n985,n986,n987);
and (n986,n863,n24);
and (n987,n867,n68);
and (n988,n987,n989);
and (n989,n811,n59);
and (n990,n986,n989);
and (n991,n992,n993);
and (n992,n751,n105);
and (n993,n772,n157);
or (n994,n995,n1007,n1010);
and (n995,n996,n1006);
or (n996,n997,n1003,n1005);
and (n997,n998,n1001);
and (n998,n999,n1000);
and (n999,n811,n105);
and (n1000,n751,n157);
xor (n1001,n1002,n989);
xor (n1002,n986,n987);
and (n1003,n1001,n1004);
xor (n1004,n992,n993);
and (n1005,n998,n1004);
xor (n1006,n984,n991);
and (n1007,n1006,n1008);
xor (n1008,n1009,n963);
xor (n1009,n955,n960);
and (n1010,n996,n1008);
and (n1011,n994,n1012);
xor (n1012,n1013,n969);
xor (n1013,n953,n966);
and (n1014,n983,n1012);
and (n1015,n1016,n1017);
xor (n1016,n979,n981);
or (n1017,n1018,n1043);
and (n1018,n1019,n1021);
xor (n1019,n1020,n1012);
xor (n1020,n983,n994);
or (n1021,n1022,n1039,n1042);
and (n1022,n1023,n1029);
and (n1023,n1024,n1028);
nor (n1024,n1025,n1027);
not (n1025,n1026);
xor (n1026,n240,n563);
and (n1027,n17,n1026);
and (n1028,n957,n20);
or (n1029,n1030,n1036,n1038);
and (n1030,n1031,n1034);
and (n1031,n1032,n1033);
and (n1032,n867,n59);
xor (n1033,n999,n1000);
xor (n1034,n1035,n1004);
xor (n1035,n998,n1001);
and (n1036,n1034,n1037);
xor (n1037,n1024,n1028);
and (n1038,n1031,n1037);
and (n1039,n1029,n1040);
xor (n1040,n1041,n1008);
xor (n1041,n996,n1006);
and (n1042,n1023,n1040);
and (n1043,n1044,n1045);
xor (n1044,n1019,n1021);
or (n1045,n1046,n1077);
and (n1046,n1047,n1049);
xor (n1047,n1048,n1040);
xor (n1048,n1023,n1029);
or (n1049,n1050,n1073,n1076);
and (n1050,n1051,n1058);
or (n1051,n1052,n1055,n1057);
and (n1052,n1053,n1054);
and (n1053,n1026,n20);
and (n1054,n957,n24);
and (n1055,n1054,n1056);
and (n1056,n863,n68);
and (n1057,n1053,n1056);
or (n1058,n1059,n1070,n1072);
and (n1059,n1060,n1068);
or (n1060,n1061,n1064,n1067);
and (n1061,n1062,n1063);
and (n1062,n863,n105);
and (n1063,n867,n157);
and (n1064,n1065,n1066);
and (n1065,n867,n105);
and (n1066,n811,n157);
and (n1067,n1061,n1066);
xor (n1068,n1069,n1056);
xor (n1069,n1053,n1054);
and (n1070,n1068,n1071);
xor (n1071,n1032,n1033);
and (n1072,n1060,n1071);
and (n1073,n1058,n1074);
xor (n1074,n1075,n1037);
xor (n1075,n1031,n1034);
and (n1076,n1051,n1074);
and (n1077,n1078,n1079);
xor (n1078,n1047,n1049);
or (n1079,n1080,n1108);
and (n1080,n1081,n1083);
xor (n1081,n1082,n1074);
xor (n1082,n1051,n1058);
or (n1083,n1084,n1104,n1107);
and (n1084,n1085,n1088);
and (n1085,n1086,n1087);
and (n1086,n957,n68);
and (n1087,n863,n59);
or (n1088,n1089,n1100,n1103);
and (n1089,n1090,n1099);
or (n1090,n1091,n1096,n1098);
and (n1091,n1092,n1095);
and (n1092,n1093,n1094);
and (n1093,n957,n105);
and (n1094,n863,n157);
and (n1095,n957,n59);
and (n1096,n1095,n1097);
xor (n1097,n1062,n1063);
and (n1098,n1092,n1097);
xor (n1099,n1086,n1087);
and (n1100,n1099,n1101);
xor (n1101,n1102,n1066);
xor (n1102,n1061,n1065);
and (n1103,n1090,n1101);
and (n1104,n1088,n1105);
xor (n1105,n1106,n1071);
xor (n1106,n1060,n1068);
and (n1107,n1085,n1105);
and (n1108,n1109,n1110);
xor (n1109,n1081,n1083);
or (n1110,n1111,n1133);
and (n1111,n1112,n1114);
xor (n1112,n1113,n1105);
xor (n1113,n1085,n1088);
and (n1114,n1115,n1131);
or (n1115,n1116,n1127,n1130);
and (n1116,n1117,n1126);
or (n1117,n1118,n1123,n1125);
and (n1118,n1119,n1122);
and (n1119,n1120,n1121);
and (n1120,n1026,n105);
and (n1121,n957,n157);
and (n1122,n1026,n59);
and (n1123,n1122,n1124);
xor (n1124,n1093,n1094);
and (n1125,n1119,n1124);
and (n1126,n1026,n68);
and (n1127,n1126,n1128);
xor (n1128,n1129,n1097);
xor (n1129,n1092,n1095);
and (n1130,n1117,n1128);
xor (n1131,n1132,n1101);
xor (n1132,n1090,n1099);
and (n1133,n1134,n1135);
xor (n1134,n1112,n1114);
and (n1135,n1136,n1137);
and (n1136,n1026,n24);
xor (n1137,n1115,n1131);
endmodule
