module top (out,n14,n15,n18,n24,n25,n30,n34,n42,n48
        ,n52,n58,n68,n77,n78,n84,n89,n95,n103,n105
        ,n111,n121,n134,n142,n148,n156,n161,n166,n172,n180
        ,n185,n393,n426);
output out;
input n14;
input n15;
input n18;
input n24;
input n25;
input n30;
input n34;
input n42;
input n48;
input n52;
input n58;
input n68;
input n77;
input n78;
input n84;
input n89;
input n95;
input n103;
input n105;
input n111;
input n121;
input n134;
input n142;
input n148;
input n156;
input n161;
input n166;
input n172;
input n180;
input n185;
input n393;
input n426;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n16;
wire n17;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
xor (out,n0,n848);
xor (n0,n1,n438);
xor (n1,n2,n342);
or (n2,n3,n341);
and (n3,n4,n290);
xor (n4,n5,n197);
xor (n5,n6,n125);
xor (n6,n7,n61);
xor (n7,n8,n37);
xor (n8,n9,n19);
nor (n9,n10,n17);
not (n10,n11);
nand (n11,n12,n16);
or (n12,n13,n15);
not (n13,n14);
nand (n16,n13,n15);
not (n17,n18);
nand (n19,n20,n31);
or (n20,n21,n28);
nor (n21,n22,n26);
and (n22,n23,n25);
not (n23,n24);
and (n26,n27,n24);
not (n27,n25);
nand (n28,n24,n29);
not (n29,n30);
or (n31,n32,n29);
nor (n32,n33,n35);
and (n33,n34,n23);
and (n35,n36,n24);
not (n36,n34);
nand (n37,n38,n55);
or (n38,n39,n50);
nand (n39,n40,n45);
nor (n40,n41,n43);
and (n41,n23,n42);
and (n43,n24,n44);
not (n44,n42);
nand (n45,n46,n49);
or (n46,n47,n42);
not (n47,n48);
nand (n49,n47,n42);
nor (n50,n51,n53);
and (n51,n47,n52);
and (n53,n54,n48);
not (n54,n52);
or (n55,n40,n56);
nor (n56,n57,n59);
and (n57,n58,n47);
and (n59,n60,n48);
not (n60,n58);
or (n61,n62,n124);
and (n62,n63,n98);
xor (n63,n64,n72);
nand (n64,n65,n71);
or (n65,n39,n66);
nor (n66,n67,n69);
and (n67,n47,n68);
and (n69,n70,n48);
not (n70,n68);
or (n71,n40,n50);
nand (n72,n73,n92);
or (n73,n74,n87);
nand (n74,n75,n82);
or (n75,n76,n79);
and (n76,n77,n78);
and (n79,n80,n81);
not (n80,n77);
not (n81,n78);
nor (n82,n83,n85);
and (n83,n84,n78);
and (n85,n86,n81);
not (n86,n84);
nor (n87,n88,n90);
and (n88,n89,n86);
and (n90,n91,n84);
not (n91,n89);
or (n92,n75,n93);
nor (n93,n94,n96);
and (n94,n95,n86);
and (n96,n97,n84);
not (n97,n95);
nand (n98,n99,n118);
or (n99,n100,n108);
not (n100,n101);
nand (n101,n102,n106);
or (n102,n103,n104);
not (n104,n105);
or (n106,n107,n105);
not (n107,n103);
nand (n108,n109,n114);
nor (n109,n110,n112);
and (n110,n111,n103);
and (n112,n113,n107);
not (n113,n111);
not (n114,n115);
nor (n115,n116,n117);
and (n116,n84,n111);
and (n117,n86,n113);
or (n118,n119,n114);
nor (n119,n120,n122);
and (n120,n107,n121);
and (n122,n103,n123);
not (n123,n121);
and (n124,n64,n72);
or (n125,n126,n196);
and (n126,n127,n175);
xor (n127,n128,n151);
nand (n128,n129,n145);
or (n129,n130,n140);
nand (n130,n131,n136);
not (n131,n132);
nand (n132,n133,n135);
or (n133,n47,n134);
nand (n135,n134,n47);
nor (n136,n137,n139);
and (n137,n80,n138);
not (n138,n134);
and (n139,n77,n134);
nor (n140,n141,n143);
and (n141,n142,n80);
and (n143,n144,n77);
not (n144,n142);
or (n145,n146,n131);
nor (n146,n147,n149);
and (n147,n148,n80);
and (n149,n150,n77);
not (n150,n148);
nand (n151,n152,n169);
or (n152,n153,n164);
nand (n153,n154,n159);
or (n154,n155,n157);
and (n155,n156,n103);
and (n157,n158,n107);
not (n158,n156);
nand (n159,n160,n162);
or (n160,n158,n161);
or (n162,n163,n156);
not (n163,n161);
nor (n164,n165,n167);
and (n165,n166,n163);
and (n167,n168,n161);
not (n168,n166);
or (n169,n170,n154);
nor (n170,n171,n173);
and (n171,n172,n163);
and (n173,n174,n161);
not (n174,n172);
nand (n175,n176,n188);
or (n176,n177,n183);
not (n177,n178);
nor (n178,n179,n181);
and (n179,n180,n161);
and (n181,n182,n163);
not (n182,n180);
nor (n183,n184,n186);
and (n184,n185,n13);
and (n186,n187,n14);
not (n187,n185);
or (n188,n189,n193);
or (n189,n190,n178);
nor (n190,n191,n192);
and (n191,n13,n180);
and (n192,n182,n14);
nor (n193,n194,n195);
and (n194,n14,n17);
and (n195,n13,n18);
and (n196,n128,n151);
xor (n197,n198,n246);
xor (n198,n199,n226);
xor (n199,n200,n213);
xor (n200,n201,n207);
nand (n201,n202,n203);
or (n202,n153,n170);
or (n203,n204,n154);
nor (n204,n205,n206);
and (n205,n163,n105);
and (n206,n161,n104);
nand (n207,n208,n209);
or (n208,n189,n183);
or (n209,n210,n177);
nor (n210,n211,n212);
and (n211,n166,n13);
and (n212,n168,n14);
and (n213,n214,n220);
nand (n214,n215,n219);
or (n215,n216,n28);
nor (n216,n217,n218);
and (n217,n23,n58);
and (n218,n60,n24);
or (n219,n21,n29);
nor (n220,n221,n13);
nor (n221,n222,n225);
and (n222,n163,n223);
not (n223,n224);
and (n224,n18,n180);
and (n225,n182,n17);
xor (n226,n227,n240);
xor (n227,n228,n234);
nand (n228,n229,n230);
or (n229,n74,n93);
or (n230,n231,n75);
nor (n231,n232,n233);
and (n232,n142,n86);
and (n233,n144,n84);
nand (n234,n235,n236);
or (n235,n108,n119);
or (n236,n237,n114);
nor (n237,n238,n239);
and (n238,n107,n89);
and (n239,n103,n91);
nand (n240,n241,n245);
or (n241,n131,n242);
nor (n242,n243,n244);
and (n243,n68,n80);
and (n244,n70,n77);
or (n245,n130,n146);
or (n246,n247,n289);
and (n247,n248,n267);
xor (n248,n249,n250);
xor (n249,n214,n220);
or (n250,n251,n266);
and (n251,n252,n260);
xor (n252,n253,n254);
nor (n253,n177,n17);
nand (n254,n255,n259);
or (n255,n256,n28);
nor (n256,n257,n258);
and (n257,n23,n52);
and (n258,n54,n24);
or (n259,n216,n29);
nand (n260,n261,n262);
or (n261,n40,n66);
or (n262,n39,n263);
nor (n263,n264,n265);
and (n264,n148,n47);
and (n265,n150,n48);
and (n266,n253,n254);
or (n267,n268,n288);
and (n268,n269,n282);
xor (n269,n270,n276);
nand (n270,n271,n275);
or (n271,n74,n272);
nor (n272,n273,n274);
and (n273,n121,n86);
and (n274,n123,n84);
or (n275,n87,n75);
nand (n276,n277,n278);
or (n277,n114,n100);
or (n278,n108,n279);
nor (n279,n280,n281);
and (n280,n107,n172);
and (n281,n103,n174);
nand (n282,n283,n284);
or (n283,n154,n164);
or (n284,n153,n285);
nor (n285,n286,n287);
and (n286,n185,n163);
and (n287,n187,n161);
and (n288,n270,n276);
and (n289,n249,n250);
or (n290,n291,n340);
and (n291,n292,n295);
xor (n292,n293,n294);
xor (n293,n127,n175);
xor (n294,n63,n98);
or (n295,n296,n339);
and (n296,n297,n317);
xor (n297,n298,n304);
nand (n298,n299,n303);
or (n299,n130,n300);
nor (n300,n301,n302);
and (n301,n95,n80);
and (n302,n97,n77);
or (n303,n131,n140);
and (n304,n305,n311);
nand (n305,n306,n310);
or (n306,n307,n28);
nor (n307,n308,n309);
and (n308,n68,n23);
and (n309,n70,n24);
or (n310,n256,n29);
nor (n311,n312,n163);
nor (n312,n313,n316);
and (n313,n107,n314);
not (n314,n315);
and (n315,n18,n156);
and (n316,n158,n17);
or (n317,n318,n338);
and (n318,n319,n332);
xor (n319,n320,n326);
nand (n320,n321,n325);
or (n321,n39,n322);
nor (n322,n323,n324);
and (n323,n142,n47);
and (n324,n144,n48);
or (n325,n40,n263);
nand (n326,n327,n331);
or (n327,n74,n328);
nor (n328,n329,n330);
and (n329,n105,n86);
and (n330,n104,n84);
or (n331,n272,n75);
nand (n332,n333,n337);
or (n333,n108,n334);
nor (n334,n335,n336);
and (n335,n166,n107);
and (n336,n168,n103);
or (n337,n279,n114);
and (n338,n320,n326);
and (n339,n298,n304);
and (n340,n293,n294);
and (n341,n5,n197);
xor (n342,n343,n376);
xor (n343,n344,n373);
xor (n344,n345,n352);
xor (n345,n346,n349);
or (n346,n347,n348);
and (n347,n227,n240);
and (n348,n228,n234);
or (n349,n350,n351);
and (n350,n200,n213);
and (n351,n201,n207);
xor (n352,n353,n366);
xor (n353,n354,n360);
nand (n354,n355,n356);
or (n355,n108,n237);
or (n356,n357,n114);
nor (n357,n358,n359);
and (n358,n107,n95);
and (n359,n103,n97);
nand (n360,n361,n362);
or (n361,n130,n242);
or (n362,n131,n363);
nor (n363,n364,n365);
and (n364,n52,n80);
and (n365,n54,n77);
nand (n366,n367,n372);
or (n367,n154,n368);
not (n368,n369);
nand (n369,n370,n371);
or (n370,n123,n161);
or (n371,n163,n121);
or (n372,n153,n204);
or (n373,n374,n375);
and (n374,n198,n246);
and (n375,n199,n226);
xor (n376,n377,n412);
xor (n377,n378,n409);
xor (n378,n379,n403);
xor (n379,n380,n386);
nand (n380,n381,n382);
or (n381,n39,n56);
or (n382,n40,n383);
nor (n383,n384,n385);
and (n384,n47,n25);
and (n385,n27,n48);
nand (n386,n387,n399);
or (n387,n388,n396);
not (n388,n389);
nor (n389,n11,n390);
nor (n390,n391,n394);
and (n391,n392,n15);
not (n392,n393);
and (n394,n395,n393);
not (n395,n15);
nor (n396,n397,n398);
and (n397,n393,n17);
and (n398,n392,n18);
or (n399,n400,n10);
nor (n400,n401,n402);
and (n401,n185,n392);
and (n402,n187,n393);
nand (n403,n404,n408);
or (n404,n405,n75);
nor (n405,n406,n407);
and (n406,n148,n86);
and (n407,n150,n84);
or (n408,n74,n231);
or (n409,n410,n411);
and (n410,n6,n125);
and (n411,n7,n61);
xor (n412,n413,n435);
xor (n413,n414,n420);
nand (n414,n415,n416);
or (n415,n189,n210);
or (n416,n417,n177);
nor (n417,n418,n419);
and (n418,n172,n13);
and (n419,n174,n14);
xor (n420,n421,n429);
nand (n421,n422,n423);
or (n422,n32,n28);
or (n423,n424,n29);
nor (n424,n425,n427);
and (n425,n426,n23);
and (n427,n428,n24);
not (n428,n426);
nor (n429,n430,n392);
nor (n430,n431,n434);
and (n431,n13,n432);
not (n432,n433);
and (n433,n18,n15);
and (n434,n395,n17);
or (n435,n436,n437);
and (n436,n8,n37);
and (n437,n9,n19);
or (n438,n439,n847);
and (n439,n440,n471);
xor (n440,n441,n470);
or (n441,n442,n469);
and (n442,n443,n468);
xor (n443,n444,n467);
or (n444,n445,n466);
and (n445,n446,n449);
xor (n446,n447,n448);
xor (n447,n252,n260);
xor (n448,n269,n282);
or (n449,n450,n465);
and (n450,n451,n464);
xor (n451,n452,n458);
nand (n452,n453,n457);
or (n453,n153,n454);
nor (n454,n455,n456);
and (n455,n161,n17);
and (n456,n163,n18);
or (n457,n285,n154);
nand (n458,n459,n463);
or (n459,n130,n460);
nor (n460,n461,n462);
and (n461,n89,n80);
and (n462,n91,n77);
or (n463,n300,n131);
xor (n464,n305,n311);
and (n465,n452,n458);
and (n466,n447,n448);
xor (n467,n248,n267);
xor (n468,n292,n295);
and (n469,n444,n467);
xor (n470,n4,n290);
nand (n471,n472,n844,n846);
or (n472,n473,n839);
nand (n473,n474,n828);
or (n474,n475,n827);
and (n475,n476,n597);
xor (n476,n477,n582);
or (n477,n478,n581);
and (n478,n479,n547);
xor (n479,n480,n502);
xor (n480,n481,n496);
xor (n481,n482,n489);
nand (n482,n483,n488);
or (n483,n74,n484);
not (n484,n485);
nor (n485,n486,n487);
and (n486,n86,n174);
and (n487,n172,n84);
or (n488,n328,n75);
nand (n489,n490,n495);
or (n490,n491,n108);
not (n491,n492);
nand (n492,n493,n494);
or (n493,n187,n103);
or (n494,n185,n107);
or (n495,n334,n114);
nand (n496,n497,n501);
or (n497,n130,n498);
nor (n498,n499,n500);
and (n499,n121,n80);
and (n500,n123,n77);
or (n501,n131,n460);
or (n502,n503,n546);
and (n503,n504,n526);
xor (n504,n505,n511);
nand (n505,n506,n510);
or (n506,n130,n507);
nor (n507,n508,n509);
and (n508,n105,n80);
and (n509,n104,n77);
or (n510,n498,n131);
xor (n511,n512,n518);
nor (n512,n513,n107);
nor (n513,n514,n517);
and (n514,n515,n86);
not (n515,n516);
and (n516,n18,n111);
and (n517,n113,n17);
nand (n518,n519,n522);
or (n519,n28,n520);
not (n520,n521);
xnor (n521,n142,n23);
or (n522,n523,n29);
nor (n523,n524,n525);
and (n524,n23,n148);
and (n525,n150,n24);
or (n526,n527,n545);
and (n527,n528,n536);
xor (n528,n529,n530);
nor (n529,n114,n17);
nand (n530,n531,n532);
or (n531,n29,n520);
or (n532,n533,n28);
nor (n533,n534,n535);
and (n534,n23,n95);
and (n535,n97,n24);
nand (n536,n537,n541);
or (n537,n74,n538);
nor (n538,n539,n540);
and (n539,n185,n86);
and (n540,n187,n84);
or (n541,n542,n75);
nor (n542,n543,n544);
and (n543,n166,n86);
and (n544,n168,n84);
and (n545,n529,n530);
and (n546,n505,n511);
xor (n547,n548,n562);
xor (n548,n549,n550);
and (n549,n512,n518);
xor (n550,n551,n556);
xor (n551,n552,n553);
nor (n552,n154,n17);
nand (n553,n554,n555);
or (n554,n523,n28);
or (n555,n307,n29);
nand (n556,n557,n561);
or (n557,n39,n558);
nor (n558,n559,n560);
and (n559,n95,n47);
and (n560,n97,n48);
or (n561,n40,n322);
or (n562,n563,n580);
and (n563,n564,n574);
xor (n564,n565,n571);
nand (n565,n566,n570);
or (n566,n39,n567);
nor (n567,n568,n569);
and (n568,n47,n89);
and (n569,n91,n48);
or (n570,n558,n40);
nand (n571,n572,n573);
or (n572,n75,n484);
or (n573,n542,n74);
nand (n574,n575,n576);
or (n575,n114,n491);
or (n576,n108,n577);
nor (n577,n578,n579);
and (n578,n103,n17);
and (n579,n107,n18);
and (n580,n565,n571);
and (n581,n480,n502);
xor (n582,n583,n588);
xor (n583,n584,n585);
xor (n584,n319,n332);
or (n585,n586,n587);
and (n586,n548,n562);
and (n587,n549,n550);
xor (n588,n589,n596);
xor (n589,n590,n593);
or (n590,n591,n592);
and (n591,n551,n556);
and (n592,n552,n553);
or (n593,n594,n595);
and (n594,n481,n496);
and (n595,n482,n489);
xor (n596,n451,n464);
or (n597,n598,n826);
and (n598,n599,n636);
xor (n599,n600,n635);
or (n600,n601,n634);
and (n601,n602,n633);
xor (n602,n603,n632);
or (n603,n604,n631);
and (n604,n605,n618);
xor (n605,n606,n612);
nand (n606,n607,n611);
or (n607,n39,n608);
nor (n608,n609,n610);
and (n609,n121,n47);
and (n610,n48,n123);
or (n611,n567,n40);
nand (n612,n613,n617);
or (n613,n130,n614);
nor (n614,n615,n616);
and (n615,n172,n80);
and (n616,n174,n77);
or (n617,n507,n131);
and (n618,n619,n625);
nor (n619,n620,n86);
nor (n620,n621,n624);
and (n621,n622,n80);
not (n622,n623);
and (n623,n18,n78);
and (n624,n81,n17);
nand (n625,n626,n630);
or (n626,n627,n28);
nor (n627,n628,n629);
and (n628,n23,n89);
and (n629,n91,n24);
or (n630,n533,n29);
and (n631,n606,n612);
xor (n632,n564,n574);
xor (n633,n504,n526);
and (n634,n603,n632);
xor (n635,n479,n547);
nand (n636,n637,n823,n825);
or (n637,n638,n696);
nand (n638,n639,n691);
not (n639,n640);
nor (n640,n641,n667);
xor (n641,n642,n666);
xor (n642,n643,n665);
or (n643,n644,n664);
and (n644,n645,n658);
xor (n645,n646,n652);
nand (n646,n647,n651);
or (n647,n74,n648);
nor (n648,n649,n650);
and (n649,n84,n17);
and (n650,n86,n18);
or (n651,n538,n75);
nand (n652,n653,n657);
or (n653,n654,n39);
nor (n654,n655,n656);
and (n655,n48,n104);
and (n656,n47,n105);
or (n657,n608,n40);
nand (n658,n659,n663);
or (n659,n130,n660);
nor (n660,n661,n662);
and (n661,n166,n80);
and (n662,n168,n77);
or (n663,n614,n131);
and (n664,n646,n652);
xor (n665,n528,n536);
xor (n666,n605,n618);
or (n667,n668,n690);
and (n668,n669,n689);
xor (n669,n670,n671);
xor (n670,n619,n625);
or (n671,n672,n688);
and (n672,n673,n682);
xor (n673,n674,n675);
nor (n674,n75,n17);
nand (n675,n676,n681);
or (n676,n677,n28);
not (n677,n678);
nand (n678,n679,n680);
or (n679,n24,n123);
nand (n680,n123,n24);
or (n681,n627,n29);
nand (n682,n683,n687);
or (n683,n39,n684);
nor (n684,n685,n686);
and (n685,n47,n172);
and (n686,n48,n174);
or (n687,n654,n40);
and (n688,n674,n675);
xor (n689,n645,n658);
and (n690,n670,n671);
or (n691,n692,n693);
xor (n692,n602,n633);
or (n693,n694,n695);
and (n694,n642,n666);
and (n695,n643,n665);
nor (n696,n697,n822);
and (n697,n698,n817);
or (n698,n699,n816);
and (n699,n700,n741);
xor (n700,n701,n734);
or (n701,n702,n733);
and (n702,n703,n719);
xor (n703,n704,n710);
nand (n704,n705,n709);
or (n705,n39,n706);
nor (n706,n707,n708);
and (n707,n48,n168);
and (n708,n47,n166);
or (n709,n684,n40);
or (n710,n711,n715);
nor (n711,n712,n131);
nor (n712,n713,n714);
and (n713,n80,n185);
and (n714,n77,n187);
nor (n715,n130,n716);
nor (n716,n717,n718);
and (n717,n77,n17);
and (n718,n80,n18);
xor (n719,n720,n726);
nor (n720,n721,n80);
nor (n721,n722,n725);
and (n722,n723,n47);
not (n723,n724);
and (n724,n18,n134);
and (n725,n138,n17);
nand (n726,n727,n732);
or (n727,n28,n728);
not (n728,n729);
nand (n729,n730,n731);
or (n730,n23,n105);
nand (n731,n105,n23);
nand (n732,n678,n30);
and (n733,n704,n710);
xor (n734,n735,n740);
xor (n735,n736,n739);
nand (n736,n737,n738);
or (n737,n130,n712);
or (n738,n660,n131);
and (n739,n720,n726);
xor (n740,n673,n682);
or (n741,n742,n815);
and (n742,n743,n763);
xor (n743,n744,n762);
or (n744,n745,n761);
and (n745,n746,n755);
xor (n746,n747,n748);
and (n747,n132,n18);
nand (n748,n749,n754);
or (n749,n28,n750);
not (n750,n751);
nand (n751,n752,n753);
or (n752,n24,n174);
nand (n753,n174,n24);
nand (n754,n729,n30);
nand (n755,n756,n760);
or (n756,n39,n757);
nor (n757,n758,n759);
and (n758,n47,n185);
and (n759,n48,n187);
or (n760,n706,n40);
and (n761,n747,n748);
xor (n762,n703,n719);
or (n763,n764,n814);
and (n764,n765,n782);
xor (n765,n766,n781);
and (n766,n767,n773);
and (n767,n768,n48);
nand (n768,n769,n772);
nand (n769,n770,n23);
not (n770,n771);
and (n771,n18,n42);
nand (n772,n44,n17);
nand (n773,n774,n775);
or (n774,n29,n750);
nand (n775,n776,n780);
not (n776,n777);
nor (n777,n778,n779);
and (n778,n168,n24);
and (n779,n166,n23);
not (n780,n28);
xor (n781,n746,n755);
or (n782,n783,n813);
and (n783,n784,n792);
xor (n784,n785,n791);
nand (n785,n786,n790);
or (n786,n39,n787);
nor (n787,n788,n789);
and (n788,n48,n17);
and (n789,n47,n18);
or (n790,n757,n40);
xor (n791,n767,n773);
or (n792,n793,n812);
and (n793,n794,n802);
xor (n794,n795,n796);
nor (n795,n40,n17);
nand (n796,n797,n801);
or (n797,n798,n28);
or (n798,n799,n800);
and (n799,n23,n187);
and (n800,n185,n24);
or (n801,n777,n29);
nor (n802,n803,n810);
nor (n803,n804,n806);
and (n804,n805,n30);
not (n805,n798);
and (n806,n807,n780);
nand (n807,n808,n809);
or (n808,n23,n18);
or (n809,n24,n17);
or (n810,n23,n811);
and (n811,n18,n30);
and (n812,n795,n796);
and (n813,n785,n791);
and (n814,n766,n781);
and (n815,n744,n762);
and (n816,n701,n734);
or (n817,n818,n819);
xor (n818,n669,n689);
or (n819,n820,n821);
and (n820,n735,n740);
and (n821,n736,n739);
and (n822,n818,n819);
nand (n823,n691,n824);
and (n824,n641,n667);
nand (n825,n692,n693);
and (n826,n600,n635);
and (n827,n477,n582);
or (n828,n829,n836);
xor (n829,n830,n835);
xor (n830,n831,n832);
xor (n831,n297,n317);
or (n832,n833,n834);
and (n833,n589,n596);
and (n834,n590,n593);
xor (n835,n446,n449);
or (n836,n837,n838);
and (n837,n583,n588);
and (n838,n584,n585);
nor (n839,n840,n841);
xor (n840,n443,n468);
or (n841,n842,n843);
and (n842,n830,n835);
and (n843,n831,n832);
or (n844,n839,n845);
nand (n845,n829,n836);
nand (n846,n840,n841);
and (n847,n441,n470);
buf (n848,n849);
xor (n849,n850,n1472);
xor (n850,n851,n1470);
xor (n851,n852,n1469);
xor (n852,n853,n1460);
xor (n853,n854,n1459);
xor (n854,n855,n1445);
xor (n855,n856,n1444);
xor (n856,n857,n1423);
xor (n857,n858,n1422);
xor (n858,n859,n1396);
xor (n859,n860,n1395);
xor (n860,n861,n1362);
xor (n861,n862,n1361);
xor (n862,n863,n1323);
xor (n863,n864,n1322);
xor (n864,n865,n1278);
xor (n865,n866,n1277);
xor (n866,n867,n1227);
xor (n867,n868,n1226);
xor (n868,n869,n1169);
xor (n869,n870,n1168);
xor (n870,n871,n1106);
xor (n871,n872,n1105);
xor (n872,n873,n1036);
xor (n873,n874,n1035);
xor (n874,n875,n961);
xor (n875,n876,n960);
xor (n876,n877,n880);
xor (n877,n878,n879);
and (n878,n426,n30);
and (n879,n34,n24);
or (n880,n881,n884);
and (n881,n882,n883);
and (n882,n34,n30);
and (n883,n25,n24);
and (n884,n885,n886);
xor (n885,n882,n883);
or (n886,n887,n890);
and (n887,n888,n889);
and (n888,n25,n30);
and (n889,n58,n24);
and (n890,n891,n892);
xor (n891,n888,n889);
or (n892,n893,n896);
and (n893,n894,n895);
and (n894,n58,n30);
and (n895,n52,n24);
and (n896,n897,n898);
xor (n897,n894,n895);
or (n898,n899,n902);
and (n899,n900,n901);
and (n900,n52,n30);
and (n901,n68,n24);
and (n902,n903,n904);
xor (n903,n900,n901);
or (n904,n905,n908);
and (n905,n906,n907);
and (n906,n68,n30);
and (n907,n148,n24);
and (n908,n909,n910);
xor (n909,n906,n907);
or (n910,n911,n914);
and (n911,n912,n913);
and (n912,n148,n30);
and (n913,n142,n24);
and (n914,n915,n916);
xor (n915,n912,n913);
or (n916,n917,n920);
and (n917,n918,n919);
and (n918,n142,n30);
and (n919,n95,n24);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
and (n924,n95,n30);
and (n925,n89,n24);
and (n926,n927,n928);
xor (n927,n924,n925);
or (n928,n929,n932);
and (n929,n930,n931);
and (n930,n89,n30);
and (n931,n121,n24);
and (n932,n933,n934);
xor (n933,n930,n931);
or (n934,n935,n938);
and (n935,n936,n937);
and (n936,n121,n30);
and (n937,n105,n24);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
and (n942,n105,n30);
and (n943,n172,n24);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
and (n948,n172,n30);
and (n949,n166,n24);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n955);
and (n953,n954,n800);
and (n954,n166,n30);
and (n955,n956,n957);
xor (n956,n954,n800);
and (n957,n958,n959);
and (n958,n185,n30);
and (n959,n18,n24);
and (n960,n25,n42);
or (n961,n962,n965);
and (n962,n963,n964);
xor (n963,n885,n886);
and (n964,n58,n42);
and (n965,n966,n967);
xor (n966,n963,n964);
or (n967,n968,n971);
and (n968,n969,n970);
xor (n969,n891,n892);
and (n970,n52,n42);
and (n971,n972,n973);
xor (n972,n969,n970);
or (n973,n974,n977);
and (n974,n975,n976);
xor (n975,n897,n898);
and (n976,n68,n42);
and (n977,n978,n979);
xor (n978,n975,n976);
or (n979,n980,n983);
and (n980,n981,n982);
xor (n981,n903,n904);
and (n982,n148,n42);
and (n983,n984,n985);
xor (n984,n981,n982);
or (n985,n986,n989);
and (n986,n987,n988);
xor (n987,n909,n910);
and (n988,n142,n42);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
xor (n993,n915,n916);
and (n994,n95,n42);
and (n995,n996,n997);
xor (n996,n993,n994);
or (n997,n998,n1001);
and (n998,n999,n1000);
xor (n999,n921,n922);
and (n1000,n89,n42);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n927,n928);
and (n1006,n121,n42);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1013);
and (n1010,n1011,n1012);
xor (n1011,n933,n934);
and (n1012,n105,n42);
and (n1013,n1014,n1015);
xor (n1014,n1011,n1012);
or (n1015,n1016,n1019);
and (n1016,n1017,n1018);
xor (n1017,n939,n940);
and (n1018,n172,n42);
and (n1019,n1020,n1021);
xor (n1020,n1017,n1018);
or (n1021,n1022,n1025);
and (n1022,n1023,n1024);
xor (n1023,n945,n946);
and (n1024,n166,n42);
and (n1025,n1026,n1027);
xor (n1026,n1023,n1024);
or (n1027,n1028,n1031);
and (n1028,n1029,n1030);
xor (n1029,n951,n952);
and (n1030,n185,n42);
and (n1031,n1032,n1033);
xor (n1032,n1029,n1030);
and (n1033,n1034,n771);
xor (n1034,n956,n957);
and (n1035,n58,n48);
or (n1036,n1037,n1040);
and (n1037,n1038,n1039);
xor (n1038,n966,n967);
and (n1039,n52,n48);
and (n1040,n1041,n1042);
xor (n1041,n1038,n1039);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n972,n973);
and (n1045,n68,n48);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n978,n979);
and (n1051,n148,n48);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n984,n985);
and (n1057,n142,n48);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
or (n1060,n1061,n1064);
and (n1061,n1062,n1063);
xor (n1062,n990,n991);
and (n1063,n95,n48);
and (n1064,n1065,n1066);
xor (n1065,n1062,n1063);
or (n1066,n1067,n1070);
and (n1067,n1068,n1069);
xor (n1068,n996,n997);
and (n1069,n89,n48);
and (n1070,n1071,n1072);
xor (n1071,n1068,n1069);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1002,n1003);
and (n1075,n121,n48);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1008,n1009);
and (n1081,n105,n48);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
xor (n1086,n1014,n1015);
and (n1087,n172,n48);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
xor (n1092,n1020,n1021);
and (n1093,n166,n48);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
or (n1096,n1097,n1100);
and (n1097,n1098,n1099);
xor (n1098,n1026,n1027);
and (n1099,n185,n48);
and (n1100,n1101,n1102);
xor (n1101,n1098,n1099);
and (n1102,n1103,n1104);
xor (n1103,n1032,n1033);
and (n1104,n18,n48);
and (n1105,n52,n134);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1041,n1042);
and (n1109,n68,n134);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1047,n1048);
and (n1115,n148,n134);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1053,n1054);
and (n1121,n142,n134);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1059,n1060);
and (n1127,n95,n134);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1065,n1066);
and (n1133,n89,n134);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1071,n1072);
and (n1139,n121,n134);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1077,n1078);
and (n1145,n105,n134);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1083,n1084);
and (n1151,n172,n134);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1089,n1090);
and (n1157,n166,n134);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1095,n1096);
and (n1163,n185,n134);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
and (n1166,n1167,n724);
xor (n1167,n1101,n1102);
and (n1168,n68,n77);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1111,n1112);
and (n1172,n148,n77);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1117,n1118);
and (n1178,n142,n77);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1123,n1124);
and (n1184,n95,n77);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1129,n1130);
and (n1190,n89,n77);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1135,n1136);
and (n1196,n121,n77);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1203);
and (n1200,n1201,n1202);
xor (n1201,n1141,n1142);
and (n1202,n105,n77);
and (n1203,n1204,n1205);
xor (n1204,n1201,n1202);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1147,n1148);
and (n1208,n172,n77);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1153,n1154);
and (n1214,n166,n77);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1159,n1160);
and (n1220,n185,n77);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
and (n1223,n1224,n1225);
xor (n1224,n1165,n1166);
and (n1225,n18,n77);
and (n1226,n148,n78);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1174,n1175);
and (n1230,n142,n78);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1180,n1181);
and (n1236,n95,n78);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1186,n1187);
and (n1242,n89,n78);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1192,n1193);
and (n1248,n121,n78);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1198,n1199);
and (n1254,n105,n78);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1204,n1205);
and (n1260,n172,n78);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1210,n1211);
and (n1266,n166,n78);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1216,n1217);
and (n1272,n185,n78);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
and (n1275,n1276,n623);
xor (n1276,n1222,n1223);
and (n1277,n142,n84);
or (n1278,n1279,n1282);
and (n1279,n1280,n1281);
xor (n1280,n1232,n1233);
and (n1281,n95,n84);
and (n1282,n1283,n1284);
xor (n1283,n1280,n1281);
or (n1284,n1285,n1288);
and (n1285,n1286,n1287);
xor (n1286,n1238,n1239);
and (n1287,n89,n84);
and (n1288,n1289,n1290);
xor (n1289,n1286,n1287);
or (n1290,n1291,n1294);
and (n1291,n1292,n1293);
xor (n1292,n1244,n1245);
and (n1293,n121,n84);
and (n1294,n1295,n1296);
xor (n1295,n1292,n1293);
or (n1296,n1297,n1300);
and (n1297,n1298,n1299);
xor (n1298,n1250,n1251);
and (n1299,n105,n84);
and (n1300,n1301,n1302);
xor (n1301,n1298,n1299);
or (n1302,n1303,n1305);
and (n1303,n1304,n487);
xor (n1304,n1256,n1257);
and (n1305,n1306,n1307);
xor (n1306,n1304,n487);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1262,n1263);
and (n1310,n166,n84);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1268,n1269);
and (n1316,n185,n84);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
and (n1319,n1320,n1321);
xor (n1320,n1274,n1275);
and (n1321,n18,n84);
and (n1322,n95,n111);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1283,n1284);
and (n1326,n89,n111);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1289,n1290);
and (n1332,n121,n111);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
or (n1335,n1336,n1339);
and (n1336,n1337,n1338);
xor (n1337,n1295,n1296);
and (n1338,n105,n111);
and (n1339,n1340,n1341);
xor (n1340,n1337,n1338);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1301,n1302);
and (n1344,n172,n111);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1351);
and (n1348,n1349,n1350);
xor (n1349,n1306,n1307);
and (n1350,n166,n111);
and (n1351,n1352,n1353);
xor (n1352,n1349,n1350);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1312,n1313);
and (n1356,n185,n111);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
and (n1359,n1360,n516);
xor (n1360,n1318,n1319);
and (n1361,n89,n103);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1328,n1329);
and (n1365,n121,n103);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1334,n1335);
and (n1371,n105,n103);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1340,n1341);
and (n1377,n172,n103);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1346,n1347);
and (n1383,n166,n103);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1352,n1353);
and (n1389,n185,n103);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
and (n1392,n1393,n1394);
xor (n1393,n1358,n1359);
and (n1394,n18,n103);
and (n1395,n121,n156);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1367,n1368);
and (n1399,n105,n156);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1373,n1374);
and (n1405,n172,n156);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1379,n1380);
and (n1411,n166,n156);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1385,n1386);
and (n1417,n185,n156);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
and (n1420,n1421,n315);
xor (n1421,n1391,n1392);
and (n1422,n105,n161);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1401,n1402);
and (n1426,n172,n161);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1407,n1408);
and (n1432,n166,n161);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1413,n1414);
and (n1438,n185,n161);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
and (n1441,n1442,n1443);
xor (n1442,n1419,n1420);
and (n1443,n18,n161);
and (n1444,n172,n180);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1428,n1429);
and (n1448,n166,n180);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1434,n1435);
and (n1454,n185,n180);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
and (n1457,n1458,n224);
xor (n1458,n1440,n1441);
and (n1459,n166,n14);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1450,n1451);
and (n1463,n185,n14);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
and (n1466,n1467,n1468);
xor (n1467,n1456,n1457);
and (n1468,n18,n14);
and (n1469,n185,n15);
and (n1470,n1471,n433);
xor (n1471,n1465,n1466);
and (n1472,n18,n393);
endmodule
