module top (out,n3,n13,n15,n16,n18,n20,n21,n26,n33
        ,n39,n42,n43,n55,n56,n62,n63,n80,n82,n83
        ,n92,n93,n95,n96,n106,n116,n134,n140,n153,n159
        ,n178,n184);
output out;
input n3;
input n13;
input n15;
input n16;
input n18;
input n20;
input n21;
input n26;
input n33;
input n39;
input n42;
input n43;
input n55;
input n56;
input n62;
input n63;
input n80;
input n82;
input n83;
input n92;
input n93;
input n95;
input n96;
input n106;
input n116;
input n134;
input n140;
input n153;
input n159;
input n178;
input n184;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n17;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n94;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
xor (out,n0,n589);
nand (n0,n1,n64);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
xor (n5,n6,n60);
xor (n6,n7,n57);
xor (n7,n8,n53);
xor (n8,n9,n44);
xor (n9,n10,n40);
xor (n10,n11,n22);
xor (n11,n12,n17);
and (n12,n13,n14);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n3);
and (s0n14,notn14,n15);
and (s1n14,n3,n16);
and (n17,n18,n19);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n3);
and (s0n19,notn19,n20);
and (s1n19,n3,n21);
or (n22,n23,n27);
and (n23,n24,n25);
and (n24,n18,n14);
and (n25,n26,n19);
and (n27,n28,n29);
xor (n28,n24,n25);
or (n29,n30,n34);
and (n30,n31,n32);
and (n31,n26,n14);
and (n32,n33,n19);
and (n34,n35,n36);
xor (n35,n31,n32);
and (n36,n37,n38);
and (n37,n33,n14);
and (n38,n39,n19);
and (n40,n26,n41);
wire s0n41,s1n41,notn41;
or (n41,s0n41,s1n41);
not(notn41,n3);
and (s0n41,notn41,n42);
and (s1n41,n3,n43);
or (n44,n45,n48);
and (n45,n46,n47);
xor (n46,n28,n29);
and (n47,n33,n41);
and (n48,n49,n50);
xor (n49,n46,n47);
and (n50,n51,n52);
xor (n51,n35,n36);
and (n52,n39,n41);
and (n53,n33,n54);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n3);
and (s0n54,notn54,n55);
and (s1n54,n3,n56);
and (n57,n58,n59);
xor (n58,n49,n50);
and (n59,n39,n54);
and (n60,n39,n61);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n3);
and (s0n61,notn61,n62);
and (s1n61,n3,n63);
nand (n64,n65,n2);
nand (n65,n66,n588);
or (n66,n67,n293);
not (n67,n68);
nand (n68,n69,n292);
nand (n69,n70,n262);
not (n70,n71);
xor (n71,n72,n222);
xor (n72,n73,n143);
xor (n73,n74,n121);
xor (n74,n75,n110);
nand (n75,n76,n102);
or (n76,n77,n87);
not (n77,n78);
nor (n78,n79,n84);
and (n79,n80,n81);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n3);
and (s0n81,notn81,n82);
and (s1n81,n3,n83);
and (n84,n85,n86);
not (n85,n80);
not (n86,n81);
nand (n87,n88,n99);
nor (n88,n89,n97);
and (n89,n90,n94);
not (n90,n91);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n3);
and (s0n91,notn91,n92);
and (s1n91,n3,n93);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n3);
and (s0n94,notn94,n95);
and (s1n94,n3,n96);
and (n97,n91,n98);
not (n98,n94);
nand (n99,n100,n101);
or (n100,n90,n81);
nand (n101,n81,n90);
nand (n102,n103,n109);
not (n103,n104);
nor (n104,n105,n107);
and (n105,n86,n106);
and (n107,n81,n108);
not (n108,n106);
not (n109,n88);
nor (n110,n111,n117);
nand (n111,n81,n112);
not (n112,n113);
wire s0n113,s1n113,notn113;
or (n113,s0n113,s1n113);
not(notn113,n3);
and (s0n113,notn113,1'b0);
and (s1n113,n3,n115);
and (n115,n116,n83);
nor (n117,n118,n120);
and (n118,n113,n119);
not (n119,n13);
and (n120,n112,n13);
nand (n121,n122,n137);
or (n122,n123,n132);
nand (n123,n124,n129);
not (n124,n125);
nand (n125,n126,n128);
or (n126,n127,n54);
not (n127,n61);
nand (n128,n54,n127);
nand (n129,n130,n131);
or (n130,n127,n94);
nand (n131,n94,n127);
nor (n132,n133,n135);
and (n133,n98,n134);
and (n135,n94,n136);
not (n136,n134);
or (n137,n124,n138);
nor (n138,n139,n141);
and (n139,n98,n140);
and (n141,n94,n142);
not (n142,n140);
xor (n143,n144,n200);
xor (n144,n145,n187);
xor (n145,n146,n163);
nand (n146,n147,n156);
or (n147,n148,n151);
not (n148,n149);
nor (n149,n150,n14);
not (n150,n19);
nor (n151,n152,n154);
and (n152,n150,n153);
and (n154,n19,n155);
not (n155,n153);
or (n156,n157,n162);
nor (n157,n158,n160);
and (n158,n150,n159);
and (n160,n19,n161);
not (n161,n159);
not (n162,n14);
nand (n163,n164,n181);
or (n164,n165,n175);
not (n165,n166);
and (n166,n167,n171);
nand (n167,n168,n170);
or (n168,n169,n54);
not (n169,n41);
nand (n170,n54,n169);
not (n171,n172);
nand (n172,n173,n174);
or (n173,n169,n19);
nand (n174,n19,n169);
nor (n175,n176,n179);
and (n176,n177,n178);
not (n177,n54);
and (n179,n54,n180);
not (n180,n178);
or (n181,n182,n171);
nor (n182,n183,n185);
and (n183,n177,n184);
and (n185,n54,n186);
not (n186,n184);
and (n187,n188,n194);
nand (n188,n189,n193);
or (n189,n148,n190);
nor (n190,n191,n192);
and (n191,n150,n184);
and (n192,n19,n186);
or (n193,n151,n162);
nand (n194,n195,n199);
or (n195,n165,n196);
nor (n196,n197,n198);
and (n197,n177,n140);
and (n198,n54,n142);
or (n199,n171,n175);
or (n200,n201,n221);
and (n201,n202,n215);
xor (n202,n203,n210);
nand (n203,n204,n209);
or (n204,n205,n87);
not (n205,n206);
nor (n206,n207,n208);
and (n207,n13,n81);
and (n208,n119,n86);
nand (n209,n109,n78);
nor (n210,n111,n211);
nor (n211,n212,n214);
and (n212,n113,n213);
not (n213,n18);
and (n214,n112,n18);
nand (n215,n216,n220);
or (n216,n123,n217);
nor (n217,n218,n219);
and (n218,n98,n106);
and (n219,n94,n108);
or (n220,n124,n132);
and (n221,n203,n210);
or (n222,n223,n261);
and (n223,n224,n239);
xor (n224,n225,n226);
xor (n225,n188,n194);
and (n226,n227,n233);
nand (n227,n228,n232);
or (n228,n148,n229);
nor (n229,n230,n231);
and (n230,n150,n178);
and (n231,n19,n180);
or (n232,n190,n162);
nand (n233,n234,n238);
or (n234,n165,n235);
nor (n235,n236,n237);
and (n236,n177,n134);
and (n237,n54,n136);
or (n238,n196,n171);
or (n239,n240,n260);
and (n240,n241,n254);
xor (n241,n242,n249);
nand (n242,n243,n248);
or (n243,n244,n87);
not (n244,n245);
nor (n245,n246,n247);
and (n246,n18,n81);
and (n247,n213,n86);
nand (n248,n109,n206);
nor (n249,n111,n250);
nor (n250,n251,n253);
and (n251,n113,n252);
not (n252,n26);
and (n253,n112,n26);
nand (n254,n255,n259);
or (n255,n123,n256);
nor (n256,n257,n258);
and (n257,n98,n80);
and (n258,n94,n85);
or (n259,n124,n217);
and (n260,n242,n249);
and (n261,n225,n226);
not (n262,n263);
or (n263,n264,n291);
and (n264,n265,n268);
xor (n265,n266,n267);
xor (n266,n202,n215);
xor (n267,n224,n239);
and (n268,n269,n270);
xor (n269,n227,n233);
or (n270,n271,n290);
and (n271,n272,n284);
xor (n272,n273,n279);
nand (n273,n274,n278);
or (n274,n275,n87);
nor (n275,n276,n277);
and (n276,n26,n86);
and (n277,n252,n81);
nand (n278,n245,n109);
nor (n279,n111,n280);
nor (n280,n281,n283);
and (n281,n113,n282);
not (n282,n33);
and (n283,n112,n33);
nand (n284,n285,n289);
or (n285,n148,n286);
nor (n286,n287,n288);
and (n287,n150,n140);
and (n288,n19,n142);
or (n289,n229,n162);
and (n290,n273,n279);
and (n291,n266,n267);
nand (n292,n71,n263);
not (n293,n294);
nand (n294,n295,n447,n587);
nand (n295,n296,n440);
nand (n296,n297,n439);
or (n297,n298,n428);
nor (n298,n299,n427);
and (n299,n300,n399);
not (n300,n301);
nor (n301,n302,n382);
or (n302,n303,n381);
and (n303,n304,n352);
xor (n304,n305,n339);
or (n305,n306,n338);
and (n306,n307,n329);
xor (n307,n308,n319);
nand (n308,n309,n315);
or (n309,n310,n87);
not (n310,n311);
nand (n311,n312,n313);
or (n312,n86,n39);
or (n313,n81,n314);
not (n314,n39);
or (n315,n88,n316);
nor (n316,n317,n318);
and (n317,n33,n86);
and (n318,n282,n81);
nand (n319,n320,n325);
or (n320,n321,n165);
not (n321,n322);
nand (n322,n323,n324);
or (n323,n54,n119);
or (n324,n177,n13);
nand (n325,n172,n326);
nor (n326,n327,n328);
and (n327,n80,n54);
and (n328,n85,n177);
nand (n329,n330,n334);
or (n330,n123,n331);
nor (n331,n332,n333);
and (n332,n98,n26);
and (n333,n94,n252);
or (n334,n124,n335);
nor (n335,n336,n337);
and (n336,n98,n18);
and (n337,n94,n213);
and (n338,n308,n319);
xor (n339,n340,n349);
xor (n340,n341,n343);
and (n341,n342,n39);
not (n342,n111);
nand (n343,n344,n348);
or (n344,n148,n345);
nor (n345,n346,n347);
and (n346,n136,n19);
and (n347,n134,n150);
or (n348,n286,n162);
nand (n349,n350,n351);
or (n350,n87,n316);
or (n351,n88,n275);
xor (n352,n353,n367);
xor (n353,n354,n361);
nand (n354,n355,n357);
or (n355,n165,n356);
not (n356,n326);
or (n357,n171,n358);
nor (n358,n359,n360);
and (n359,n177,n106);
and (n360,n54,n108);
nand (n361,n362,n363);
or (n362,n123,n335);
or (n363,n124,n364);
nor (n364,n365,n366);
and (n365,n98,n13);
and (n366,n94,n119);
and (n367,n368,n373);
nor (n368,n369,n86);
nor (n369,n370,n372);
and (n370,n98,n371);
nand (n371,n91,n39);
and (n372,n90,n314);
nand (n373,n374,n379);
or (n374,n375,n148);
not (n375,n376);
nor (n376,n377,n378);
and (n377,n106,n19);
and (n378,n108,n150);
nand (n379,n380,n14);
not (n380,n345);
and (n381,n305,n339);
xor (n382,n383,n388);
xor (n383,n384,n385);
xor (n384,n272,n284);
or (n385,n386,n387);
and (n386,n353,n367);
and (n387,n354,n361);
xor (n388,n389,n396);
xor (n389,n390,n393);
nand (n390,n391,n392);
or (n391,n123,n364);
or (n392,n124,n256);
nand (n393,n394,n395);
or (n394,n165,n358);
or (n395,n235,n171);
or (n396,n397,n398);
and (n397,n340,n349);
and (n398,n341,n343);
not (n399,n400);
nand (n400,n401,n402);
xor (n401,n304,n352);
or (n402,n403,n426);
and (n403,n404,n425);
xor (n404,n405,n406);
xor (n405,n368,n373);
or (n406,n407,n424);
and (n407,n408,n417);
xor (n408,n409,n410);
and (n409,n109,n39);
nand (n410,n411,n412);
or (n411,n162,n375);
nand (n412,n413,n149);
not (n413,n414);
nor (n414,n415,n416);
and (n415,n80,n150);
and (n416,n85,n19);
nand (n417,n418,n423);
or (n418,n419,n165);
not (n419,n420);
nor (n420,n421,n422);
and (n421,n18,n54);
and (n422,n177,n213);
nand (n423,n172,n322);
and (n424,n409,n410);
xor (n425,n307,n329);
and (n426,n405,n406);
and (n427,n302,n382);
nor (n428,n429,n436);
xor (n429,n430,n433);
xor (n430,n431,n432);
xor (n431,n241,n254);
xor (n432,n269,n270);
or (n433,n434,n435);
and (n434,n389,n396);
and (n435,n390,n393);
or (n436,n437,n438);
and (n437,n383,n388);
and (n438,n384,n385);
nand (n439,n429,n436);
nand (n440,n441,n443);
not (n441,n442);
xor (n442,n265,n268);
not (n443,n444);
or (n444,n445,n446);
and (n445,n430,n433);
and (n446,n431,n432);
nand (n447,n440,n448,n586);
nor (n448,n449,n583);
nor (n449,n450,n581);
and (n450,n451,n576);
or (n451,n452,n575);
and (n452,n453,n494);
xor (n453,n454,n487);
or (n454,n455,n486);
and (n455,n456,n475);
xor (n456,n457,n464);
nand (n457,n458,n463);
or (n458,n459,n165);
not (n459,n460);
nor (n460,n461,n462);
and (n461,n252,n177);
and (n462,n26,n54);
nand (n463,n172,n420);
nand (n464,n465,n470);
or (n465,n466,n124);
not (n466,n467);
nor (n467,n468,n469);
and (n468,n33,n94);
and (n469,n282,n98);
nand (n470,n471,n472);
not (n471,n123);
nand (n472,n473,n474);
or (n473,n98,n39);
or (n474,n94,n314);
xor (n475,n476,n480);
and (n476,n477,n94);
nand (n477,n478,n479);
or (n478,n54,n60);
or (n479,n61,n39);
nand (n480,n481,n485);
or (n481,n148,n482);
nor (n482,n483,n484);
and (n483,n150,n13);
and (n484,n19,n119);
or (n485,n414,n162);
and (n486,n457,n464);
xor (n487,n488,n493);
xor (n488,n489,n492);
nand (n489,n490,n491);
or (n490,n466,n123);
or (n491,n124,n331);
and (n492,n476,n480);
xor (n493,n408,n417);
or (n494,n495,n574);
and (n495,n496,n515);
xor (n496,n497,n514);
or (n497,n498,n513);
and (n498,n499,n507);
xor (n499,n500,n501);
and (n500,n125,n39);
nand (n501,n502,n506);
or (n502,n503,n165);
not (n503,n504);
nor (n504,n53,n505);
and (n505,n282,n177);
nand (n506,n460,n172);
nand (n507,n508,n512);
or (n508,n148,n509);
not (n509,n510);
nor (n510,n511,n17);
and (n511,n213,n150);
or (n512,n482,n162);
and (n513,n500,n501);
xor (n514,n456,n475);
or (n515,n516,n573);
and (n516,n517,n572);
xor (n517,n518,n531);
nor (n518,n519,n527);
not (n519,n520);
nand (n520,n521,n526);
or (n521,n522,n148);
not (n522,n523);
nand (n523,n524,n525);
or (n524,n252,n19);
nand (n525,n19,n252);
nand (n526,n510,n14);
nand (n527,n528,n54);
nand (n528,n529,n530);
or (n529,n19,n52);
or (n530,n41,n39);
nand (n531,n532,n570);
or (n532,n533,n556);
not (n533,n534);
nand (n534,n535,n555);
or (n535,n536,n545);
nor (n536,n537,n544);
nand (n537,n538,n543);
or (n538,n539,n148);
not (n539,n540);
nand (n540,n541,n542);
or (n541,n282,n19);
nand (n542,n19,n282);
nand (n543,n523,n14);
nor (n544,n171,n314);
nand (n545,n546,n553);
nand (n546,n547,n552);
or (n547,n548,n148);
not (n548,n549);
nand (n549,n550,n551);
or (n550,n150,n39);
or (n551,n19,n314);
nand (n552,n540,n14);
nor (n553,n554,n150);
and (n554,n39,n14);
nand (n555,n537,n544);
not (n556,n557);
nand (n557,n558,n566);
not (n558,n559);
nand (n559,n560,n565);
or (n560,n561,n165);
not (n561,n562);
nand (n562,n563,n564);
or (n563,n177,n39);
or (n564,n54,n314);
nand (n565,n172,n504);
nor (n566,n567,n569);
and (n567,n519,n568);
not (n568,n527);
and (n569,n520,n527);
nand (n570,n571,n559);
not (n571,n566);
xor (n572,n499,n507);
and (n573,n518,n531);
and (n574,n497,n514);
and (n575,n454,n487);
or (n576,n577,n578);
xor (n577,n404,n425);
or (n578,n579,n580);
and (n579,n488,n493);
and (n580,n489,n492);
not (n581,n582);
nand (n582,n577,n578);
nand (n583,n584,n300);
not (n584,n585);
nor (n585,n401,n402);
not (n586,n428);
nand (n587,n442,n444);
or (n588,n294,n68);
wire s0n589,s1n589,notn589;
or (n589,s0n589,s1n589);
not(notn589,n3);
and (s0n589,notn589,n590);
and (s1n589,n3,n5);
xor (n590,n591,n911);
xor (n591,n592,n931);
xor (n592,n593,n906);
xor (n593,n594,n924);
xor (n594,n595,n900);
xor (n595,n596,n912);
xor (n596,n597,n894);
xor (n597,n598,n891);
xor (n598,n599,n890);
xor (n599,n600,n865);
xor (n600,n601,n79);
xor (n601,n602,n832);
xor (n602,n603,n831);
xor (n603,n604,n793);
xor (n604,n605,n792);
xor (n605,n606,n749);
xor (n606,n607,n748);
xor (n607,n608,n706);
xor (n608,n609,n705);
xor (n609,n610,n660);
xor (n610,n611,n659);
xor (n611,n612,n615);
xor (n612,n613,n614);
and (n613,n159,n14);
and (n614,n153,n19);
or (n615,n616,n619);
and (n616,n617,n618);
and (n617,n153,n14);
and (n618,n184,n19);
and (n619,n620,n621);
xor (n620,n617,n618);
or (n621,n622,n625);
and (n622,n623,n624);
and (n623,n184,n14);
and (n624,n178,n19);
and (n625,n626,n627);
xor (n626,n623,n624);
or (n627,n628,n631);
and (n628,n629,n630);
and (n629,n178,n14);
and (n630,n140,n19);
and (n631,n632,n633);
xor (n632,n629,n630);
or (n633,n634,n637);
and (n634,n635,n636);
and (n635,n140,n14);
and (n636,n134,n19);
and (n637,n638,n639);
xor (n638,n635,n636);
or (n639,n640,n642);
and (n640,n641,n377);
and (n641,n134,n14);
and (n642,n643,n644);
xor (n643,n641,n377);
or (n644,n645,n648);
and (n645,n646,n647);
and (n646,n106,n14);
and (n647,n80,n19);
and (n648,n649,n650);
xor (n649,n646,n647);
or (n650,n651,n654);
and (n651,n652,n653);
and (n652,n80,n14);
and (n653,n13,n19);
and (n654,n655,n656);
xor (n655,n652,n653);
or (n656,n657,n658);
and (n657,n12,n17);
and (n658,n11,n22);
and (n659,n184,n41);
or (n660,n661,n664);
and (n661,n662,n663);
xor (n662,n620,n621);
and (n663,n178,n41);
and (n664,n665,n666);
xor (n665,n662,n663);
or (n666,n667,n670);
and (n667,n668,n669);
xor (n668,n626,n627);
and (n669,n140,n41);
and (n670,n671,n672);
xor (n671,n668,n669);
or (n672,n673,n676);
and (n673,n674,n675);
xor (n674,n632,n633);
and (n675,n134,n41);
and (n676,n677,n678);
xor (n677,n674,n675);
or (n678,n679,n682);
and (n679,n680,n681);
xor (n680,n638,n639);
and (n681,n106,n41);
and (n682,n683,n684);
xor (n683,n680,n681);
or (n684,n685,n688);
and (n685,n686,n687);
xor (n686,n643,n644);
and (n687,n80,n41);
and (n688,n689,n690);
xor (n689,n686,n687);
or (n690,n691,n694);
and (n691,n692,n693);
xor (n692,n649,n650);
and (n693,n13,n41);
and (n694,n695,n696);
xor (n695,n692,n693);
or (n696,n697,n700);
and (n697,n698,n699);
xor (n698,n655,n656);
and (n699,n18,n41);
and (n700,n701,n702);
xor (n701,n698,n699);
or (n702,n703,n704);
and (n703,n10,n40);
and (n704,n9,n44);
and (n705,n178,n54);
or (n706,n707,n710);
and (n707,n708,n709);
xor (n708,n665,n666);
and (n709,n140,n54);
and (n710,n711,n712);
xor (n711,n708,n709);
or (n712,n713,n716);
and (n713,n714,n715);
xor (n714,n671,n672);
and (n715,n134,n54);
and (n716,n717,n718);
xor (n717,n714,n715);
or (n718,n719,n722);
and (n719,n720,n721);
xor (n720,n677,n678);
and (n721,n106,n54);
and (n722,n723,n724);
xor (n723,n720,n721);
or (n724,n725,n727);
and (n725,n726,n327);
xor (n726,n683,n684);
and (n727,n728,n729);
xor (n728,n726,n327);
or (n729,n730,n733);
and (n730,n731,n732);
xor (n731,n689,n690);
and (n732,n13,n54);
and (n733,n734,n735);
xor (n734,n731,n732);
or (n735,n736,n738);
and (n736,n737,n421);
xor (n737,n695,n696);
and (n738,n739,n740);
xor (n739,n737,n421);
or (n740,n741,n743);
and (n741,n742,n462);
xor (n742,n701,n702);
and (n743,n744,n745);
xor (n744,n742,n462);
or (n745,n746,n747);
and (n746,n8,n53);
and (n747,n7,n57);
and (n748,n140,n61);
or (n749,n750,n753);
and (n750,n751,n752);
xor (n751,n711,n712);
and (n752,n134,n61);
and (n753,n754,n755);
xor (n754,n751,n752);
or (n755,n756,n759);
and (n756,n757,n758);
xor (n757,n717,n718);
and (n758,n106,n61);
and (n759,n760,n761);
xor (n760,n757,n758);
or (n761,n762,n765);
and (n762,n763,n764);
xor (n763,n723,n724);
and (n764,n80,n61);
and (n765,n766,n767);
xor (n766,n763,n764);
or (n767,n768,n771);
and (n768,n769,n770);
xor (n769,n728,n729);
and (n770,n13,n61);
and (n771,n772,n773);
xor (n772,n769,n770);
or (n773,n774,n777);
and (n774,n775,n776);
xor (n775,n734,n735);
and (n776,n18,n61);
and (n777,n778,n779);
xor (n778,n775,n776);
or (n779,n780,n783);
and (n780,n781,n782);
xor (n781,n739,n740);
and (n782,n26,n61);
and (n783,n784,n785);
xor (n784,n781,n782);
or (n785,n786,n789);
and (n786,n787,n788);
xor (n787,n744,n745);
and (n788,n33,n61);
and (n789,n790,n791);
xor (n790,n787,n788);
and (n791,n6,n60);
and (n792,n134,n94);
or (n793,n794,n797);
and (n794,n795,n796);
xor (n795,n754,n755);
and (n796,n106,n94);
and (n797,n798,n799);
xor (n798,n795,n796);
or (n799,n800,n803);
and (n800,n801,n802);
xor (n801,n760,n761);
and (n802,n80,n94);
and (n803,n804,n805);
xor (n804,n801,n802);
or (n805,n806,n809);
and (n806,n807,n808);
xor (n807,n766,n767);
and (n808,n13,n94);
and (n809,n810,n811);
xor (n810,n807,n808);
or (n811,n812,n815);
and (n812,n813,n814);
xor (n813,n772,n773);
and (n814,n18,n94);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n821);
and (n818,n819,n820);
xor (n819,n778,n779);
and (n820,n26,n94);
and (n821,n822,n823);
xor (n822,n819,n820);
or (n823,n824,n826);
and (n824,n825,n468);
xor (n825,n784,n785);
and (n826,n827,n828);
xor (n827,n825,n468);
and (n828,n829,n830);
xor (n829,n790,n791);
and (n830,n39,n94);
and (n831,n106,n91);
or (n832,n833,n836);
and (n833,n834,n835);
xor (n834,n798,n799);
and (n835,n80,n91);
and (n836,n837,n838);
xor (n837,n834,n835);
or (n838,n839,n842);
and (n839,n840,n841);
xor (n840,n804,n805);
and (n841,n13,n91);
and (n842,n843,n844);
xor (n843,n840,n841);
or (n844,n845,n848);
and (n845,n846,n847);
xor (n846,n810,n811);
and (n847,n18,n91);
and (n848,n849,n850);
xor (n849,n846,n847);
or (n850,n851,n854);
and (n851,n852,n853);
xor (n852,n816,n817);
and (n853,n26,n91);
and (n854,n855,n856);
xor (n855,n852,n853);
or (n856,n857,n860);
and (n857,n858,n859);
xor (n858,n822,n823);
and (n859,n33,n91);
and (n860,n861,n862);
xor (n861,n858,n859);
and (n862,n863,n864);
xor (n863,n827,n828);
not (n864,n371);
or (n865,n866,n868);
and (n866,n867,n207);
xor (n867,n837,n838);
and (n868,n869,n870);
xor (n869,n867,n207);
or (n870,n871,n873);
and (n871,n872,n246);
xor (n872,n843,n844);
and (n873,n874,n875);
xor (n874,n872,n246);
or (n875,n876,n879);
and (n876,n877,n878);
xor (n877,n849,n850);
and (n878,n26,n81);
and (n879,n880,n881);
xor (n880,n877,n878);
or (n881,n882,n885);
and (n882,n883,n884);
xor (n883,n855,n856);
and (n884,n33,n81);
and (n885,n886,n887);
xor (n886,n883,n884);
and (n887,n888,n889);
xor (n888,n861,n862);
and (n889,n39,n81);
and (n890,n13,n113);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n869,n870);
and (n894,n18,n113);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n874,n875);
and (n900,n26,n113);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n880,n881);
and (n906,n33,n113);
and (n907,n908,n909);
xor (n908,n905,n906);
and (n909,n910,n911);
xor (n910,n886,n887);
and (n911,n39,n113);
or (n912,n913,n915);
and (n913,n914,n900);
xor (n914,n896,n897);
and (n915,n916,n917);
xor (n916,n914,n900);
or (n917,n918,n920);
and (n918,n919,n906);
xor (n919,n902,n903);
and (n920,n921,n922);
xor (n921,n919,n906);
and (n922,n923,n911);
xor (n923,n908,n909);
or (n924,n925,n927);
and (n925,n926,n906);
xor (n926,n916,n917);
and (n927,n928,n929);
xor (n928,n926,n906);
and (n929,n930,n911);
xor (n930,n921,n922);
and (n931,n932,n911);
xor (n932,n928,n929);
endmodule
