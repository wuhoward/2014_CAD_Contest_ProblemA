module top (out,n20,n21,n28,n29,n40,n47,n49,n56,n57
        ,n67,n75,n80,n86,n92,n102,n104,n110,n119,n124
        ,n134,n145,n154,n159,n189,n194,n221,n280,n301,n302
        ,n332,n431,n500,n560,n645,n1617,n1618,n1621);
output out;
input n20;
input n21;
input n28;
input n29;
input n40;
input n47;
input n49;
input n56;
input n57;
input n67;
input n75;
input n80;
input n86;
input n92;
input n102;
input n104;
input n110;
input n119;
input n124;
input n134;
input n145;
input n154;
input n159;
input n189;
input n194;
input n221;
input n280;
input n301;
input n302;
input n332;
input n431;
input n500;
input n560;
input n645;
input n1617;
input n1618;
input n1621;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1619;
wire n1620;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
xor (out,n0,n1622);
nand (n0,n1,n1619);
or (n1,n2,n1615);
not (n2,n3);
nor (n3,n4,n1612);
and (n4,n5,n447);
nor (n5,n6,n446);
and (n6,n7,n382);
xor (n7,n8,n286);
xor (n8,n9,n182);
xor (n9,n10,n163);
xor (n10,n11,n95);
or (n11,n12,n94);
and (n12,n13,n69);
xor (n13,n14,n42);
nand (n14,n15,n35);
or (n15,n16,n24);
not (n16,n17);
nand (n17,n18,n22);
or (n18,n19,n21);
not (n19,n20);
or (n22,n20,n23);
not (n23,n21);
nand (n24,n25,n32);
nor (n25,n26,n30);
and (n26,n27,n29);
not (n27,n28);
and (n30,n28,n31);
not (n31,n29);
nor (n32,n33,n34);
and (n33,n27,n23);
and (n34,n28,n21);
nand (n35,n36,n37);
not (n36,n25);
nor (n37,n38,n41);
and (n38,n23,n39);
not (n39,n40);
and (n41,n40,n21);
nand (n42,n43,n63);
or (n43,n44,n51);
not (n44,n45);
nand (n45,n46,n50);
or (n46,n47,n48);
not (n48,n49);
nand (n50,n48,n47);
not (n51,n52);
nor (n52,n53,n59);
nand (n53,n54,n58);
or (n54,n55,n57);
not (n55,n56);
nand (n58,n55,n57);
nor (n59,n60,n61);
and (n60,n48,n57);
and (n61,n49,n62);
not (n62,n57);
nand (n63,n53,n64);
nor (n64,n65,n68);
and (n65,n66,n48);
not (n66,n67);
and (n68,n67,n49);
nand (n69,n70,n88);
or (n70,n71,n82);
nand (n71,n72,n77);
not (n72,n73);
nand (n73,n74,n76);
or (n74,n23,n75);
nand (n76,n75,n23);
nand (n77,n78,n81);
or (n78,n75,n79);
not (n79,n80);
nand (n81,n79,n75);
not (n82,n83);
nor (n83,n84,n87);
and (n84,n85,n79);
not (n85,n86);
and (n87,n86,n80);
or (n88,n72,n89);
nor (n89,n90,n93);
and (n90,n91,n80);
not (n91,n92);
and (n93,n92,n79);
and (n94,n14,n42);
or (n95,n96,n162);
and (n96,n97,n137);
xor (n97,n98,n113);
nand (n98,n99,n110);
or (n99,n100,n106);
nand (n100,n101,n105);
or (n101,n102,n103);
not (n103,n104);
nand (n105,n102,n103);
nor (n106,n100,n107);
nor (n107,n108,n111);
and (n108,n109,n110);
not (n109,n102);
and (n111,n102,n112);
not (n112,n110);
nand (n113,n114,n130);
or (n114,n115,n121);
not (n115,n116);
nor (n116,n117,n120);
and (n117,n118,n55);
not (n118,n119);
and (n120,n119,n56);
nand (n121,n122,n126);
nand (n122,n123,n125);
or (n123,n124,n55);
nand (n125,n55,n124);
not (n126,n127);
nand (n127,n128,n129);
or (n128,n112,n124);
nand (n129,n124,n112);
nand (n130,n131,n127);
not (n131,n132);
nor (n132,n133,n135);
and (n133,n55,n134);
and (n135,n56,n136);
not (n136,n134);
nand (n137,n138,n156);
or (n138,n139,n150);
not (n139,n140);
and (n140,n141,n147);
not (n141,n142);
nand (n142,n143,n146);
or (n143,n144,n49);
not (n144,n145);
nand (n146,n49,n144);
nand (n147,n148,n149);
nand (n148,n29,n144);
nand (n149,n145,n31);
not (n150,n151);
nor (n151,n152,n155);
and (n152,n153,n31);
not (n153,n154);
and (n155,n154,n29);
or (n156,n141,n157);
nor (n157,n158,n160);
and (n158,n31,n159);
and (n160,n29,n161);
not (n161,n159);
and (n162,n98,n113);
xor (n163,n164,n179);
xor (n164,n165,n172);
nand (n165,n166,n168);
or (n166,n24,n167);
not (n167,n37);
or (n168,n169,n25);
nor (n169,n170,n171);
and (n170,n154,n23);
and (n171,n21,n153);
nand (n172,n173,n178);
or (n173,n174,n72);
not (n174,n175);
nor (n175,n176,n177);
and (n176,n20,n80);
and (n177,n19,n79);
or (n178,n71,n89);
nand (n179,n180,n181);
or (n180,n121,n132);
or (n181,n126,n55);
xor (n182,n183,n257);
xor (n183,n184,n215);
xor (n184,n185,n206);
xor (n185,n186,n198);
nand (n186,n187,n197);
or (n187,n188,n190);
not (n188,n189);
not (n190,n191);
nor (n191,n192,n196);
nand (n192,n193,n195);
or (n193,n79,n194);
nand (n195,n194,n79);
not (n196,n194);
nand (n197,n192,n86);
nand (n198,n199,n200);
or (n199,n139,n157);
or (n200,n141,n201);
not (n201,n202);
nor (n202,n203,n205);
and (n203,n204,n31);
not (n204,n47);
and (n205,n47,n29);
not (n206,n207);
nand (n207,n208,n210);
or (n208,n209,n51);
not (n209,n64);
nand (n210,n211,n53);
not (n211,n212);
nor (n212,n213,n214);
and (n213,n118,n49);
and (n214,n119,n48);
or (n215,n216,n256);
and (n216,n217,n231);
xor (n217,n218,n224);
nand (n218,n219,n222);
or (n219,n220,n190);
not (n220,n221);
or (n222,n223,n188);
not (n223,n192);
not (n224,n225);
nor (n225,n226,n230);
and (n226,n106,n227);
nor (n227,n228,n229);
and (n228,n136,n112);
and (n229,n134,n110);
and (n230,n100,n110);
or (n231,n232,n255);
and (n232,n233,n248);
xor (n233,n234,n241);
nand (n234,n235,n240);
or (n235,n236,n121);
not (n236,n237);
nor (n237,n238,n239);
and (n238,n66,n55);
and (n239,n67,n56);
nand (n240,n127,n116);
nand (n241,n242,n247);
or (n242,n243,n139);
not (n243,n244);
nor (n244,n245,n246);
and (n245,n39,n31);
and (n246,n40,n29);
nand (n247,n142,n151);
nand (n248,n249,n250);
or (n249,n16,n25);
nand (n250,n251,n252);
not (n251,n24);
nor (n252,n253,n254);
and (n253,n91,n23);
and (n254,n92,n21);
and (n255,n234,n241);
and (n256,n218,n224);
or (n257,n258,n285);
and (n258,n259,n284);
xor (n259,n260,n283);
or (n260,n261,n282);
and (n261,n262,n277);
xor (n262,n263,n270);
nand (n263,n264,n269);
or (n264,n265,n51);
not (n265,n266);
nor (n266,n267,n268);
and (n267,n161,n48);
and (n268,n159,n49);
nand (n269,n53,n45);
nand (n270,n271,n276);
or (n271,n272,n71);
not (n272,n273);
nor (n273,n274,n275);
and (n274,n188,n79);
and (n275,n189,n80);
nand (n276,n73,n83);
nand (n277,n278,n281);
or (n278,n279,n190);
not (n279,n280);
nand (n281,n192,n221);
and (n282,n263,n270);
xor (n283,n13,n69);
xor (n284,n97,n137);
and (n285,n260,n283);
or (n286,n287,n381);
and (n287,n288,n350);
xor (n288,n289,n290);
xor (n289,n217,n231);
or (n290,n291,n349);
and (n291,n292,n326);
xor (n292,n225,n293);
or (n293,n294,n325);
and (n294,n295,n318);
xor (n295,n296,n310);
nand (n296,n297,n104);
or (n297,n298,n304);
nand (n298,n299,n303);
or (n299,n300,n302);
not (n300,n301);
nand (n303,n302,n300);
not (n304,n305);
nand (n305,n306,n307);
not (n306,n298);
nand (n307,n308,n309);
or (n308,n300,n104);
nand (n309,n300,n104);
nand (n310,n311,n317);
or (n311,n312,n316);
not (n312,n313);
nand (n313,n314,n315);
or (n314,n119,n112);
nand (n315,n112,n119);
not (n316,n106);
nand (n317,n227,n100);
nand (n318,n319,n324);
or (n319,n320,n51);
not (n320,n321);
nor (n321,n322,n323);
and (n322,n153,n48);
and (n323,n154,n49);
nand (n324,n53,n266);
and (n325,n296,n310);
or (n326,n327,n348);
and (n327,n328,n341);
xor (n328,n329,n334);
nand (n329,n330,n333);
or (n330,n331,n190);
not (n331,n332);
nand (n333,n192,n280);
nand (n334,n335,n340);
or (n335,n336,n139);
not (n336,n337);
nor (n337,n338,n339);
and (n338,n19,n31);
and (n339,n20,n29);
nand (n340,n142,n244);
nand (n341,n342,n343);
or (n342,n236,n126);
or (n343,n121,n344);
not (n344,n345);
nor (n345,n346,n347);
and (n346,n204,n55);
and (n347,n47,n56);
and (n348,n329,n334);
and (n349,n225,n293);
or (n350,n351,n380);
and (n351,n352,n355);
xor (n352,n353,n354);
xor (n353,n262,n277);
xor (n354,n233,n248);
or (n355,n356,n379);
and (n356,n357,n372);
xor (n357,n358,n365);
nand (n358,n359,n364);
or (n359,n360,n24);
not (n360,n361);
nor (n361,n362,n363);
and (n362,n23,n85);
and (n363,n86,n21);
nand (n364,n36,n252);
nand (n365,n366,n371);
or (n366,n367,n71);
not (n367,n368);
nor (n368,n369,n370);
and (n369,n220,n79);
and (n370,n221,n80);
nand (n371,n73,n273);
not (n372,n373);
nor (n373,n374,n378);
and (n374,n304,n375);
nor (n375,n376,n377);
and (n376,n136,n103);
and (n377,n134,n104);
nor (n378,n306,n103);
and (n379,n358,n365);
and (n380,n353,n354);
and (n381,n289,n290);
or (n382,n383,n445);
and (n383,n384,n387);
xor (n384,n385,n386);
xor (n385,n259,n284);
xor (n386,n288,n350);
or (n387,n388,n444);
and (n388,n389,n443);
xor (n389,n390,n391);
xor (n390,n292,n326);
or (n391,n392,n442);
and (n392,n393,n441);
xor (n393,n394,n418);
or (n394,n395,n417);
and (n395,n396,n411);
xor (n396,n397,n404);
nand (n397,n398,n403);
or (n398,n399,n139);
not (n399,n400);
nand (n400,n401,n402);
or (n401,n92,n31);
nand (n402,n31,n92);
nand (n403,n337,n142);
nand (n404,n405,n410);
or (n405,n406,n121);
not (n406,n407);
nor (n407,n408,n409);
and (n408,n161,n55);
and (n409,n159,n56);
nand (n410,n127,n345);
nand (n411,n412,n413);
or (n412,n25,n360);
or (n413,n24,n414);
nor (n414,n415,n416);
and (n415,n189,n23);
and (n416,n21,n188);
and (n417,n397,n404);
or (n418,n419,n440);
and (n419,n420,n433);
xor (n420,n421,n428);
nand (n421,n422,n427);
or (n422,n423,n316);
not (n423,n424);
nor (n424,n425,n426);
and (n425,n66,n112);
and (n426,n67,n110);
nand (n427,n100,n313);
nand (n428,n429,n432);
or (n429,n430,n190);
not (n430,n431);
nand (n432,n192,n332);
nand (n433,n434,n439);
or (n434,n435,n51);
not (n435,n436);
nor (n436,n437,n438);
and (n437,n39,n48);
and (n438,n40,n49);
nand (n439,n53,n321);
and (n440,n421,n428);
xor (n441,n295,n318);
and (n442,n394,n418);
xor (n443,n352,n355);
and (n444,n390,n391);
and (n445,n385,n386);
nor (n446,n7,n382);
nand (n447,n448,n1611);
or (n448,n449,n572);
nor (n449,n450,n451);
xor (n450,n384,n387);
or (n451,n452,n571);
and (n452,n453,n480);
xor (n453,n454,n479);
or (n454,n455,n478);
and (n455,n456,n459);
xor (n456,n457,n458);
xor (n457,n328,n341);
xor (n458,n357,n372);
or (n459,n460,n477);
and (n460,n461,n469);
xor (n461,n462,n373);
nand (n462,n463,n468);
or (n463,n464,n71);
not (n464,n465);
nor (n465,n466,n467);
and (n466,n279,n79);
and (n467,n280,n80);
nand (n468,n73,n368);
nand (n469,n470,n302);
nor (n470,n471,n476);
and (n471,n472,n473);
not (n472,n121);
nand (n473,n474,n475);
or (n474,n154,n55);
nand (n475,n55,n154);
and (n476,n127,n407);
and (n477,n462,n373);
and (n478,n457,n458);
xor (n479,n389,n443);
or (n480,n481,n570);
and (n481,n482,n534);
xor (n482,n483,n484);
xor (n483,n393,n441);
or (n484,n485,n533);
and (n485,n486,n532);
xor (n486,n487,n509);
or (n487,n488,n508);
and (n488,n489,n502);
xor (n489,n490,n497);
nand (n490,n491,n496);
or (n491,n492,n71);
not (n492,n493);
nand (n493,n494,n495);
or (n494,n331,n80);
nand (n495,n80,n331);
nand (n496,n465,n73);
nand (n497,n498,n501);
or (n498,n499,n190);
not (n499,n500);
nand (n501,n192,n431);
nand (n502,n503,n505);
or (n503,n504,n306);
not (n504,n375);
or (n505,n305,n506);
not (n506,n507);
xor (n507,n118,n103);
and (n508,n490,n497);
or (n509,n510,n531);
and (n510,n511,n525);
xor (n511,n512,n519);
nand (n512,n513,n518);
or (n513,n514,n51);
not (n514,n515);
nor (n515,n516,n517);
and (n516,n19,n48);
and (n517,n20,n49);
nand (n518,n53,n436);
nand (n519,n520,n524);
or (n520,n521,n316);
nor (n521,n522,n523);
and (n522,n204,n110);
and (n523,n47,n112);
nand (n524,n424,n100);
nand (n525,n526,n530);
or (n526,n139,n527);
nor (n527,n528,n529);
and (n528,n85,n29);
and (n529,n86,n31);
or (n530,n141,n399);
and (n531,n512,n519);
xor (n532,n396,n411);
and (n533,n487,n509);
or (n534,n535,n569);
and (n535,n536,n539);
xor (n536,n537,n538);
xor (n537,n420,n433);
xor (n538,n461,n469);
and (n539,n540,n563);
or (n540,n541,n562);
and (n541,n542,n557);
xor (n542,n543,n550);
nand (n543,n544,n549);
or (n544,n545,n121);
not (n545,n546);
nor (n546,n547,n548);
and (n547,n39,n55);
and (n548,n40,n56);
nand (n549,n473,n127);
nand (n550,n551,n556);
or (n551,n552,n71);
not (n552,n553);
nand (n553,n554,n555);
or (n554,n431,n79);
nand (n555,n431,n79);
nand (n556,n73,n493);
nand (n557,n558,n561);
or (n558,n559,n190);
not (n559,n560);
nand (n561,n192,n500);
and (n562,n543,n550);
nand (n563,n564,n568);
or (n564,n24,n565);
nor (n565,n566,n567);
and (n566,n23,n221);
and (n567,n21,n220);
or (n568,n25,n414);
and (n569,n537,n538);
and (n570,n483,n484);
and (n571,n454,n479);
not (n572,n573);
nand (n573,n574,n1606);
or (n574,n575,n750);
not (n575,n576);
nor (n576,n577,n657);
nor (n577,n578,n579);
xor (n578,n453,n480);
or (n579,n580,n656);
and (n580,n581,n584);
xor (n581,n582,n583);
xor (n582,n456,n459);
xor (n583,n482,n534);
or (n584,n585,n655);
and (n585,n586,n619);
xor (n586,n587,n588);
xor (n587,n486,n532);
or (n588,n589,n618);
and (n589,n590,n616);
xor (n590,n591,n615);
or (n591,n592,n614);
and (n592,n593,n608);
xor (n593,n594,n601);
nand (n594,n595,n600);
or (n595,n596,n305);
not (n596,n597);
nor (n597,n598,n599);
and (n598,n66,n103);
and (n599,n67,n104);
nand (n600,n298,n507);
nand (n601,n602,n607);
or (n602,n603,n51);
not (n603,n604);
nor (n604,n605,n606);
and (n605,n91,n48);
and (n606,n92,n49);
nand (n607,n53,n515);
nand (n608,n609,n612);
or (n609,n316,n610);
not (n610,n611);
xor (n611,n161,n112);
or (n612,n521,n613);
not (n613,n100);
and (n614,n594,n601);
xor (n615,n511,n525);
nand (n616,n617,n469);
or (n617,n302,n470);
and (n618,n591,n615);
or (n619,n620,n654);
and (n620,n621,n653);
xor (n621,n622,n623);
xor (n622,n489,n502);
or (n623,n624,n652);
and (n624,n625,n641);
xor (n625,n626,n634);
nand (n626,n627,n632);
or (n627,n628,n139);
not (n628,n629);
nand (n629,n630,n631);
or (n630,n29,n188);
or (n631,n31,n189);
nand (n632,n633,n142);
not (n633,n527);
nand (n634,n635,n640);
or (n635,n636,n24);
not (n636,n637);
nand (n637,n638,n639);
or (n638,n21,n279);
or (n639,n23,n280);
or (n640,n25,n565);
nand (n641,n642,n651);
or (n642,n643,n646);
nand (n643,n644,n302);
not (n644,n645);
not (n646,n647);
nor (n647,n648,n650);
and (n648,n136,n649);
not (n649,n302);
and (n650,n134,n302);
or (n651,n649,n644);
and (n652,n626,n634);
xor (n653,n563,n540);
and (n654,n622,n623);
and (n655,n587,n588);
and (n656,n582,n583);
nor (n657,n658,n659);
xor (n658,n581,n584);
or (n659,n660,n749);
and (n660,n661,n748);
xor (n661,n662,n663);
xor (n662,n536,n539);
or (n663,n664,n747);
and (n664,n665,n746);
xor (n665,n666,n739);
or (n666,n667,n738);
and (n667,n668,n712);
xor (n668,n669,n687);
or (n669,n670,n686);
and (n670,n671,n679);
xor (n671,n672,n673);
and (n672,n192,n560);
nand (n673,n674,n678);
or (n674,n643,n675);
nor (n675,n676,n677);
and (n676,n118,n302);
and (n677,n119,n649);
nand (n678,n647,n645);
nand (n679,n680,n685);
or (n680,n681,n305);
not (n681,n682);
nor (n682,n683,n684);
and (n683,n204,n103);
and (n684,n47,n104);
nand (n685,n298,n597);
and (n686,n672,n673);
or (n687,n688,n711);
and (n688,n689,n704);
xor (n689,n690,n697);
nand (n690,n691,n696);
or (n691,n692,n316);
not (n692,n693);
nor (n693,n694,n695);
and (n694,n153,n112);
and (n695,n154,n110);
nand (n696,n611,n100);
nand (n697,n698,n699);
or (n698,n141,n628);
nand (n699,n700,n140);
not (n700,n701);
nor (n701,n702,n703);
and (n702,n221,n31);
and (n703,n220,n29);
nand (n704,n705,n706);
or (n705,n636,n25);
nand (n706,n707,n251);
not (n707,n708);
nor (n708,n709,n710);
and (n709,n332,n23);
and (n710,n21,n331);
and (n711,n690,n697);
or (n712,n713,n737);
and (n713,n714,n729);
xor (n714,n715,n722);
nand (n715,n716,n721);
or (n716,n717,n71);
not (n717,n718);
nor (n718,n719,n720);
and (n719,n499,n79);
and (n720,n500,n80);
nand (n721,n553,n73);
nand (n722,n723,n728);
or (n723,n724,n121);
not (n724,n725);
nand (n725,n726,n727);
or (n726,n56,n19);
or (n727,n55,n20);
nand (n728,n127,n546);
nand (n729,n730,n735);
or (n730,n51,n731);
not (n731,n732);
nor (n732,n733,n734);
and (n733,n85,n48);
and (n734,n86,n49);
or (n735,n736,n603);
not (n736,n53);
and (n737,n715,n722);
and (n738,n669,n687);
or (n739,n740,n745);
and (n740,n741,n744);
xor (n741,n742,n743);
xor (n742,n542,n557);
xor (n743,n593,n608);
xor (n744,n625,n641);
and (n745,n742,n743);
xor (n746,n590,n616);
and (n747,n666,n739);
xor (n748,n586,n619);
and (n749,n662,n663);
not (n750,n751);
nand (n751,n752,n1591);
or (n752,n753,n1521);
not (n753,n754);
nand (n754,n755,n1508);
or (n755,n756,n1209);
not (n756,n757);
nand (n757,n758,n1198,n1208);
nand (n758,n759,n986,n1064);
nor (n759,n760,n924);
not (n760,n761);
or (n761,n762,n887);
xor (n762,n763,n847);
xor (n763,n764,n794);
xor (n764,n765,n785);
xor (n765,n766,n776);
nand (n766,n767,n772);
or (n767,n768,n51);
not (n768,n769);
nor (n769,n770,n771);
and (n770,n499,n48);
and (n771,n500,n49);
nand (n772,n53,n773);
nand (n773,n774,n775);
or (n774,n49,n430);
or (n775,n48,n431);
nand (n776,n777,n781);
or (n777,n778,n643);
nor (n778,n779,n780);
and (n779,n649,n20);
and (n780,n302,n19);
or (n781,n782,n644);
nor (n782,n783,n784);
and (n783,n649,n40);
and (n784,n302,n39);
nand (n785,n786,n790);
or (n786,n316,n787);
nor (n787,n788,n789);
and (n788,n112,n221);
and (n789,n110,n220);
or (n790,n791,n613);
nor (n791,n792,n793);
and (n792,n112,n189);
and (n793,n110,n188);
or (n794,n795,n846);
and (n795,n796,n821);
xor (n796,n797,n803);
nand (n797,n798,n802);
or (n798,n316,n799);
nor (n799,n800,n801);
and (n800,n112,n280);
and (n801,n110,n279);
or (n802,n613,n787);
xor (n803,n804,n810);
and (n804,n805,n49);
nand (n805,n806,n807);
or (n806,n560,n57);
nand (n807,n808,n55);
not (n808,n809);
and (n809,n560,n57);
nand (n810,n811,n816);
or (n811,n812,n306);
not (n812,n813);
nand (n813,n814,n815);
or (n814,n104,n85);
or (n815,n103,n86);
nand (n816,n817,n304);
not (n817,n818);
nor (n818,n819,n820);
and (n819,n103,n189);
and (n820,n104,n188);
or (n821,n822,n845);
and (n822,n823,n835);
xor (n823,n824,n825);
and (n824,n53,n560);
nand (n825,n826,n831);
or (n826,n644,n827);
not (n827,n828);
nor (n828,n829,n830);
and (n829,n91,n649);
and (n830,n92,n302);
or (n831,n832,n643);
nor (n832,n833,n834);
and (n833,n649,n86);
and (n834,n302,n85);
nand (n835,n836,n840);
or (n836,n121,n837);
nor (n837,n838,n839);
and (n838,n55,n500);
and (n839,n56,n499);
or (n840,n126,n841);
not (n841,n842);
nor (n842,n843,n844);
and (n843,n431,n56);
and (n844,n430,n55);
and (n845,n824,n825);
and (n846,n797,n803);
xor (n847,n848,n870);
xor (n848,n849,n850);
and (n849,n804,n810);
or (n850,n851,n869);
and (n851,n852,n866);
xor (n852,n853,n859);
nand (n853,n854,n855);
or (n854,n841,n121);
nand (n855,n127,n856);
nor (n856,n857,n858);
and (n857,n331,n55);
and (n858,n332,n56);
nand (n859,n860,n865);
or (n860,n861,n51);
not (n861,n862);
nand (n862,n863,n864);
or (n863,n48,n560);
or (n864,n559,n49);
nand (n865,n53,n769);
nand (n866,n867,n868);
or (n867,n643,n827);
or (n868,n778,n644);
and (n869,n853,n859);
xor (n870,n871,n879);
xor (n871,n872,n873);
and (n872,n142,n560);
nand (n873,n874,n875);
or (n874,n812,n305);
nand (n875,n298,n876);
nand (n876,n877,n878);
or (n877,n104,n91);
or (n878,n103,n92);
nand (n879,n880,n882);
or (n880,n881,n121);
not (n881,n856);
nand (n882,n883,n127);
not (n883,n884);
nor (n884,n885,n886);
and (n885,n55,n280);
and (n886,n56,n279);
or (n887,n888,n923);
and (n888,n889,n922);
xor (n889,n890,n891);
xor (n890,n852,n866);
or (n891,n892,n921);
and (n892,n893,n906);
xor (n893,n894,n900);
nand (n894,n895,n899);
or (n895,n305,n896);
nor (n896,n897,n898);
and (n897,n103,n221);
and (n898,n104,n220);
or (n899,n306,n818);
nand (n900,n901,n905);
or (n901,n316,n902);
nor (n902,n903,n904);
and (n903,n112,n332);
and (n904,n110,n331);
or (n905,n799,n613);
and (n906,n907,n914);
nor (n907,n908,n55);
nor (n908,n909,n912);
and (n909,n910,n112);
not (n910,n911);
and (n911,n560,n124);
and (n912,n559,n913);
not (n913,n124);
nand (n914,n915,n920);
or (n915,n916,n643);
not (n916,n917);
nor (n917,n918,n919);
and (n918,n188,n649);
and (n919,n189,n302);
or (n920,n832,n644);
and (n921,n894,n900);
xor (n922,n796,n821);
and (n923,n890,n891);
nand (n924,n925,n980);
not (n925,n926);
nor (n926,n927,n955);
xor (n927,n928,n954);
xor (n928,n929,n953);
or (n929,n930,n952);
and (n930,n931,n946);
xor (n931,n932,n940);
nand (n932,n933,n938);
or (n933,n934,n121);
not (n934,n935);
nand (n935,n936,n937);
or (n936,n55,n560);
or (n937,n56,n559);
nand (n938,n939,n127);
not (n939,n837);
nand (n940,n941,n945);
or (n941,n305,n942);
nor (n942,n943,n944);
and (n943,n103,n280);
and (n944,n104,n279);
or (n945,n896,n306);
nand (n946,n947,n951);
or (n947,n316,n948);
nor (n948,n949,n950);
and (n949,n112,n431);
and (n950,n110,n430);
or (n951,n902,n613);
and (n952,n932,n940);
xor (n953,n823,n835);
xor (n954,n893,n906);
or (n955,n956,n979);
and (n956,n957,n978);
xor (n957,n958,n959);
xor (n958,n907,n914);
or (n959,n960,n977);
and (n960,n961,n970);
xor (n961,n962,n963);
and (n962,n127,n560);
nand (n963,n964,n969);
or (n964,n643,n965);
not (n965,n966);
nor (n966,n967,n968);
and (n967,n221,n302);
and (n968,n220,n649);
nand (n969,n917,n645);
nand (n970,n971,n976);
or (n971,n305,n972);
not (n972,n973);
nor (n973,n974,n975);
and (n974,n331,n103);
and (n975,n332,n104);
or (n976,n306,n942);
and (n977,n962,n963);
xor (n978,n931,n946);
and (n979,n958,n959);
not (n980,n981);
nor (n981,n982,n983);
xor (n982,n889,n922);
or (n983,n984,n985);
and (n984,n928,n954);
and (n985,n929,n953);
nand (n986,n987,n1060);
not (n987,n988);
xor (n988,n989,n1057);
xor (n989,n990,n1027);
xor (n990,n991,n1009);
xor (n991,n992,n1003);
nand (n992,n993,n998);
or (n993,n994,n141);
not (n994,n995);
nand (n995,n996,n997);
or (n996,n29,n499);
or (n997,n31,n500);
nand (n998,n999,n140);
not (n999,n1000);
nor (n1000,n1001,n1002);
and (n1001,n559,n29);
and (n1002,n31,n560);
nand (n1003,n1004,n1005);
or (n1004,n316,n791);
or (n1005,n613,n1006);
nor (n1006,n1007,n1008);
and (n1007,n112,n86);
and (n1008,n110,n85);
nand (n1009,n1010,n1026);
or (n1010,n1011,n1018);
not (n1011,n1012);
nand (n1012,n1013,n29);
nand (n1013,n1014,n1015);
or (n1014,n560,n145);
nand (n1015,n1016,n48);
not (n1016,n1017);
and (n1017,n560,n145);
not (n1018,n1019);
nand (n1019,n1020,n1022);
or (n1020,n1021,n305);
not (n1021,n876);
nand (n1022,n298,n1023);
nor (n1023,n1024,n1025);
and (n1024,n19,n103);
and (n1025,n20,n104);
or (n1026,n1019,n1012);
xor (n1027,n1028,n1035);
xor (n1028,n1029,n1032);
or (n1029,n1030,n1031);
and (n1030,n871,n879);
and (n1031,n872,n873);
or (n1032,n1033,n1034);
and (n1033,n765,n785);
and (n1034,n766,n776);
xor (n1035,n1036,n1050);
xor (n1036,n1037,n1043);
nand (n1037,n1038,n1039);
or (n1038,n121,n884);
or (n1039,n1040,n126);
nor (n1040,n1041,n1042);
and (n1041,n55,n221);
and (n1042,n56,n220);
nand (n1043,n1044,n1049);
or (n1044,n1045,n736);
not (n1045,n1046);
nand (n1046,n1047,n1048);
or (n1047,n331,n49);
or (n1048,n48,n332);
nand (n1049,n52,n773);
nand (n1050,n1051,n1052);
or (n1051,n782,n643);
or (n1052,n1053,n644);
not (n1053,n1054);
nor (n1054,n1055,n1056);
and (n1055,n153,n649);
and (n1056,n154,n302);
or (n1057,n1058,n1059);
and (n1058,n848,n870);
and (n1059,n849,n850);
not (n1060,n1061);
or (n1061,n1062,n1063);
and (n1062,n763,n847);
and (n1063,n764,n794);
or (n1064,n1065,n1197);
and (n1065,n1066,n1094);
xor (n1066,n1067,n1093);
or (n1067,n1068,n1092);
and (n1068,n1069,n1091);
xor (n1069,n1070,n1077);
nand (n1070,n1071,n1076);
or (n1071,n316,n1072);
not (n1072,n1073);
nor (n1073,n1074,n1075);
and (n1074,n500,n110);
and (n1075,n499,n112);
or (n1076,n948,n613);
and (n1077,n1078,n1084);
nor (n1078,n1079,n112);
nor (n1079,n1080,n1083);
and (n1080,n1081,n103);
not (n1081,n1082);
and (n1082,n560,n102);
and (n1083,n559,n109);
nand (n1084,n1085,n1086);
or (n1085,n644,n965);
nand (n1086,n1087,n1090);
nand (n1087,n1088,n1089);
or (n1088,n280,n649);
nand (n1089,n649,n280);
not (n1090,n643);
xor (n1091,n961,n970);
and (n1092,n1070,n1077);
xor (n1093,n957,n978);
or (n1094,n1095,n1196);
and (n1095,n1096,n1115);
xor (n1096,n1097,n1114);
or (n1097,n1098,n1113);
and (n1098,n1099,n1112);
xor (n1099,n1100,n1105);
nand (n1100,n1101,n1104);
or (n1101,n1102,n305);
not (n1102,n1103);
xor (n1103,n430,n103);
nand (n1104,n298,n973);
nand (n1105,n1106,n1111);
or (n1106,n1107,n316);
not (n1107,n1108);
nand (n1108,n1109,n1110);
or (n1109,n112,n560);
or (n1110,n559,n110);
nand (n1111,n1073,n100);
xor (n1112,n1078,n1084);
and (n1113,n1100,n1105);
xor (n1114,n1069,n1091);
or (n1115,n1116,n1195);
and (n1116,n1117,n1139);
xor (n1117,n1118,n1138);
or (n1118,n1119,n1137);
and (n1119,n1120,n1129);
xor (n1120,n1121,n1122);
and (n1121,n100,n560);
nand (n1122,n1123,n1128);
or (n1123,n1124,n305);
not (n1124,n1125);
nor (n1125,n1126,n1127);
and (n1126,n499,n103);
and (n1127,n500,n104);
nand (n1128,n298,n1103);
nand (n1129,n1130,n1135);
or (n1130,n643,n1131);
not (n1131,n1132);
nand (n1132,n1133,n1134);
or (n1133,n332,n649);
nand (n1134,n649,n332);
or (n1135,n1136,n644);
not (n1136,n1087);
and (n1137,n1121,n1122);
xor (n1138,n1099,n1112);
nand (n1139,n1140,n1194);
or (n1140,n1141,n1156);
nor (n1141,n1142,n1143);
xor (n1142,n1120,n1129);
nor (n1143,n1144,n1151);
not (n1144,n1145);
nand (n1145,n1146,n1150);
or (n1146,n643,n1147);
nor (n1147,n1148,n1149);
and (n1148,n430,n302);
and (n1149,n431,n649);
nand (n1150,n1132,n645);
nand (n1151,n1152,n104);
nand (n1152,n1153,n1155);
or (n1153,n1154,n302);
and (n1154,n560,n301);
or (n1155,n560,n301);
nor (n1156,n1157,n1193);
and (n1157,n1158,n1169);
nand (n1158,n1159,n1163);
nor (n1159,n1160,n1161);
and (n1160,n1151,n1145);
and (n1161,n1162,n1144);
not (n1162,n1151);
nor (n1163,n1164,n1168);
and (n1164,n304,n1165);
nand (n1165,n1166,n1167);
or (n1166,n103,n560);
or (n1167,n559,n104);
and (n1168,n298,n1125);
nand (n1169,n1170,n1192);
or (n1170,n1171,n1186);
not (n1171,n1172);
nor (n1172,n1173,n1184);
not (n1173,n1174);
nand (n1174,n1175,n1180);
or (n1175,n644,n1176);
not (n1176,n1177);
nor (n1177,n1178,n1179);
and (n1178,n499,n649);
and (n1179,n500,n302);
nand (n1180,n1181,n1090);
nor (n1181,n1182,n1183);
and (n1182,n559,n649);
and (n1183,n560,n302);
nand (n1184,n1185,n302);
nand (n1185,n560,n645);
not (n1186,n1187);
nand (n1187,n1188,n1191);
nor (n1188,n1189,n1190);
nor (n1189,n1176,n643);
nor (n1190,n1147,n644);
nand (n1191,n560,n298);
or (n1192,n1188,n1191);
nor (n1193,n1163,n1159);
nand (n1194,n1142,n1143);
and (n1195,n1118,n1138);
and (n1196,n1097,n1114);
and (n1197,n1067,n1093);
nand (n1198,n1199,n986);
or (n1199,n1200,n1202);
not (n1200,n1201);
nand (n1201,n762,n887);
not (n1202,n1203);
nand (n1203,n761,n1204);
nand (n1204,n1205,n1207);
or (n1205,n981,n1206);
nand (n1206,n927,n955);
nand (n1207,n982,n983);
nand (n1208,n988,n1061);
not (n1209,n1210);
nor (n1210,n1211,n1471);
nor (n1211,n1212,n1448);
xor (n1212,n1213,n1368);
xor (n1213,n1214,n1285);
xor (n1214,n1215,n1265);
xor (n1215,n1216,n1250);
or (n1216,n1217,n1249);
and (n1217,n1218,n1238);
xor (n1218,n1219,n1229);
nand (n1219,n1220,n1225);
or (n1220,n1221,n121);
not (n1221,n1222);
nor (n1222,n1223,n1224);
and (n1223,n86,n56);
and (n1224,n85,n55);
nand (n1225,n127,n1226);
nor (n1226,n1227,n1228);
and (n1227,n91,n55);
and (n1228,n92,n56);
nand (n1229,n1230,n1234);
or (n1230,n51,n1231);
nor (n1231,n1232,n1233);
and (n1232,n220,n49);
and (n1233,n221,n48);
nand (n1234,n53,n1235);
nor (n1235,n1236,n1237);
and (n1236,n188,n48);
and (n1237,n189,n49);
nand (n1238,n1239,n1244);
or (n1239,n613,n1240);
not (n1240,n1241);
nand (n1241,n1242,n1243);
or (n1242,n110,n39);
or (n1243,n112,n40);
nand (n1244,n1245,n106);
not (n1245,n1246);
nor (n1246,n1247,n1248);
and (n1247,n112,n20);
and (n1248,n110,n19);
and (n1249,n1219,n1229);
xor (n1250,n1251,n1259);
xor (n1251,n1252,n1256);
nand (n1252,n1253,n1255);
or (n1253,n1254,n51);
not (n1254,n1235);
nand (n1255,n53,n732);
nand (n1256,n1257,n1258);
or (n1257,n1240,n316);
nand (n1258,n100,n693);
nand (n1259,n1260,n1264);
or (n1260,n139,n1261);
nor (n1261,n1262,n1263);
and (n1262,n31,n280);
and (n1263,n29,n279);
or (n1264,n141,n701);
xor (n1265,n1266,n1281);
xor (n1266,n1267,n1274);
nand (n1267,n1268,n1273);
or (n1268,n1269,n305);
not (n1269,n1270);
nor (n1270,n1271,n1272);
and (n1271,n161,n103);
and (n1272,n159,n104);
nand (n1273,n682,n298);
nand (n1274,n1275,n1280);
or (n1275,n1276,n71);
not (n1276,n1277);
nand (n1277,n1278,n1279);
or (n1278,n79,n560);
or (n1279,n80,n559);
nand (n1280,n718,n73);
nand (n1281,n1282,n1283);
or (n1282,n724,n126);
or (n1283,n121,n1284);
not (n1284,n1226);
or (n1285,n1286,n1367);
and (n1286,n1287,n1324);
xor (n1287,n1288,n1289);
xor (n1288,n1218,n1238);
xor (n1289,n1290,n1308);
xor (n1290,n1291,n1298);
nand (n1291,n1292,n1296);
or (n1292,n1293,n139);
nor (n1293,n1294,n1295);
and (n1294,n331,n29);
and (n1295,n332,n31);
nand (n1296,n1297,n142);
not (n1297,n1261);
nand (n1298,n1299,n1303);
or (n1299,n24,n1300);
nor (n1300,n1301,n1302);
and (n1301,n23,n500);
and (n1302,n21,n499);
nand (n1303,n1304,n36);
not (n1304,n1305);
nor (n1305,n1306,n1307);
and (n1306,n23,n431);
and (n1307,n21,n430);
and (n1308,n1309,n1314);
nor (n1309,n1310,n23);
nor (n1310,n1311,n1313);
and (n1311,n1312,n31);
nand (n1312,n560,n28);
and (n1313,n559,n27);
nand (n1314,n1315,n1320);
or (n1315,n643,n1316);
not (n1316,n1317);
nor (n1317,n1318,n1319);
and (n1318,n161,n649);
and (n1319,n159,n302);
nand (n1320,n1321,n645);
nor (n1321,n1322,n1323);
and (n1322,n204,n649);
and (n1323,n47,n302);
or (n1324,n1325,n1366);
and (n1325,n1326,n1347);
xor (n1326,n1327,n1328);
xor (n1327,n1309,n1314);
or (n1328,n1329,n1346);
and (n1329,n1330,n1339);
xor (n1330,n1331,n1332);
and (n1331,n36,n560);
nand (n1332,n1333,n1335);
or (n1333,n1334,n305);
not (n1334,n1023);
nand (n1335,n298,n1336);
nor (n1336,n1337,n1338);
and (n1337,n39,n103);
and (n1338,n40,n104);
nand (n1339,n1340,n1345);
or (n1340,n1341,n126);
not (n1341,n1342);
nand (n1342,n1343,n1344);
or (n1343,n56,n188);
or (n1344,n55,n189);
or (n1345,n121,n1040);
and (n1346,n1331,n1332);
or (n1347,n1348,n1365);
and (n1348,n1349,n1359);
xor (n1349,n1350,n1356);
nand (n1350,n1351,n1352);
or (n1351,n1045,n51);
nand (n1352,n1353,n53);
nor (n1353,n1354,n1355);
and (n1354,n279,n48);
and (n1355,n280,n49);
nand (n1356,n1357,n1358);
or (n1357,n644,n1316);
nand (n1358,n1054,n1090);
nand (n1359,n1360,n1361);
or (n1360,n994,n139);
nand (n1361,n1362,n142);
nor (n1362,n1363,n1364);
and (n1363,n430,n31);
and (n1364,n431,n29);
and (n1365,n1350,n1356);
and (n1366,n1327,n1328);
and (n1367,n1288,n1289);
xor (n1368,n1369,n1408);
xor (n1369,n1370,n1373);
or (n1370,n1371,n1372);
and (n1371,n1290,n1308);
and (n1372,n1291,n1298);
xor (n1373,n1374,n1392);
xor (n1374,n1375,n1378);
nand (n1375,n1376,n1377);
or (n1376,n24,n1305);
or (n1377,n25,n708);
xor (n1378,n1379,n1385);
nor (n1379,n1380,n79);
nor (n1380,n1381,n1383);
and (n1381,n1382,n23);
nand (n1382,n560,n75);
and (n1383,n559,n1384);
not (n1384,n75);
nand (n1385,n1386,n1391);
or (n1386,n1387,n643);
not (n1387,n1388);
nor (n1388,n1389,n1390);
and (n1389,n66,n649);
and (n1390,n67,n302);
or (n1391,n675,n644);
or (n1392,n1393,n1407);
and (n1393,n1394,n1400);
xor (n1394,n1395,n1396);
and (n1395,n73,n560);
nand (n1396,n1397,n1399);
or (n1397,n643,n1398);
not (n1398,n1321);
nand (n1399,n1388,n645);
nand (n1400,n1401,n1406);
or (n1401,n305,n1402);
not (n1402,n1403);
nor (n1403,n1404,n1405);
and (n1404,n103,n153);
and (n1405,n154,n104);
or (n1406,n306,n1269);
and (n1407,n1395,n1396);
or (n1408,n1409,n1447);
and (n1409,n1410,n1446);
xor (n1410,n1411,n1426);
or (n1411,n1412,n1425);
and (n1412,n1413,n1421);
xor (n1413,n1414,n1418);
nand (n1414,n1415,n1417);
or (n1415,n1416,n305);
not (n1416,n1336);
nand (n1417,n1403,n298);
nand (n1418,n1419,n1420);
or (n1419,n1341,n121);
nand (n1420,n127,n1222);
nand (n1421,n1422,n1424);
or (n1422,n51,n1423);
not (n1423,n1353);
or (n1424,n736,n1231);
and (n1425,n1414,n1418);
or (n1426,n1427,n1445);
and (n1427,n1428,n1439);
xor (n1428,n1429,n1435);
nand (n1429,n1430,n1434);
or (n1430,n316,n1431);
nor (n1431,n1432,n1433);
and (n1432,n92,n112);
and (n1433,n91,n110);
or (n1434,n1246,n613);
nand (n1435,n1436,n1438);
or (n1436,n139,n1437);
not (n1437,n1362);
or (n1438,n1293,n141);
nand (n1439,n1440,n1444);
or (n1440,n24,n1441);
nor (n1441,n1442,n1443);
and (n1442,n559,n21);
and (n1443,n560,n23);
or (n1444,n1300,n25);
and (n1445,n1429,n1435);
xor (n1446,n1394,n1400);
and (n1447,n1411,n1426);
or (n1448,n1449,n1470);
and (n1449,n1450,n1453);
xor (n1450,n1451,n1452);
xor (n1451,n1410,n1446);
xor (n1452,n1287,n1324);
or (n1453,n1454,n1469);
and (n1454,n1455,n1458);
xor (n1455,n1456,n1457);
xor (n1456,n1428,n1439);
xor (n1457,n1413,n1421);
or (n1458,n1459,n1468);
and (n1459,n1460,n1465);
xor (n1460,n1461,n1464);
nand (n1461,n1462,n1463);
or (n1462,n316,n1006);
or (n1463,n1431,n613);
nor (n1464,n1018,n1012);
or (n1465,n1466,n1467);
and (n1466,n1036,n1050);
and (n1467,n1037,n1043);
and (n1468,n1461,n1464);
and (n1469,n1456,n1457);
and (n1470,n1451,n1452);
nand (n1471,n1472,n1501);
nor (n1472,n1473,n1496);
nor (n1473,n1474,n1487);
xor (n1474,n1475,n1486);
xor (n1475,n1476,n1477);
xor (n1476,n1326,n1347);
or (n1477,n1478,n1485);
and (n1478,n1479,n1482);
xor (n1479,n1480,n1481);
xor (n1480,n1349,n1359);
xor (n1481,n1330,n1339);
or (n1482,n1483,n1484);
and (n1483,n991,n1009);
and (n1484,n992,n1003);
and (n1485,n1480,n1481);
xor (n1486,n1455,n1458);
or (n1487,n1488,n1495);
and (n1488,n1489,n1494);
xor (n1489,n1490,n1491);
xor (n1490,n1460,n1465);
or (n1491,n1492,n1493);
and (n1492,n1028,n1035);
and (n1493,n1029,n1032);
xor (n1494,n1479,n1482);
and (n1495,n1490,n1491);
nor (n1496,n1497,n1500);
or (n1497,n1498,n1499);
and (n1498,n989,n1057);
and (n1499,n990,n1027);
xor (n1500,n1489,n1494);
nand (n1501,n1502,n1504);
not (n1502,n1503);
xor (n1503,n1450,n1453);
not (n1504,n1505);
or (n1505,n1506,n1507);
and (n1506,n1475,n1486);
and (n1507,n1476,n1477);
nor (n1508,n1509,n1520);
and (n1509,n1510,n1519);
nand (n1510,n1511,n1518);
or (n1511,n1512,n1513);
not (n1512,n1501);
not (n1513,n1514);
nand (n1514,n1515,n1517);
or (n1515,n1473,n1516);
nand (n1516,n1497,n1500);
nand (n1517,n1474,n1487);
nand (n1518,n1503,n1505);
not (n1519,n1211);
and (n1520,n1212,n1448);
not (n1521,n1522);
and (n1522,n1523,n1574);
nor (n1523,n1524,n1555);
nor (n1524,n1525,n1526);
xor (n1525,n661,n748);
or (n1526,n1527,n1554);
and (n1527,n1528,n1553);
xor (n1528,n1529,n1530);
xor (n1529,n621,n653);
or (n1530,n1531,n1552);
and (n1531,n1532,n1545);
xor (n1532,n1533,n1544);
or (n1533,n1534,n1543);
and (n1534,n1535,n1540);
xor (n1535,n1536,n1537);
and (n1536,n1379,n1385);
or (n1537,n1538,n1539);
and (n1538,n1266,n1281);
and (n1539,n1267,n1274);
or (n1540,n1541,n1542);
and (n1541,n1251,n1259);
and (n1542,n1252,n1256);
and (n1543,n1536,n1537);
xor (n1544,n668,n712);
or (n1545,n1546,n1551);
and (n1546,n1547,n1550);
xor (n1547,n1548,n1549);
xor (n1548,n689,n704);
xor (n1549,n671,n679);
xor (n1550,n714,n729);
and (n1551,n1548,n1549);
and (n1552,n1533,n1544);
xor (n1553,n665,n746);
and (n1554,n1529,n1530);
nor (n1555,n1556,n1557);
xor (n1556,n1528,n1553);
or (n1557,n1558,n1573);
and (n1558,n1559,n1572);
xor (n1559,n1560,n1561);
xor (n1560,n741,n744);
or (n1561,n1562,n1571);
and (n1562,n1563,n1568);
xor (n1563,n1564,n1567);
or (n1564,n1565,n1566);
and (n1565,n1374,n1392);
and (n1566,n1375,n1378);
xor (n1567,n1535,n1540);
or (n1568,n1569,n1570);
and (n1569,n1215,n1265);
and (n1570,n1216,n1250);
and (n1571,n1564,n1567);
xor (n1572,n1532,n1545);
and (n1573,n1560,n1561);
nor (n1574,n1575,n1586);
nor (n1575,n1576,n1577);
xor (n1576,n1559,n1572);
or (n1577,n1578,n1585);
and (n1578,n1579,n1584);
xor (n1579,n1580,n1581);
xor (n1580,n1547,n1550);
or (n1581,n1582,n1583);
and (n1582,n1369,n1408);
and (n1583,n1370,n1373);
xor (n1584,n1563,n1568);
and (n1585,n1580,n1581);
nor (n1586,n1587,n1588);
xor (n1587,n1579,n1584);
or (n1588,n1589,n1590);
and (n1589,n1213,n1368);
and (n1590,n1214,n1285);
not (n1591,n1592);
nand (n1592,n1593,n1600);
or (n1593,n1594,n1599);
not (n1594,n1595);
nor (n1595,n1596,n1575);
and (n1596,n1597,n1598);
nand (n1597,n1576,n1577);
nand (n1598,n1587,n1588);
not (n1599,n1523);
nor (n1600,n1601,n1605);
and (n1601,n1602,n1603);
not (n1602,n1524);
not (n1603,n1604);
nand (n1604,n1556,n1557);
and (n1605,n1525,n1526);
not (n1606,n1607);
nor (n1607,n1608,n577);
and (n1608,n1609,n1610);
nand (n1609,n579,n578);
nand (n1610,n658,n659);
nand (n1611,n450,n451);
and (n1612,n1613,n1614);
not (n1613,n5);
not (n1614,n447);
nand (n1615,n1616,n1618);
not (n1616,n1617);
nand (n1619,n1620,n1621);
nor (n1620,n1618,n1617);
wire s0n1622,s1n1622,notn1622;
or (n1622,s0n1622,s1n1622);
not(notn1622,n1617);
and (s0n1622,notn1622,n1623);
and (s1n1622,n1617,1'b0);
wire s0n1623,s1n1623,notn1623;
or (n1623,s0n1623,s1n1623);
not(notn1623,n1618);
and (s0n1623,notn1623,n1621);
and (s1n1623,n1618,n1624);
xor (n1624,n1625,n2801);
xor (n1625,n1626,n2800);
xor (n1626,n1627,n2760);
xor (n1627,n1628,n2759);
xor (n1628,n1629,n2708);
xor (n1629,n1630,n2707);
xor (n1630,n1631,n2652);
xor (n1631,n1632,n41);
xor (n1632,n1633,n2589);
xor (n1633,n1634,n2588);
xor (n1634,n1635,n2523);
xor (n1635,n1636,n2522);
xor (n1636,n1637,n2448);
xor (n1637,n1638,n2447);
xor (n1638,n1639,n2375);
xor (n1639,n1640,n68);
xor (n1640,n1641,n2289);
xor (n1641,n1642,n2288);
xor (n1642,n1643,n2204);
xor (n1643,n1644,n2203);
or (n1644,n1645,n2109);
and (n1645,n1646,n2108);
or (n1646,n1647,n2016);
and (n1647,n1648,n229);
or (n1648,n1649,n1922);
and (n1649,n1650,n1921);
or (n1650,n1651,n1834);
and (n1651,n1652,n377);
or (n1652,n1653,n1740);
and (n1653,n1654,n1739);
and (n1654,n650,n1655);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
and (n1657,n134,n645);
and (n1658,n119,n302);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1664);
and (n1662,n1663,n1390);
and (n1663,n119,n645);
and (n1664,n1665,n1666);
xor (n1665,n1663,n1390);
or (n1666,n1667,n1669);
and (n1667,n1668,n1323);
and (n1668,n67,n645);
and (n1669,n1670,n1671);
xor (n1670,n1668,n1323);
or (n1671,n1672,n1674);
and (n1672,n1673,n1319);
and (n1673,n47,n645);
and (n1674,n1675,n1676);
xor (n1675,n1673,n1319);
or (n1676,n1677,n1679);
and (n1677,n1678,n1056);
and (n1678,n159,n645);
and (n1679,n1680,n1681);
xor (n1680,n1678,n1056);
or (n1681,n1682,n1685);
and (n1682,n1683,n1684);
and (n1683,n154,n645);
and (n1684,n40,n302);
and (n1685,n1686,n1687);
xor (n1686,n1683,n1684);
or (n1687,n1688,n1691);
and (n1688,n1689,n1690);
and (n1689,n40,n645);
and (n1690,n20,n302);
and (n1691,n1692,n1693);
xor (n1692,n1689,n1690);
or (n1693,n1694,n1696);
and (n1694,n1695,n830);
and (n1695,n20,n645);
and (n1696,n1697,n1698);
xor (n1697,n1695,n830);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
and (n1700,n92,n645);
and (n1701,n86,n302);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1707);
and (n1705,n1706,n919);
and (n1706,n86,n645);
and (n1707,n1708,n1709);
xor (n1708,n1706,n919);
or (n1709,n1710,n1712);
and (n1710,n1711,n967);
and (n1711,n189,n645);
and (n1712,n1713,n1714);
xor (n1713,n1711,n967);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
and (n1716,n221,n645);
and (n1717,n280,n302);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
and (n1722,n280,n645);
and (n1723,n332,n302);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
and (n1728,n332,n645);
and (n1729,n431,n302);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1735);
and (n1733,n1734,n1179);
and (n1734,n431,n645);
and (n1735,n1736,n1737);
xor (n1736,n1734,n1179);
and (n1737,n1738,n1183);
and (n1738,n500,n645);
and (n1739,n134,n301);
and (n1740,n1741,n1742);
xor (n1741,n1654,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n650,n1655);
and (n1745,n119,n301);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1660,n1661);
and (n1751,n67,n301);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1665,n1666);
and (n1757,n47,n301);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1670,n1671);
and (n1763,n159,n301);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1675,n1676);
and (n1769,n154,n301);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
or (n1772,n1773,n1776);
and (n1773,n1774,n1775);
xor (n1774,n1680,n1681);
and (n1775,n40,n301);
and (n1776,n1777,n1778);
xor (n1777,n1774,n1775);
or (n1778,n1779,n1782);
and (n1779,n1780,n1781);
xor (n1780,n1686,n1687);
and (n1781,n20,n301);
and (n1782,n1783,n1784);
xor (n1783,n1780,n1781);
or (n1784,n1785,n1788);
and (n1785,n1786,n1787);
xor (n1786,n1692,n1693);
and (n1787,n92,n301);
and (n1788,n1789,n1790);
xor (n1789,n1786,n1787);
or (n1790,n1791,n1794);
and (n1791,n1792,n1793);
xor (n1792,n1697,n1698);
and (n1793,n86,n301);
and (n1794,n1795,n1796);
xor (n1795,n1792,n1793);
or (n1796,n1797,n1800);
and (n1797,n1798,n1799);
xor (n1798,n1703,n1704);
and (n1799,n189,n301);
and (n1800,n1801,n1802);
xor (n1801,n1798,n1799);
or (n1802,n1803,n1806);
and (n1803,n1804,n1805);
xor (n1804,n1708,n1709);
and (n1805,n221,n301);
and (n1806,n1807,n1808);
xor (n1807,n1804,n1805);
or (n1808,n1809,n1812);
and (n1809,n1810,n1811);
xor (n1810,n1713,n1714);
and (n1811,n280,n301);
and (n1812,n1813,n1814);
xor (n1813,n1810,n1811);
or (n1814,n1815,n1818);
and (n1815,n1816,n1817);
xor (n1816,n1719,n1720);
and (n1817,n332,n301);
and (n1818,n1819,n1820);
xor (n1819,n1816,n1817);
or (n1820,n1821,n1824);
and (n1821,n1822,n1823);
xor (n1822,n1725,n1726);
and (n1823,n431,n301);
and (n1824,n1825,n1826);
xor (n1825,n1822,n1823);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1731,n1732);
and (n1829,n500,n301);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
and (n1832,n1833,n1154);
xor (n1833,n1736,n1737);
and (n1834,n1835,n1836);
xor (n1835,n1652,n377);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1741,n1742);
and (n1839,n119,n104);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1845);
and (n1843,n1844,n599);
xor (n1844,n1747,n1748);
and (n1845,n1846,n1847);
xor (n1846,n1844,n599);
or (n1847,n1848,n1850);
and (n1848,n1849,n684);
xor (n1849,n1753,n1754);
and (n1850,n1851,n1852);
xor (n1851,n1849,n684);
or (n1852,n1853,n1855);
and (n1853,n1854,n1272);
xor (n1854,n1759,n1760);
and (n1855,n1856,n1857);
xor (n1856,n1854,n1272);
or (n1857,n1858,n1860);
and (n1858,n1859,n1405);
xor (n1859,n1765,n1766);
and (n1860,n1861,n1862);
xor (n1861,n1859,n1405);
or (n1862,n1863,n1865);
and (n1863,n1864,n1338);
xor (n1864,n1771,n1772);
and (n1865,n1866,n1867);
xor (n1866,n1864,n1338);
or (n1867,n1868,n1870);
and (n1868,n1869,n1025);
xor (n1869,n1777,n1778);
and (n1870,n1871,n1872);
xor (n1871,n1869,n1025);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1783,n1784);
and (n1875,n92,n104);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1789,n1790);
and (n1881,n86,n104);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1795,n1796);
and (n1887,n189,n104);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1801,n1802);
and (n1893,n221,n104);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1807,n1808);
and (n1899,n280,n104);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1905);
and (n1903,n1904,n975);
xor (n1904,n1813,n1814);
and (n1905,n1906,n1907);
xor (n1906,n1904,n975);
or (n1907,n1908,n1911);
and (n1908,n1909,n1910);
xor (n1909,n1819,n1820);
and (n1910,n431,n104);
and (n1911,n1912,n1913);
xor (n1912,n1909,n1910);
or (n1913,n1914,n1916);
and (n1914,n1915,n1127);
xor (n1915,n1825,n1826);
and (n1916,n1917,n1918);
xor (n1917,n1915,n1127);
and (n1918,n1919,n1920);
xor (n1919,n1831,n1832);
and (n1920,n560,n104);
and (n1921,n134,n102);
and (n1922,n1923,n1924);
xor (n1923,n1650,n1921);
or (n1924,n1925,n1928);
and (n1925,n1926,n1927);
xor (n1926,n1835,n1836);
and (n1927,n119,n102);
and (n1928,n1929,n1930);
xor (n1929,n1926,n1927);
or (n1930,n1931,n1934);
and (n1931,n1932,n1933);
xor (n1932,n1841,n1842);
and (n1933,n67,n102);
and (n1934,n1935,n1936);
xor (n1935,n1932,n1933);
or (n1936,n1937,n1940);
and (n1937,n1938,n1939);
xor (n1938,n1846,n1847);
and (n1939,n47,n102);
and (n1940,n1941,n1942);
xor (n1941,n1938,n1939);
or (n1942,n1943,n1946);
and (n1943,n1944,n1945);
xor (n1944,n1851,n1852);
and (n1945,n159,n102);
and (n1946,n1947,n1948);
xor (n1947,n1944,n1945);
or (n1948,n1949,n1952);
and (n1949,n1950,n1951);
xor (n1950,n1856,n1857);
and (n1951,n154,n102);
and (n1952,n1953,n1954);
xor (n1953,n1950,n1951);
or (n1954,n1955,n1958);
and (n1955,n1956,n1957);
xor (n1956,n1861,n1862);
and (n1957,n40,n102);
and (n1958,n1959,n1960);
xor (n1959,n1956,n1957);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
xor (n1962,n1866,n1867);
and (n1963,n20,n102);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
xor (n1968,n1871,n1872);
and (n1969,n92,n102);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
xor (n1974,n1877,n1878);
and (n1975,n86,n102);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
xor (n1980,n1883,n1884);
and (n1981,n189,n102);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
xor (n1986,n1889,n1890);
and (n1987,n221,n102);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
or (n1990,n1991,n1994);
and (n1991,n1992,n1993);
xor (n1992,n1895,n1896);
and (n1993,n280,n102);
and (n1994,n1995,n1996);
xor (n1995,n1992,n1993);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
xor (n1998,n1901,n1902);
and (n1999,n332,n102);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2006);
and (n2003,n2004,n2005);
xor (n2004,n1906,n1907);
and (n2005,n431,n102);
and (n2006,n2007,n2008);
xor (n2007,n2004,n2005);
or (n2008,n2009,n2012);
and (n2009,n2010,n2011);
xor (n2010,n1912,n1913);
and (n2011,n500,n102);
and (n2012,n2013,n2014);
xor (n2013,n2010,n2011);
and (n2014,n2015,n1082);
xor (n2015,n1917,n1918);
and (n2016,n2017,n2018);
xor (n2017,n1648,n229);
or (n2018,n2019,n2022);
and (n2019,n2020,n2021);
xor (n2020,n1923,n1924);
and (n2021,n119,n110);
and (n2022,n2023,n2024);
xor (n2023,n2020,n2021);
or (n2024,n2025,n2027);
and (n2025,n2026,n426);
xor (n2026,n1929,n1930);
and (n2027,n2028,n2029);
xor (n2028,n2026,n426);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1935,n1936);
and (n2032,n47,n110);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1941,n1942);
and (n2038,n159,n110);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
or (n2041,n2042,n2044);
and (n2042,n2043,n695);
xor (n2043,n1947,n1948);
and (n2044,n2045,n2046);
xor (n2045,n2043,n695);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1953,n1954);
and (n2049,n40,n110);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
or (n2052,n2053,n2056);
and (n2053,n2054,n2055);
xor (n2054,n1959,n1960);
and (n2055,n20,n110);
and (n2056,n2057,n2058);
xor (n2057,n2054,n2055);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n1965,n1966);
and (n2061,n92,n110);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n1971,n1972);
and (n2067,n86,n110);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2074);
and (n2071,n2072,n2073);
xor (n2072,n1977,n1978);
and (n2073,n189,n110);
and (n2074,n2075,n2076);
xor (n2075,n2072,n2073);
or (n2076,n2077,n2080);
and (n2077,n2078,n2079);
xor (n2078,n1983,n1984);
and (n2079,n221,n110);
and (n2080,n2081,n2082);
xor (n2081,n2078,n2079);
or (n2082,n2083,n2086);
and (n2083,n2084,n2085);
xor (n2084,n1989,n1990);
and (n2085,n280,n110);
and (n2086,n2087,n2088);
xor (n2087,n2084,n2085);
or (n2088,n2089,n2092);
and (n2089,n2090,n2091);
xor (n2090,n1995,n1996);
and (n2091,n332,n110);
and (n2092,n2093,n2094);
xor (n2093,n2090,n2091);
or (n2094,n2095,n2098);
and (n2095,n2096,n2097);
xor (n2096,n2001,n2002);
and (n2097,n431,n110);
and (n2098,n2099,n2100);
xor (n2099,n2096,n2097);
or (n2100,n2101,n2103);
and (n2101,n2102,n1074);
xor (n2102,n2007,n2008);
and (n2103,n2104,n2105);
xor (n2104,n2102,n1074);
and (n2105,n2106,n2107);
xor (n2106,n2013,n2014);
and (n2107,n560,n110);
and (n2108,n134,n124);
and (n2109,n2110,n2111);
xor (n2110,n1646,n2108);
or (n2111,n2112,n2115);
and (n2112,n2113,n2114);
xor (n2113,n2017,n2018);
and (n2114,n119,n124);
and (n2115,n2116,n2117);
xor (n2116,n2113,n2114);
or (n2117,n2118,n2121);
and (n2118,n2119,n2120);
xor (n2119,n2023,n2024);
and (n2120,n67,n124);
and (n2121,n2122,n2123);
xor (n2122,n2119,n2120);
or (n2123,n2124,n2127);
and (n2124,n2125,n2126);
xor (n2125,n2028,n2029);
and (n2126,n47,n124);
and (n2127,n2128,n2129);
xor (n2128,n2125,n2126);
or (n2129,n2130,n2133);
and (n2130,n2131,n2132);
xor (n2131,n2034,n2035);
and (n2132,n159,n124);
and (n2133,n2134,n2135);
xor (n2134,n2131,n2132);
or (n2135,n2136,n2139);
and (n2136,n2137,n2138);
xor (n2137,n2040,n2041);
and (n2138,n154,n124);
and (n2139,n2140,n2141);
xor (n2140,n2137,n2138);
or (n2141,n2142,n2145);
and (n2142,n2143,n2144);
xor (n2143,n2045,n2046);
and (n2144,n40,n124);
and (n2145,n2146,n2147);
xor (n2146,n2143,n2144);
or (n2147,n2148,n2151);
and (n2148,n2149,n2150);
xor (n2149,n2051,n2052);
and (n2150,n20,n124);
and (n2151,n2152,n2153);
xor (n2152,n2149,n2150);
or (n2153,n2154,n2157);
and (n2154,n2155,n2156);
xor (n2155,n2057,n2058);
and (n2156,n92,n124);
and (n2157,n2158,n2159);
xor (n2158,n2155,n2156);
or (n2159,n2160,n2163);
and (n2160,n2161,n2162);
xor (n2161,n2063,n2064);
and (n2162,n86,n124);
and (n2163,n2164,n2165);
xor (n2164,n2161,n2162);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2069,n2070);
and (n2168,n189,n124);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2075,n2076);
and (n2174,n221,n124);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
or (n2177,n2178,n2181);
and (n2178,n2179,n2180);
xor (n2179,n2081,n2082);
and (n2180,n280,n124);
and (n2181,n2182,n2183);
xor (n2182,n2179,n2180);
or (n2183,n2184,n2187);
and (n2184,n2185,n2186);
xor (n2185,n2087,n2088);
and (n2186,n332,n124);
and (n2187,n2188,n2189);
xor (n2188,n2185,n2186);
or (n2189,n2190,n2193);
and (n2190,n2191,n2192);
xor (n2191,n2093,n2094);
and (n2192,n431,n124);
and (n2193,n2194,n2195);
xor (n2194,n2191,n2192);
or (n2195,n2196,n2199);
and (n2196,n2197,n2198);
xor (n2197,n2099,n2100);
and (n2198,n500,n124);
and (n2199,n2200,n2201);
xor (n2200,n2197,n2198);
and (n2201,n2202,n911);
xor (n2202,n2104,n2105);
and (n2203,n134,n56);
or (n2204,n2205,n2207);
and (n2205,n2206,n120);
xor (n2206,n2110,n2111);
and (n2207,n2208,n2209);
xor (n2208,n2206,n120);
or (n2209,n2210,n2212);
and (n2210,n2211,n239);
xor (n2211,n2116,n2117);
and (n2212,n2213,n2214);
xor (n2213,n2211,n239);
or (n2214,n2215,n2217);
and (n2215,n2216,n347);
xor (n2216,n2122,n2123);
and (n2217,n2218,n2219);
xor (n2218,n2216,n347);
or (n2219,n2220,n2222);
and (n2220,n2221,n409);
xor (n2221,n2128,n2129);
and (n2222,n2223,n2224);
xor (n2223,n2221,n409);
or (n2224,n2225,n2228);
and (n2225,n2226,n2227);
xor (n2226,n2134,n2135);
and (n2227,n154,n56);
and (n2228,n2229,n2230);
xor (n2229,n2226,n2227);
or (n2230,n2231,n2233);
and (n2231,n2232,n548);
xor (n2232,n2140,n2141);
and (n2233,n2234,n2235);
xor (n2234,n2232,n548);
or (n2235,n2236,n2239);
and (n2236,n2237,n2238);
xor (n2237,n2146,n2147);
and (n2238,n20,n56);
and (n2239,n2240,n2241);
xor (n2240,n2237,n2238);
or (n2241,n2242,n2244);
and (n2242,n2243,n1228);
xor (n2243,n2152,n2153);
and (n2244,n2245,n2246);
xor (n2245,n2243,n1228);
or (n2246,n2247,n2249);
and (n2247,n2248,n1223);
xor (n2248,n2158,n2159);
and (n2249,n2250,n2251);
xor (n2250,n2248,n1223);
or (n2251,n2252,n2255);
and (n2252,n2253,n2254);
xor (n2253,n2164,n2165);
and (n2254,n189,n56);
and (n2255,n2256,n2257);
xor (n2256,n2253,n2254);
or (n2257,n2258,n2261);
and (n2258,n2259,n2260);
xor (n2259,n2170,n2171);
and (n2260,n221,n56);
and (n2261,n2262,n2263);
xor (n2262,n2259,n2260);
or (n2263,n2264,n2267);
and (n2264,n2265,n2266);
xor (n2265,n2176,n2177);
and (n2266,n280,n56);
and (n2267,n2268,n2269);
xor (n2268,n2265,n2266);
or (n2269,n2270,n2272);
and (n2270,n2271,n858);
xor (n2271,n2182,n2183);
and (n2272,n2273,n2274);
xor (n2273,n2271,n858);
or (n2274,n2275,n2277);
and (n2275,n2276,n843);
xor (n2276,n2188,n2189);
and (n2277,n2278,n2279);
xor (n2278,n2276,n843);
or (n2279,n2280,n2283);
and (n2280,n2281,n2282);
xor (n2281,n2194,n2195);
and (n2282,n500,n56);
and (n2283,n2284,n2285);
xor (n2284,n2281,n2282);
and (n2285,n2286,n2287);
xor (n2286,n2200,n2201);
and (n2287,n560,n56);
and (n2288,n119,n57);
or (n2289,n2290,n2293);
and (n2290,n2291,n2292);
xor (n2291,n2208,n2209);
and (n2292,n67,n57);
and (n2293,n2294,n2295);
xor (n2294,n2291,n2292);
or (n2295,n2296,n2299);
and (n2296,n2297,n2298);
xor (n2297,n2213,n2214);
and (n2298,n47,n57);
and (n2299,n2300,n2301);
xor (n2300,n2297,n2298);
or (n2301,n2302,n2305);
and (n2302,n2303,n2304);
xor (n2303,n2218,n2219);
and (n2304,n159,n57);
and (n2305,n2306,n2307);
xor (n2306,n2303,n2304);
or (n2307,n2308,n2311);
and (n2308,n2309,n2310);
xor (n2309,n2223,n2224);
and (n2310,n154,n57);
and (n2311,n2312,n2313);
xor (n2312,n2309,n2310);
or (n2313,n2314,n2317);
and (n2314,n2315,n2316);
xor (n2315,n2229,n2230);
and (n2316,n40,n57);
and (n2317,n2318,n2319);
xor (n2318,n2315,n2316);
or (n2319,n2320,n2323);
and (n2320,n2321,n2322);
xor (n2321,n2234,n2235);
and (n2322,n20,n57);
and (n2323,n2324,n2325);
xor (n2324,n2321,n2322);
or (n2325,n2326,n2329);
and (n2326,n2327,n2328);
xor (n2327,n2240,n2241);
and (n2328,n92,n57);
and (n2329,n2330,n2331);
xor (n2330,n2327,n2328);
or (n2331,n2332,n2335);
and (n2332,n2333,n2334);
xor (n2333,n2245,n2246);
and (n2334,n86,n57);
and (n2335,n2336,n2337);
xor (n2336,n2333,n2334);
or (n2337,n2338,n2341);
and (n2338,n2339,n2340);
xor (n2339,n2250,n2251);
and (n2340,n189,n57);
and (n2341,n2342,n2343);
xor (n2342,n2339,n2340);
or (n2343,n2344,n2347);
and (n2344,n2345,n2346);
xor (n2345,n2256,n2257);
and (n2346,n221,n57);
and (n2347,n2348,n2349);
xor (n2348,n2345,n2346);
or (n2349,n2350,n2353);
and (n2350,n2351,n2352);
xor (n2351,n2262,n2263);
and (n2352,n280,n57);
and (n2353,n2354,n2355);
xor (n2354,n2351,n2352);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2268,n2269);
and (n2358,n332,n57);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2273,n2274);
and (n2364,n431,n57);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2278,n2279);
and (n2370,n500,n57);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
and (n2373,n2374,n809);
xor (n2374,n2284,n2285);
or (n2375,n2376,n2379);
and (n2376,n2377,n2378);
xor (n2377,n2294,n2295);
and (n2378,n47,n49);
and (n2379,n2380,n2381);
xor (n2380,n2377,n2378);
or (n2381,n2382,n2384);
and (n2382,n2383,n268);
xor (n2383,n2300,n2301);
and (n2384,n2385,n2386);
xor (n2385,n2383,n268);
or (n2386,n2387,n2389);
and (n2387,n2388,n323);
xor (n2388,n2306,n2307);
and (n2389,n2390,n2391);
xor (n2390,n2388,n323);
or (n2391,n2392,n2394);
and (n2392,n2393,n438);
xor (n2393,n2312,n2313);
and (n2394,n2395,n2396);
xor (n2395,n2393,n438);
or (n2396,n2397,n2399);
and (n2397,n2398,n517);
xor (n2398,n2318,n2319);
and (n2399,n2400,n2401);
xor (n2400,n2398,n517);
or (n2401,n2402,n2404);
and (n2402,n2403,n606);
xor (n2403,n2324,n2325);
and (n2404,n2405,n2406);
xor (n2405,n2403,n606);
or (n2406,n2407,n2409);
and (n2407,n2408,n734);
xor (n2408,n2330,n2331);
and (n2409,n2410,n2411);
xor (n2410,n2408,n734);
or (n2411,n2412,n2414);
and (n2412,n2413,n1237);
xor (n2413,n2336,n2337);
and (n2414,n2415,n2416);
xor (n2415,n2413,n1237);
or (n2416,n2417,n2420);
and (n2417,n2418,n2419);
xor (n2418,n2342,n2343);
and (n2419,n221,n49);
and (n2420,n2421,n2422);
xor (n2421,n2418,n2419);
or (n2422,n2423,n2425);
and (n2423,n2424,n1355);
xor (n2424,n2348,n2349);
and (n2425,n2426,n2427);
xor (n2426,n2424,n1355);
or (n2427,n2428,n2431);
and (n2428,n2429,n2430);
xor (n2429,n2354,n2355);
and (n2430,n332,n49);
and (n2431,n2432,n2433);
xor (n2432,n2429,n2430);
or (n2433,n2434,n2437);
and (n2434,n2435,n2436);
xor (n2435,n2360,n2361);
and (n2436,n431,n49);
and (n2437,n2438,n2439);
xor (n2438,n2435,n2436);
or (n2439,n2440,n2442);
and (n2440,n2441,n771);
xor (n2441,n2366,n2367);
and (n2442,n2443,n2444);
xor (n2443,n2441,n771);
and (n2444,n2445,n2446);
xor (n2445,n2372,n2373);
and (n2446,n560,n49);
and (n2447,n47,n145);
or (n2448,n2449,n2452);
and (n2449,n2450,n2451);
xor (n2450,n2380,n2381);
and (n2451,n159,n145);
and (n2452,n2453,n2454);
xor (n2453,n2450,n2451);
or (n2454,n2455,n2458);
and (n2455,n2456,n2457);
xor (n2456,n2385,n2386);
and (n2457,n154,n145);
and (n2458,n2459,n2460);
xor (n2459,n2456,n2457);
or (n2460,n2461,n2464);
and (n2461,n2462,n2463);
xor (n2462,n2390,n2391);
and (n2463,n40,n145);
and (n2464,n2465,n2466);
xor (n2465,n2462,n2463);
or (n2466,n2467,n2470);
and (n2467,n2468,n2469);
xor (n2468,n2395,n2396);
and (n2469,n20,n145);
and (n2470,n2471,n2472);
xor (n2471,n2468,n2469);
or (n2472,n2473,n2476);
and (n2473,n2474,n2475);
xor (n2474,n2400,n2401);
and (n2475,n92,n145);
and (n2476,n2477,n2478);
xor (n2477,n2474,n2475);
or (n2478,n2479,n2482);
and (n2479,n2480,n2481);
xor (n2480,n2405,n2406);
and (n2481,n86,n145);
and (n2482,n2483,n2484);
xor (n2483,n2480,n2481);
or (n2484,n2485,n2488);
and (n2485,n2486,n2487);
xor (n2486,n2410,n2411);
and (n2487,n189,n145);
and (n2488,n2489,n2490);
xor (n2489,n2486,n2487);
or (n2490,n2491,n2494);
and (n2491,n2492,n2493);
xor (n2492,n2415,n2416);
and (n2493,n221,n145);
and (n2494,n2495,n2496);
xor (n2495,n2492,n2493);
or (n2496,n2497,n2500);
and (n2497,n2498,n2499);
xor (n2498,n2421,n2422);
and (n2499,n280,n145);
and (n2500,n2501,n2502);
xor (n2501,n2498,n2499);
or (n2502,n2503,n2506);
and (n2503,n2504,n2505);
xor (n2504,n2426,n2427);
and (n2505,n332,n145);
and (n2506,n2507,n2508);
xor (n2507,n2504,n2505);
or (n2508,n2509,n2512);
and (n2509,n2510,n2511);
xor (n2510,n2432,n2433);
and (n2511,n431,n145);
and (n2512,n2513,n2514);
xor (n2513,n2510,n2511);
or (n2514,n2515,n2518);
and (n2515,n2516,n2517);
xor (n2516,n2438,n2439);
and (n2517,n500,n145);
and (n2518,n2519,n2520);
xor (n2519,n2516,n2517);
and (n2520,n2521,n1017);
xor (n2521,n2443,n2444);
and (n2522,n159,n29);
or (n2523,n2524,n2526);
and (n2524,n2525,n155);
xor (n2525,n2453,n2454);
and (n2526,n2527,n2528);
xor (n2527,n2525,n155);
or (n2528,n2529,n2531);
and (n2529,n2530,n246);
xor (n2530,n2459,n2460);
and (n2531,n2532,n2533);
xor (n2532,n2530,n246);
or (n2533,n2534,n2536);
and (n2534,n2535,n339);
xor (n2535,n2465,n2466);
and (n2536,n2537,n2538);
xor (n2537,n2535,n339);
or (n2538,n2539,n2542);
and (n2539,n2540,n2541);
xor (n2540,n2471,n2472);
and (n2541,n92,n29);
and (n2542,n2543,n2544);
xor (n2543,n2540,n2541);
or (n2544,n2545,n2548);
and (n2545,n2546,n2547);
xor (n2546,n2477,n2478);
and (n2547,n86,n29);
and (n2548,n2549,n2550);
xor (n2549,n2546,n2547);
or (n2550,n2551,n2554);
and (n2551,n2552,n2553);
xor (n2552,n2483,n2484);
and (n2553,n189,n29);
and (n2554,n2555,n2556);
xor (n2555,n2552,n2553);
or (n2556,n2557,n2560);
and (n2557,n2558,n2559);
xor (n2558,n2489,n2490);
and (n2559,n221,n29);
and (n2560,n2561,n2562);
xor (n2561,n2558,n2559);
or (n2562,n2563,n2566);
and (n2563,n2564,n2565);
xor (n2564,n2495,n2496);
and (n2565,n280,n29);
and (n2566,n2567,n2568);
xor (n2567,n2564,n2565);
or (n2568,n2569,n2572);
and (n2569,n2570,n2571);
xor (n2570,n2501,n2502);
and (n2571,n332,n29);
and (n2572,n2573,n2574);
xor (n2573,n2570,n2571);
or (n2574,n2575,n2577);
and (n2575,n2576,n1364);
xor (n2576,n2507,n2508);
and (n2577,n2578,n2579);
xor (n2578,n2576,n1364);
or (n2579,n2580,n2583);
and (n2580,n2581,n2582);
xor (n2581,n2513,n2514);
and (n2582,n500,n29);
and (n2583,n2584,n2585);
xor (n2584,n2581,n2582);
and (n2585,n2586,n2587);
xor (n2586,n2519,n2520);
and (n2587,n560,n29);
and (n2588,n154,n28);
or (n2589,n2590,n2593);
and (n2590,n2591,n2592);
xor (n2591,n2527,n2528);
and (n2592,n40,n28);
and (n2593,n2594,n2595);
xor (n2594,n2591,n2592);
or (n2595,n2596,n2599);
and (n2596,n2597,n2598);
xor (n2597,n2532,n2533);
and (n2598,n20,n28);
and (n2599,n2600,n2601);
xor (n2600,n2597,n2598);
or (n2601,n2602,n2605);
and (n2602,n2603,n2604);
xor (n2603,n2537,n2538);
and (n2604,n92,n28);
and (n2605,n2606,n2607);
xor (n2606,n2603,n2604);
or (n2607,n2608,n2611);
and (n2608,n2609,n2610);
xor (n2609,n2543,n2544);
and (n2610,n86,n28);
and (n2611,n2612,n2613);
xor (n2612,n2609,n2610);
or (n2613,n2614,n2617);
and (n2614,n2615,n2616);
xor (n2615,n2549,n2550);
and (n2616,n189,n28);
and (n2617,n2618,n2619);
xor (n2618,n2615,n2616);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
xor (n2621,n2555,n2556);
and (n2622,n221,n28);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
xor (n2627,n2561,n2562);
and (n2628,n280,n28);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
xor (n2633,n2567,n2568);
and (n2634,n332,n28);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
xor (n2639,n2573,n2574);
and (n2640,n431,n28);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
or (n2643,n2644,n2647);
and (n2644,n2645,n2646);
xor (n2645,n2578,n2579);
and (n2646,n500,n28);
and (n2647,n2648,n2649);
xor (n2648,n2645,n2646);
and (n2649,n2650,n2651);
xor (n2650,n2584,n2585);
not (n2651,n1312);
or (n2652,n2653,n2656);
and (n2653,n2654,n2655);
xor (n2654,n2594,n2595);
and (n2655,n20,n21);
and (n2656,n2657,n2658);
xor (n2657,n2654,n2655);
or (n2658,n2659,n2661);
and (n2659,n2660,n254);
xor (n2660,n2600,n2601);
and (n2661,n2662,n2663);
xor (n2662,n2660,n254);
or (n2663,n2664,n2666);
and (n2664,n2665,n363);
xor (n2665,n2606,n2607);
and (n2666,n2667,n2668);
xor (n2667,n2665,n363);
or (n2668,n2669,n2672);
and (n2669,n2670,n2671);
xor (n2670,n2612,n2613);
and (n2671,n189,n21);
and (n2672,n2673,n2674);
xor (n2673,n2670,n2671);
or (n2674,n2675,n2678);
and (n2675,n2676,n2677);
xor (n2676,n2618,n2619);
and (n2677,n221,n21);
and (n2678,n2679,n2680);
xor (n2679,n2676,n2677);
or (n2680,n2681,n2684);
and (n2681,n2682,n2683);
xor (n2682,n2624,n2625);
and (n2683,n280,n21);
and (n2684,n2685,n2686);
xor (n2685,n2682,n2683);
or (n2686,n2687,n2690);
and (n2687,n2688,n2689);
xor (n2688,n2630,n2631);
and (n2689,n332,n21);
and (n2690,n2691,n2692);
xor (n2691,n2688,n2689);
or (n2692,n2693,n2696);
and (n2693,n2694,n2695);
xor (n2694,n2636,n2637);
and (n2695,n431,n21);
and (n2696,n2697,n2698);
xor (n2697,n2694,n2695);
or (n2698,n2699,n2702);
and (n2699,n2700,n2701);
xor (n2700,n2642,n2643);
and (n2701,n500,n21);
and (n2702,n2703,n2704);
xor (n2703,n2700,n2701);
and (n2704,n2705,n2706);
xor (n2705,n2648,n2649);
and (n2706,n560,n21);
and (n2707,n20,n75);
or (n2708,n2709,n2712);
and (n2709,n2710,n2711);
xor (n2710,n2657,n2658);
and (n2711,n92,n75);
and (n2712,n2713,n2714);
xor (n2713,n2710,n2711);
or (n2714,n2715,n2718);
and (n2715,n2716,n2717);
xor (n2716,n2662,n2663);
and (n2717,n86,n75);
and (n2718,n2719,n2720);
xor (n2719,n2716,n2717);
or (n2720,n2721,n2724);
and (n2721,n2722,n2723);
xor (n2722,n2667,n2668);
and (n2723,n189,n75);
and (n2724,n2725,n2726);
xor (n2725,n2722,n2723);
or (n2726,n2727,n2730);
and (n2727,n2728,n2729);
xor (n2728,n2673,n2674);
and (n2729,n221,n75);
and (n2730,n2731,n2732);
xor (n2731,n2728,n2729);
or (n2732,n2733,n2736);
and (n2733,n2734,n2735);
xor (n2734,n2679,n2680);
and (n2735,n280,n75);
and (n2736,n2737,n2738);
xor (n2737,n2734,n2735);
or (n2738,n2739,n2742);
and (n2739,n2740,n2741);
xor (n2740,n2685,n2686);
and (n2741,n332,n75);
and (n2742,n2743,n2744);
xor (n2743,n2740,n2741);
or (n2744,n2745,n2748);
and (n2745,n2746,n2747);
xor (n2746,n2691,n2692);
and (n2747,n431,n75);
and (n2748,n2749,n2750);
xor (n2749,n2746,n2747);
or (n2750,n2751,n2754);
and (n2751,n2752,n2753);
xor (n2752,n2697,n2698);
and (n2753,n500,n75);
and (n2754,n2755,n2756);
xor (n2755,n2752,n2753);
and (n2756,n2757,n2758);
xor (n2757,n2703,n2704);
not (n2758,n1382);
and (n2759,n92,n80);
or (n2760,n2761,n2763);
and (n2761,n2762,n87);
xor (n2762,n2713,n2714);
and (n2763,n2764,n2765);
xor (n2764,n2762,n87);
or (n2765,n2766,n2768);
and (n2766,n2767,n275);
xor (n2767,n2719,n2720);
and (n2768,n2769,n2770);
xor (n2769,n2767,n275);
or (n2770,n2771,n2773);
and (n2771,n2772,n370);
xor (n2772,n2725,n2726);
and (n2773,n2774,n2775);
xor (n2774,n2772,n370);
or (n2775,n2776,n2778);
and (n2776,n2777,n467);
xor (n2777,n2731,n2732);
and (n2778,n2779,n2780);
xor (n2779,n2777,n467);
or (n2780,n2781,n2784);
and (n2781,n2782,n2783);
xor (n2782,n2737,n2738);
and (n2783,n332,n80);
and (n2784,n2785,n2786);
xor (n2785,n2782,n2783);
or (n2786,n2787,n2790);
and (n2787,n2788,n2789);
xor (n2788,n2743,n2744);
and (n2789,n431,n80);
and (n2790,n2791,n2792);
xor (n2791,n2788,n2789);
or (n2792,n2793,n2795);
and (n2793,n2794,n720);
xor (n2794,n2749,n2750);
and (n2795,n2796,n2797);
xor (n2796,n2794,n720);
and (n2797,n2798,n2799);
xor (n2798,n2755,n2756);
and (n2799,n560,n80);
and (n2800,n86,n194);
or (n2801,n2802,n2805);
and (n2802,n2803,n2804);
xor (n2803,n2764,n2765);
and (n2804,n189,n194);
and (n2805,n2806,n2807);
xor (n2806,n2803,n2804);
or (n2807,n2808,n2811);
and (n2808,n2809,n2810);
xor (n2809,n2769,n2770);
and (n2810,n221,n194);
and (n2811,n2812,n2813);
xor (n2812,n2809,n2810);
or (n2813,n2814,n2817);
and (n2814,n2815,n2816);
xor (n2815,n2774,n2775);
and (n2816,n280,n194);
and (n2817,n2818,n2819);
xor (n2818,n2815,n2816);
or (n2819,n2820,n2823);
and (n2820,n2821,n2822);
xor (n2821,n2779,n2780);
and (n2822,n332,n194);
and (n2823,n2824,n2825);
xor (n2824,n2821,n2822);
or (n2825,n2826,n2829);
and (n2826,n2827,n2828);
xor (n2827,n2785,n2786);
and (n2828,n431,n194);
and (n2829,n2830,n2831);
xor (n2830,n2827,n2828);
or (n2831,n2832,n2835);
and (n2832,n2833,n2834);
xor (n2833,n2791,n2792);
and (n2834,n500,n194);
and (n2835,n2836,n2837);
xor (n2836,n2833,n2834);
and (n2837,n2838,n2839);
xor (n2838,n2796,n2797);
and (n2839,n560,n194);
endmodule
