module top (out,n18,n19,n25,n30,n36,n43,n44,n53,n54
        ,n62,n71,n78,n84,n93,n99,n103,n110,n130,n170
        ,n184);
output out;
input n18;
input n19;
input n25;
input n30;
input n36;
input n43;
input n44;
input n53;
input n54;
input n62;
input n71;
input n78;
input n84;
input n93;
input n99;
input n103;
input n110;
input n130;
input n170;
input n184;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
xor (out,n0,n388);
nand (n0,n1,n387);
or (n1,n2,n217);
not (n2,n3);
nand (n3,n4,n216);
nand (n4,n5,n153);
not (n5,n6);
or (n6,n7,n152);
and (n7,n8,n122);
xor (n8,n9,n88);
or (n9,n10,n87);
and (n10,n11,n65);
xor (n11,n12,n38);
nand (n12,n13,n32);
or (n13,n14,n27);
nand (n14,n15,n22);
nor (n15,n16,n20);
and (n16,n17,n19);
not (n17,n18);
and (n20,n18,n21);
not (n21,n19);
nand (n22,n23,n26);
or (n23,n19,n24);
not (n24,n25);
nand (n26,n24,n19);
nor (n27,n28,n31);
and (n28,n29,n25);
not (n29,n30);
and (n31,n30,n24);
or (n32,n33,n15);
or (n33,n34,n37);
and (n34,n35,n24);
not (n35,n36);
and (n37,n36,n25);
nand (n38,n39,n59);
or (n39,n40,n48);
not (n40,n41);
nor (n41,n42,n45);
and (n42,n43,n44);
and (n45,n46,n47);
not (n46,n43);
not (n47,n44);
nand (n48,n49,n56);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n54);
not (n52,n53);
nand (n55,n52,n54);
nand (n56,n57,n58);
or (n57,n52,n44);
nand (n58,n44,n52);
or (n59,n49,n60);
nor (n60,n61,n63);
and (n61,n47,n62);
and (n63,n44,n64);
not (n64,n62);
nand (n65,n66,n81);
or (n66,n67,n76);
nand (n67,n68,n73);
nor (n68,n69,n72);
and (n69,n70,n44);
not (n70,n71);
and (n72,n71,n47);
nand (n73,n74,n75);
or (n74,n71,n17);
nand (n75,n17,n71);
nor (n76,n77,n79);
and (n77,n78,n17);
and (n79,n18,n80);
not (n80,n78);
or (n81,n68,n82);
nor (n82,n83,n85);
and (n83,n84,n17);
and (n85,n18,n86);
not (n86,n84);
and (n87,n12,n38);
xor (n88,n89,n114);
xor (n89,n90,n96);
nor (n90,n91,n29);
nor (n91,n92,n94);
and (n92,n24,n93);
and (n94,n25,n95);
not (n95,n93);
nand (n96,n97,n107);
or (n97,n98,n100);
not (n98,n99);
not (n100,n101);
nor (n101,n102,n104);
and (n102,n103,n54);
and (n104,n105,n106);
not (n105,n103);
not (n106,n54);
or (n107,n108,n113);
nor (n108,n109,n111);
and (n109,n110,n106);
and (n111,n112,n54);
not (n112,n110);
nand (n113,n98,n54);
nand (n114,n115,n119);
or (n115,n15,n116);
nor (n116,n117,n118);
and (n117,n78,n24);
and (n118,n80,n25);
nand (n119,n120,n121);
not (n120,n33);
not (n121,n14);
xor (n122,n123,n138);
xor (n123,n124,n132);
nand (n124,n125,n126);
or (n125,n48,n60);
or (n126,n49,n127);
nor (n127,n128,n131);
and (n128,n129,n44);
not (n129,n130);
and (n131,n130,n47);
nand (n132,n133,n134);
or (n133,n67,n82);
or (n134,n68,n135);
nor (n135,n136,n137);
and (n136,n17,n43);
and (n137,n18,n46);
and (n138,n139,n145);
nor (n139,n140,n24);
nor (n140,n141,n144);
and (n141,n142,n17);
not (n142,n143);
and (n143,n30,n19);
and (n144,n29,n21);
nand (n145,n146,n151);
or (n146,n147,n113);
not (n147,n148);
nor (n148,n149,n150);
and (n149,n129,n106);
and (n150,n130,n54);
or (n151,n108,n98);
and (n152,n9,n88);
not (n153,n154);
xor (n154,n155,n190);
xor (n155,n156,n187);
xor (n156,n157,n179);
xor (n157,n158,n164);
nand (n158,n159,n160);
or (n159,n14,n116);
or (n160,n161,n15);
nor (n161,n162,n163);
and (n162,n24,n84);
and (n163,n25,n86);
nand (n164,n165,n175);
or (n165,n166,n172);
nand (n166,n91,n167);
nand (n167,n168,n171);
or (n168,n169,n93);
not (n169,n170);
nand (n171,n169,n93);
nor (n172,n173,n174);
and (n173,n29,n170);
and (n174,n30,n169);
or (n175,n176,n91);
nor (n176,n177,n178);
and (n177,n36,n169);
and (n178,n35,n170);
nand (n179,n180,n181);
or (n180,n113,n100);
or (n181,n182,n98);
nor (n182,n183,n185);
and (n183,n184,n106);
and (n185,n186,n54);
not (n186,n184);
or (n187,n188,n189);
and (n188,n123,n138);
and (n189,n124,n132);
xor (n190,n191,n213);
xor (n191,n192,n198);
nand (n192,n193,n194);
or (n193,n67,n135);
or (n194,n68,n195);
nor (n195,n196,n197);
and (n196,n17,n62);
and (n197,n18,n64);
xor (n198,n199,n204);
nor (n199,n200,n169);
nor (n200,n201,n203);
and (n201,n202,n24);
nand (n202,n30,n93);
and (n203,n29,n95);
nand (n204,n205,n210);
or (n205,n49,n206);
not (n206,n207);
nand (n207,n208,n209);
or (n208,n44,n112);
or (n209,n47,n110);
nand (n210,n211,n212);
not (n211,n127);
not (n212,n48);
or (n213,n214,n215);
and (n214,n89,n114);
and (n215,n90,n96);
nand (n216,n154,n6);
not (n217,n218);
nand (n218,n219,n386);
or (n219,n220,n381);
not (n220,n221);
or (n221,n222,n380);
and (n222,n223,n272);
xor (n223,n224,n265);
or (n224,n225,n264);
and (n225,n226,n250);
xor (n226,n227,n233);
nand (n227,n228,n232);
or (n228,n67,n229);
nor (n229,n230,n231);
and (n230,n17,n36);
and (n231,n18,n35);
or (n232,n76,n68);
and (n233,n234,n240);
and (n234,n235,n18);
nand (n235,n236,n237);
or (n236,n30,n71);
nand (n237,n238,n47);
not (n238,n239);
and (n239,n30,n71);
nand (n240,n241,n246);
or (n241,n98,n242);
not (n242,n243);
nor (n243,n244,n245);
and (n244,n64,n106);
and (n245,n62,n54);
or (n246,n247,n113);
nor (n247,n248,n249);
and (n248,n106,n43);
and (n249,n54,n46);
xor (n250,n251,n257);
xor (n251,n252,n254);
and (n252,n253,n30);
not (n253,n15);
nand (n254,n255,n256);
or (n255,n113,n242);
nand (n256,n148,n99);
nand (n257,n258,n263);
or (n258,n259,n48);
not (n259,n260);
nor (n260,n261,n262);
and (n261,n86,n47);
and (n262,n84,n44);
nand (n263,n41,n50);
and (n264,n227,n233);
xor (n265,n266,n271);
xor (n266,n267,n268);
xor (n267,n139,n145);
or (n268,n269,n270);
and (n269,n251,n257);
and (n270,n252,n254);
xor (n271,n11,n65);
nand (n272,n273,n379);
or (n273,n274,n374);
nor (n274,n275,n373);
and (n275,n276,n352);
nand (n276,n277,n350);
or (n277,n278,n333);
not (n278,n279);
or (n279,n280,n332);
and (n280,n281,n310);
xor (n281,n282,n291);
nand (n282,n283,n287);
or (n283,n48,n284);
nor (n284,n285,n286);
and (n285,n44,n29);
and (n286,n30,n47);
or (n287,n49,n288);
nor (n288,n289,n290);
and (n289,n35,n44);
and (n290,n36,n47);
nand (n291,n292,n309);
or (n292,n293,n299);
not (n293,n294);
nand (n294,n295,n44);
nand (n295,n296,n298);
or (n296,n297,n54);
and (n297,n30,n53);
nand (n298,n29,n52);
not (n299,n300);
nand (n300,n301,n305);
or (n301,n302,n113);
or (n302,n303,n304);
and (n303,n78,n54);
and (n304,n80,n106);
or (n305,n306,n98);
nor (n306,n307,n308);
and (n307,n86,n54);
and (n308,n84,n106);
or (n309,n300,n294);
or (n310,n311,n331);
and (n311,n312,n320);
xor (n312,n313,n314);
nor (n313,n49,n29);
nand (n314,n315,n319);
or (n315,n316,n113);
nor (n316,n317,n318);
and (n317,n35,n54);
and (n318,n36,n106);
or (n319,n302,n98);
nor (n320,n321,n329);
nor (n321,n322,n324);
and (n322,n323,n99);
not (n323,n316);
and (n324,n325,n328);
nand (n325,n326,n327);
or (n326,n29,n54);
nand (n327,n54,n29);
not (n328,n113);
or (n329,n330,n106);
and (n330,n30,n99);
and (n331,n313,n314);
and (n332,n282,n291);
not (n333,n334);
nand (n334,n335,n349);
not (n335,n336);
xor (n336,n337,n346);
xor (n337,n338,n340);
and (n338,n339,n30);
not (n339,n68);
nand (n340,n341,n342);
or (n341,n288,n48);
nand (n342,n343,n50);
nor (n343,n344,n345);
and (n344,n80,n47);
and (n345,n78,n44);
nand (n346,n347,n348);
or (n347,n306,n113);
or (n348,n247,n98);
nand (n349,n293,n300);
nand (n350,n351,n336);
not (n351,n349);
nand (n352,n353,n369);
not (n353,n354);
xor (n354,n355,n368);
xor (n355,n356,n360);
nand (n356,n357,n359);
or (n357,n358,n48);
not (n358,n343);
nand (n359,n260,n50);
nand (n360,n361,n366);
or (n361,n362,n67);
not (n362,n363);
nand (n363,n364,n365);
or (n364,n30,n17);
or (n365,n29,n18);
nand (n366,n367,n339);
not (n367,n229);
xor (n368,n234,n240);
not (n369,n370);
or (n370,n371,n372);
and (n371,n337,n346);
and (n372,n338,n340);
nor (n373,n353,n369);
nor (n374,n375,n376);
xor (n375,n226,n250);
or (n376,n377,n378);
and (n377,n355,n368);
and (n378,n356,n360);
nand (n379,n375,n376);
and (n380,n224,n265);
nor (n381,n382,n383);
xor (n382,n8,n122);
or (n383,n384,n385);
and (n384,n266,n271);
and (n385,n267,n268);
nand (n386,n382,n383);
or (n387,n218,n3);
xor (n388,n389,n595);
xor (n389,n390,n592);
xor (n390,n391,n591);
xor (n391,n392,n583);
xor (n392,n393,n582);
xor (n393,n394,n568);
xor (n394,n395,n567);
xor (n395,n396,n546);
xor (n396,n397,n545);
xor (n397,n398,n519);
xor (n398,n399,n518);
xor (n399,n400,n488);
xor (n400,n401,n487);
xor (n401,n402,n449);
xor (n402,n403,n448);
xor (n403,n404,n406);
xor (n404,n405,n102);
and (n405,n184,n99);
or (n406,n407,n410);
and (n407,n408,n409);
and (n408,n103,n99);
and (n409,n110,n54);
and (n410,n411,n412);
xor (n411,n408,n409);
or (n412,n413,n415);
and (n413,n414,n150);
and (n414,n110,n99);
and (n415,n416,n417);
xor (n416,n414,n150);
or (n417,n418,n420);
and (n418,n419,n245);
and (n419,n130,n99);
and (n420,n421,n422);
xor (n421,n419,n245);
or (n422,n423,n426);
and (n423,n424,n425);
and (n424,n62,n99);
and (n425,n43,n54);
and (n426,n427,n428);
xor (n427,n424,n425);
or (n428,n429,n432);
and (n429,n430,n431);
and (n430,n43,n99);
and (n431,n84,n54);
and (n432,n433,n434);
xor (n433,n430,n431);
or (n434,n435,n437);
and (n435,n436,n303);
and (n436,n84,n99);
and (n437,n438,n439);
xor (n438,n436,n303);
or (n439,n440,n443);
and (n440,n441,n442);
and (n441,n78,n99);
and (n442,n36,n54);
and (n443,n444,n445);
xor (n444,n441,n442);
and (n445,n446,n447);
and (n446,n36,n99);
and (n447,n30,n54);
and (n448,n110,n53);
or (n449,n450,n453);
and (n450,n451,n452);
xor (n451,n411,n412);
and (n452,n130,n53);
and (n453,n454,n455);
xor (n454,n451,n452);
or (n455,n456,n459);
and (n456,n457,n458);
xor (n457,n416,n417);
and (n458,n62,n53);
and (n459,n460,n461);
xor (n460,n457,n458);
or (n461,n462,n465);
and (n462,n463,n464);
xor (n463,n421,n422);
and (n464,n43,n53);
and (n465,n466,n467);
xor (n466,n463,n464);
or (n467,n468,n471);
and (n468,n469,n470);
xor (n469,n427,n428);
and (n470,n84,n53);
and (n471,n472,n473);
xor (n472,n469,n470);
or (n473,n474,n477);
and (n474,n475,n476);
xor (n475,n433,n434);
and (n476,n78,n53);
and (n477,n478,n479);
xor (n478,n475,n476);
or (n479,n480,n483);
and (n480,n481,n482);
xor (n481,n438,n439);
and (n482,n36,n53);
and (n483,n484,n485);
xor (n484,n481,n482);
and (n485,n486,n297);
xor (n486,n444,n445);
and (n487,n130,n44);
or (n488,n489,n492);
and (n489,n490,n491);
xor (n490,n454,n455);
and (n491,n62,n44);
and (n492,n493,n494);
xor (n493,n490,n491);
or (n494,n495,n497);
and (n495,n496,n42);
xor (n496,n460,n461);
and (n497,n498,n499);
xor (n498,n496,n42);
or (n499,n500,n502);
and (n500,n501,n262);
xor (n501,n466,n467);
and (n502,n503,n504);
xor (n503,n501,n262);
or (n504,n505,n507);
and (n505,n506,n345);
xor (n506,n472,n473);
and (n507,n508,n509);
xor (n508,n506,n345);
or (n509,n510,n513);
and (n510,n511,n512);
xor (n511,n478,n479);
and (n512,n36,n44);
and (n513,n514,n515);
xor (n514,n511,n512);
and (n515,n516,n517);
xor (n516,n484,n485);
and (n517,n30,n44);
and (n518,n62,n71);
or (n519,n520,n523);
and (n520,n521,n522);
xor (n521,n493,n494);
and (n522,n43,n71);
and (n523,n524,n525);
xor (n524,n521,n522);
or (n525,n526,n529);
and (n526,n527,n528);
xor (n527,n498,n499);
and (n528,n84,n71);
and (n529,n530,n531);
xor (n530,n527,n528);
or (n531,n532,n535);
and (n532,n533,n534);
xor (n533,n503,n504);
and (n534,n78,n71);
and (n535,n536,n537);
xor (n536,n533,n534);
or (n537,n538,n541);
and (n538,n539,n540);
xor (n539,n508,n509);
and (n540,n36,n71);
and (n541,n542,n543);
xor (n542,n539,n540);
and (n543,n544,n239);
xor (n544,n514,n515);
and (n545,n43,n18);
or (n546,n547,n550);
and (n547,n548,n549);
xor (n548,n524,n525);
and (n549,n84,n18);
and (n550,n551,n552);
xor (n551,n548,n549);
or (n552,n553,n556);
and (n553,n554,n555);
xor (n554,n530,n531);
and (n555,n78,n18);
and (n556,n557,n558);
xor (n557,n554,n555);
or (n558,n559,n562);
and (n559,n560,n561);
xor (n560,n536,n537);
and (n561,n36,n18);
and (n562,n563,n564);
xor (n563,n560,n561);
and (n564,n565,n566);
xor (n565,n542,n543);
and (n566,n30,n18);
and (n567,n84,n19);
or (n568,n569,n572);
and (n569,n570,n571);
xor (n570,n551,n552);
and (n571,n78,n19);
and (n572,n573,n574);
xor (n573,n570,n571);
or (n574,n575,n578);
and (n575,n576,n577);
xor (n576,n557,n558);
and (n577,n36,n19);
and (n578,n579,n580);
xor (n579,n576,n577);
and (n580,n581,n143);
xor (n581,n563,n564);
and (n582,n78,n25);
or (n583,n584,n586);
and (n584,n585,n37);
xor (n585,n573,n574);
and (n586,n587,n588);
xor (n587,n585,n37);
and (n588,n589,n590);
xor (n589,n579,n580);
and (n590,n30,n25);
and (n591,n36,n93);
and (n592,n593,n594);
xor (n593,n587,n588);
not (n594,n202);
and (n595,n30,n170);
endmodule
