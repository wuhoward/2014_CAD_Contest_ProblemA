module top (out,n13,n16,n17,n21,n24,n25,n35,n38,n39
        ,n43,n53,n56,n57,n61,n68,n71,n72,n76,n84
        ,n87,n88,n92,n102,n105,n106,n110,n115,n310,n372
        ,n466,n539,n624);
output out;
input n13;
input n16;
input n17;
input n21;
input n24;
input n25;
input n35;
input n38;
input n39;
input n43;
input n53;
input n56;
input n57;
input n61;
input n68;
input n71;
input n72;
input n76;
input n84;
input n87;
input n88;
input n92;
input n102;
input n105;
input n106;
input n110;
input n115;
input n310;
input n372;
input n466;
input n539;
input n624;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
xor (out,n0,n1281);
xor (n0,n1,n334);
xor (n1,n2,n268);
xor (n2,n3,n227);
or (n3,n4,n205,n226);
and (n4,n5,n176);
or (n5,n6,n147,n175);
and (n6,n7,n117);
or (n7,n8,n97,n116);
and (n8,n9,n48);
or (n9,n10,n31,n47);
and (n10,n11,n18);
not (n11,n12);
and (n12,n13,n14);
not (n14,n15);
and (n15,n16,n17);
xnor (n18,n19,n28);
not (n19,n20);
and (n20,n21,n22);
and (n22,n23,n26);
xor (n23,n24,n25);
not (n26,n27);
xor (n27,n25,n13);
and (n28,n24,n29);
not (n29,n30);
and (n30,n25,n13);
and (n31,n18,n32);
xnor (n32,n33,n44);
nor (n33,n34,n42);
and (n34,n35,n36);
and (n36,n37,n40);
xor (n37,n38,n39);
not (n40,n41);
xor (n41,n39,n24);
and (n42,n43,n41);
and (n44,n38,n45);
not (n45,n46);
and (n46,n39,n24);
and (n47,n11,n32);
or (n48,n49,n80,n96);
and (n49,n50,n65);
xnor (n50,n51,n62);
nor (n51,n52,n60);
and (n52,n53,n54);
and (n54,n55,n58);
xor (n55,n56,n57);
not (n58,n59);
xor (n59,n57,n38);
and (n60,n61,n59);
and (n62,n56,n63);
not (n63,n64);
and (n64,n57,n38);
xnor (n65,n66,n77);
nor (n66,n67,n75);
and (n67,n68,n69);
and (n69,n70,n73);
xor (n70,n71,n72);
not (n73,n74);
xor (n74,n72,n56);
and (n75,n76,n74);
and (n77,n71,n78);
not (n78,n79);
and (n79,n72,n56);
and (n80,n65,n81);
xnor (n81,n82,n93);
nor (n82,n83,n91);
and (n83,n84,n85);
and (n85,n86,n89);
xor (n86,n87,n88);
not (n89,n90);
xor (n90,n88,n71);
and (n91,n92,n90);
and (n93,n87,n94);
not (n94,n95);
and (n95,n88,n71);
and (n96,n50,n81);
and (n97,n48,n98);
and (n98,n99,n114);
xnor (n99,n100,n111);
nor (n100,n101,n109);
and (n101,n102,n103);
and (n103,n104,n107);
xor (n104,n105,n106);
not (n107,n108);
xor (n108,n106,n87);
and (n109,n110,n108);
and (n111,n105,n112);
not (n112,n113);
and (n113,n106,n87);
and (n114,n115,n105);
and (n116,n9,n98);
or (n117,n118,n143,n146);
and (n118,n119,n129);
xor (n119,n120,n125);
xor (n120,n28,n121);
xnor (n121,n122,n44);
nor (n122,n123,n124);
and (n123,n43,n36);
and (n124,n21,n41);
xnor (n125,n126,n62);
nor (n126,n127,n128);
and (n127,n61,n54);
and (n128,n35,n59);
xor (n129,n130,n139);
xor (n130,n131,n135);
xnor (n131,n132,n77);
nor (n132,n133,n134);
and (n133,n76,n69);
and (n134,n53,n74);
xnor (n135,n136,n93);
nor (n136,n137,n138);
and (n137,n92,n85);
and (n138,n68,n90);
xnor (n139,n140,n111);
nor (n140,n141,n142);
and (n141,n110,n103);
and (n142,n84,n108);
and (n143,n129,n144);
not (n144,n145);
and (n145,n102,n105);
and (n146,n119,n144);
and (n147,n117,n148);
xor (n148,n149,n165);
xor (n149,n150,n151);
and (n150,n110,n105);
xor (n151,n152,n161);
xor (n152,n153,n157);
xnor (n153,n154,n77);
nor (n154,n155,n156);
and (n155,n53,n69);
and (n156,n61,n74);
xnor (n157,n158,n93);
nor (n158,n159,n160);
and (n159,n68,n85);
and (n160,n76,n90);
xnor (n161,n162,n111);
nor (n162,n163,n164);
and (n163,n84,n103);
and (n164,n92,n108);
xor (n165,n166,n171);
xor (n166,n167,n168);
not (n167,n28);
xnor (n168,n169,n44);
not (n169,n170);
and (n170,n21,n36);
xnor (n171,n172,n62);
nor (n172,n173,n174);
and (n173,n35,n54);
and (n174,n43,n59);
and (n175,n7,n148);
xor (n176,n177,n194);
xor (n177,n178,n190);
or (n178,n179,n188,n189);
and (n179,n180,n184);
or (n180,n181,n182,n183);
and (n181,n28,n121);
and (n182,n121,n125);
and (n183,n28,n125);
or (n184,n185,n186,n187);
and (n185,n131,n135);
and (n186,n135,n139);
and (n187,n131,n139);
and (n188,n184,n145);
and (n189,n180,n145);
or (n190,n191,n192,n193);
and (n191,n150,n151);
and (n192,n151,n165);
and (n193,n150,n165);
xor (n194,n195,n204);
xor (n195,n196,n200);
xnor (n196,n197,n93);
nor (n197,n198,n199);
and (n198,n76,n85);
and (n199,n53,n90);
xnor (n200,n201,n111);
nor (n201,n202,n203);
and (n202,n92,n103);
and (n203,n68,n108);
and (n204,n84,n105);
and (n205,n176,n206);
xor (n206,n207,n217);
xor (n207,n208,n213);
xor (n208,n44,n209);
xnor (n209,n210,n62);
nor (n210,n211,n212);
and (n211,n43,n54);
and (n212,n21,n59);
xnor (n213,n214,n77);
nor (n214,n215,n216);
and (n215,n61,n69);
and (n216,n35,n74);
xnor (n217,n218,n222);
or (n218,n219,n220,n221);
and (n219,n153,n157);
and (n220,n157,n161);
and (n221,n153,n161);
or (n222,n223,n224,n225);
and (n223,n167,n168);
and (n224,n168,n171);
and (n225,n167,n171);
and (n226,n5,n206);
xor (n227,n228,n234);
xor (n228,n229,n233);
or (n229,n230,n231,n232);
and (n230,n178,n190);
and (n231,n190,n194);
and (n232,n178,n194);
and (n233,n207,n217);
xor (n234,n235,n247);
xor (n235,n236,n237);
or (n236,n218,n222);
xor (n237,n238,n243);
xor (n238,n239,n240);
not (n239,n44);
xnor (n240,n241,n62);
not (n241,n242);
and (n242,n21,n54);
xnor (n243,n244,n77);
nor (n244,n245,n246);
and (n245,n35,n69);
and (n246,n43,n74);
xor (n247,n248,n257);
xor (n248,n249,n253);
or (n249,n250,n251,n252);
and (n250,n196,n200);
and (n251,n200,n204);
and (n252,n196,n204);
or (n253,n254,n255,n256);
and (n254,n44,n209);
and (n255,n209,n213);
and (n256,n44,n213);
xor (n257,n258,n267);
xor (n258,n259,n263);
xnor (n259,n260,n93);
nor (n260,n261,n262);
and (n261,n53,n85);
and (n262,n61,n90);
xnor (n263,n264,n111);
nor (n264,n265,n266);
and (n265,n68,n103);
and (n266,n76,n108);
and (n267,n92,n105);
and (n268,n269,n332);
or (n269,n270,n328,n331);
and (n270,n271,n326);
or (n271,n272,n321,n325);
and (n272,n273,n312);
or (n273,n274,n303,n311);
and (n274,n275,n287);
or (n275,n276,n281,n286);
and (n276,n12,n277);
xnor (n277,n278,n28);
nor (n278,n279,n280);
and (n279,n43,n22);
and (n280,n21,n27);
and (n281,n277,n282);
xnor (n282,n283,n44);
nor (n283,n284,n285);
and (n284,n61,n36);
and (n285,n35,n41);
and (n286,n12,n282);
or (n287,n288,n297,n302);
and (n288,n289,n293);
xnor (n289,n290,n62);
nor (n290,n291,n292);
and (n291,n76,n54);
and (n292,n53,n59);
xnor (n293,n294,n77);
nor (n294,n295,n296);
and (n295,n92,n69);
and (n296,n68,n74);
and (n297,n293,n298);
xnor (n298,n299,n93);
nor (n299,n300,n301);
and (n300,n110,n85);
and (n301,n84,n90);
and (n302,n289,n298);
and (n303,n287,n304);
or (n304,n305,n309);
xnor (n305,n306,n111);
nor (n306,n307,n308);
and (n307,n115,n103);
and (n308,n102,n108);
and (n309,n310,n105);
and (n311,n275,n304);
or (n312,n313,n318,n320);
and (n313,n314,n316);
xor (n314,n315,n32);
xor (n315,n11,n18);
xor (n316,n317,n81);
xor (n317,n50,n65);
and (n318,n316,n319);
xor (n319,n99,n114);
and (n320,n314,n319);
and (n321,n312,n322);
xor (n322,n323,n129);
xor (n323,n145,n324);
not (n324,n119);
and (n325,n273,n322);
xor (n326,n327,n145);
xor (n327,n180,n184);
and (n328,n326,n329);
xor (n329,n330,n148);
xor (n330,n7,n117);
and (n331,n271,n329);
xor (n332,n333,n206);
xor (n333,n5,n176);
or (n334,n335,n413);
and (n335,n336,n337);
xor (n336,n269,n332);
and (n337,n338,n411);
or (n338,n339,n407,n410);
and (n339,n340,n405);
or (n340,n341,n401,n404);
and (n341,n342,n392);
or (n342,n343,n374,n391);
and (n343,n344,n360);
or (n344,n345,n354,n359);
and (n345,n346,n347);
not (n346,n17);
xnor (n347,n348,n12);
not (n348,n349);
and (n349,n21,n350);
and (n350,n351,n352);
xor (n351,n13,n16);
not (n352,n353);
xor (n353,n16,n17);
and (n354,n347,n355);
xnor (n355,n356,n28);
nor (n356,n357,n358);
and (n357,n35,n22);
and (n358,n43,n27);
and (n359,n346,n355);
or (n360,n361,n370,n373);
and (n361,n362,n366);
xnor (n362,n363,n93);
nor (n363,n364,n365);
and (n364,n102,n85);
and (n365,n110,n90);
xnor (n366,n367,n111);
nor (n367,n368,n369);
and (n368,n310,n103);
and (n369,n115,n108);
and (n370,n366,n371);
and (n371,n372,n105);
and (n373,n362,n371);
and (n374,n360,n375);
or (n375,n376,n385,n390);
and (n376,n377,n381);
xnor (n377,n378,n44);
nor (n378,n379,n380);
and (n379,n53,n36);
and (n380,n61,n41);
xnor (n381,n382,n62);
nor (n382,n383,n384);
and (n383,n68,n54);
and (n384,n76,n59);
and (n385,n381,n386);
xnor (n386,n387,n77);
nor (n387,n388,n389);
and (n388,n84,n69);
and (n389,n92,n74);
and (n390,n377,n386);
and (n391,n344,n375);
or (n392,n393,n398,n400);
and (n393,n394,n396);
xor (n394,n395,n282);
xor (n395,n12,n277);
xor (n396,n397,n298);
xor (n397,n289,n293);
and (n398,n396,n399);
xnor (n399,n305,n309);
and (n400,n394,n399);
and (n401,n392,n402);
xor (n402,n403,n319);
xor (n403,n314,n316);
and (n404,n342,n402);
xor (n405,n406,n98);
xor (n406,n9,n48);
and (n407,n405,n408);
xor (n408,n409,n322);
xor (n409,n273,n312);
and (n410,n340,n408);
xor (n411,n412,n329);
xor (n412,n271,n326);
and (n413,n414,n415);
xor (n414,n336,n337);
or (n415,n416,n488);
and (n416,n417,n418);
xor (n417,n338,n411);
and (n418,n419,n486);
or (n419,n420,n482,n485);
and (n420,n421,n480);
or (n421,n422,n474,n479);
and (n422,n423,n469);
or (n423,n424,n453,n468);
and (n424,n425,n441);
or (n425,n426,n435,n440);
and (n426,n427,n431);
xnor (n427,n428,n44);
nor (n428,n429,n430);
and (n429,n76,n36);
and (n430,n53,n41);
xnor (n431,n432,n62);
nor (n432,n433,n434);
and (n433,n92,n54);
and (n434,n68,n59);
and (n435,n431,n436);
xnor (n436,n437,n77);
nor (n437,n438,n439);
and (n438,n110,n69);
and (n439,n84,n74);
and (n440,n427,n436);
or (n441,n442,n447,n452);
and (n442,n17,n443);
xnor (n443,n444,n12);
nor (n444,n445,n446);
and (n445,n43,n350);
and (n446,n21,n353);
and (n447,n443,n448);
xnor (n448,n449,n28);
nor (n449,n450,n451);
and (n450,n61,n22);
and (n451,n35,n27);
and (n452,n17,n448);
and (n453,n441,n454);
or (n454,n455,n464,n467);
and (n455,n456,n460);
xnor (n456,n457,n93);
nor (n457,n458,n459);
and (n458,n115,n85);
and (n459,n102,n90);
xnor (n460,n461,n111);
nor (n461,n462,n463);
and (n462,n372,n103);
and (n463,n310,n108);
and (n464,n460,n465);
and (n465,n466,n105);
and (n467,n456,n465);
and (n468,n425,n454);
or (n469,n470,n472);
xor (n470,n471,n371);
xor (n471,n362,n366);
xor (n472,n473,n386);
xor (n473,n377,n381);
and (n474,n469,n475);
xor (n475,n476,n478);
xor (n476,n477,n396);
not (n477,n394);
not (n478,n399);
and (n479,n423,n475);
xor (n480,n481,n304);
xor (n481,n275,n287);
and (n482,n480,n483);
xor (n483,n484,n402);
xor (n484,n342,n392);
and (n485,n421,n483);
xor (n486,n487,n408);
xor (n487,n340,n405);
and (n488,n489,n490);
xor (n489,n417,n418);
or (n490,n491,n570);
and (n491,n492,n493);
xor (n492,n419,n486);
and (n493,n494,n568);
or (n494,n495,n564,n567);
and (n495,n496,n560);
or (n496,n497,n556,n559);
and (n497,n498,n546);
or (n498,n499,n532,n545);
and (n499,n500,n516);
or (n500,n501,n510,n515);
and (n501,n502,n506);
xnor (n502,n503,n28);
nor (n503,n504,n505);
and (n504,n53,n22);
and (n505,n61,n27);
xnor (n506,n507,n44);
nor (n507,n508,n509);
and (n508,n68,n36);
and (n509,n76,n41);
and (n510,n506,n511);
xnor (n511,n512,n62);
nor (n512,n513,n514);
and (n513,n84,n54);
and (n514,n92,n59);
and (n515,n502,n511);
or (n516,n517,n526,n531);
and (n517,n518,n522);
xnor (n518,n519,n77);
nor (n519,n520,n521);
and (n520,n102,n69);
and (n521,n110,n74);
xnor (n522,n523,n93);
nor (n523,n524,n525);
and (n524,n310,n85);
and (n525,n115,n90);
and (n526,n522,n527);
xnor (n527,n528,n111);
nor (n528,n529,n530);
and (n529,n466,n103);
and (n530,n372,n108);
and (n531,n518,n527);
and (n532,n516,n533);
and (n533,n534,n541);
xnor (n534,n535,n17);
not (n535,n536);
and (n536,n21,n537);
and (n537,n538,n540);
xor (n538,n17,n539);
not (n540,n539);
xnor (n541,n542,n12);
nor (n542,n543,n544);
and (n543,n35,n350);
and (n544,n43,n353);
and (n545,n500,n533);
or (n546,n547,n552,n555);
and (n547,n548,n550);
xor (n548,n549,n436);
xor (n549,n427,n431);
xor (n550,n551,n448);
xor (n551,n17,n443);
and (n552,n550,n553);
xor (n553,n554,n465);
xor (n554,n456,n460);
and (n555,n548,n553);
and (n556,n546,n557);
xor (n557,n558,n355);
xor (n558,n346,n347);
and (n559,n498,n557);
and (n560,n561,n563);
xor (n561,n562,n454);
xor (n562,n425,n441);
xnor (n563,n470,n472);
and (n564,n560,n565);
xor (n565,n566,n375);
xor (n566,n344,n360);
and (n567,n496,n565);
xor (n568,n569,n483);
xor (n569,n421,n480);
and (n570,n571,n572);
xor (n571,n492,n493);
or (n572,n573,n652);
and (n573,n574,n575);
xor (n574,n494,n568);
or (n575,n576,n648,n651);
and (n576,n577,n646);
or (n577,n578,n643,n645);
and (n578,n579,n641);
or (n579,n580,n637,n640);
and (n580,n581,n627);
or (n581,n582,n615,n626);
and (n582,n583,n599);
or (n583,n584,n593,n598);
and (n584,n585,n589);
xnor (n585,n586,n17);
nor (n586,n587,n588);
and (n587,n43,n537);
and (n588,n21,n539);
xnor (n589,n590,n12);
nor (n590,n591,n592);
and (n591,n61,n350);
and (n592,n35,n353);
and (n593,n589,n594);
xnor (n594,n595,n28);
nor (n595,n596,n597);
and (n596,n76,n22);
and (n597,n53,n27);
and (n598,n585,n594);
or (n599,n600,n609,n614);
and (n600,n601,n605);
xnor (n601,n602,n44);
nor (n602,n603,n604);
and (n603,n92,n36);
and (n604,n68,n41);
xnor (n605,n606,n62);
nor (n606,n607,n608);
and (n607,n110,n54);
and (n608,n84,n59);
and (n609,n605,n610);
xnor (n610,n611,n77);
nor (n611,n612,n613);
and (n612,n115,n69);
and (n613,n102,n74);
and (n614,n601,n610);
and (n615,n599,n616);
and (n616,n617,n621);
xnor (n617,n618,n93);
nor (n618,n619,n620);
and (n619,n372,n85);
and (n620,n310,n90);
xnor (n621,n622,n111);
nor (n622,n623,n625);
and (n623,n624,n103);
and (n625,n466,n108);
and (n626,n583,n616);
or (n627,n628,n633,n636);
and (n628,n629,n631);
not (n629,n630);
nand (n630,n624,n105);
xor (n631,n632,n511);
xor (n632,n502,n506);
and (n633,n631,n634);
xor (n634,n635,n527);
xor (n635,n518,n522);
and (n636,n629,n634);
and (n637,n627,n638);
xor (n638,n639,n553);
xor (n639,n548,n550);
and (n640,n581,n638);
xor (n641,n642,n557);
xor (n642,n498,n546);
and (n643,n641,n644);
xor (n644,n561,n563);
and (n645,n579,n644);
xor (n646,n647,n565);
xor (n647,n496,n560);
and (n648,n646,n649);
xor (n649,n650,n475);
xor (n650,n423,n469);
and (n651,n577,n649);
and (n652,n653,n654);
xor (n653,n574,n575);
or (n654,n655,n732);
and (n655,n656,n658);
xor (n656,n657,n649);
xor (n657,n577,n646);
and (n658,n659,n730);
or (n659,n660,n726,n729);
and (n660,n661,n721);
or (n661,n662,n718,n720);
and (n662,n663,n709);
or (n663,n664,n691,n708);
and (n664,n665,n679);
or (n665,n666,n675,n678);
and (n666,n667,n671);
xnor (n667,n668,n77);
nor (n668,n669,n670);
and (n669,n310,n69);
and (n670,n115,n74);
xnor (n671,n672,n93);
nor (n672,n673,n674);
and (n673,n466,n85);
and (n674,n372,n90);
and (n675,n671,n676);
xnor (n676,n677,n111);
nand (n677,n624,n108);
and (n678,n667,n676);
or (n679,n680,n689,n690);
and (n680,n681,n685);
xnor (n681,n682,n17);
nor (n682,n683,n684);
and (n683,n35,n537);
and (n684,n43,n539);
xnor (n685,n686,n12);
nor (n686,n687,n688);
and (n687,n53,n350);
and (n688,n61,n353);
and (n689,n685,n111);
and (n690,n681,n111);
and (n691,n679,n692);
or (n692,n693,n702,n707);
and (n693,n694,n698);
xnor (n694,n695,n28);
nor (n695,n696,n697);
and (n696,n68,n22);
and (n697,n76,n27);
xnor (n698,n699,n44);
nor (n699,n700,n701);
and (n700,n84,n36);
and (n701,n92,n41);
and (n702,n698,n703);
xnor (n703,n704,n62);
nor (n704,n705,n706);
and (n705,n102,n54);
and (n706,n110,n59);
and (n707,n694,n703);
and (n708,n665,n692);
or (n709,n710,n715,n717);
and (n710,n711,n713);
xor (n711,n712,n594);
xor (n712,n585,n589);
xor (n713,n714,n610);
xor (n714,n601,n605);
and (n715,n713,n716);
xor (n716,n617,n621);
and (n717,n711,n716);
and (n718,n709,n719);
xor (n719,n534,n541);
and (n720,n663,n719);
and (n721,n722,n724);
xor (n722,n723,n616);
xor (n723,n583,n599);
xor (n724,n725,n634);
xor (n725,n629,n631);
and (n726,n721,n727);
xor (n727,n728,n533);
xor (n728,n500,n516);
and (n729,n661,n727);
xor (n730,n731,n644);
xor (n731,n579,n641);
and (n732,n733,n734);
xor (n733,n656,n658);
or (n734,n735,n742);
and (n735,n736,n737);
xor (n736,n659,n730);
and (n737,n738,n740);
xor (n738,n739,n727);
xor (n739,n661,n721);
xor (n740,n741,n638);
xor (n741,n581,n627);
and (n742,n743,n744);
xor (n743,n736,n737);
or (n744,n745,n808);
and (n745,n746,n752);
xor (n746,n747,n750);
xor (n747,n727,n748);
xor (n748,n741,n749);
not (n749,n550);
xor (n750,n739,n751);
xnor (n751,n548,n553);
or (n752,n753,n805,n807);
and (n753,n754,n803);
or (n754,n755,n799,n802);
and (n755,n756,n794);
or (n756,n757,n790,n793);
and (n757,n758,n774);
or (n758,n759,n768,n773);
and (n759,n760,n764);
xnor (n760,n761,n17);
nor (n761,n762,n763);
and (n762,n61,n537);
and (n763,n35,n539);
xnor (n764,n765,n12);
nor (n765,n766,n767);
and (n766,n76,n350);
and (n767,n53,n353);
and (n768,n764,n769);
xnor (n769,n770,n28);
nor (n770,n771,n772);
and (n771,n92,n22);
and (n772,n68,n27);
and (n773,n760,n769);
or (n774,n775,n784,n789);
and (n775,n776,n780);
xnor (n776,n777,n44);
nor (n777,n778,n779);
and (n778,n110,n36);
and (n779,n84,n41);
xnor (n780,n781,n62);
nor (n781,n782,n783);
and (n782,n115,n54);
and (n783,n102,n59);
and (n784,n780,n785);
xnor (n785,n786,n77);
nor (n786,n787,n788);
and (n787,n372,n69);
and (n788,n310,n74);
and (n789,n776,n785);
and (n790,n774,n791);
xor (n791,n792,n676);
xor (n792,n667,n671);
and (n793,n758,n791);
and (n794,n795,n797);
xor (n795,n796,n111);
xor (n796,n681,n685);
xor (n797,n798,n703);
xor (n798,n694,n698);
and (n799,n794,n800);
xor (n800,n801,n716);
xor (n801,n711,n713);
and (n802,n756,n800);
xor (n803,n804,n719);
xor (n804,n663,n709);
and (n805,n803,n806);
xor (n806,n722,n724);
and (n807,n754,n806);
and (n808,n809,n810);
xor (n809,n746,n752);
or (n810,n811,n865);
and (n811,n812,n814);
xor (n812,n813,n806);
xor (n813,n754,n803);
or (n814,n815,n861,n864);
and (n815,n816,n859);
or (n816,n817,n856,n858);
and (n817,n818,n854);
or (n818,n819,n848,n853);
and (n819,n820,n832);
or (n820,n821,n830,n831);
and (n821,n822,n826);
xnor (n822,n823,n17);
nor (n823,n824,n825);
and (n824,n53,n537);
and (n825,n61,n539);
xnor (n826,n827,n12);
nor (n827,n828,n829);
and (n828,n68,n350);
and (n829,n76,n353);
and (n830,n826,n93);
and (n831,n822,n93);
or (n832,n833,n842,n847);
and (n833,n834,n838);
xnor (n834,n835,n28);
nor (n835,n836,n837);
and (n836,n84,n22);
and (n837,n92,n27);
xnor (n838,n839,n44);
nor (n839,n840,n841);
and (n840,n102,n36);
and (n841,n110,n41);
and (n842,n838,n843);
xnor (n843,n844,n62);
nor (n844,n845,n846);
and (n845,n310,n54);
and (n846,n115,n59);
and (n847,n834,n843);
and (n848,n832,n849);
xnor (n849,n850,n93);
nor (n850,n851,n852);
and (n851,n624,n85);
and (n852,n466,n90);
and (n853,n820,n849);
xor (n854,n855,n791);
xor (n855,n758,n774);
and (n856,n854,n857);
xor (n857,n795,n797);
and (n858,n818,n857);
xor (n859,n860,n692);
xor (n860,n665,n679);
and (n861,n859,n862);
xor (n862,n863,n800);
xor (n863,n756,n794);
and (n864,n816,n862);
and (n865,n866,n867);
xor (n866,n812,n814);
or (n867,n868,n938);
and (n868,n869,n871);
xor (n869,n870,n862);
xor (n870,n816,n859);
or (n871,n872,n934,n937);
and (n872,n873,n929);
or (n873,n874,n925,n928);
and (n874,n875,n915);
or (n875,n876,n909,n914);
and (n876,n877,n893);
or (n877,n878,n887,n892);
and (n878,n879,n883);
xnor (n879,n880,n44);
nor (n880,n881,n882);
and (n881,n115,n36);
and (n882,n102,n41);
xnor (n883,n884,n62);
nor (n884,n885,n886);
and (n885,n372,n54);
and (n886,n310,n59);
and (n887,n883,n888);
xnor (n888,n889,n77);
nor (n889,n890,n891);
and (n890,n624,n69);
and (n891,n466,n74);
and (n892,n879,n888);
or (n893,n894,n903,n908);
and (n894,n895,n899);
xnor (n895,n896,n17);
nor (n896,n897,n898);
and (n897,n76,n537);
and (n898,n53,n539);
xnor (n899,n900,n12);
nor (n900,n901,n902);
and (n901,n92,n350);
and (n902,n68,n353);
and (n903,n899,n904);
xnor (n904,n905,n28);
nor (n905,n906,n907);
and (n906,n110,n22);
and (n907,n84,n27);
and (n908,n895,n904);
and (n909,n893,n910);
xnor (n910,n911,n77);
nor (n911,n912,n913);
and (n912,n466,n69);
and (n913,n372,n74);
and (n914,n877,n910);
or (n915,n916,n921,n924);
and (n916,n917,n919);
xnor (n917,n918,n93);
nand (n918,n624,n90);
xor (n919,n920,n93);
xor (n920,n822,n826);
and (n921,n919,n922);
xor (n922,n923,n843);
xor (n923,n834,n838);
and (n924,n917,n922);
and (n925,n915,n926);
xor (n926,n927,n785);
xor (n927,n776,n780);
and (n928,n875,n926);
and (n929,n930,n932);
xor (n930,n931,n769);
xor (n931,n760,n764);
xor (n932,n933,n849);
xor (n933,n820,n832);
and (n934,n929,n935);
xor (n935,n936,n857);
xor (n936,n818,n854);
and (n937,n873,n935);
and (n938,n939,n940);
xor (n939,n869,n871);
or (n940,n941,n993);
and (n941,n942,n944);
xor (n942,n943,n935);
xor (n943,n873,n929);
or (n944,n945,n990,n992);
and (n945,n946,n988);
or (n946,n947,n984,n987);
and (n947,n948,n982);
or (n948,n949,n978,n981);
and (n949,n950,n966);
or (n950,n951,n960,n965);
and (n951,n952,n956);
xnor (n952,n953,n28);
nor (n953,n954,n955);
and (n954,n102,n22);
and (n955,n110,n27);
xnor (n956,n957,n44);
nor (n957,n958,n959);
and (n958,n310,n36);
and (n959,n115,n41);
and (n960,n956,n961);
xnor (n961,n962,n62);
nor (n962,n963,n964);
and (n963,n466,n54);
and (n964,n372,n59);
and (n965,n952,n961);
or (n966,n967,n976,n977);
and (n967,n968,n972);
xnor (n968,n969,n17);
nor (n969,n970,n971);
and (n970,n68,n537);
and (n971,n76,n539);
xnor (n972,n973,n12);
nor (n973,n974,n975);
and (n974,n84,n350);
and (n975,n92,n353);
and (n976,n972,n77);
and (n977,n968,n77);
and (n978,n966,n979);
xor (n979,n980,n888);
xor (n980,n879,n883);
and (n981,n950,n979);
xor (n982,n983,n910);
xor (n983,n877,n893);
and (n984,n982,n985);
xor (n985,n986,n922);
xor (n986,n917,n919);
and (n987,n948,n985);
xor (n988,n989,n926);
xor (n989,n875,n915);
and (n990,n988,n991);
xor (n991,n930,n932);
and (n992,n946,n991);
and (n993,n994,n995);
xor (n994,n942,n944);
or (n995,n996,n1034);
and (n996,n997,n999);
xor (n997,n998,n991);
xor (n998,n946,n988);
and (n999,n1000,n1032);
or (n1000,n1001,n1028,n1031);
and (n1001,n1002,n1026);
or (n1002,n1003,n1022,n1025);
and (n1003,n1004,n1020);
or (n1004,n1005,n1014,n1019);
and (n1005,n1006,n1010);
xnor (n1006,n1007,n17);
nor (n1007,n1008,n1009);
and (n1008,n92,n537);
and (n1009,n68,n539);
xnor (n1010,n1011,n12);
nor (n1011,n1012,n1013);
and (n1012,n110,n350);
and (n1013,n84,n353);
and (n1014,n1010,n1015);
xnor (n1015,n1016,n28);
nor (n1016,n1017,n1018);
and (n1017,n115,n22);
and (n1018,n102,n27);
and (n1019,n1006,n1015);
xnor (n1020,n1021,n77);
nand (n1021,n624,n74);
and (n1022,n1020,n1023);
xor (n1023,n1024,n961);
xor (n1024,n952,n956);
and (n1025,n1004,n1023);
xor (n1026,n1027,n904);
xor (n1027,n895,n899);
and (n1028,n1026,n1029);
xor (n1029,n1030,n979);
xor (n1030,n950,n966);
and (n1031,n1002,n1029);
xor (n1032,n1033,n985);
xor (n1033,n948,n982);
and (n1034,n1035,n1036);
xor (n1035,n997,n999);
or (n1036,n1037,n1089);
and (n1037,n1038,n1039);
xor (n1038,n1000,n1032);
and (n1039,n1040,n1087);
or (n1040,n1041,n1083,n1086);
and (n1041,n1042,n1076);
or (n1042,n1043,n1070,n1075);
and (n1043,n1044,n1058);
or (n1044,n1045,n1054,n1057);
and (n1045,n1046,n1050);
xnor (n1046,n1047,n28);
nor (n1047,n1048,n1049);
and (n1048,n310,n22);
and (n1049,n115,n27);
xnor (n1050,n1051,n44);
nor (n1051,n1052,n1053);
and (n1052,n466,n36);
and (n1053,n372,n41);
and (n1054,n1050,n1055);
xnor (n1055,n1056,n62);
nand (n1056,n624,n59);
and (n1057,n1046,n1055);
or (n1058,n1059,n1068,n1069);
and (n1059,n1060,n1064);
xnor (n1060,n1061,n17);
nor (n1061,n1062,n1063);
and (n1062,n84,n537);
and (n1063,n92,n539);
xnor (n1064,n1065,n12);
nor (n1065,n1066,n1067);
and (n1066,n102,n350);
and (n1067,n110,n353);
and (n1068,n1064,n62);
and (n1069,n1060,n62);
and (n1070,n1058,n1071);
xnor (n1071,n1072,n44);
nor (n1072,n1073,n1074);
and (n1073,n372,n36);
and (n1074,n310,n41);
and (n1075,n1044,n1071);
and (n1076,n1077,n1081);
xnor (n1077,n1078,n62);
nor (n1078,n1079,n1080);
and (n1079,n624,n54);
and (n1080,n466,n59);
xor (n1081,n1082,n1015);
xor (n1082,n1006,n1010);
and (n1083,n1076,n1084);
xor (n1084,n1085,n77);
xor (n1085,n968,n972);
and (n1086,n1042,n1084);
xor (n1087,n1088,n1029);
xor (n1088,n1002,n1026);
and (n1089,n1090,n1091);
xor (n1090,n1038,n1039);
or (n1091,n1092,n1099);
and (n1092,n1093,n1094);
xor (n1093,n1040,n1087);
and (n1094,n1095,n1097);
xor (n1095,n1096,n1023);
xor (n1096,n1004,n1020);
xor (n1097,n1098,n1084);
xor (n1098,n1042,n1076);
and (n1099,n1100,n1101);
xor (n1100,n1093,n1094);
or (n1101,n1102,n1135);
and (n1102,n1103,n1104);
xor (n1103,n1095,n1097);
or (n1104,n1105,n1132,n1134);
and (n1105,n1106,n1130);
or (n1106,n1107,n1126,n1129);
and (n1107,n1108,n1124);
or (n1108,n1109,n1118,n1123);
and (n1109,n1110,n1114);
xnor (n1110,n1111,n17);
nor (n1111,n1112,n1113);
and (n1112,n110,n537);
and (n1113,n84,n539);
xnor (n1114,n1115,n12);
nor (n1115,n1116,n1117);
and (n1116,n115,n350);
and (n1117,n102,n353);
and (n1118,n1114,n1119);
xnor (n1119,n1120,n28);
nor (n1120,n1121,n1122);
and (n1121,n372,n22);
and (n1122,n310,n27);
and (n1123,n1110,n1119);
xor (n1124,n1125,n1055);
xor (n1125,n1046,n1050);
and (n1126,n1124,n1127);
xor (n1127,n1128,n62);
xor (n1128,n1060,n1064);
and (n1129,n1108,n1127);
xor (n1130,n1131,n1071);
xor (n1131,n1044,n1058);
and (n1132,n1130,n1133);
xor (n1133,n1077,n1081);
and (n1134,n1106,n1133);
and (n1135,n1136,n1137);
xor (n1136,n1103,n1104);
or (n1137,n1138,n1171);
and (n1138,n1139,n1141);
xor (n1139,n1140,n1133);
xor (n1140,n1106,n1130);
and (n1141,n1142,n1169);
or (n1142,n1143,n1163,n1168);
and (n1143,n1144,n1156);
or (n1144,n1145,n1154,n1155);
and (n1145,n1146,n1150);
xnor (n1146,n1147,n17);
nor (n1147,n1148,n1149);
and (n1148,n102,n537);
and (n1149,n110,n539);
xnor (n1150,n1151,n12);
nor (n1151,n1152,n1153);
and (n1152,n310,n350);
and (n1153,n115,n353);
and (n1154,n1150,n44);
and (n1155,n1146,n44);
and (n1156,n1157,n1161);
xnor (n1157,n1158,n28);
nor (n1158,n1159,n1160);
and (n1159,n466,n22);
and (n1160,n372,n27);
xnor (n1161,n1162,n44);
nand (n1162,n624,n41);
and (n1163,n1156,n1164);
xnor (n1164,n1165,n44);
nor (n1165,n1166,n1167);
and (n1166,n624,n36);
and (n1167,n466,n41);
and (n1168,n1144,n1164);
xor (n1169,n1170,n1127);
xor (n1170,n1108,n1124);
and (n1171,n1172,n1173);
xor (n1172,n1139,n1141);
or (n1173,n1174,n1181);
and (n1174,n1175,n1176);
xor (n1175,n1142,n1169);
and (n1176,n1177,n1179);
xor (n1177,n1178,n1119);
xor (n1178,n1110,n1114);
xor (n1179,n1180,n1164);
xor (n1180,n1144,n1156);
and (n1181,n1182,n1183);
xor (n1182,n1175,n1176);
or (n1183,n1184,n1209);
and (n1184,n1185,n1186);
xor (n1185,n1177,n1179);
or (n1186,n1187,n1206,n1208);
and (n1187,n1188,n1204);
or (n1188,n1189,n1198,n1203);
and (n1189,n1190,n1194);
xnor (n1190,n1191,n17);
nor (n1191,n1192,n1193);
and (n1192,n115,n537);
and (n1193,n102,n539);
xnor (n1194,n1195,n12);
nor (n1195,n1196,n1197);
and (n1196,n372,n350);
and (n1197,n310,n353);
and (n1198,n1194,n1199);
xnor (n1199,n1200,n28);
nor (n1200,n1201,n1202);
and (n1201,n624,n22);
and (n1202,n466,n27);
and (n1203,n1190,n1199);
xor (n1204,n1205,n44);
xor (n1205,n1146,n1150);
and (n1206,n1204,n1207);
xor (n1207,n1157,n1161);
and (n1208,n1188,n1207);
and (n1209,n1210,n1211);
xor (n1210,n1185,n1186);
or (n1211,n1212,n1230);
and (n1212,n1213,n1215);
xor (n1213,n1214,n1207);
xor (n1214,n1188,n1204);
and (n1215,n1216,n1228);
or (n1216,n1217,n1226,n1227);
and (n1217,n1218,n1222);
xnor (n1218,n1219,n17);
nor (n1219,n1220,n1221);
and (n1220,n310,n537);
and (n1221,n115,n539);
xnor (n1222,n1223,n12);
nor (n1223,n1224,n1225);
and (n1224,n466,n350);
and (n1225,n372,n353);
and (n1226,n1222,n28);
and (n1227,n1218,n28);
xor (n1228,n1229,n1199);
xor (n1229,n1190,n1194);
and (n1230,n1231,n1232);
xor (n1231,n1213,n1215);
or (n1232,n1233,n1240);
and (n1233,n1234,n1235);
xor (n1234,n1216,n1228);
and (n1235,n1236,n1238);
xnor (n1236,n1237,n28);
nand (n1237,n624,n27);
xor (n1238,n1239,n28);
xor (n1239,n1218,n1222);
and (n1240,n1241,n1242);
xor (n1241,n1234,n1235);
or (n1242,n1243,n1254);
and (n1243,n1244,n1245);
xor (n1244,n1236,n1238);
and (n1245,n1246,n1250);
xnor (n1246,n1247,n17);
nor (n1247,n1248,n1249);
and (n1248,n372,n537);
and (n1249,n310,n539);
xnor (n1250,n1251,n12);
nor (n1251,n1252,n1253);
and (n1252,n624,n350);
and (n1253,n466,n353);
and (n1254,n1255,n1256);
xor (n1255,n1244,n1245);
or (n1256,n1257,n1264);
and (n1257,n1258,n1259);
xor (n1258,n1246,n1250);
and (n1259,n1260,n12);
xnor (n1260,n1261,n17);
nor (n1261,n1262,n1263);
and (n1262,n466,n537);
and (n1263,n372,n539);
and (n1264,n1265,n1266);
xor (n1265,n1258,n1259);
or (n1266,n1267,n1271);
and (n1267,n1268,n1270);
xnor (n1268,n1269,n12);
nand (n1269,n624,n353);
xor (n1270,n1260,n12);
and (n1271,n1272,n1273);
xor (n1272,n1268,n1270);
and (n1273,n1274,n1278);
xnor (n1274,n1275,n17);
nor (n1275,n1276,n1277);
and (n1276,n624,n537);
and (n1277,n466,n539);
and (n1278,n1279,n17);
xnor (n1279,n1280,n17);
nand (n1280,n624,n539);
xor (n1281,n1282,n1377);
xor (n1282,n1283,n1346);
xor (n1283,n1284,n1332);
xor (n1284,n1285,n1302);
or (n1285,n1286,n1292,n1301);
and (n1286,n1287,n1291);
or (n1287,n1288,n184);
or (n1288,n1289,n182,n1290);
and (n1289,n167,n121);
and (n1290,n167,n125);
not (n1291,n207);
and (n1292,n1291,n1293);
xor (n1293,n1294,n194);
xor (n1294,n1295,n1298);
or (n1295,n220,n1296,n1297);
and (n1296,n161,n150);
and (n1297,n157,n150);
or (n1298,n224,n1299,n1300);
and (n1299,n171,n153);
and (n1300,n168,n153);
and (n1301,n1287,n1293);
or (n1302,n1303,n1328,n1331);
and (n1303,n1304,n1324);
or (n1304,n1305,n1320,n1323);
and (n1305,n1306,n1316);
or (n1306,n1307,n1314,n1315);
and (n1307,n1308,n1311);
or (n1308,n31,n1309,n1310);
and (n1309,n32,n50);
and (n1310,n18,n50);
or (n1311,n80,n1312,n1313);
and (n1312,n81,n99);
and (n1313,n65,n99);
and (n1314,n1311,n114);
and (n1315,n1308,n114);
or (n1316,n1317,n1318,n1319);
and (n1317,n145,n324);
and (n1318,n324,n129);
and (n1319,n145,n129);
and (n1320,n1316,n1321);
xor (n1321,n1322,n150);
xor (n1322,n157,n161);
and (n1323,n1306,n1321);
and (n1324,n1325,n1327);
xor (n1325,n1326,n153);
xor (n1326,n168,n171);
xnor (n1327,n1288,n184);
and (n1328,n1324,n1329);
xor (n1329,n1330,n1293);
xor (n1330,n1287,n1291);
and (n1331,n1304,n1329);
xor (n1332,n1333,n1340);
xor (n1333,n1334,n1338);
or (n1334,n1335,n1336,n1337);
and (n1335,n1295,n1298);
and (n1336,n1298,n194);
and (n1337,n1295,n194);
xor (n1338,n1339,n259);
xor (n1339,n240,n243);
xor (n1340,n1341,n1345);
xor (n1341,n249,n1342);
or (n1342,n1343,n255,n1344);
and (n1343,n239,n209);
and (n1344,n239,n213);
xnor (n1345,n263,n267);
and (n1346,n1347,n1375);
or (n1347,n1348,n1372,n1374);
and (n1348,n1349,n1370);
or (n1349,n1350,n1368,n1369);
and (n1350,n1351,n1359);
or (n1351,n1352,n1356,n1358);
and (n1352,n1353,n287);
or (n1353,n1354,n281,n1355);
and (n1354,n11,n277);
and (n1355,n11,n282);
and (n1356,n287,n1357);
and (n1357,n305,n309);
and (n1358,n1353,n1357);
or (n1359,n1360,n1365,n1367);
and (n1360,n1361,n1363);
xor (n1361,n1362,n50);
xor (n1362,n18,n32);
xor (n1363,n1364,n99);
xor (n1364,n65,n81);
and (n1365,n1363,n1366);
not (n1366,n114);
and (n1367,n1361,n1366);
and (n1368,n1359,n322);
and (n1369,n1351,n322);
xor (n1370,n1371,n1321);
xor (n1371,n1306,n1316);
and (n1372,n1370,n1373);
xor (n1373,n1325,n1327);
and (n1374,n1349,n1373);
xor (n1375,n1376,n1329);
xor (n1376,n1304,n1324);
or (n1377,n1378,n1412);
and (n1378,n1379,n1380);
xor (n1379,n1347,n1375);
and (n1380,n1381,n1410);
or (n1381,n1382,n1406,n1409);
and (n1382,n1383,n1404);
or (n1383,n1384,n1400,n1403);
and (n1384,n1385,n1396);
or (n1385,n1386,n1393,n1395);
and (n1386,n1387,n1390);
or (n1387,n354,n1388,n1389);
and (n1388,n355,n377);
and (n1389,n347,n377);
or (n1390,n385,n1391,n1392);
and (n1391,n386,n362);
and (n1392,n381,n362);
and (n1393,n1390,n1394);
or (n1394,n366,n371);
and (n1395,n1387,n1394);
or (n1396,n1397,n1398,n1399);
and (n1397,n477,n396);
and (n1398,n396,n478);
and (n1399,n477,n478);
and (n1400,n1396,n1401);
xor (n1401,n1402,n1366);
xor (n1402,n1361,n1363);
and (n1403,n1385,n1401);
xor (n1404,n1405,n114);
xor (n1405,n1308,n1311);
and (n1406,n1404,n1407);
xor (n1407,n1408,n322);
xor (n1408,n1351,n1359);
and (n1409,n1383,n1407);
xor (n1410,n1411,n1373);
xor (n1411,n1349,n1370);
and (n1412,n1413,n1414);
xor (n1413,n1379,n1380);
or (n1414,n1415,n1447);
and (n1415,n1416,n1417);
xor (n1416,n1381,n1410);
and (n1417,n1418,n1445);
or (n1418,n1419,n1441,n1444);
and (n1419,n1420,n1439);
or (n1420,n1421,n1437,n1438);
and (n1421,n1422,n1428);
or (n1422,n1423,n1427,n468);
and (n1423,n425,n1424);
or (n1424,n1425,n447,n1426);
and (n1425,n346,n443);
and (n1426,n346,n448);
and (n1427,n1424,n454);
or (n1428,n1429,n1434,n1436);
and (n1429,n1430,n1432);
xor (n1430,n1431,n377);
xor (n1431,n347,n355);
xor (n1432,n1433,n362);
xor (n1433,n381,n386);
and (n1434,n1432,n1435);
xnor (n1435,n366,n371);
and (n1436,n1430,n1435);
and (n1437,n1428,n475);
and (n1438,n1422,n475);
xor (n1439,n1440,n1357);
xor (n1440,n1353,n287);
and (n1441,n1439,n1442);
xor (n1442,n1443,n1401);
xor (n1443,n1385,n1396);
and (n1444,n1420,n1442);
xor (n1445,n1446,n1407);
xor (n1446,n1383,n1404);
and (n1447,n1448,n1449);
xor (n1448,n1416,n1417);
or (n1449,n1450,n1470);
and (n1450,n1451,n1452);
xor (n1451,n1418,n1445);
and (n1452,n1453,n1468);
or (n1453,n1454,n1464,n1467);
and (n1454,n1455,n1462);
or (n1455,n1456,n1458,n1461);
and (n1456,n498,n1457);
or (n1457,n548,n553);
and (n1458,n1457,n1459);
xor (n1459,n1460,n1435);
xor (n1460,n1430,n1432);
and (n1461,n498,n1459);
xor (n1462,n1463,n1394);
xor (n1463,n1387,n1390);
and (n1464,n1462,n1465);
xor (n1465,n1466,n475);
xor (n1466,n1422,n1428);
and (n1467,n1455,n1465);
xor (n1468,n1469,n1442);
xor (n1469,n1420,n1439);
and (n1470,n1471,n1472);
xor (n1471,n1451,n1452);
or (n1472,n1473,n1489);
and (n1473,n1474,n1475);
xor (n1474,n1453,n1468);
and (n1475,n1476,n1487);
or (n1476,n1477,n1483,n1486);
and (n1477,n1478,n1481);
or (n1478,n580,n1479,n1480);
and (n1479,n627,n749);
and (n1480,n581,n749);
xor (n1481,n1482,n454);
xor (n1482,n425,n1424);
and (n1483,n1481,n1484);
xor (n1484,n1485,n1459);
xor (n1485,n498,n1457);
and (n1486,n1478,n1484);
xor (n1487,n1488,n1465);
xor (n1488,n1455,n1462);
and (n1489,n1490,n1491);
xor (n1490,n1474,n1475);
or (n1491,n1492,n1500);
and (n1492,n1493,n1494);
xor (n1493,n1476,n1487);
and (n1494,n1495,n1498);
or (n1495,n660,n1496,n1497);
and (n1496,n721,n751);
and (n1497,n661,n751);
xor (n1498,n1499,n1484);
xor (n1499,n1478,n1481);
and (n1500,n1501,n1502);
xor (n1501,n1493,n1494);
or (n1502,n1503,n742);
and (n1503,n1504,n1505);
xor (n1504,n1495,n1498);
or (n1505,n1506,n1507,n1508);
and (n1506,n727,n748);
and (n1507,n748,n750);
and (n1508,n727,n750);
endmodule
