module top (out,n3,n37,n38,n43,n45,n53,n62,n63,n69
        ,n76,n81,n91,n92,n97,n102,n108,n119,n120,n126
        ,n131,n138,n147,n156,n163,n173,n174,n179,n180,n192
        ,n196,n203,n217,n223,n229,n230,n234,n240,n249,n251
        ,n257,n267,n278,n280,n288,n297,n306,n307,n314,n323
        ,n335,n358,n360,n368,n376,n384,n385,n392,n403,n416
        ,n452,n460,n490,n496,n517,n556,n3518,n3519,n3528,n3529
        ,n3537,n3545,n3546,n3554,n3566,n3573,n3575,n3581,n3586,n3592
        ,n3602,n3603,n3611,n3615,n3622,n3624,n3632,n3633,n3641,n3650
        ,n3651,n3657,n3659,n3670,n3680,n3687,n3695,n3704,n3723,n3732
        ,n3733,n3741,n3756,n3763,n3774,n3783,n3790,n3800,n3806,n3808
        ,n3820,n3828,n3837,n3843,n3866,n3867,n3929,n3935,n3952,n3959
        ,n4025,n4032,n4342,n4350,n4384,n4406,n4413,n4423,n5233,n5241
        ,n7034,n7036,n7042,n7049,n7055,n7064,n7065,n7072,n7078,n7084
        ,n7091,n7093,n7102,n7109,n7120,n7123,n7124,n7129,n7134,n7146
        ,n7147,n7154,n7165,n7173,n7174,n7180,n7181,n7194,n7204,n7205
        ,n7212,n7223,n7232,n7237,n7242,n7251,n7253,n7261,n7270,n7289
        ,n7308,n7330,n7339,n7355,n7366,n7378,n7383,n7385,n7391,n7463
        ,n7471,n7479,n7483,n7497,n7527,n7558,n7595,n7745,n7753,n7758
        ,n7853,n7859,n7867,n7917,n10462,n10471,n10472,n10476,n10477,n10481
        ,n10482,n10485,n10487,n10504,n10511,n10512,n10516,n10517,n10519,n10521
        ,n10524,n10535,n10536,n10541,n10543,n10548,n10549,n10553,n10554,n10571
        ,n10572,n10577,n10578,n10581,n10582,n10585,n10586,n10607,n10609,n10612
        ,n10613,n10622,n10623,n10628,n10629,n10635,n10637,n10638,n10644,n10646
        ,n10649,n10650,n10661,n10662,n10665,n10666,n10669,n10670,n10674,n10675
        ,n10690,n10691,n10696,n10697,n10700,n10701,n10704,n10705,n10714,n10715
        ,n10717);
output out;
input n3;
input n37;
input n38;
input n43;
input n45;
input n53;
input n62;
input n63;
input n69;
input n76;
input n81;
input n91;
input n92;
input n97;
input n102;
input n108;
input n119;
input n120;
input n126;
input n131;
input n138;
input n147;
input n156;
input n163;
input n173;
input n174;
input n179;
input n180;
input n192;
input n196;
input n203;
input n217;
input n223;
input n229;
input n230;
input n234;
input n240;
input n249;
input n251;
input n257;
input n267;
input n278;
input n280;
input n288;
input n297;
input n306;
input n307;
input n314;
input n323;
input n335;
input n358;
input n360;
input n368;
input n376;
input n384;
input n385;
input n392;
input n403;
input n416;
input n452;
input n460;
input n490;
input n496;
input n517;
input n556;
input n3518;
input n3519;
input n3528;
input n3529;
input n3537;
input n3545;
input n3546;
input n3554;
input n3566;
input n3573;
input n3575;
input n3581;
input n3586;
input n3592;
input n3602;
input n3603;
input n3611;
input n3615;
input n3622;
input n3624;
input n3632;
input n3633;
input n3641;
input n3650;
input n3651;
input n3657;
input n3659;
input n3670;
input n3680;
input n3687;
input n3695;
input n3704;
input n3723;
input n3732;
input n3733;
input n3741;
input n3756;
input n3763;
input n3774;
input n3783;
input n3790;
input n3800;
input n3806;
input n3808;
input n3820;
input n3828;
input n3837;
input n3843;
input n3866;
input n3867;
input n3929;
input n3935;
input n3952;
input n3959;
input n4025;
input n4032;
input n4342;
input n4350;
input n4384;
input n4406;
input n4413;
input n4423;
input n5233;
input n5241;
input n7034;
input n7036;
input n7042;
input n7049;
input n7055;
input n7064;
input n7065;
input n7072;
input n7078;
input n7084;
input n7091;
input n7093;
input n7102;
input n7109;
input n7120;
input n7123;
input n7124;
input n7129;
input n7134;
input n7146;
input n7147;
input n7154;
input n7165;
input n7173;
input n7174;
input n7180;
input n7181;
input n7194;
input n7204;
input n7205;
input n7212;
input n7223;
input n7232;
input n7237;
input n7242;
input n7251;
input n7253;
input n7261;
input n7270;
input n7289;
input n7308;
input n7330;
input n7339;
input n7355;
input n7366;
input n7378;
input n7383;
input n7385;
input n7391;
input n7463;
input n7471;
input n7479;
input n7483;
input n7497;
input n7527;
input n7558;
input n7595;
input n7745;
input n7753;
input n7758;
input n7853;
input n7859;
input n7867;
input n7917;
input n10462;
input n10471;
input n10472;
input n10476;
input n10477;
input n10481;
input n10482;
input n10485;
input n10487;
input n10504;
input n10511;
input n10512;
input n10516;
input n10517;
input n10519;
input n10521;
input n10524;
input n10535;
input n10536;
input n10541;
input n10543;
input n10548;
input n10549;
input n10553;
input n10554;
input n10571;
input n10572;
input n10577;
input n10578;
input n10581;
input n10582;
input n10585;
input n10586;
input n10607;
input n10609;
input n10612;
input n10613;
input n10622;
input n10623;
input n10628;
input n10629;
input n10635;
input n10637;
input n10638;
input n10644;
input n10646;
input n10649;
input n10650;
input n10661;
input n10662;
input n10665;
input n10666;
input n10669;
input n10670;
input n10674;
input n10675;
input n10690;
input n10691;
input n10696;
input n10697;
input n10700;
input n10701;
input n10704;
input n10705;
input n10714;
input n10715;
input n10717;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n175;
wire n176;
wire n177;
wire n178;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n231;
wire n232;
wire n233;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n250;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3574;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3612;
wire n3613;
wire n3614;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3623;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3658;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3807;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7035;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7092;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7121;
wire n7122;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7252;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7384;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7480;
wire n7481;
wire n7482;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10449;
wire n10450;
wire n10451;
wire n10452;
wire n10453;
wire n10454;
wire n10455;
wire n10456;
wire n10457;
wire n10458;
wire n10459;
wire n10460;
wire n10461;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10467;
wire n10468;
wire n10469;
wire n10470;
wire n10473;
wire n10474;
wire n10475;
wire n10478;
wire n10479;
wire n10480;
wire n10483;
wire n10484;
wire n10486;
wire n10488;
wire n10489;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10505;
wire n10506;
wire n10507;
wire n10508;
wire n10509;
wire n10510;
wire n10513;
wire n10514;
wire n10515;
wire n10518;
wire n10520;
wire n10522;
wire n10523;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10537;
wire n10538;
wire n10539;
wire n10540;
wire n10542;
wire n10544;
wire n10545;
wire n10546;
wire n10547;
wire n10550;
wire n10551;
wire n10552;
wire n10555;
wire n10556;
wire n10557;
wire n10558;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10566;
wire n10567;
wire n10568;
wire n10569;
wire n10570;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10579;
wire n10580;
wire n10583;
wire n10584;
wire n10587;
wire n10588;
wire n10589;
wire n10590;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10602;
wire n10603;
wire n10604;
wire n10605;
wire n10606;
wire n10608;
wire n10610;
wire n10611;
wire n10614;
wire n10615;
wire n10616;
wire n10617;
wire n10618;
wire n10619;
wire n10620;
wire n10621;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10636;
wire n10639;
wire n10640;
wire n10641;
wire n10642;
wire n10643;
wire n10645;
wire n10647;
wire n10648;
wire n10651;
wire n10652;
wire n10653;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10663;
wire n10664;
wire n10667;
wire n10668;
wire n10671;
wire n10672;
wire n10673;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10683;
wire n10684;
wire n10685;
wire n10686;
wire n10687;
wire n10688;
wire n10689;
wire n10692;
wire n10693;
wire n10694;
wire n10695;
wire n10698;
wire n10699;
wire n10702;
wire n10703;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10716;
wire n10718;
wire n10719;
wire n10720;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10729;
wire n10730;
wire n10731;
wire n10732;
wire n10733;
wire n10734;
wire n10735;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10747;
wire n10748;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10766;
wire n10767;
wire n10768;
wire n10769;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10780;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10793;
wire n10794;
wire n10795;
wire n10796;
wire n10797;
wire n10798;
wire n10799;
wire n10800;
wire n10801;
wire n10802;
wire n10803;
wire n10804;
wire n10805;
wire n10806;
wire n10807;
wire n10808;
wire n10809;
wire n10810;
wire n10811;
wire n10812;
wire n10813;
wire n10814;
wire n10815;
wire n10816;
wire n10817;
wire n10818;
wire n10819;
wire n10820;
wire n10821;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10831;
wire n10832;
wire n10833;
wire n10834;
wire n10835;
wire n10836;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10842;
wire n10843;
wire n10844;
wire n10845;
wire n10846;
wire n10847;
wire n10848;
wire n10849;
wire n10850;
wire n10851;
wire n10852;
wire n10853;
wire n10854;
wire n10855;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n10869;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10877;
wire n10878;
wire n10879;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n10890;
wire n10891;
wire n10892;
wire n10893;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10899;
wire n10900;
wire n10901;
wire n10902;
wire n10903;
wire n10904;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10917;
wire n10918;
wire n10919;
wire n10920;
wire n10921;
wire n10922;
wire n10923;
wire n10924;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10930;
wire n10931;
wire n10932;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10937;
wire n10938;
wire n10939;
wire n10940;
wire n10941;
wire n10942;
wire n10943;
wire n10944;
wire n10945;
wire n10946;
wire n10947;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10963;
wire n10964;
wire n10965;
wire n10966;
wire n10967;
wire n10968;
wire n10969;
wire n10970;
wire n10971;
wire n10972;
wire n10973;
wire n10974;
wire n10975;
wire n10976;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10986;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10992;
wire n10993;
wire n10994;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11006;
wire n11007;
wire n11008;
wire n11009;
wire n11010;
wire n11011;
wire n11012;
wire n11013;
wire n11014;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n11020;
wire n11021;
wire n11022;
wire n11023;
wire n11024;
wire n11025;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11030;
wire n11031;
wire n11032;
wire n11033;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11038;
wire n11039;
wire n11040;
wire n11041;
wire n11042;
wire n11043;
wire n11044;
wire n11045;
wire n11046;
wire n11047;
wire n11048;
wire n11049;
wire n11050;
wire n11051;
wire n11052;
wire n11053;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n11058;
wire n11059;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11071;
wire n11072;
wire n11073;
wire n11074;
wire n11075;
wire n11076;
wire n11077;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11087;
wire n11088;
wire n11089;
wire n11090;
wire n11091;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11097;
wire n11098;
wire n11099;
wire n11100;
wire n11101;
wire n11102;
wire n11103;
wire n11104;
wire n11105;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11114;
wire n11115;
wire n11116;
wire n11117;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11132;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11145;
wire n11146;
wire n11147;
wire n11148;
wire n11149;
wire n11150;
wire n11151;
wire n11152;
wire n11153;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n11160;
wire n11161;
wire n11162;
wire n11163;
wire n11164;
wire n11165;
wire n11166;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11180;
wire n11181;
wire n11182;
wire n11183;
wire n11184;
wire n11185;
wire n11186;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11228;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11239;
wire n11240;
wire n11241;
wire n11242;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11247;
wire n11248;
wire n11249;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11260;
wire n11261;
wire n11262;
wire n11263;
wire n11264;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11273;
wire n11274;
wire n11275;
wire n11276;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11292;
wire n11293;
wire n11294;
wire n11295;
wire n11296;
wire n11297;
wire n11298;
wire n11299;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11338;
wire n11339;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11346;
wire n11347;
wire n11348;
wire n11349;
wire n11350;
wire n11351;
wire n11352;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11396;
wire n11397;
wire n11398;
wire n11399;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n11450;
wire n11451;
wire n11452;
wire n11453;
wire n11454;
wire n11455;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11460;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11469;
wire n11470;
wire n11471;
wire n11472;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11493;
wire n11494;
wire n11495;
wire n11496;
wire n11497;
wire n11498;
wire n11499;
wire n11500;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11506;
wire n11507;
wire n11508;
wire n11509;
wire n11510;
wire n11511;
wire n11512;
wire n11513;
wire n11514;
wire n11515;
wire n11516;
wire n11517;
wire n11518;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11525;
wire n11526;
wire n11527;
wire n11528;
wire n11529;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11563;
wire n11564;
wire n11565;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11578;
wire n11579;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11588;
wire n11589;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11597;
wire n11598;
wire n11599;
wire n11600;
wire n11601;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11607;
wire n11608;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11623;
wire n11624;
wire n11625;
wire n11626;
wire n11627;
wire n11628;
wire n11629;
wire n11630;
wire n11631;
wire n11632;
wire n11633;
wire n11634;
wire n11635;
wire n11636;
wire n11637;
wire n11638;
wire n11639;
wire n11640;
wire n11641;
wire n11642;
wire n11643;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11649;
wire n11650;
wire n11651;
wire n11652;
wire n11653;
wire n11654;
wire n11655;
wire n11656;
wire n11657;
wire n11658;
wire n11659;
wire n11660;
wire n11661;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11666;
wire n11667;
wire n11668;
wire n11669;
wire n11670;
wire n11671;
wire n11672;
wire n11673;
wire n11674;
wire n11675;
wire n11676;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11689;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11728;
wire n11729;
wire n11730;
wire n11731;
wire n11732;
wire n11733;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11757;
wire n11758;
wire n11759;
wire n11760;
wire n11761;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11766;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11771;
wire n11772;
wire n11773;
wire n11774;
wire n11775;
wire n11776;
wire n11777;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11789;
wire n11790;
wire n11791;
wire n11792;
wire n11793;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11798;
wire n11799;
wire n11800;
wire n11801;
wire n11802;
wire n11803;
wire n11804;
wire n11805;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11813;
wire n11814;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11835;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11840;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11850;
wire n11851;
wire n11852;
wire n11853;
wire n11854;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11869;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11874;
wire n11875;
wire n11876;
wire n11877;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11887;
wire n11888;
wire n11889;
wire n11890;
wire n11891;
wire n11892;
wire n11893;
wire n11894;
wire n11895;
wire n11896;
wire n11897;
wire n11898;
wire n11899;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11907;
wire n11908;
wire n11909;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11925;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11936;
wire n11937;
wire n11938;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11949;
wire n11950;
wire n11951;
wire n11952;
wire n11953;
wire n11954;
wire n11955;
wire n11956;
wire n11957;
wire n11958;
wire n11959;
wire n11960;
wire n11961;
wire n11962;
wire n11963;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11988;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11996;
wire n11997;
wire n11998;
wire n11999;
wire n12000;
wire n12001;
wire n12002;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12007;
wire n12008;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12024;
wire n12025;
wire n12026;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12043;
wire n12044;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12049;
wire n12050;
wire n12051;
wire n12052;
wire n12053;
wire n12054;
wire n12055;
wire n12056;
wire n12057;
wire n12058;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12067;
wire n12068;
wire n12069;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12076;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12081;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12095;
wire n12096;
wire n12097;
wire n12098;
wire n12099;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12122;
wire n12123;
wire n12124;
wire n12125;
wire n12126;
wire n12127;
wire n12128;
wire n12129;
wire n12130;
wire n12131;
wire n12132;
wire n12133;
wire n12134;
wire n12135;
wire n12136;
wire n12137;
wire n12138;
wire n12139;
wire n12140;
wire n12141;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12146;
wire n12147;
wire n12148;
wire n12149;
wire n12150;
wire n12151;
wire n12152;
wire n12153;
wire n12154;
wire n12155;
wire n12156;
wire n12157;
wire n12158;
wire n12159;
wire n12160;
wire n12161;
wire n12162;
wire n12163;
wire n12164;
wire n12165;
wire n12166;
wire n12167;
wire n12168;
wire n12169;
wire n12170;
wire n12171;
wire n12172;
wire n12173;
wire n12174;
wire n12175;
wire n12176;
wire n12177;
wire n12178;
wire n12179;
wire n12180;
wire n12181;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12189;
wire n12190;
wire n12191;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n12200;
wire n12201;
wire n12202;
wire n12203;
wire n12204;
wire n12205;
wire n12206;
wire n12207;
wire n12208;
wire n12209;
wire n12210;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12228;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12233;
wire n12234;
wire n12235;
wire n12236;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12244;
wire n12245;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12255;
wire n12256;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12266;
wire n12267;
wire n12268;
wire n12269;
wire n12270;
wire n12271;
wire n12272;
wire n12273;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12281;
wire n12282;
wire n12283;
wire n12284;
wire n12285;
wire n12286;
wire n12287;
wire n12288;
wire n12289;
wire n12290;
wire n12291;
wire n12292;
wire n12293;
wire n12294;
wire n12295;
wire n12296;
wire n12297;
wire n12298;
wire n12299;
wire n12300;
wire n12301;
wire n12302;
wire n12303;
wire n12304;
wire n12305;
wire n12306;
wire n12307;
wire n12308;
wire n12309;
wire n12310;
wire n12311;
wire n12312;
wire n12313;
wire n12314;
wire n12315;
wire n12316;
wire n12317;
wire n12318;
wire n12319;
wire n12320;
wire n12321;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12326;
wire n12327;
wire n12328;
wire n12329;
wire n12330;
wire n12331;
wire n12332;
wire n12333;
wire n12334;
wire n12335;
wire n12336;
wire n12337;
wire n12338;
wire n12339;
wire n12340;
wire n12341;
wire n12342;
wire n12343;
wire n12344;
wire n12345;
wire n12346;
wire n12347;
wire n12348;
wire n12349;
wire n12350;
wire n12351;
wire n12352;
wire n12353;
wire n12354;
wire n12355;
wire n12356;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n12370;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12389;
wire n12390;
wire n12391;
wire n12392;
wire n12393;
wire n12394;
wire n12395;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n12400;
wire n12401;
wire n12402;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12409;
wire n12410;
wire n12411;
wire n12412;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12417;
wire n12418;
wire n12419;
wire n12420;
wire n12421;
wire n12422;
wire n12423;
wire n12424;
wire n12425;
wire n12426;
wire n12427;
wire n12428;
wire n12429;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12440;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12455;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12479;
wire n12480;
wire n12481;
wire n12482;
wire n12483;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12494;
wire n12495;
wire n12496;
wire n12497;
wire n12498;
wire n12499;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12519;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12527;
wire n12528;
wire n12529;
wire n12530;
wire n12531;
wire n12532;
wire n12533;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12558;
wire n12559;
wire n12560;
wire n12561;
wire n12562;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12582;
wire n12583;
wire n12584;
wire n12585;
wire n12586;
wire n12587;
wire n12588;
wire n12589;
wire n12590;
wire n12591;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n12600;
wire n12601;
wire n12602;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12632;
wire n12633;
wire n12634;
wire n12635;
wire n12636;
wire n12637;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12649;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12665;
wire n12666;
wire n12667;
wire n12668;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12673;
wire n12674;
wire n12675;
wire n12676;
wire n12677;
wire n12678;
wire n12679;
wire n12680;
wire n12681;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12725;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12743;
wire n12744;
wire n12745;
wire n12746;
wire n12747;
wire n12748;
wire n12749;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12754;
wire n12755;
wire n12756;
wire n12757;
wire n12758;
wire n12759;
wire n12760;
wire n12761;
wire n12762;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12772;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12777;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12813;
wire n12814;
wire n12815;
wire n12816;
wire n12817;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12825;
wire n12826;
wire n12827;
wire n12828;
wire n12829;
wire n12830;
wire n12831;
wire n12832;
wire n12833;
wire n12834;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12842;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12865;
wire n12866;
wire n12867;
wire n12868;
wire n12869;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12874;
wire n12875;
wire n12876;
wire n12877;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12946;
wire n12947;
wire n12948;
wire n12949;
wire n12950;
wire n12951;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12985;
wire n12986;
wire n12987;
wire n12988;
wire n12989;
wire n12990;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13004;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13042;
wire n13043;
wire n13044;
wire n13045;
wire n13046;
wire n13047;
wire n13048;
wire n13049;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13086;
wire n13087;
wire n13088;
wire n13089;
wire n13090;
wire n13091;
wire n13092;
wire n13093;
wire n13094;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n13100;
wire n13101;
wire n13102;
wire n13103;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13135;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13140;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13176;
wire n13177;
wire n13178;
wire n13179;
wire n13180;
wire n13181;
wire n13182;
wire n13183;
wire n13184;
wire n13185;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13198;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13221;
wire n13222;
wire n13223;
wire n13224;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13261;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13276;
wire n13277;
wire n13278;
wire n13279;
wire n13280;
wire n13281;
wire n13282;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13303;
wire n13304;
wire n13305;
wire n13306;
wire n13307;
wire n13308;
wire n13309;
wire n13310;
wire n13311;
wire n13312;
wire n13313;
wire n13314;
wire n13315;
wire n13316;
wire n13317;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13365;
wire n13366;
wire n13367;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13394;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13404;
wire n13405;
wire n13406;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13425;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n13480;
wire n13481;
wire n13482;
wire n13483;
wire n13484;
wire n13485;
wire n13486;
wire n13487;
wire n13488;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13513;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n13530;
wire n13531;
wire n13532;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13550;
wire n13551;
wire n13552;
wire n13553;
wire n13554;
wire n13555;
wire n13556;
wire n13557;
wire n13558;
wire n13559;
wire n13560;
wire n13561;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13566;
wire n13567;
wire n13568;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13584;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13597;
wire n13598;
wire n13599;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13608;
wire n13609;
wire n13610;
wire n13611;
wire n13612;
wire n13613;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13618;
wire n13619;
wire n13620;
wire n13621;
wire n13622;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n13630;
wire n13631;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13636;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13667;
wire n13668;
wire n13669;
wire n13670;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n13680;
wire n13681;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13692;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13697;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13715;
wire n13716;
wire n13717;
wire n13718;
wire n13719;
wire n13720;
wire n13721;
wire n13722;
wire n13723;
wire n13724;
wire n13725;
wire n13726;
wire n13727;
wire n13728;
wire n13729;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13741;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13746;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13765;
wire n13766;
wire n13767;
wire n13768;
wire n13769;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13791;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13796;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n13820;
wire n13821;
wire n13822;
wire n13823;
wire n13824;
wire n13825;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13831;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13840;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13845;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13851;
wire n13852;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13868;
wire n13869;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13877;
wire n13878;
wire n13879;
wire n13880;
wire n13881;
wire n13882;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13887;
wire n13888;
wire n13889;
wire n13890;
wire n13891;
wire n13892;
wire n13893;
wire n13894;
wire n13895;
wire n13896;
wire n13897;
wire n13898;
wire n13899;
wire n13900;
wire n13901;
wire n13902;
wire n13903;
wire n13904;
wire n13905;
wire n13906;
wire n13907;
wire n13908;
wire n13909;
wire n13910;
wire n13911;
wire n13912;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13919;
wire n13920;
wire n13921;
wire n13922;
wire n13923;
wire n13924;
wire n13925;
wire n13926;
wire n13927;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13934;
wire n13935;
wire n13936;
wire n13937;
wire n13938;
wire n13939;
wire n13940;
wire n13941;
wire n13942;
wire n13943;
wire n13944;
wire n13945;
wire n13946;
wire n13947;
wire n13948;
wire n13949;
wire n13950;
wire n13951;
wire n13952;
wire n13953;
wire n13954;
wire n13955;
wire n13956;
wire n13957;
wire n13958;
wire n13959;
wire n13960;
wire n13961;
wire n13962;
wire n13963;
wire n13964;
wire n13965;
wire n13966;
wire n13967;
wire n13968;
wire n13969;
wire n13970;
wire n13971;
wire n13972;
wire n13973;
wire n13974;
wire n13975;
wire n13976;
wire n13977;
wire n13978;
wire n13979;
wire n13980;
wire n13981;
wire n13982;
wire n13983;
wire n13984;
wire n13985;
wire n13986;
wire n13987;
wire n13988;
wire n13989;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13997;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14002;
wire n14003;
wire n14004;
wire n14005;
wire n14006;
wire n14007;
wire n14008;
wire n14009;
wire n14010;
wire n14011;
wire n14012;
wire n14013;
wire n14014;
wire n14015;
wire n14016;
wire n14017;
wire n14018;
wire n14019;
wire n14020;
wire n14021;
wire n14022;
wire n14023;
wire n14024;
wire n14025;
wire n14026;
wire n14027;
wire n14028;
wire n14029;
wire n14030;
wire n14031;
wire n14032;
wire n14033;
wire n14034;
wire n14035;
wire n14036;
wire n14037;
wire n14038;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14043;
wire n14044;
wire n14045;
wire n14046;
wire n14047;
wire n14048;
wire n14049;
wire n14050;
wire n14051;
wire n14052;
wire n14053;
wire n14054;
wire n14055;
wire n14056;
wire n14057;
wire n14058;
wire n14059;
wire n14060;
wire n14061;
wire n14062;
wire n14063;
wire n14064;
wire n14065;
wire n14066;
wire n14067;
wire n14068;
wire n14069;
wire n14070;
wire n14071;
wire n14072;
wire n14073;
wire n14074;
wire n14075;
wire n14076;
wire n14077;
wire n14078;
wire n14079;
wire n14080;
wire n14081;
wire n14082;
wire n14083;
wire n14084;
wire n14085;
wire n14086;
wire n14087;
wire n14088;
wire n14089;
wire n14090;
wire n14091;
wire n14092;
wire n14093;
wire n14094;
wire n14095;
wire n14096;
wire n14097;
wire n14098;
wire n14099;
wire n14100;
wire n14101;
wire n14102;
wire n14103;
wire n14104;
wire n14105;
wire n14106;
wire n14107;
wire n14108;
wire n14109;
wire n14110;
wire n14111;
wire n14112;
wire n14113;
wire n14114;
wire n14115;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14121;
wire n14122;
wire n14123;
wire n14124;
wire n14125;
wire n14126;
wire n14127;
wire n14128;
wire n14129;
wire n14130;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14135;
wire n14136;
wire n14137;
wire n14138;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14146;
wire n14147;
wire n14148;
wire n14149;
wire n14150;
wire n14151;
wire n14152;
wire n14153;
wire n14154;
wire n14155;
wire n14156;
wire n14157;
wire n14158;
wire n14159;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14164;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14170;
wire n14171;
wire n14172;
wire n14173;
wire n14174;
wire n14175;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14192;
wire n14193;
wire n14194;
wire n14195;
wire n14196;
wire n14197;
wire n14198;
wire n14199;
wire n14200;
wire n14201;
wire n14202;
wire n14203;
wire n14204;
wire n14205;
wire n14206;
wire n14207;
wire n14208;
wire n14209;
wire n14210;
wire n14211;
wire n14212;
wire n14213;
wire n14214;
wire n14215;
wire n14216;
wire n14217;
wire n14218;
wire n14219;
wire n14220;
wire n14221;
wire n14222;
wire n14223;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14233;
wire n14234;
wire n14235;
wire n14236;
wire n14237;
wire n14238;
wire n14239;
wire n14240;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n14250;
wire n14251;
wire n14252;
wire n14253;
wire n14254;
wire n14255;
wire n14256;
wire n14257;
wire n14258;
wire n14259;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14265;
wire n14266;
wire n14267;
wire n14268;
wire n14269;
wire n14270;
wire n14271;
wire n14272;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14278;
wire n14279;
wire n14280;
wire n14281;
wire n14282;
wire n14283;
wire n14284;
wire n14285;
wire n14286;
wire n14287;
wire n14288;
wire n14289;
wire n14290;
wire n14291;
wire n14292;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n14300;
wire n14301;
wire n14302;
wire n14303;
wire n14304;
wire n14305;
wire n14306;
wire n14307;
wire n14308;
wire n14309;
wire n14310;
wire n14311;
wire n14312;
wire n14313;
wire n14314;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14320;
wire n14321;
wire n14322;
wire n14323;
wire n14324;
wire n14325;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14332;
wire n14333;
wire n14334;
wire n14335;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14341;
wire n14342;
wire n14343;
wire n14344;
wire n14345;
wire n14346;
wire n14347;
wire n14348;
wire n14349;
wire n14350;
wire n14351;
wire n14352;
wire n14353;
wire n14354;
wire n14355;
wire n14356;
wire n14357;
wire n14358;
wire n14359;
wire n14360;
wire n14361;
wire n14362;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14369;
wire n14370;
wire n14371;
wire n14372;
wire n14373;
wire n14374;
wire n14375;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14390;
wire n14391;
wire n14392;
wire n14393;
wire n14394;
wire n14395;
wire n14396;
wire n14397;
wire n14398;
wire n14399;
wire n14400;
wire n14401;
wire n14402;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14407;
wire n14408;
wire n14409;
wire n14410;
wire n14411;
wire n14412;
wire n14413;
wire n14414;
wire n14415;
wire n14416;
wire n14417;
wire n14418;
wire n14419;
wire n14420;
wire n14421;
wire n14422;
wire n14423;
wire n14424;
wire n14425;
wire n14426;
wire n14427;
wire n14428;
wire n14429;
wire n14430;
wire n14431;
wire n14432;
wire n14433;
wire n14434;
wire n14435;
wire n14436;
wire n14437;
wire n14438;
wire n14439;
wire n14440;
wire n14441;
wire n14442;
wire n14443;
wire n14444;
wire n14445;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14453;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n14460;
wire n14461;
wire n14462;
wire n14463;
wire n14464;
wire n14465;
wire n14466;
wire n14467;
wire n14468;
wire n14469;
wire n14470;
wire n14471;
wire n14472;
wire n14473;
wire n14474;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14480;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14486;
wire n14487;
wire n14488;
wire n14489;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14501;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14507;
wire n14508;
wire n14509;
wire n14510;
wire n14511;
wire n14512;
wire n14513;
wire n14514;
wire n14515;
wire n14516;
wire n14517;
wire n14518;
wire n14519;
wire n14520;
wire n14521;
wire n14522;
wire n14523;
wire n14524;
wire n14525;
wire n14526;
wire n14527;
wire n14528;
wire n14529;
wire n14530;
wire n14531;
wire n14532;
wire n14533;
wire n14534;
wire n14535;
wire n14536;
wire n14537;
wire n14538;
wire n14539;
wire n14540;
wire n14541;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14546;
wire n14547;
wire n14548;
wire n14549;
wire n14550;
wire n14551;
wire n14552;
wire n14553;
wire n14554;
wire n14555;
wire n14556;
wire n14557;
wire n14558;
wire n14559;
wire n14560;
wire n14561;
wire n14562;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14568;
wire n14569;
wire n14570;
wire n14571;
wire n14572;
wire n14573;
wire n14574;
wire n14575;
wire n14576;
wire n14577;
wire n14578;
wire n14579;
wire n14580;
wire n14581;
wire n14582;
wire n14583;
wire n14584;
wire n14585;
wire n14586;
wire n14587;
wire n14588;
wire n14589;
wire n14590;
wire n14591;
wire n14592;
wire n14593;
wire n14594;
wire n14595;
wire n14596;
wire n14597;
wire n14598;
wire n14599;
wire n14600;
wire n14601;
wire n14602;
wire n14603;
wire n14604;
wire n14605;
wire n14606;
wire n14607;
wire n14608;
wire n14609;
wire n14610;
wire n14611;
wire n14612;
wire n14613;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14618;
wire n14619;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14624;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n14640;
wire n14641;
wire n14642;
wire n14643;
wire n14644;
wire n14645;
wire n14646;
wire n14647;
wire n14648;
wire n14649;
wire n14650;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14657;
wire n14658;
wire n14659;
wire n14660;
wire n14661;
wire n14662;
wire n14663;
wire n14664;
wire n14665;
wire n14666;
wire n14667;
wire n14668;
wire n14669;
wire n14670;
wire n14671;
wire n14672;
wire n14673;
wire n14674;
wire n14675;
wire n14676;
wire n14677;
wire n14678;
wire n14679;
wire n14680;
wire n14681;
wire n14682;
wire n14683;
wire n14684;
wire n14685;
wire n14686;
wire n14687;
wire n14688;
wire n14689;
wire n14690;
wire n14691;
wire n14692;
wire n14693;
wire n14694;
wire n14695;
wire n14696;
wire n14697;
wire n14698;
wire n14699;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14707;
wire n14708;
wire n14709;
wire n14710;
wire n14711;
wire n14712;
wire n14713;
wire n14714;
wire n14715;
wire n14716;
wire n14717;
wire n14718;
wire n14719;
wire n14720;
wire n14721;
wire n14722;
wire n14723;
wire n14724;
wire n14725;
wire n14726;
wire n14727;
wire n14728;
wire n14729;
wire n14730;
wire n14731;
wire n14732;
wire n14733;
wire n14734;
wire n14735;
wire n14736;
wire n14737;
wire n14738;
wire n14739;
wire n14740;
wire n14741;
wire n14742;
wire n14743;
wire n14744;
wire n14745;
wire n14746;
wire n14747;
wire n14748;
wire n14749;
wire n14750;
wire n14751;
wire n14752;
wire n14753;
wire n14754;
wire n14755;
wire n14756;
wire n14757;
wire n14758;
wire n14759;
wire n14760;
wire n14761;
wire n14762;
wire n14763;
wire n14764;
wire n14765;
wire n14766;
wire n14767;
wire n14768;
wire n14769;
wire n14770;
wire n14771;
wire n14772;
wire n14773;
wire n14774;
wire n14775;
wire n14776;
wire n14777;
wire n14778;
wire n14779;
wire n14780;
wire n14781;
wire n14782;
wire n14783;
wire n14784;
wire n14785;
wire n14786;
wire n14787;
wire n14788;
wire n14789;
wire n14790;
wire n14791;
wire n14792;
wire n14793;
wire n14794;
wire n14795;
wire n14796;
wire n14797;
wire n14798;
wire n14799;
wire n14800;
wire n14801;
wire n14802;
wire n14803;
wire n14804;
wire n14805;
wire n14806;
wire n14807;
wire n14808;
wire n14809;
wire n14810;
wire n14811;
wire n14812;
wire n14813;
wire n14814;
wire n14815;
wire n14816;
wire n14817;
wire n14818;
wire n14819;
wire n14820;
wire n14821;
wire n14822;
wire n14823;
wire n14824;
wire n14825;
wire n14826;
wire n14827;
wire n14828;
wire n14829;
wire n14830;
wire n14831;
wire n14832;
wire n14833;
wire n14834;
wire n14835;
wire n14836;
wire n14837;
wire n14838;
wire n14839;
wire n14840;
wire n14841;
wire n14842;
wire n14843;
wire n14844;
wire n14845;
wire n14846;
wire n14847;
wire n14848;
wire n14849;
wire n14850;
wire n14851;
wire n14852;
wire n14853;
wire n14854;
wire n14855;
wire n14856;
wire n14857;
wire n14858;
wire n14859;
wire n14860;
wire n14861;
wire n14862;
wire n14863;
wire n14864;
wire n14865;
wire n14866;
wire n14867;
wire n14868;
wire n14869;
wire n14870;
wire n14871;
wire n14872;
wire n14873;
wire n14874;
wire n14875;
wire n14876;
wire n14877;
wire n14878;
wire n14879;
wire n14880;
wire n14881;
wire n14882;
wire n14883;
wire n14884;
wire n14885;
wire n14886;
wire n14887;
wire n14888;
wire n14889;
wire n14890;
wire n14891;
wire n14892;
wire n14893;
wire n14894;
wire n14895;
wire n14896;
wire n14897;
wire n14898;
wire n14899;
wire n14900;
wire n14901;
wire n14902;
wire n14903;
wire n14904;
wire n14905;
wire n14906;
wire n14907;
wire n14908;
wire n14909;
wire n14910;
wire n14911;
wire n14912;
wire n14913;
wire n14914;
wire n14915;
wire n14916;
wire n14917;
wire n14918;
wire n14919;
wire n14920;
wire n14921;
wire n14922;
wire n14923;
wire n14924;
wire n14925;
wire n14926;
wire n14927;
wire n14928;
wire n14929;
wire n14930;
wire n14931;
wire n14932;
wire n14933;
wire n14934;
wire n14935;
wire n14936;
wire n14937;
wire n14938;
wire n14939;
wire n14940;
wire n14941;
wire n14942;
wire n14943;
wire n14944;
wire n14945;
wire n14946;
wire n14947;
wire n14948;
wire n14949;
wire n14950;
wire n14951;
wire n14952;
wire n14953;
wire n14954;
wire n14955;
wire n14956;
wire n14957;
wire n14958;
wire n14959;
wire n14960;
wire n14961;
wire n14962;
wire n14963;
wire n14964;
wire n14965;
wire n14966;
wire n14967;
wire n14968;
wire n14969;
wire n14970;
wire n14971;
wire n14972;
wire n14973;
wire n14974;
wire n14975;
wire n14976;
wire n14977;
wire n14978;
wire n14979;
wire n14980;
wire n14981;
wire n14982;
wire n14983;
wire n14984;
wire n14985;
wire n14986;
wire n14987;
wire n14988;
wire n14989;
wire n14990;
wire n14991;
wire n14992;
wire n14993;
wire n14994;
wire n14995;
wire n14996;
wire n14997;
wire n14998;
wire n14999;
wire n15000;
wire n15001;
wire n15002;
wire n15003;
wire n15004;
wire n15005;
wire n15006;
wire n15007;
wire n15008;
wire n15009;
wire n15010;
wire n15011;
wire n15012;
wire n15013;
wire n15014;
wire n15015;
wire n15016;
wire n15017;
wire n15018;
wire n15019;
wire n15020;
wire n15021;
wire n15022;
wire n15023;
wire n15024;
wire n15025;
wire n15026;
wire n15027;
wire n15028;
wire n15029;
wire n15030;
wire n15031;
wire n15032;
wire n15033;
wire n15034;
wire n15035;
wire n15036;
wire n15037;
wire n15038;
wire n15039;
wire n15040;
wire n15041;
wire n15042;
wire n15043;
wire n15044;
wire n15045;
wire n15046;
wire n15047;
wire n15048;
wire n15049;
wire n15050;
wire n15051;
wire n15052;
wire n15053;
wire n15054;
wire n15055;
wire n15056;
wire n15057;
wire n15058;
wire n15059;
wire n15060;
wire n15061;
wire n15062;
wire n15063;
wire n15064;
wire n15065;
wire n15066;
wire n15067;
wire n15068;
wire n15069;
wire n15070;
wire n15071;
wire n15072;
wire n15073;
wire n15074;
wire n15075;
wire n15076;
wire n15077;
wire n15078;
wire n15079;
wire n15080;
wire n15081;
wire n15082;
wire n15083;
wire n15084;
wire n15085;
wire n15086;
wire n15087;
wire n15088;
wire n15089;
wire n15090;
wire n15091;
wire n15092;
wire n15093;
wire n15094;
wire n15095;
wire n15096;
wire n15097;
wire n15098;
wire n15099;
wire n15100;
wire n15101;
wire n15102;
wire n15103;
wire n15104;
wire n15105;
wire n15106;
wire n15107;
wire n15108;
wire n15109;
wire n15110;
wire n15111;
wire n15112;
wire n15113;
wire n15114;
wire n15115;
wire n15116;
wire n15117;
wire n15118;
wire n15119;
wire n15120;
wire n15121;
wire n15122;
wire n15123;
wire n15124;
wire n15125;
wire n15126;
wire n15127;
wire n15128;
wire n15129;
wire n15130;
wire n15131;
wire n15132;
wire n15133;
wire n15134;
wire n15135;
wire n15136;
wire n15137;
wire n15138;
wire n15139;
wire n15140;
wire n15141;
wire n15142;
wire n15143;
wire n15144;
wire n15145;
wire n15146;
wire n15147;
wire n15148;
wire n15149;
wire n15150;
wire n15151;
wire n15152;
wire n15153;
wire n15154;
wire n15155;
wire n15156;
wire n15157;
wire n15158;
wire n15159;
wire n15160;
wire n15161;
wire n15162;
wire n15163;
wire n15164;
wire n15165;
wire n15166;
wire n15167;
wire n15168;
wire n15169;
wire n15170;
wire n15171;
wire n15172;
wire n15173;
wire n15174;
wire n15175;
wire n15176;
wire n15177;
wire n15178;
wire n15179;
wire n15180;
wire n15181;
wire n15182;
wire n15183;
wire n15184;
wire n15185;
wire n15186;
wire n15187;
wire n15188;
wire n15189;
wire n15190;
wire n15191;
wire n15192;
wire n15193;
wire n15194;
wire n15195;
wire n15196;
wire n15197;
wire n15198;
wire n15199;
wire n15200;
wire n15201;
wire n15202;
wire n15203;
wire n15204;
wire n15205;
wire n15206;
wire n15207;
wire n15208;
wire n15209;
wire n15210;
wire n15211;
wire n15212;
wire n15213;
wire n15214;
wire n15215;
wire n15216;
wire n15217;
wire n15218;
wire n15219;
wire n15220;
wire n15221;
wire n15222;
wire n15223;
wire n15224;
wire n15225;
wire n15226;
wire n15227;
wire n15228;
wire n15229;
wire n15230;
wire n15231;
wire n15232;
wire n15233;
wire n15234;
wire n15235;
wire n15236;
wire n15237;
wire n15238;
wire n15239;
wire n15240;
wire n15241;
wire n15242;
wire n15243;
wire n15244;
wire n15245;
wire n15246;
wire n15247;
wire n15248;
wire n15249;
wire n15250;
wire n15251;
wire n15252;
wire n15253;
wire n15254;
wire n15255;
wire n15256;
wire n15257;
wire n15258;
wire n15259;
wire n15260;
wire n15261;
wire n15262;
wire n15263;
wire n15264;
wire n15265;
wire n15266;
wire n15267;
wire n15268;
wire n15269;
wire n15270;
wire n15271;
wire n15272;
wire n15273;
wire n15274;
wire n15275;
wire n15276;
wire n15277;
wire n15278;
wire n15279;
wire n15280;
wire n15281;
wire n15282;
wire n15283;
wire n15284;
wire n15285;
wire n15286;
wire n15287;
wire n15288;
wire n15289;
wire n15290;
wire n15291;
wire n15292;
wire n15293;
wire n15294;
wire n15295;
wire n15296;
wire n15297;
wire n15298;
wire n15299;
wire n15300;
wire n15301;
wire n15302;
wire n15303;
wire n15304;
wire n15305;
wire n15306;
wire n15307;
wire n15308;
wire n15309;
wire n15310;
wire n15311;
wire n15312;
wire n15313;
wire n15314;
wire n15315;
wire n15316;
wire n15317;
wire n15318;
wire n15319;
wire n15320;
wire n15321;
wire n15322;
wire n15323;
wire n15324;
wire n15325;
wire n15326;
wire n15327;
wire n15328;
wire n15329;
wire n15330;
wire n15331;
wire n15332;
wire n15333;
wire n15334;
wire n15335;
wire n15336;
wire n15337;
wire n15338;
wire n15339;
wire n15340;
wire n15341;
wire n15342;
wire n15343;
wire n15344;
wire n15345;
wire n15346;
wire n15347;
wire n15348;
wire n15349;
wire n15350;
wire n15351;
wire n15352;
wire n15353;
wire n15354;
wire n15355;
wire n15356;
wire n15357;
wire n15358;
wire n15359;
wire n15360;
wire n15361;
wire n15362;
wire n15363;
wire n15364;
wire n15365;
wire n15366;
wire n15367;
wire n15368;
wire n15369;
wire n15370;
wire n15371;
wire n15372;
wire n15373;
wire n15374;
wire n15375;
wire n15376;
wire n15377;
wire n15378;
wire n15379;
wire n15380;
wire n15381;
wire n15382;
wire n15383;
wire n15384;
wire n15385;
wire n15386;
wire n15387;
wire n15388;
wire n15389;
wire n15390;
wire n15391;
wire n15392;
wire n15393;
wire n15394;
wire n15395;
wire n15396;
wire n15397;
wire n15398;
wire n15399;
wire n15400;
wire n15401;
wire n15402;
wire n15403;
wire n15404;
wire n15405;
wire n15406;
wire n15407;
wire n15408;
wire n15409;
wire n15410;
wire n15411;
wire n15412;
wire n15413;
wire n15414;
wire n15415;
wire n15416;
wire n15417;
wire n15418;
wire n15419;
wire n15420;
wire n15421;
wire n15422;
wire n15423;
wire n15424;
wire n15425;
wire n15426;
wire n15427;
wire n15428;
wire n15429;
wire n15430;
wire n15431;
wire n15432;
wire n15433;
wire n15434;
wire n15435;
wire n15436;
wire n15437;
wire n15438;
wire n15439;
wire n15440;
wire n15441;
wire n15442;
wire n15443;
wire n15444;
wire n15445;
wire n15446;
wire n15447;
wire n15448;
wire n15449;
wire n15450;
wire n15451;
wire n15452;
wire n15453;
wire n15454;
wire n15455;
wire n15456;
wire n15457;
wire n15458;
wire n15459;
wire n15460;
wire n15461;
wire n15462;
wire n15463;
wire n15464;
wire n15465;
wire n15466;
wire n15467;
wire n15468;
wire n15469;
wire n15470;
wire n15471;
wire n15472;
wire n15473;
wire n15474;
wire n15475;
wire n15476;
wire n15477;
wire n15478;
wire n15479;
wire n15480;
wire n15481;
wire n15482;
wire n15483;
wire n15484;
wire n15485;
wire n15486;
wire n15487;
wire n15488;
wire n15489;
wire n15490;
wire n15491;
wire n15492;
wire n15493;
wire n15494;
wire n15495;
wire n15496;
wire n15497;
wire n15498;
wire n15499;
wire n15500;
wire n15501;
wire n15502;
wire n15503;
wire n15504;
wire n15505;
wire n15506;
wire n15507;
wire n15508;
wire n15509;
wire n15510;
wire n15511;
wire n15512;
wire n15513;
wire n15514;
wire n15515;
wire n15516;
wire n15517;
wire n15518;
wire n15519;
wire n15520;
wire n15521;
wire n15522;
wire n15523;
wire n15524;
wire n15525;
wire n15526;
wire n15527;
wire n15528;
wire n15529;
wire n15530;
wire n15531;
wire n15532;
wire n15533;
wire n15534;
wire n15535;
wire n15536;
wire n15537;
wire n15538;
wire n15539;
wire n15540;
wire n15541;
wire n15542;
wire n15543;
wire n15544;
wire n15545;
wire n15546;
wire n15547;
wire n15548;
wire n15549;
wire n15550;
wire n15551;
wire n15552;
wire n15553;
wire n15554;
wire n15555;
wire n15556;
wire n15557;
wire n15558;
wire n15559;
wire n15560;
wire n15561;
wire n15562;
wire n15563;
wire n15564;
wire n15565;
wire n15566;
wire n15567;
wire n15568;
wire n15569;
wire n15570;
wire n15571;
wire n15572;
wire n15573;
wire n15574;
wire n15575;
wire n15576;
wire n15577;
wire n15578;
wire n15579;
wire n15580;
wire n15581;
wire n15582;
wire n15583;
wire n15584;
wire n15585;
wire n15586;
wire n15587;
wire n15588;
wire n15589;
wire n15590;
wire n15591;
wire n15592;
wire n15593;
wire n15594;
wire n15595;
wire n15596;
wire n15597;
wire n15598;
wire n15599;
wire n15600;
wire n15601;
wire n15602;
wire n15603;
wire n15604;
wire n15605;
wire n15606;
wire n15607;
wire n15608;
wire n15609;
wire n15610;
wire n15611;
wire n15612;
wire n15613;
wire n15614;
wire n15615;
wire n15616;
wire n15617;
wire n15618;
wire n15619;
wire n15620;
wire n15621;
wire n15622;
wire n15623;
wire n15624;
wire n15625;
wire n15626;
wire n15627;
wire n15628;
wire n15629;
wire n15630;
wire n15631;
wire n15632;
wire n15633;
wire n15634;
wire n15635;
wire n15636;
wire n15637;
wire n15638;
wire n15639;
wire n15640;
wire n15641;
wire n15642;
wire n15643;
wire n15644;
wire n15645;
wire n15646;
wire n15647;
wire n15648;
wire n15649;
wire n15650;
wire n15651;
wire n15652;
wire n15653;
wire n15654;
wire n15655;
wire n15656;
wire n15657;
wire n15658;
wire n15659;
wire n15660;
wire n15661;
wire n15662;
wire n15663;
wire n15664;
wire n15665;
wire n15666;
wire n15667;
wire n15668;
wire n15669;
wire n15670;
wire n15671;
wire n15672;
wire n15673;
wire n15674;
wire n15675;
wire n15676;
wire n15677;
wire n15678;
wire n15679;
wire n15680;
wire n15681;
wire n15682;
wire n15683;
wire n15684;
wire n15685;
wire n15686;
wire n15687;
wire n15688;
wire n15689;
wire n15690;
wire n15691;
wire n15692;
wire n15693;
wire n15694;
wire n15695;
wire n15696;
wire n15697;
wire n15698;
wire n15699;
wire n15700;
wire n15701;
wire n15702;
wire n15703;
wire n15704;
wire n15705;
wire n15706;
wire n15707;
wire n15708;
wire n15709;
wire n15710;
wire n15711;
wire n15712;
wire n15713;
wire n15714;
wire n15715;
wire n15716;
wire n15717;
wire n15718;
wire n15719;
wire n15720;
wire n15721;
wire n15722;
wire n15723;
wire n15724;
wire n15725;
wire n15726;
wire n15727;
wire n15728;
wire n15729;
wire n15730;
wire n15731;
wire n15732;
wire n15733;
wire n15734;
wire n15735;
wire n15736;
wire n15737;
wire n15738;
wire n15739;
wire n15740;
wire n15741;
wire n15742;
wire n15743;
wire n15744;
wire n15745;
wire n15746;
wire n15747;
wire n15748;
wire n15749;
wire n15750;
wire n15751;
wire n15752;
wire n15753;
wire n15754;
wire n15755;
wire n15756;
wire n15757;
wire n15758;
wire n15759;
wire n15760;
wire n15761;
wire n15762;
wire n15763;
wire n15764;
wire n15765;
wire n15766;
wire n15767;
wire n15768;
wire n15769;
wire n15770;
wire n15771;
wire n15772;
wire n15773;
wire n15774;
wire n15775;
wire n15776;
wire n15777;
wire n15778;
wire n15779;
wire n15780;
wire n15781;
wire n15782;
wire n15783;
wire n15784;
wire n15785;
wire n15786;
wire n15787;
wire n15788;
wire n15789;
wire n15790;
wire n15791;
wire n15792;
wire n15793;
wire n15794;
wire n15795;
wire n15796;
wire n15797;
wire n15798;
wire n15799;
wire n15800;
wire n15801;
wire n15802;
wire n15803;
wire n15804;
wire n15805;
wire n15806;
wire n15807;
wire n15808;
wire n15809;
wire n15810;
wire n15811;
wire n15812;
wire n15813;
wire n15814;
wire n15815;
wire n15816;
wire n15817;
wire n15818;
wire n15819;
wire n15820;
wire n15821;
wire n15822;
wire n15823;
wire n15824;
wire n15825;
wire n15826;
wire n15827;
wire n15828;
wire n15829;
wire n15830;
wire n15831;
wire n15832;
wire n15833;
wire n15834;
wire n15835;
wire n15836;
wire n15837;
wire n15838;
wire n15839;
wire n15840;
wire n15841;
wire n15842;
wire n15843;
wire n15844;
wire n15845;
wire n15846;
wire n15847;
wire n15848;
wire n15849;
wire n15850;
wire n15851;
wire n15852;
wire n15853;
wire n15854;
wire n15855;
wire n15856;
wire n15857;
wire n15858;
wire n15859;
wire n15860;
wire n15861;
wire n15862;
wire n15863;
wire n15864;
wire n15865;
wire n15866;
wire n15867;
wire n15868;
wire n15869;
wire n15870;
wire n15871;
wire n15872;
wire n15873;
wire n15874;
wire n15875;
wire n15876;
wire n15877;
wire n15878;
wire n15879;
wire n15880;
wire n15881;
wire n15882;
wire n15883;
wire n15884;
wire n15885;
wire n15886;
wire n15887;
wire n15888;
wire n15889;
wire n15890;
wire n15891;
wire n15892;
wire n15893;
wire n15894;
wire n15895;
wire n15896;
wire n15897;
wire n15898;
wire n15899;
wire n15900;
wire n15901;
wire n15902;
wire n15903;
wire n15904;
wire n15905;
wire n15906;
wire n15907;
wire n15908;
wire n15909;
wire n15910;
wire n15911;
wire n15912;
wire n15913;
wire n15914;
wire n15915;
wire n15916;
wire n15917;
wire n15918;
wire n15919;
wire n15920;
wire n15921;
wire n15922;
wire n15923;
wire n15924;
wire n15925;
wire n15926;
wire n15927;
wire n15928;
wire n15929;
wire n15930;
wire n15931;
wire n15932;
wire n15933;
wire n15934;
wire n15935;
wire n15936;
wire n15937;
wire n15938;
wire n15939;
wire n15940;
wire n15941;
wire n15942;
wire n15943;
wire n15944;
wire n15945;
wire n15946;
wire n15947;
wire n15948;
wire n15949;
wire n15950;
wire n15951;
wire n15952;
wire n15953;
wire n15954;
wire n15955;
wire n15956;
wire n15957;
wire n15958;
wire n15959;
wire n15960;
wire n15961;
wire n15962;
wire n15963;
wire n15964;
wire n15965;
wire n15966;
wire n15967;
wire n15968;
wire n15969;
wire n15970;
wire n15971;
wire n15972;
wire n15973;
wire n15974;
wire n15975;
wire n15976;
wire n15977;
wire n15978;
wire n15979;
wire n15980;
wire n15981;
wire n15982;
wire n15983;
wire n15984;
wire n15985;
wire n15986;
wire n15987;
wire n15988;
wire n15989;
wire n15990;
wire n15991;
wire n15992;
wire n15993;
wire n15994;
wire n15995;
wire n15996;
wire n15997;
wire n15998;
wire n15999;
wire n16000;
wire n16001;
wire n16002;
wire n16003;
wire n16004;
wire n16005;
wire n16006;
wire n16007;
wire n16008;
wire n16009;
wire n16010;
wire n16011;
wire n16012;
wire n16013;
wire n16014;
wire n16015;
wire n16016;
wire n16017;
wire n16018;
wire n16019;
wire n16020;
wire n16021;
wire n16022;
wire n16023;
wire n16024;
wire n16025;
wire n16026;
wire n16027;
wire n16028;
wire n16029;
wire n16030;
wire n16031;
wire n16032;
wire n16033;
wire n16034;
wire n16035;
wire n16036;
wire n16037;
wire n16038;
wire n16039;
wire n16040;
wire n16041;
wire n16042;
wire n16043;
wire n16044;
wire n16045;
wire n16046;
wire n16047;
wire n16048;
wire n16049;
wire n16050;
wire n16051;
wire n16052;
wire n16053;
wire n16054;
wire n16055;
wire n16056;
wire n16057;
wire n16058;
wire n16059;
wire n16060;
wire n16061;
wire n16062;
wire n16063;
wire n16064;
wire n16065;
wire n16066;
wire n16067;
wire n16068;
wire n16069;
wire n16070;
wire n16071;
wire n16072;
wire n16073;
wire n16074;
wire n16075;
wire n16076;
wire n16077;
wire n16078;
wire n16079;
wire n16080;
wire n16081;
wire n16082;
wire n16083;
wire n16084;
wire n16085;
wire n16086;
wire n16087;
wire n16088;
wire n16089;
wire n16090;
wire n16091;
wire n16092;
wire n16093;
wire n16094;
wire n16095;
wire n16096;
wire n16097;
wire n16098;
wire n16099;
wire n16100;
wire n16101;
wire n16102;
wire n16103;
wire n16104;
wire n16105;
wire n16106;
wire n16107;
wire n16108;
wire n16109;
wire n16110;
wire n16111;
wire n16112;
wire n16113;
wire n16114;
wire n16115;
wire n16116;
wire n16117;
wire n16118;
wire n16119;
wire n16120;
wire n16121;
wire n16122;
wire n16123;
wire n16124;
wire n16125;
wire n16126;
wire n16127;
wire n16128;
wire n16129;
wire n16130;
wire n16131;
wire n16132;
wire n16133;
wire n16134;
wire n16135;
wire n16136;
wire n16137;
wire n16138;
wire n16139;
wire n16140;
wire n16141;
wire n16142;
wire n16143;
wire n16144;
wire n16145;
wire n16146;
wire n16147;
wire n16148;
wire n16149;
wire n16150;
wire n16151;
wire n16152;
wire n16153;
wire n16154;
wire n16155;
wire n16156;
wire n16157;
wire n16158;
wire n16159;
wire n16160;
wire n16161;
wire n16162;
wire n16163;
wire n16164;
wire n16165;
wire n16166;
wire n16167;
wire n16168;
wire n16169;
wire n16170;
wire n16171;
wire n16172;
wire n16173;
wire n16174;
wire n16175;
wire n16176;
wire n16177;
wire n16178;
wire n16179;
wire n16180;
wire n16181;
wire n16182;
wire n16183;
wire n16184;
wire n16185;
wire n16186;
wire n16187;
wire n16188;
wire n16189;
wire n16190;
wire n16191;
wire n16192;
wire n16193;
wire n16194;
wire n16195;
wire n16196;
wire n16197;
wire n16198;
wire n16199;
wire n16200;
wire n16201;
wire n16202;
wire n16203;
wire n16204;
wire n16205;
wire n16206;
wire n16207;
wire n16208;
wire n16209;
wire n16210;
wire n16211;
wire n16212;
wire n16213;
wire n16214;
wire n16215;
wire n16216;
wire n16217;
wire n16218;
wire n16219;
wire n16220;
wire n16221;
wire n16222;
wire n16223;
wire n16224;
wire n16225;
wire n16226;
wire n16227;
wire n16228;
wire n16229;
wire n16230;
wire n16231;
wire n16232;
wire n16233;
wire n16234;
wire n16235;
wire n16236;
wire n16237;
wire n16238;
wire n16239;
wire n16240;
wire n16241;
wire n16242;
wire n16243;
wire n16244;
wire n16245;
wire n16246;
wire n16247;
wire n16248;
wire n16249;
wire n16250;
wire n16251;
wire n16252;
wire n16253;
wire n16254;
wire n16255;
wire n16256;
wire n16257;
wire n16258;
wire n16259;
wire n16260;
wire n16261;
wire n16262;
wire n16263;
wire n16264;
wire n16265;
wire n16266;
wire n16267;
wire n16268;
wire n16269;
wire n16270;
wire n16271;
wire n16272;
wire n16273;
wire n16274;
wire n16275;
wire n16276;
wire n16277;
wire n16278;
wire n16279;
wire n16280;
wire n16281;
wire n16282;
wire n16283;
wire n16284;
wire n16285;
wire n16286;
wire n16287;
wire n16288;
wire n16289;
wire n16290;
wire n16291;
wire n16292;
wire n16293;
wire n16294;
wire n16295;
wire n16296;
wire n16297;
wire n16298;
wire n16299;
wire n16300;
wire n16301;
wire n16302;
wire n16303;
wire n16304;
wire n16305;
wire n16306;
wire n16307;
wire n16308;
wire n16309;
wire n16310;
wire n16311;
wire n16312;
wire n16313;
wire n16314;
wire n16315;
wire n16316;
wire n16317;
wire n16318;
wire n16319;
wire n16320;
wire n16321;
wire n16322;
wire n16323;
wire n16324;
wire n16325;
wire n16326;
wire n16327;
wire n16328;
wire n16329;
wire n16330;
wire n16331;
wire n16332;
wire n16333;
wire n16334;
wire n16335;
wire n16336;
wire n16337;
wire n16338;
wire n16339;
wire n16340;
wire n16341;
wire n16342;
wire n16343;
wire n16344;
wire n16345;
wire n16346;
wire n16347;
wire n16348;
wire n16349;
wire n16350;
wire n16351;
wire n16352;
wire n16353;
wire n16354;
wire n16355;
wire n16356;
wire n16357;
wire n16358;
wire n16359;
wire n16360;
wire n16361;
wire n16362;
wire n16363;
wire n16364;
wire n16365;
wire n16366;
wire n16367;
wire n16368;
wire n16369;
wire n16370;
wire n16371;
wire n16372;
wire n16373;
wire n16374;
wire n16375;
wire n16376;
wire n16377;
wire n16378;
wire n16379;
wire n16380;
wire n16381;
wire n16382;
wire n16383;
wire n16384;
wire n16385;
wire n16386;
wire n16387;
wire n16388;
wire n16389;
wire n16390;
wire n16391;
wire n16392;
wire n16393;
wire n16394;
wire n16395;
wire n16396;
wire n16397;
wire n16398;
wire n16399;
wire n16400;
wire n16401;
wire n16402;
wire n16403;
wire n16404;
wire n16405;
wire n16406;
wire n16407;
wire n16408;
wire n16409;
wire n16410;
wire n16411;
wire n16412;
wire n16413;
wire n16414;
wire n16415;
wire n16416;
wire n16417;
wire n16418;
wire n16419;
wire n16420;
wire n16421;
wire n16422;
wire n16423;
wire n16424;
wire n16425;
wire n16426;
wire n16427;
wire n16428;
wire n16429;
wire n16430;
wire n16431;
wire n16432;
wire n16433;
wire n16434;
wire n16435;
wire n16436;
wire n16437;
wire n16438;
wire n16439;
wire n16440;
wire n16441;
wire n16442;
wire n16443;
wire n16444;
wire n16445;
wire n16446;
wire n16447;
wire n16448;
wire n16449;
wire n16450;
wire n16451;
wire n16452;
wire n16453;
wire n16454;
wire n16455;
wire n16456;
wire n16457;
wire n16458;
wire n16459;
wire n16460;
wire n16461;
wire n16462;
wire n16463;
wire n16464;
wire n16465;
wire n16466;
wire n16467;
wire n16468;
wire n16469;
wire n16470;
wire n16471;
wire n16472;
wire n16473;
wire n16474;
wire n16475;
wire n16476;
wire n16477;
wire n16478;
wire n16479;
wire n16480;
wire n16481;
wire n16482;
wire n16483;
wire n16484;
wire n16485;
wire n16486;
wire n16487;
wire n16488;
wire n16489;
wire n16490;
wire n16491;
wire n16492;
wire n16493;
wire n16494;
wire n16495;
wire n16496;
wire n16497;
wire n16498;
wire n16499;
wire n16500;
wire n16501;
wire n16502;
wire n16503;
wire n16504;
wire n16505;
wire n16506;
wire n16507;
wire n16508;
wire n16509;
wire n16510;
wire n16511;
wire n16512;
wire n16513;
wire n16514;
wire n16515;
wire n16516;
wire n16517;
wire n16518;
wire n16519;
wire n16520;
wire n16521;
wire n16522;
wire n16523;
wire n16524;
wire n16525;
wire n16526;
wire n16527;
wire n16528;
wire n16529;
wire n16530;
wire n16531;
wire n16532;
wire n16533;
wire n16534;
wire n16535;
wire n16536;
wire n16537;
wire n16538;
wire n16539;
wire n16540;
wire n16541;
wire n16542;
wire n16543;
wire n16544;
wire n16545;
wire n16546;
wire n16547;
wire n16548;
wire n16549;
wire n16550;
wire n16551;
wire n16552;
wire n16553;
wire n16554;
wire n16555;
wire n16556;
wire n16557;
wire n16558;
wire n16559;
wire n16560;
wire n16561;
wire n16562;
wire n16563;
wire n16564;
wire n16565;
wire n16566;
wire n16567;
wire n16568;
wire n16569;
wire n16570;
wire n16571;
wire n16572;
wire n16573;
wire n16574;
wire n16575;
wire n16576;
wire n16577;
wire n16578;
wire n16579;
wire n16580;
wire n16581;
wire n16582;
wire n16583;
wire n16584;
wire n16585;
wire n16586;
wire n16587;
wire n16588;
wire n16589;
wire n16590;
wire n16591;
wire n16592;
wire n16593;
wire n16594;
wire n16595;
wire n16596;
wire n16597;
wire n16598;
wire n16599;
wire n16600;
wire n16601;
wire n16602;
wire n16603;
wire n16604;
wire n16605;
wire n16606;
wire n16607;
wire n16608;
wire n16609;
wire n16610;
wire n16611;
wire n16612;
wire n16613;
wire n16614;
wire n16615;
wire n16616;
wire n16617;
wire n16618;
wire n16619;
wire n16620;
wire n16621;
wire n16622;
wire n16623;
wire n16624;
wire n16625;
wire n16626;
wire n16627;
wire n16628;
wire n16629;
wire n16630;
wire n16631;
wire n16632;
wire n16633;
wire n16634;
wire n16635;
wire n16636;
wire n16637;
wire n16638;
wire n16639;
wire n16640;
wire n16641;
wire n16642;
wire n16643;
wire n16644;
wire n16645;
wire n16646;
wire n16647;
wire n16648;
wire n16649;
wire n16650;
wire n16651;
wire n16652;
wire n16653;
wire n16654;
wire n16655;
wire n16656;
wire n16657;
wire n16658;
wire n16659;
wire n16660;
wire n16661;
wire n16662;
wire n16663;
wire n16664;
wire n16665;
wire n16666;
wire n16667;
wire n16668;
wire n16669;
wire n16670;
wire n16671;
wire n16672;
wire n16673;
wire n16674;
wire n16675;
wire n16676;
wire n16677;
wire n16678;
wire n16679;
wire n16680;
wire n16681;
wire n16682;
wire n16683;
wire n16684;
wire n16685;
wire n16686;
wire n16687;
wire n16688;
wire n16689;
wire n16690;
wire n16691;
wire n16692;
wire n16693;
wire n16694;
wire n16695;
wire n16696;
wire n16697;
wire n16698;
wire n16699;
wire n16700;
wire n16701;
wire n16702;
wire n16703;
wire n16704;
wire n16705;
wire n16706;
wire n16707;
wire n16708;
wire n16709;
wire n16710;
wire n16711;
wire n16712;
wire n16713;
wire n16714;
wire n16715;
wire n16716;
wire n16717;
wire n16718;
wire n16719;
wire n16720;
wire n16721;
wire n16722;
wire n16723;
wire n16724;
wire n16725;
wire n16726;
wire n16727;
wire n16728;
wire n16729;
wire n16730;
wire n16731;
wire n16732;
wire n16733;
wire n16734;
wire n16735;
wire n16736;
wire n16737;
wire n16738;
wire n16739;
wire n16740;
wire n16741;
wire n16742;
wire n16743;
wire n16744;
wire n16745;
wire n16746;
wire n16747;
wire n16748;
wire n16749;
wire n16750;
wire n16751;
wire n16752;
wire n16753;
wire n16754;
wire n16755;
wire n16756;
wire n16757;
wire n16758;
wire n16759;
wire n16760;
wire n16761;
wire n16762;
wire n16763;
wire n16764;
wire n16765;
wire n16766;
wire n16767;
wire n16768;
wire n16769;
wire n16770;
wire n16771;
wire n16772;
wire n16773;
wire n16774;
wire n16775;
wire n16776;
wire n16777;
wire n16778;
wire n16779;
wire n16780;
wire n16781;
wire n16782;
wire n16783;
wire n16784;
wire n16785;
wire n16786;
wire n16787;
wire n16788;
wire n16789;
wire n16790;
wire n16791;
wire n16792;
wire n16793;
wire n16794;
wire n16795;
wire n16796;
wire n16797;
wire n16798;
wire n16799;
wire n16800;
wire n16801;
wire n16802;
wire n16803;
wire n16804;
wire n16805;
wire n16806;
wire n16807;
wire n16808;
wire n16809;
wire n16810;
wire n16811;
wire n16812;
wire n16813;
wire n16814;
wire n16815;
wire n16816;
wire n16817;
wire n16818;
wire n16819;
wire n16820;
wire n16821;
wire n16822;
wire n16823;
wire n16824;
wire n16825;
wire n16826;
wire n16827;
wire n16828;
wire n16829;
wire n16830;
wire n16831;
wire n16832;
wire n16833;
wire n16834;
wire n16835;
wire n16836;
wire n16837;
wire n16838;
wire n16839;
wire n16840;
wire n16841;
wire n16842;
wire n16843;
wire n16844;
wire n16845;
wire n16846;
wire n16847;
wire n16848;
wire n16849;
wire n16850;
wire n16851;
wire n16852;
wire n16853;
wire n16854;
wire n16855;
wire n16856;
wire n16857;
wire n16858;
wire n16859;
wire n16860;
wire n16861;
wire n16862;
wire n16863;
wire n16864;
wire n16865;
wire n16866;
wire n16867;
wire n16868;
wire n16869;
wire n16870;
wire n16871;
wire n16872;
wire n16873;
wire n16874;
wire n16875;
wire n16876;
wire n16877;
wire n16878;
wire n16879;
wire n16880;
wire n16881;
wire n16882;
wire n16883;
wire n16884;
wire n16885;
wire n16886;
wire n16887;
wire n16888;
wire n16889;
wire n16890;
wire n16891;
wire n16892;
wire n16893;
wire n16894;
wire n16895;
wire n16896;
wire n16897;
wire n16898;
wire n16899;
wire n16900;
wire n16901;
wire n16902;
wire n16903;
wire n16904;
wire n16905;
wire n16906;
wire n16907;
wire n16908;
wire n16909;
wire n16910;
wire n16911;
wire n16912;
wire n16913;
wire n16914;
wire n16915;
wire n16916;
wire n16917;
wire n16918;
wire n16919;
wire n16920;
wire n16921;
wire n16922;
wire n16923;
wire n16924;
wire n16925;
wire n16926;
wire n16927;
wire n16928;
wire n16929;
wire n16930;
wire n16931;
wire n16932;
wire n16933;
wire n16934;
wire n16935;
wire n16936;
wire n16937;
wire n16938;
wire n16939;
wire n16940;
wire n16941;
wire n16942;
wire n16943;
wire n16944;
wire n16945;
wire n16946;
wire n16947;
wire n16948;
wire n16949;
wire n16950;
wire n16951;
wire n16952;
wire n16953;
wire n16954;
wire n16955;
wire n16956;
wire n16957;
wire n16958;
wire n16959;
wire n16960;
wire n16961;
wire n16962;
wire n16963;
wire n16964;
wire n16965;
wire n16966;
wire n16967;
wire n16968;
wire n16969;
wire n16970;
wire n16971;
wire n16972;
wire n16973;
wire n16974;
wire n16975;
wire n16976;
wire n16977;
wire n16978;
wire n16979;
wire n16980;
wire n16981;
wire n16982;
wire n16983;
wire n16984;
wire n16985;
wire n16986;
wire n16987;
wire n16988;
wire n16989;
wire n16990;
wire n16991;
wire n16992;
wire n16993;
wire n16994;
wire n16995;
wire n16996;
wire n16997;
wire n16998;
wire n16999;
wire n17000;
wire n17001;
wire n17002;
wire n17003;
wire n17004;
wire n17005;
wire n17006;
wire n17007;
wire n17008;
wire n17009;
wire n17010;
wire n17011;
wire n17012;
wire n17013;
wire n17014;
wire n17015;
wire n17016;
wire n17017;
wire n17018;
wire n17019;
wire n17020;
wire n17021;
wire n17022;
wire n17023;
wire n17024;
wire n17025;
wire n17026;
wire n17027;
wire n17028;
wire n17029;
wire n17030;
wire n17031;
wire n17032;
wire n17033;
wire n17034;
wire n17035;
wire n17036;
wire n17037;
wire n17038;
wire n17039;
wire n17040;
wire n17041;
wire n17042;
wire n17043;
wire n17044;
wire n17045;
wire n17046;
wire n17047;
wire n17048;
wire n17049;
wire n17050;
wire n17051;
wire n17052;
wire n17053;
wire n17054;
wire n17055;
wire n17056;
wire n17057;
wire n17058;
wire n17059;
wire n17060;
wire n17061;
wire n17062;
wire n17063;
wire n17064;
wire n17065;
wire n17066;
wire n17067;
wire n17068;
wire n17069;
wire n17070;
wire n17071;
wire n17072;
wire n17073;
wire n17074;
wire n17075;
wire n17076;
wire n17077;
wire n17078;
wire n17079;
wire n17080;
wire n17081;
wire n17082;
wire n17083;
wire n17084;
wire n17085;
wire n17086;
wire n17087;
wire n17088;
wire n17089;
wire n17090;
wire n17091;
wire n17092;
wire n17093;
wire n17094;
wire n17095;
wire n17096;
wire n17097;
wire n17098;
wire n17099;
wire n17100;
wire n17101;
wire n17102;
wire n17103;
wire n17104;
wire n17105;
wire n17106;
wire n17107;
wire n17108;
wire n17109;
wire n17110;
wire n17111;
wire n17112;
wire n17113;
wire n17114;
wire n17115;
wire n17116;
wire n17117;
wire n17118;
wire n17119;
wire n17120;
wire n17121;
wire n17122;
wire n17123;
wire n17124;
wire n17125;
wire n17126;
wire n17127;
wire n17128;
wire n17129;
wire n17130;
wire n17131;
wire n17132;
wire n17133;
wire n17134;
wire n17135;
wire n17136;
wire n17137;
wire n17138;
wire n17139;
wire n17140;
wire n17141;
wire n17142;
wire n17143;
wire n17144;
wire n17145;
wire n17146;
wire n17147;
wire n17148;
wire n17149;
wire n17150;
wire n17151;
wire n17152;
wire n17153;
wire n17154;
wire n17155;
wire n17156;
wire n17157;
wire n17158;
wire n17159;
wire n17160;
wire n17161;
wire n17162;
wire n17163;
wire n17164;
wire n17165;
wire n17166;
wire n17167;
wire n17168;
wire n17169;
wire n17170;
wire n17171;
wire n17172;
wire n17173;
wire n17174;
wire n17175;
wire n17176;
wire n17177;
wire n17178;
wire n17179;
wire n17180;
wire n17181;
wire n17182;
wire n17183;
wire n17184;
wire n17185;
wire n17186;
wire n17187;
wire n17188;
wire n17189;
wire n17190;
wire n17191;
wire n17192;
wire n17193;
wire n17194;
wire n17195;
wire n17196;
wire n17197;
wire n17198;
wire n17199;
wire n17200;
wire n17201;
wire n17202;
wire n17203;
wire n17204;
wire n17205;
wire n17206;
wire n17207;
wire n17208;
wire n17209;
wire n17210;
wire n17211;
wire n17212;
wire n17213;
wire n17214;
wire n17215;
wire n17216;
wire n17217;
wire n17218;
wire n17219;
wire n17220;
wire n17221;
wire n17222;
wire n17223;
wire n17224;
wire n17225;
wire n17226;
wire n17227;
wire n17228;
wire n17229;
wire n17230;
wire n17231;
wire n17232;
wire n17233;
wire n17234;
wire n17235;
wire n17236;
wire n17237;
wire n17238;
wire n17239;
wire n17240;
wire n17241;
wire n17242;
wire n17243;
wire n17244;
wire n17245;
wire n17246;
wire n17247;
wire n17248;
wire n17249;
wire n17250;
wire n17251;
wire n17252;
wire n17253;
wire n17254;
wire n17255;
wire n17256;
wire n17257;
wire n17258;
wire n17259;
wire n17260;
wire n17261;
wire n17262;
wire n17263;
wire n17264;
wire n17265;
wire n17266;
wire n17267;
wire n17268;
wire n17269;
wire n17270;
wire n17271;
wire n17272;
wire n17273;
wire n17274;
wire n17275;
wire n17276;
wire n17277;
wire n17278;
wire n17279;
wire n17280;
wire n17281;
wire n17282;
wire n17283;
wire n17284;
wire n17285;
wire n17286;
wire n17287;
wire n17288;
wire n17289;
wire n17290;
wire n17291;
wire n17292;
wire n17293;
wire n17294;
wire n17295;
wire n17296;
wire n17297;
wire n17298;
wire n17299;
wire n17300;
wire n17301;
wire n17302;
wire n17303;
wire n17304;
wire n17305;
wire n17306;
wire n17307;
wire n17308;
wire n17309;
wire n17310;
wire n17311;
wire n17312;
wire n17313;
wire n17314;
wire n17315;
wire n17316;
wire n17317;
wire n17318;
wire n17319;
wire n17320;
wire n17321;
wire n17322;
wire n17323;
wire n17324;
wire n17325;
wire n17326;
wire n17327;
wire n17328;
wire n17329;
wire n17330;
wire n17331;
wire n17332;
wire n17333;
wire n17334;
wire n17335;
wire n17336;
wire n17337;
wire n17338;
wire n17339;
wire n17340;
wire n17341;
wire n17342;
wire n17343;
wire n17344;
wire n17345;
wire n17346;
wire n17347;
wire n17348;
wire n17349;
wire n17350;
wire n17351;
wire n17352;
wire n17353;
wire n17354;
wire n17355;
wire n17356;
wire n17357;
wire n17358;
wire n17359;
wire n17360;
wire n17361;
wire n17362;
wire n17363;
wire n17364;
wire n17365;
wire n17366;
wire n17367;
wire n17368;
wire n17369;
wire n17370;
wire n17371;
wire n17372;
wire n17373;
wire n17374;
wire n17375;
wire n17376;
wire n17377;
wire n17378;
wire n17379;
wire n17380;
wire n17381;
wire n17382;
wire n17383;
wire n17384;
wire n17385;
wire n17386;
wire n17387;
wire n17388;
wire n17389;
wire n17390;
wire n17391;
wire n17392;
wire n17393;
wire n17394;
wire n17395;
wire n17396;
wire n17397;
wire n17398;
wire n17399;
wire n17400;
wire n17401;
wire n17402;
wire n17403;
wire n17404;
wire n17405;
wire n17406;
wire n17407;
wire n17408;
wire n17409;
wire n17410;
wire n17411;
wire n17412;
wire n17413;
wire n17414;
wire n17415;
wire n17416;
wire n17417;
wire n17418;
wire n17419;
wire n17420;
wire n17421;
wire n17422;
wire n17423;
wire n17424;
wire n17425;
wire n17426;
wire n17427;
wire n17428;
wire n17429;
wire n17430;
wire n17431;
wire n17432;
wire n17433;
wire n17434;
wire n17435;
wire n17436;
wire n17437;
wire n17438;
wire n17439;
wire n17440;
wire n17441;
wire n17442;
wire n17443;
wire n17444;
wire n17445;
wire n17446;
wire n17447;
wire n17448;
wire n17449;
wire n17450;
wire n17451;
wire n17452;
wire n17453;
wire n17454;
wire n17455;
wire n17456;
wire n17457;
wire n17458;
wire n17459;
wire n17460;
wire n17461;
wire n17462;
wire n17463;
wire n17464;
wire n17465;
wire n17466;
wire n17467;
wire n17468;
wire n17469;
wire n17470;
wire n17471;
wire n17472;
wire n17473;
wire n17474;
wire n17475;
wire n17476;
wire n17477;
wire n17478;
wire n17479;
wire n17480;
wire n17481;
wire n17482;
wire n17483;
wire n17484;
wire n17485;
wire n17486;
wire n17487;
wire n17488;
wire n17489;
wire n17490;
wire n17491;
wire n17492;
wire n17493;
wire n17494;
wire n17495;
wire n17496;
wire n17497;
wire n17498;
wire n17499;
wire n17500;
wire n17501;
wire n17502;
wire n17503;
wire n17504;
wire n17505;
wire n17506;
wire n17507;
wire n17508;
wire n17509;
wire n17510;
wire n17511;
wire n17512;
wire n17513;
wire n17514;
wire n17515;
wire n17516;
wire n17517;
wire n17518;
wire n17519;
wire n17520;
wire n17521;
wire n17522;
wire n17523;
wire n17524;
wire n17525;
wire n17526;
wire n17527;
wire n17528;
wire n17529;
wire n17530;
wire n17531;
wire n17532;
wire n17533;
wire n17534;
wire n17535;
wire n17536;
wire n17537;
wire n17538;
wire n17539;
wire n17540;
wire n17541;
wire n17542;
wire n17543;
wire n17544;
wire n17545;
wire n17546;
wire n17547;
wire n17548;
wire n17549;
wire n17550;
wire n17551;
wire n17552;
wire n17553;
wire n17554;
wire n17555;
wire n17556;
wire n17557;
wire n17558;
wire n17559;
wire n17560;
wire n17561;
wire n17562;
wire n17563;
wire n17564;
wire n17565;
wire n17566;
wire n17567;
wire n17568;
wire n17569;
wire n17570;
wire n17571;
wire n17572;
wire n17573;
wire n17574;
wire n17575;
wire n17576;
wire n17577;
wire n17578;
wire n17579;
wire n17580;
wire n17581;
wire n17582;
wire n17583;
wire n17584;
wire n17585;
wire n17586;
wire n17587;
wire n17588;
wire n17589;
wire n17590;
wire n17591;
wire n17592;
wire n17593;
wire n17594;
wire n17595;
wire n17596;
wire n17597;
wire n17598;
wire n17599;
wire n17600;
wire n17601;
wire n17602;
wire n17603;
wire n17604;
wire n17605;
wire n17606;
wire n17607;
wire n17608;
wire n17609;
wire n17610;
wire n17611;
wire n17612;
wire n17613;
wire n17614;
wire n17615;
wire n17616;
wire n17617;
wire n17618;
wire n17619;
wire n17620;
wire n17621;
wire n17622;
wire n17623;
wire n17624;
wire n17625;
wire n17626;
wire n17627;
wire n17628;
wire n17629;
wire n17630;
wire n17631;
wire n17632;
wire n17633;
wire n17634;
wire n17635;
wire n17636;
wire n17637;
wire n17638;
wire n17639;
wire n17640;
wire n17641;
wire n17642;
wire n17643;
wire n17644;
wire n17645;
wire n17646;
wire n17647;
wire n17648;
wire n17649;
wire n17650;
wire n17651;
wire n17652;
wire n17653;
wire n17654;
wire n17655;
wire n17656;
wire n17657;
wire n17658;
wire n17659;
wire n17660;
wire n17661;
wire n17662;
wire n17663;
wire n17664;
wire n17665;
wire n17666;
wire n17667;
wire n17668;
wire n17669;
wire n17670;
wire n17671;
wire n17672;
wire n17673;
wire n17674;
wire n17675;
wire n17676;
wire n17677;
wire n17678;
wire n17679;
wire n17680;
wire n17681;
wire n17682;
wire n17683;
wire n17684;
wire n17685;
wire n17686;
wire n17687;
wire n17688;
wire n17689;
wire n17690;
wire n17691;
wire n17692;
wire n17693;
wire n17694;
wire n17695;
wire n17696;
wire n17697;
wire n17698;
wire n17699;
wire n17700;
wire n17701;
wire n17702;
wire n17703;
wire n17704;
wire n17705;
wire n17706;
wire n17707;
wire n17708;
wire n17709;
wire n17710;
wire n17711;
wire n17712;
wire n17713;
wire n17714;
wire n17715;
wire n17716;
wire n17717;
wire n17718;
wire n17719;
wire n17720;
wire n17721;
wire n17722;
wire n17723;
wire n17724;
wire n17725;
wire n17726;
wire n17727;
wire n17728;
wire n17729;
wire n17730;
wire n17731;
wire n17732;
wire n17733;
wire n17734;
wire n17735;
wire n17736;
wire n17737;
wire n17738;
wire n17739;
wire n17740;
wire n17741;
wire n17742;
wire n17743;
wire n17744;
wire n17745;
wire n17746;
wire n17747;
wire n17748;
wire n17749;
wire n17750;
wire n17751;
wire n17752;
wire n17753;
wire n17754;
wire n17755;
wire n17756;
wire n17757;
wire n17758;
wire n17759;
wire n17760;
wire n17761;
wire n17762;
wire n17763;
wire n17764;
wire n17765;
wire n17766;
wire n17767;
wire n17768;
wire n17769;
wire n17770;
wire n17771;
wire n17772;
wire n17773;
wire n17774;
wire n17775;
wire n17776;
wire n17777;
wire n17778;
wire n17779;
wire n17780;
wire n17781;
wire n17782;
wire n17783;
wire n17784;
wire n17785;
wire n17786;
wire n17787;
wire n17788;
wire n17789;
wire n17790;
wire n17791;
wire n17792;
wire n17793;
wire n17794;
wire n17795;
wire n17796;
wire n17797;
wire n17798;
wire n17799;
wire n17800;
wire n17801;
wire n17802;
wire n17803;
wire n17804;
wire n17805;
wire n17806;
wire n17807;
wire n17808;
wire n17809;
wire n17810;
wire n17811;
wire n17812;
wire n17813;
wire n17814;
wire n17815;
wire n17816;
wire n17817;
wire n17818;
wire n17819;
wire n17820;
wire n17821;
wire n17822;
wire n17823;
wire n17824;
wire n17825;
wire n17826;
wire n17827;
wire n17828;
wire n17829;
wire n17830;
wire n17831;
wire n17832;
wire n17833;
wire n17834;
wire n17835;
wire n17836;
wire n17837;
wire n17838;
wire n17839;
wire n17840;
wire n17841;
wire n17842;
wire n17843;
wire n17844;
wire n17845;
wire n17846;
wire n17847;
wire n17848;
wire n17849;
wire n17850;
wire n17851;
wire n17852;
wire n17853;
wire n17854;
wire n17855;
wire n17856;
wire n17857;
wire n17858;
wire n17859;
wire n17860;
wire n17861;
wire n17862;
wire n17863;
wire n17864;
wire n17865;
wire n17866;
wire n17867;
wire n17868;
wire n17869;
wire n17870;
wire n17871;
wire n17872;
wire n17873;
wire n17874;
wire n17875;
wire n17876;
wire n17877;
wire n17878;
wire n17879;
wire n17880;
wire n17881;
wire n17882;
wire n17883;
wire n17884;
wire n17885;
wire n17886;
wire n17887;
wire n17888;
wire n17889;
wire n17890;
wire n17891;
wire n17892;
wire n17893;
wire n17894;
wire n17895;
wire n17896;
wire n17897;
wire n17898;
wire n17899;
wire n17900;
wire n17901;
wire n17902;
wire n17903;
wire n17904;
wire n17905;
wire n17906;
wire n17907;
wire n17908;
wire n17909;
wire n17910;
wire n17911;
wire n17912;
wire n17913;
wire n17914;
wire n17915;
wire n17916;
wire n17917;
wire n17918;
wire n17919;
wire n17920;
wire n17921;
wire n17922;
wire n17923;
wire n17924;
wire n17925;
wire n17926;
wire n17927;
wire n17928;
wire n17929;
wire n17930;
wire n17931;
wire n17932;
wire n17933;
wire n17934;
wire n17935;
wire n17936;
wire n17937;
wire n17938;
wire n17939;
wire n17940;
wire n17941;
wire n17942;
wire n17943;
wire n17944;
wire n17945;
wire n17946;
wire n17947;
wire n17948;
wire n17949;
wire n17950;
wire n17951;
wire n17952;
wire n17953;
wire n17954;
wire n17955;
wire n17956;
wire n17957;
wire n17958;
wire n17959;
wire n17960;
wire n17961;
wire n17962;
wire n17963;
wire n17964;
wire n17965;
wire n17966;
wire n17967;
wire n17968;
wire n17969;
wire n17970;
wire n17971;
wire n17972;
wire n17973;
wire n17974;
wire n17975;
wire n17976;
wire n17977;
wire n17978;
wire n17979;
wire n17980;
wire n17981;
wire n17982;
wire n17983;
wire n17984;
wire n17985;
wire n17986;
wire n17987;
wire n17988;
wire n17989;
wire n17990;
wire n17991;
wire n17992;
wire n17993;
wire n17994;
wire n17995;
wire n17996;
wire n17997;
wire n17998;
wire n17999;
wire n18000;
wire n18001;
wire n18002;
wire n18003;
wire n18004;
wire n18005;
wire n18006;
wire n18007;
wire n18008;
wire n18009;
wire n18010;
wire n18011;
wire n18012;
wire n18013;
wire n18014;
wire n18015;
wire n18016;
wire n18017;
wire n18018;
wire n18019;
wire n18020;
wire n18021;
wire n18022;
wire n18023;
wire n18024;
wire n18025;
wire n18026;
wire n18027;
wire n18028;
wire n18029;
wire n18030;
wire n18031;
wire n18032;
wire n18033;
wire n18034;
wire n18035;
wire n18036;
wire n18037;
wire n18038;
wire n18039;
wire n18040;
wire n18041;
wire n18042;
wire n18043;
wire n18044;
wire n18045;
wire n18046;
wire n18047;
wire n18048;
wire n18049;
wire n18050;
wire n18051;
wire n18052;
wire n18053;
wire n18054;
wire n18055;
wire n18056;
wire n18057;
wire n18058;
wire n18059;
wire n18060;
wire n18061;
wire n18062;
wire n18063;
wire n18064;
wire n18065;
wire n18066;
wire n18067;
wire n18068;
wire n18069;
wire n18070;
wire n18071;
wire n18072;
wire n18073;
wire n18074;
wire n18075;
wire n18076;
wire n18077;
wire n18078;
wire n18079;
wire n18080;
wire n18081;
wire n18082;
wire n18083;
wire n18084;
wire n18085;
wire n18086;
wire n18087;
wire n18088;
wire n18089;
wire n18090;
wire n18091;
wire n18092;
wire n18093;
wire n18094;
wire n18095;
wire n18096;
wire n18097;
wire n18098;
wire n18099;
wire n18100;
wire n18101;
wire n18102;
wire n18103;
wire n18104;
wire n18105;
wire n18106;
wire n18107;
wire n18108;
wire n18109;
wire n18110;
wire n18111;
wire n18112;
wire n18113;
wire n18114;
wire n18115;
wire n18116;
wire n18117;
wire n18118;
wire n18119;
wire n18120;
wire n18121;
wire n18122;
wire n18123;
wire n18124;
wire n18125;
wire n18126;
wire n18127;
wire n18128;
wire n18129;
wire n18130;
wire n18131;
wire n18132;
wire n18133;
wire n18134;
wire n18135;
wire n18136;
wire n18137;
wire n18138;
wire n18139;
wire n18140;
wire n18141;
wire n18142;
wire n18143;
wire n18144;
wire n18145;
wire n18146;
wire n18147;
wire n18148;
wire n18149;
wire n18150;
wire n18151;
wire n18152;
wire n18153;
wire n18154;
wire n18155;
wire n18156;
wire n18157;
wire n18158;
wire n18159;
wire n18160;
wire n18161;
wire n18162;
wire n18163;
wire n18164;
wire n18165;
wire n18166;
wire n18167;
wire n18168;
wire n18169;
wire n18170;
wire n18171;
wire n18172;
wire n18173;
wire n18174;
wire n18175;
wire n18176;
wire n18177;
wire n18178;
wire n18179;
wire n18180;
wire n18181;
wire n18182;
wire n18183;
wire n18184;
wire n18185;
wire n18186;
wire n18187;
wire n18188;
wire n18189;
wire n18190;
wire n18191;
wire n18192;
wire n18193;
wire n18194;
wire n18195;
wire n18196;
wire n18197;
wire n18198;
wire n18199;
wire n18200;
wire n18201;
wire n18202;
wire n18203;
wire n18204;
wire n18205;
wire n18206;
wire n18207;
wire n18208;
wire n18209;
wire n18210;
wire n18211;
wire n18212;
wire n18213;
wire n18214;
wire n18215;
wire n18216;
wire n18217;
wire n18218;
wire n18219;
wire n18220;
wire n18221;
wire n18222;
wire n18223;
wire n18224;
wire n18225;
wire n18226;
wire n18227;
wire n18228;
wire n18229;
wire n18230;
wire n18231;
wire n18232;
wire n18233;
wire n18234;
wire n18235;
wire n18236;
wire n18237;
wire n18238;
wire n18239;
wire n18240;
wire n18241;
wire n18242;
wire n18243;
wire n18244;
wire n18245;
wire n18246;
wire n18247;
wire n18248;
wire n18249;
wire n18250;
wire n18251;
wire n18252;
wire n18253;
wire n18254;
wire n18255;
wire n18256;
wire n18257;
wire n18258;
wire n18259;
wire n18260;
wire n18261;
wire n18262;
wire n18263;
wire n18264;
wire n18265;
wire n18266;
wire n18267;
wire n18268;
wire n18269;
wire n18270;
wire n18271;
wire n18272;
wire n18273;
wire n18274;
wire n18275;
wire n18276;
wire n18277;
wire n18278;
wire n18279;
wire n18280;
wire n18281;
wire n18282;
wire n18283;
wire n18284;
wire n18285;
wire n18286;
wire n18287;
wire n18288;
wire n18289;
wire n18290;
wire n18291;
wire n18292;
wire n18293;
wire n18294;
wire n18295;
wire n18296;
wire n18297;
wire n18298;
wire n18299;
wire n18300;
wire n18301;
wire n18302;
wire n18303;
wire n18304;
wire n18305;
wire n18306;
wire n18307;
wire n18308;
wire n18309;
wire n18310;
wire n18311;
wire n18312;
wire n18313;
wire n18314;
wire n18315;
wire n18316;
wire n18317;
wire n18318;
wire n18319;
wire n18320;
wire n18321;
wire n18322;
wire n18323;
wire n18324;
wire n18325;
wire n18326;
wire n18327;
wire n18328;
wire n18329;
wire n18330;
wire n18331;
wire n18332;
wire n18333;
wire n18334;
wire n18335;
wire n18336;
wire n18337;
wire n18338;
wire n18339;
wire n18340;
wire n18341;
wire n18342;
wire n18343;
wire n18344;
wire n18345;
wire n18346;
wire n18347;
wire n18348;
wire n18349;
wire n18350;
wire n18351;
wire n18352;
wire n18353;
wire n18354;
wire n18355;
wire n18356;
wire n18357;
wire n18358;
wire n18359;
wire n18360;
wire n18361;
wire n18362;
wire n18363;
wire n18364;
wire n18365;
wire n18366;
wire n18367;
wire n18368;
wire n18369;
wire n18370;
wire n18371;
wire n18372;
wire n18373;
wire n18374;
wire n18375;
wire n18376;
wire n18377;
wire n18378;
wire n18379;
wire n18380;
wire n18381;
wire n18382;
wire n18383;
wire n18384;
wire n18385;
wire n18386;
wire n18387;
wire n18388;
wire n18389;
wire n18390;
wire n18391;
wire n18392;
wire n18393;
wire n18394;
wire n18395;
wire n18396;
wire n18397;
wire n18398;
wire n18399;
wire n18400;
wire n18401;
wire n18402;
wire n18403;
wire n18404;
wire n18405;
wire n18406;
wire n18407;
wire n18408;
wire n18409;
wire n18410;
wire n18411;
wire n18412;
wire n18413;
wire n18414;
wire n18415;
wire n18416;
wire n18417;
wire n18418;
wire n18419;
wire n18420;
wire n18421;
wire n18422;
wire n18423;
wire n18424;
wire n18425;
wire n18426;
wire n18427;
wire n18428;
wire n18429;
wire n18430;
wire n18431;
wire n18432;
wire n18433;
wire n18434;
wire n18435;
wire n18436;
wire n18437;
wire n18438;
wire n18439;
wire n18440;
wire n18441;
wire n18442;
wire n18443;
wire n18444;
wire n18445;
wire n18446;
wire n18447;
wire n18448;
wire n18449;
wire n18450;
wire n18451;
wire n18452;
wire n18453;
wire n18454;
wire n18455;
wire n18456;
wire n18457;
wire n18458;
wire n18459;
wire n18460;
wire n18461;
wire n18462;
wire n18463;
wire n18464;
wire n18465;
wire n18466;
wire n18467;
wire n18468;
wire n18469;
wire n18470;
wire n18471;
wire n18472;
wire n18473;
wire n18474;
wire n18475;
wire n18476;
wire n18477;
wire n18478;
wire n18479;
wire n18480;
wire n18481;
wire n18482;
wire n18483;
wire n18484;
wire n18485;
wire n18486;
wire n18487;
wire n18488;
wire n18489;
wire n18490;
wire n18491;
wire n18492;
wire n18493;
wire n18494;
wire n18495;
wire n18496;
wire n18497;
wire n18498;
wire n18499;
wire n18500;
wire n18501;
wire n18502;
wire n18503;
wire n18504;
wire n18505;
wire n18506;
wire n18507;
wire n18508;
wire n18509;
wire n18510;
wire n18511;
wire n18512;
wire n18513;
wire n18514;
wire n18515;
wire n18516;
wire n18517;
wire n18518;
wire n18519;
wire n18520;
wire n18521;
wire n18522;
wire n18523;
wire n18524;
wire n18525;
wire n18526;
wire n18527;
wire n18528;
wire n18529;
wire n18530;
wire n18531;
wire n18532;
wire n18533;
wire n18534;
wire n18535;
wire n18536;
wire n18537;
wire n18538;
wire n18539;
wire n18540;
wire n18541;
wire n18542;
wire n18543;
wire n18544;
wire n18545;
wire n18546;
wire n18547;
wire n18548;
wire n18549;
wire n18550;
wire n18551;
wire n18552;
wire n18553;
wire n18554;
wire n18555;
wire n18556;
wire n18557;
wire n18558;
wire n18559;
wire n18560;
wire n18561;
wire n18562;
wire n18563;
wire n18564;
wire n18565;
wire n18566;
wire n18567;
wire n18568;
wire n18569;
wire n18570;
wire n18571;
wire n18572;
wire n18573;
wire n18574;
wire n18575;
wire n18576;
wire n18577;
wire n18578;
wire n18579;
wire n18580;
wire n18581;
wire n18582;
wire n18583;
wire n18584;
wire n18585;
wire n18586;
wire n18587;
wire n18588;
wire n18589;
wire n18590;
wire n18591;
wire n18592;
wire n18593;
wire n18594;
wire n18595;
wire n18596;
wire n18597;
wire n18598;
wire n18599;
wire n18600;
wire n18601;
wire n18602;
wire n18603;
wire n18604;
wire n18605;
wire n18606;
wire n18607;
wire n18608;
wire n18609;
wire n18610;
wire n18611;
wire n18612;
wire n18613;
wire n18614;
wire n18615;
wire n18616;
wire n18617;
wire n18618;
wire n18619;
wire n18620;
wire n18621;
wire n18622;
wire n18623;
wire n18624;
wire n18625;
wire n18626;
wire n18627;
wire n18628;
wire n18629;
wire n18630;
wire n18631;
wire n18632;
wire n18633;
wire n18634;
wire n18635;
wire n18636;
wire n18637;
wire n18638;
wire n18639;
wire n18640;
wire n18641;
wire n18642;
wire n18643;
wire n18644;
wire n18645;
wire n18646;
wire n18647;
wire n18648;
wire n18649;
wire n18650;
wire n18651;
wire n18652;
wire n18653;
wire n18654;
wire n18655;
wire n18656;
wire n18657;
wire n18658;
wire n18659;
wire n18660;
wire n18661;
wire n18662;
wire n18663;
wire n18664;
wire n18665;
wire n18666;
wire n18667;
wire n18668;
wire n18669;
wire n18670;
wire n18671;
wire n18672;
wire n18673;
wire n18674;
wire n18675;
wire n18676;
wire n18677;
wire n18678;
wire n18679;
wire n18680;
wire n18681;
wire n18682;
wire n18683;
wire n18684;
wire n18685;
wire n18686;
wire n18687;
wire n18688;
wire n18689;
wire n18690;
wire n18691;
wire n18692;
wire n18693;
wire n18694;
wire n18695;
wire n18696;
wire n18697;
wire n18698;
wire n18699;
wire n18700;
wire n18701;
wire n18702;
wire n18703;
wire n18704;
wire n18705;
wire n18706;
wire n18707;
wire n18708;
wire n18709;
wire n18710;
wire n18711;
wire n18712;
wire n18713;
wire n18714;
wire n18715;
wire n18716;
wire n18717;
wire n18718;
wire n18719;
wire n18720;
wire n18721;
wire n18722;
wire n18723;
wire n18724;
wire n18725;
wire n18726;
wire n18727;
wire n18728;
wire n18729;
wire n18730;
wire n18731;
wire n18732;
wire n18733;
wire n18734;
wire n18735;
wire n18736;
wire n18737;
wire n18738;
wire n18739;
wire n18740;
wire n18741;
wire n18742;
wire n18743;
wire n18744;
wire n18745;
wire n18746;
wire n18747;
wire n18748;
wire n18749;
wire n18750;
wire n18751;
wire n18752;
wire n18753;
wire n18754;
wire n18755;
wire n18756;
wire n18757;
wire n18758;
wire n18759;
wire n18760;
wire n18761;
wire n18762;
wire n18763;
wire n18764;
wire n18765;
wire n18766;
wire n18767;
wire n18768;
wire n18769;
wire n18770;
wire n18771;
wire n18772;
wire n18773;
wire n18774;
wire n18775;
wire n18776;
wire n18777;
wire n18778;
wire n18779;
wire n18780;
wire n18781;
wire n18782;
wire n18783;
wire n18784;
wire n18785;
wire n18786;
wire n18787;
wire n18788;
wire n18789;
wire n18790;
wire n18791;
wire n18792;
wire n18793;
wire n18794;
wire n18795;
wire n18796;
wire n18797;
wire n18798;
wire n18799;
wire n18800;
wire n18801;
wire n18802;
wire n18803;
wire n18804;
wire n18805;
wire n18806;
wire n18807;
wire n18808;
wire n18809;
wire n18810;
wire n18811;
wire n18812;
wire n18813;
wire n18814;
wire n18815;
wire n18816;
wire n18817;
wire n18818;
wire n18819;
wire n18820;
wire n18821;
wire n18822;
wire n18823;
wire n18824;
wire n18825;
wire n18826;
wire n18827;
wire n18828;
wire n18829;
wire n18830;
wire n18831;
wire n18832;
wire n18833;
wire n18834;
wire n18835;
wire n18836;
wire n18837;
wire n18838;
wire n18839;
wire n18840;
wire n18841;
wire n18842;
wire n18843;
wire n18844;
wire n18845;
wire n18846;
wire n18847;
wire n18848;
wire n18849;
wire n18850;
wire n18851;
wire n18852;
wire n18853;
wire n18854;
wire n18855;
wire n18856;
wire n18857;
wire n18858;
wire n18859;
wire n18860;
wire n18861;
wire n18862;
wire n18863;
wire n18864;
wire n18865;
wire n18866;
wire n18867;
wire n18868;
wire n18869;
wire n18870;
wire n18871;
wire n18872;
wire n18873;
wire n18874;
wire n18875;
wire n18876;
wire n18877;
wire n18878;
wire n18879;
wire n18880;
wire n18881;
wire n18882;
wire n18883;
wire n18884;
wire n18885;
wire n18886;
wire n18887;
wire n18888;
wire n18889;
wire n18890;
wire n18891;
wire n18892;
wire n18893;
wire n18894;
wire n18895;
wire n18896;
wire n18897;
wire n18898;
wire n18899;
wire n18900;
wire n18901;
wire n18902;
wire n18903;
wire n18904;
wire n18905;
wire n18906;
wire n18907;
wire n18908;
wire n18909;
wire n18910;
wire n18911;
wire n18912;
wire n18913;
wire n18914;
wire n18915;
wire n18916;
wire n18917;
wire n18918;
wire n18919;
wire n18920;
wire n18921;
wire n18922;
wire n18923;
wire n18924;
wire n18925;
wire n18926;
wire n18927;
wire n18928;
wire n18929;
wire n18930;
wire n18931;
wire n18932;
wire n18933;
wire n18934;
wire n18935;
wire n18936;
wire n18937;
wire n18938;
wire n18939;
wire n18940;
wire n18941;
wire n18942;
wire n18943;
wire n18944;
wire n18945;
wire n18946;
wire n18947;
wire n18948;
wire n18949;
wire n18950;
wire n18951;
wire n18952;
wire n18953;
wire n18954;
wire n18955;
wire n18956;
wire n18957;
wire n18958;
wire n18959;
wire n18960;
wire n18961;
wire n18962;
wire n18963;
wire n18964;
wire n18965;
wire n18966;
wire n18967;
wire n18968;
wire n18969;
wire n18970;
wire n18971;
wire n18972;
wire n18973;
wire n18974;
wire n18975;
wire n18976;
wire n18977;
wire n18978;
wire n18979;
wire n18980;
wire n18981;
wire n18982;
wire n18983;
wire n18984;
wire n18985;
wire n18986;
wire n18987;
wire n18988;
wire n18989;
wire n18990;
wire n18991;
wire n18992;
wire n18993;
wire n18994;
wire n18995;
wire n18996;
wire n18997;
wire n18998;
wire n18999;
wire n19000;
wire n19001;
wire n19002;
wire n19003;
wire n19004;
wire n19005;
wire n19006;
wire n19007;
wire n19008;
wire n19009;
wire n19010;
wire n19011;
wire n19012;
wire n19013;
wire n19014;
wire n19015;
wire n19016;
wire n19017;
wire n19018;
wire n19019;
wire n19020;
wire n19021;
wire n19022;
wire n19023;
wire n19024;
wire n19025;
wire n19026;
wire n19027;
wire n19028;
wire n19029;
wire n19030;
wire n19031;
wire n19032;
wire n19033;
wire n19034;
wire n19035;
wire n19036;
wire n19037;
wire n19038;
wire n19039;
wire n19040;
wire n19041;
wire n19042;
wire n19043;
wire n19044;
wire n19045;
wire n19046;
wire n19047;
wire n19048;
wire n19049;
wire n19050;
wire n19051;
wire n19052;
wire n19053;
wire n19054;
wire n19055;
wire n19056;
wire n19057;
wire n19058;
wire n19059;
wire n19060;
wire n19061;
wire n19062;
wire n19063;
wire n19064;
wire n19065;
wire n19066;
wire n19067;
wire n19068;
wire n19069;
wire n19070;
wire n19071;
wire n19072;
wire n19073;
wire n19074;
wire n19075;
wire n19076;
wire n19077;
wire n19078;
wire n19079;
wire n19080;
wire n19081;
wire n19082;
wire n19083;
wire n19084;
wire n19085;
wire n19086;
wire n19087;
wire n19088;
wire n19089;
wire n19090;
wire n19091;
wire n19092;
wire n19093;
wire n19094;
wire n19095;
wire n19096;
wire n19097;
wire n19098;
wire n19099;
wire n19100;
wire n19101;
wire n19102;
wire n19103;
wire n19104;
wire n19105;
wire n19106;
wire n19107;
wire n19108;
wire n19109;
wire n19110;
wire n19111;
wire n19112;
wire n19113;
wire n19114;
wire n19115;
wire n19116;
wire n19117;
wire n19118;
wire n19119;
wire n19120;
wire n19121;
wire n19122;
wire n19123;
wire n19124;
wire n19125;
wire n19126;
wire n19127;
wire n19128;
wire n19129;
wire n19130;
wire n19131;
wire n19132;
wire n19133;
wire n19134;
wire n19135;
wire n19136;
wire n19137;
wire n19138;
wire n19139;
wire n19140;
wire n19141;
wire n19142;
wire n19143;
wire n19144;
wire n19145;
wire n19146;
wire n19147;
wire n19148;
wire n19149;
wire n19150;
wire n19151;
wire n19152;
wire n19153;
wire n19154;
wire n19155;
wire n19156;
wire n19157;
wire n19158;
wire n19159;
wire n19160;
wire n19161;
wire n19162;
wire n19163;
wire n19164;
wire n19165;
wire n19166;
wire n19167;
wire n19168;
wire n19169;
wire n19170;
wire n19171;
wire n19172;
wire n19173;
wire n19174;
wire n19175;
wire n19176;
wire n19177;
wire n19178;
wire n19179;
wire n19180;
wire n19181;
wire n19182;
wire n19183;
wire n19184;
wire n19185;
wire n19186;
wire n19187;
wire n19188;
wire n19189;
wire n19190;
wire n19191;
wire n19192;
wire n19193;
wire n19194;
wire n19195;
wire n19196;
wire n19197;
wire n19198;
wire n19199;
wire n19200;
wire n19201;
wire n19202;
wire n19203;
wire n19204;
wire n19205;
wire n19206;
wire n19207;
wire n19208;
wire n19209;
wire n19210;
wire n19211;
wire n19212;
wire n19213;
wire n19214;
wire n19215;
wire n19216;
wire n19217;
wire n19218;
wire n19219;
wire n19220;
wire n19221;
wire n19222;
wire n19223;
wire n19224;
wire n19225;
wire n19226;
wire n19227;
wire n19228;
wire n19229;
wire n19230;
wire n19231;
wire n19232;
wire n19233;
wire n19234;
wire n19235;
wire n19236;
wire n19237;
wire n19238;
wire n19239;
wire n19240;
wire n19241;
wire n19242;
wire n19243;
wire n19244;
wire n19245;
wire n19246;
wire n19247;
wire n19248;
wire n19249;
wire n19250;
wire n19251;
wire n19252;
wire n19253;
wire n19254;
wire n19255;
wire n19256;
wire n19257;
wire n19258;
wire n19259;
wire n19260;
wire n19261;
wire n19262;
wire n19263;
wire n19264;
wire n19265;
wire n19266;
wire n19267;
wire n19268;
wire n19269;
wire n19270;
wire n19271;
wire n19272;
wire n19273;
wire n19274;
wire n19275;
wire n19276;
wire n19277;
wire n19278;
wire n19279;
wire n19280;
wire n19281;
wire n19282;
wire n19283;
wire n19284;
wire n19285;
wire n19286;
wire n19287;
wire n19288;
wire n19289;
wire n19290;
wire n19291;
wire n19292;
wire n19293;
wire n19294;
wire n19295;
wire n19296;
wire n19297;
wire n19298;
wire n19299;
wire n19300;
wire n19301;
wire n19302;
wire n19303;
wire n19304;
wire n19305;
wire n19306;
wire n19307;
wire n19308;
wire n19309;
wire n19310;
wire n19311;
wire n19312;
wire n19313;
wire n19314;
wire n19315;
wire n19316;
wire n19317;
wire n19318;
wire n19319;
wire n19320;
wire n19321;
wire n19322;
wire n19323;
wire n19324;
wire n19325;
wire n19326;
wire n19327;
wire n19328;
wire n19329;
wire n19330;
wire n19331;
wire n19332;
wire n19333;
wire n19334;
wire n19335;
wire n19336;
wire n19337;
wire n19338;
wire n19339;
wire n19340;
wire n19341;
wire n19342;
wire n19343;
wire n19344;
wire n19345;
wire n19346;
wire n19347;
wire n19348;
wire n19349;
wire n19350;
wire n19351;
wire n19352;
wire n19353;
wire n19354;
wire n19355;
wire n19356;
wire n19357;
wire n19358;
wire n19359;
wire n19360;
wire n19361;
wire n19362;
wire n19363;
wire n19364;
wire n19365;
wire n19366;
wire n19367;
wire n19368;
wire n19369;
wire n19370;
wire n19371;
wire n19372;
wire n19373;
wire n19374;
wire n19375;
wire n19376;
wire n19377;
wire n19378;
wire n19379;
wire n19380;
wire n19381;
wire n19382;
wire n19383;
wire n19384;
wire n19385;
wire n19386;
wire n19387;
wire n19388;
wire n19389;
wire n19390;
wire n19391;
wire n19392;
wire n19393;
wire n19394;
wire n19395;
wire n19396;
wire n19397;
wire n19398;
wire n19399;
wire n19400;
wire n19401;
wire n19402;
wire n19403;
wire n19404;
wire n19405;
wire n19406;
wire n19407;
wire n19408;
wire n19409;
wire n19410;
wire n19411;
wire n19412;
wire n19413;
wire n19414;
wire n19415;
wire n19416;
wire n19417;
wire n19418;
wire n19419;
wire n19420;
wire n19421;
wire n19422;
wire n19423;
wire n19424;
wire n19425;
wire n19426;
wire n19427;
wire n19428;
wire n19429;
wire n19430;
wire n19431;
wire n19432;
wire n19433;
wire n19434;
wire n19435;
wire n19436;
wire n19437;
wire n19438;
wire n19439;
wire n19440;
wire n19441;
wire n19442;
wire n19443;
wire n19444;
wire n19445;
wire n19446;
wire n19447;
wire n19448;
wire n19449;
wire n19450;
wire n19451;
wire n19452;
wire n19453;
wire n19454;
wire n19455;
wire n19456;
wire n19457;
wire n19458;
wire n19459;
wire n19460;
wire n19461;
wire n19462;
wire n19463;
wire n19464;
wire n19465;
wire n19466;
wire n19467;
wire n19468;
wire n19469;
wire n19470;
wire n19471;
wire n19472;
wire n19473;
wire n19474;
wire n19475;
wire n19476;
wire n19477;
wire n19478;
wire n19479;
wire n19480;
wire n19481;
wire n19482;
wire n19483;
wire n19484;
wire n19485;
wire n19486;
wire n19487;
wire n19488;
wire n19489;
wire n19490;
wire n19491;
wire n19492;
wire n19493;
wire n19494;
wire n19495;
wire n19496;
wire n19497;
wire n19498;
wire n19499;
wire n19500;
wire n19501;
wire n19502;
wire n19503;
wire n19504;
wire n19505;
wire n19506;
wire n19507;
wire n19508;
wire n19509;
wire n19510;
wire n19511;
wire n19512;
wire n19513;
wire n19514;
wire n19515;
wire n19516;
wire n19517;
wire n19518;
wire n19519;
wire n19520;
wire n19521;
wire n19522;
wire n19523;
wire n19524;
wire n19525;
wire n19526;
wire n19527;
wire n19528;
wire n19529;
wire n19530;
wire n19531;
wire n19532;
wire n19533;
wire n19534;
wire n19535;
wire n19536;
wire n19537;
wire n19538;
wire n19539;
wire n19540;
wire n19541;
wire n19542;
wire n19543;
wire n19544;
wire n19545;
wire n19546;
wire n19547;
wire n19548;
wire n19549;
wire n19550;
wire n19551;
wire n19552;
wire n19553;
wire n19554;
wire n19555;
wire n19556;
wire n19557;
wire n19558;
wire n19559;
wire n19560;
wire n19561;
wire n19562;
wire n19563;
wire n19564;
wire n19565;
wire n19566;
wire n19567;
wire n19568;
wire n19569;
wire n19570;
wire n19571;
wire n19572;
wire n19573;
wire n19574;
wire n19575;
wire n19576;
wire n19577;
wire n19578;
wire n19579;
wire n19580;
wire n19581;
wire n19582;
wire n19583;
wire n19584;
wire n19585;
wire n19586;
wire n19587;
wire n19588;
wire n19589;
wire n19590;
wire n19591;
wire n19592;
wire n19593;
wire n19594;
wire n19595;
wire n19596;
wire n19597;
wire n19598;
wire n19599;
wire n19600;
wire n19601;
wire n19602;
wire n19603;
wire n19604;
wire n19605;
wire n19606;
wire n19607;
wire n19608;
wire n19609;
wire n19610;
wire n19611;
wire n19612;
wire n19613;
wire n19614;
wire n19615;
wire n19616;
wire n19617;
wire n19618;
wire n19619;
wire n19620;
wire n19621;
wire n19622;
wire n19623;
wire n19624;
wire n19625;
wire n19626;
wire n19627;
wire n19628;
wire n19629;
wire n19630;
wire n19631;
wire n19632;
wire n19633;
wire n19634;
wire n19635;
wire n19636;
wire n19637;
wire n19638;
wire n19639;
wire n19640;
wire n19641;
wire n19642;
wire n19643;
wire n19644;
wire n19645;
wire n19646;
wire n19647;
wire n19648;
wire n19649;
wire n19650;
wire n19651;
wire n19652;
wire n19653;
wire n19654;
wire n19655;
wire n19656;
wire n19657;
wire n19658;
wire n19659;
wire n19660;
wire n19661;
wire n19662;
wire n19663;
wire n19664;
wire n19665;
wire n19666;
wire n19667;
wire n19668;
wire n19669;
wire n19670;
wire n19671;
wire n19672;
wire n19673;
wire n19674;
wire n19675;
wire n19676;
wire n19677;
wire n19678;
wire n19679;
wire n19680;
wire n19681;
wire n19682;
wire n19683;
wire n19684;
wire n19685;
wire n19686;
wire n19687;
wire n19688;
wire n19689;
wire n19690;
wire n19691;
wire n19692;
wire n19693;
wire n19694;
wire n19695;
wire n19696;
wire n19697;
wire n19698;
wire n19699;
wire n19700;
wire n19701;
wire n19702;
wire n19703;
wire n19704;
wire n19705;
wire n19706;
wire n19707;
wire n19708;
wire n19709;
wire n19710;
wire n19711;
wire n19712;
wire n19713;
wire n19714;
wire n19715;
wire n19716;
wire n19717;
wire n19718;
wire n19719;
wire n19720;
wire n19721;
wire n19722;
wire n19723;
wire n19724;
wire n19725;
wire n19726;
wire n19727;
wire n19728;
wire n19729;
wire n19730;
wire n19731;
wire n19732;
wire n19733;
wire n19734;
wire n19735;
wire n19736;
wire n19737;
wire n19738;
wire n19739;
wire n19740;
wire n19741;
wire n19742;
wire n19743;
wire n19744;
wire n19745;
wire n19746;
wire n19747;
wire n19748;
wire n19749;
wire n19750;
wire n19751;
wire n19752;
wire n19753;
wire n19754;
wire n19755;
wire n19756;
wire n19757;
wire n19758;
wire n19759;
wire n19760;
wire n19761;
wire n19762;
wire n19763;
wire n19764;
wire n19765;
wire n19766;
wire n19767;
wire n19768;
wire n19769;
wire n19770;
wire n19771;
wire n19772;
wire n19773;
wire n19774;
wire n19775;
wire n19776;
wire n19777;
wire n19778;
wire n19779;
wire n19780;
wire n19781;
wire n19782;
wire n19783;
wire n19784;
wire n19785;
wire n19786;
wire n19787;
wire n19788;
wire n19789;
wire n19790;
wire n19791;
wire n19792;
wire n19793;
wire n19794;
wire n19795;
wire n19796;
wire n19797;
wire n19798;
wire n19799;
wire n19800;
wire n19801;
wire n19802;
wire n19803;
wire n19804;
wire n19805;
wire n19806;
wire n19807;
wire n19808;
wire n19809;
wire n19810;
wire n19811;
wire n19812;
wire n19813;
wire n19814;
wire n19815;
wire n19816;
wire n19817;
wire n19818;
wire n19819;
wire n19820;
wire n19821;
wire n19822;
wire n19823;
wire n19824;
wire n19825;
wire n19826;
wire n19827;
wire n19828;
wire n19829;
wire n19830;
wire n19831;
wire n19832;
wire n19833;
wire n19834;
wire n19835;
wire n19836;
wire n19837;
wire n19838;
wire n19839;
wire n19840;
wire n19841;
wire n19842;
wire n19843;
wire n19844;
wire n19845;
wire n19846;
wire n19847;
wire n19848;
wire n19849;
wire n19850;
wire n19851;
wire n19852;
wire n19853;
wire n19854;
wire n19855;
wire n19856;
wire n19857;
wire n19858;
wire n19859;
wire n19860;
wire n19861;
wire n19862;
wire n19863;
wire n19864;
wire n19865;
wire n19866;
wire n19867;
wire n19868;
wire n19869;
wire n19870;
wire n19871;
wire n19872;
wire n19873;
wire n19874;
wire n19875;
wire n19876;
wire n19877;
wire n19878;
wire n19879;
wire n19880;
wire n19881;
wire n19882;
wire n19883;
wire n19884;
wire n19885;
wire n19886;
wire n19887;
wire n19888;
wire n19889;
wire n19890;
wire n19891;
wire n19892;
wire n19893;
wire n19894;
wire n19895;
wire n19896;
wire n19897;
wire n19898;
wire n19899;
wire n19900;
wire n19901;
wire n19902;
wire n19903;
wire n19904;
wire n19905;
wire n19906;
wire n19907;
wire n19908;
wire n19909;
wire n19910;
wire n19911;
wire n19912;
wire n19913;
wire n19914;
wire n19915;
wire n19916;
wire n19917;
wire n19918;
wire n19919;
wire n19920;
wire n19921;
wire n19922;
wire n19923;
wire n19924;
wire n19925;
wire n19926;
wire n19927;
wire n19928;
wire n19929;
wire n19930;
wire n19931;
wire n19932;
wire n19933;
wire n19934;
wire n19935;
wire n19936;
wire n19937;
wire n19938;
wire n19939;
wire n19940;
wire n19941;
wire n19942;
wire n19943;
wire n19944;
wire n19945;
wire n19946;
wire n19947;
wire n19948;
wire n19949;
wire n19950;
wire n19951;
wire n19952;
wire n19953;
wire n19954;
wire n19955;
wire n19956;
wire n19957;
wire n19958;
wire n19959;
wire n19960;
wire n19961;
wire n19962;
wire n19963;
wire n19964;
wire n19965;
wire n19966;
wire n19967;
wire n19968;
wire n19969;
wire n19970;
wire n19971;
wire n19972;
wire n19973;
wire n19974;
wire n19975;
wire n19976;
wire n19977;
wire n19978;
wire n19979;
wire n19980;
wire n19981;
wire n19982;
wire n19983;
wire n19984;
wire n19985;
wire n19986;
wire n19987;
wire n19988;
wire n19989;
wire n19990;
wire n19991;
wire n19992;
wire n19993;
wire n19994;
wire n19995;
wire n19996;
wire n19997;
wire n19998;
wire n19999;
wire n20000;
wire n20001;
wire n20002;
wire n20003;
wire n20004;
wire n20005;
wire n20006;
wire n20007;
wire n20008;
wire n20009;
wire n20010;
wire n20011;
wire n20012;
wire n20013;
wire n20014;
wire n20015;
wire n20016;
wire n20017;
wire n20018;
wire n20019;
wire n20020;
wire n20021;
wire n20022;
wire n20023;
wire n20024;
wire n20025;
wire n20026;
wire n20027;
wire n20028;
wire n20029;
wire n20030;
wire n20031;
wire n20032;
wire n20033;
wire n20034;
wire n20035;
wire n20036;
wire n20037;
wire n20038;
wire n20039;
wire n20040;
wire n20041;
wire n20042;
wire n20043;
wire n20044;
wire n20045;
wire n20046;
wire n20047;
wire n20048;
wire n20049;
wire n20050;
wire n20051;
wire n20052;
wire n20053;
wire n20054;
wire n20055;
wire n20056;
wire n20057;
wire n20058;
wire n20059;
wire n20060;
wire n20061;
wire n20062;
wire n20063;
wire n20064;
wire n20065;
wire n20066;
wire n20067;
wire n20068;
wire n20069;
wire n20070;
wire n20071;
wire n20072;
wire n20073;
wire n20074;
wire n20075;
wire n20076;
wire n20077;
wire n20078;
wire n20079;
wire n20080;
wire n20081;
wire n20082;
wire n20083;
wire n20084;
wire n20085;
wire n20086;
wire n20087;
wire n20088;
wire n20089;
wire n20090;
wire n20091;
wire n20092;
wire n20093;
wire n20094;
wire n20095;
wire n20096;
wire n20097;
wire n20098;
wire n20099;
wire n20100;
wire n20101;
wire n20102;
wire n20103;
wire n20104;
wire n20105;
wire n20106;
wire n20107;
wire n20108;
wire n20109;
wire n20110;
wire n20111;
wire n20112;
wire n20113;
wire n20114;
wire n20115;
wire n20116;
wire n20117;
wire n20118;
wire n20119;
wire n20120;
wire n20121;
wire n20122;
wire n20123;
wire n20124;
wire n20125;
wire n20126;
wire n20127;
wire n20128;
wire n20129;
wire n20130;
wire n20131;
wire n20132;
wire n20133;
wire n20134;
wire n20135;
wire n20136;
wire n20137;
wire n20138;
wire n20139;
wire n20140;
wire n20141;
wire n20142;
wire n20143;
wire n20144;
wire n20145;
wire n20146;
wire n20147;
wire n20148;
wire n20149;
wire n20150;
wire n20151;
wire n20152;
wire n20153;
wire n20154;
wire n20155;
wire n20156;
wire n20157;
wire n20158;
wire n20159;
wire n20160;
wire n20161;
wire n20162;
wire n20163;
wire n20164;
wire n20165;
wire n20166;
wire n20167;
wire n20168;
wire n20169;
wire n20170;
wire n20171;
wire n20172;
wire n20173;
wire n20174;
wire n20175;
wire n20176;
wire n20177;
wire n20178;
wire n20179;
wire n20180;
wire n20181;
wire n20182;
wire n20183;
wire n20184;
wire n20185;
wire n20186;
wire n20187;
wire n20188;
wire n20189;
wire n20190;
wire n20191;
wire n20192;
wire n20193;
wire n20194;
wire n20195;
wire n20196;
wire n20197;
wire n20198;
wire n20199;
wire n20200;
wire n20201;
wire n20202;
wire n20203;
wire n20204;
wire n20205;
wire n20206;
wire n20207;
wire n20208;
wire n20209;
wire n20210;
wire n20211;
wire n20212;
wire n20213;
wire n20214;
wire n20215;
wire n20216;
wire n20217;
wire n20218;
wire n20219;
wire n20220;
wire n20221;
wire n20222;
wire n20223;
wire n20224;
wire n20225;
wire n20226;
wire n20227;
wire n20228;
wire n20229;
wire n20230;
wire n20231;
wire n20232;
wire n20233;
wire n20234;
wire n20235;
wire n20236;
wire n20237;
wire n20238;
wire n20239;
wire n20240;
wire n20241;
wire n20242;
wire n20243;
wire n20244;
wire n20245;
wire n20246;
wire n20247;
wire n20248;
wire n20249;
wire n20250;
wire n20251;
wire n20252;
wire n20253;
wire n20254;
wire n20255;
wire n20256;
wire n20257;
wire n20258;
wire n20259;
wire n20260;
wire n20261;
wire n20262;
wire n20263;
wire n20264;
wire n20265;
wire n20266;
wire n20267;
wire n20268;
wire n20269;
wire n20270;
wire n20271;
wire n20272;
wire n20273;
wire n20274;
wire n20275;
wire n20276;
wire n20277;
wire n20278;
wire n20279;
wire n20280;
wire n20281;
wire n20282;
wire n20283;
wire n20284;
wire n20285;
wire n20286;
wire n20287;
wire n20288;
wire n20289;
wire n20290;
wire n20291;
wire n20292;
wire n20293;
wire n20294;
wire n20295;
wire n20296;
wire n20297;
wire n20298;
wire n20299;
wire n20300;
wire n20301;
wire n20302;
wire n20303;
wire n20304;
wire n20305;
wire n20306;
wire n20307;
wire n20308;
wire n20309;
wire n20310;
wire n20311;
wire n20312;
wire n20313;
wire n20314;
wire n20315;
wire n20316;
wire n20317;
wire n20318;
wire n20319;
wire n20320;
wire n20321;
wire n20322;
wire n20323;
wire n20324;
wire n20325;
wire n20326;
wire n20327;
wire n20328;
wire n20329;
wire n20330;
wire n20331;
wire n20332;
wire n20333;
wire n20334;
wire n20335;
wire n20336;
wire n20337;
wire n20338;
wire n20339;
wire n20340;
wire n20341;
wire n20342;
wire n20343;
wire n20344;
wire n20345;
wire n20346;
wire n20347;
wire n20348;
wire n20349;
wire n20350;
wire n20351;
wire n20352;
wire n20353;
wire n20354;
wire n20355;
wire n20356;
wire n20357;
wire n20358;
wire n20359;
wire n20360;
wire n20361;
wire n20362;
wire n20363;
wire n20364;
wire n20365;
wire n20366;
wire n20367;
wire n20368;
wire n20369;
wire n20370;
wire n20371;
wire n20372;
wire n20373;
wire n20374;
wire n20375;
wire n20376;
wire n20377;
wire n20378;
wire n20379;
wire n20380;
wire n20381;
wire n20382;
wire n20383;
wire n20384;
wire n20385;
wire n20386;
wire n20387;
wire n20388;
wire n20389;
wire n20390;
wire n20391;
wire n20392;
wire n20393;
wire n20394;
wire n20395;
wire n20396;
wire n20397;
wire n20398;
wire n20399;
wire n20400;
wire n20401;
wire n20402;
wire n20403;
wire n20404;
wire n20405;
wire n20406;
wire n20407;
wire n20408;
wire n20409;
wire n20410;
wire n20411;
wire n20412;
wire n20413;
wire n20414;
wire n20415;
wire n20416;
wire n20417;
wire n20418;
wire n20419;
wire n20420;
wire n20421;
wire n20422;
wire n20423;
wire n20424;
wire n20425;
wire n20426;
wire n20427;
wire n20428;
wire n20429;
wire n20430;
wire n20431;
wire n20432;
wire n20433;
wire n20434;
wire n20435;
wire n20436;
wire n20437;
wire n20438;
wire n20439;
wire n20440;
wire n20441;
wire n20442;
wire n20443;
wire n20444;
wire n20445;
wire n20446;
wire n20447;
wire n20448;
wire n20449;
wire n20450;
wire n20451;
wire n20452;
wire n20453;
wire n20454;
wire n20455;
wire n20456;
wire n20457;
wire n20458;
wire n20459;
wire n20460;
wire n20461;
wire n20462;
wire n20463;
wire n20464;
wire n20465;
wire n20466;
wire n20467;
wire n20468;
wire n20469;
wire n20470;
wire n20471;
wire n20472;
wire n20473;
wire n20474;
wire n20475;
wire n20476;
wire n20477;
wire n20478;
wire n20479;
wire n20480;
wire n20481;
wire n20482;
wire n20483;
wire n20484;
wire n20485;
wire n20486;
wire n20487;
wire n20488;
wire n20489;
wire n20490;
wire n20491;
wire n20492;
wire n20493;
wire n20494;
wire n20495;
wire n20496;
wire n20497;
wire n20498;
wire n20499;
wire n20500;
wire n20501;
wire n20502;
wire n20503;
wire n20504;
wire n20505;
wire n20506;
wire n20507;
wire n20508;
wire n20509;
wire n20510;
wire n20511;
wire n20512;
wire n20513;
wire n20514;
wire n20515;
wire n20516;
wire n20517;
wire n20518;
wire n20519;
wire n20520;
wire n20521;
wire n20522;
wire n20523;
wire n20524;
wire n20525;
wire n20526;
wire n20527;
wire n20528;
wire n20529;
wire n20530;
wire n20531;
wire n20532;
wire n20533;
wire n20534;
wire n20535;
wire n20536;
wire n20537;
wire n20538;
wire n20539;
wire n20540;
wire n20541;
wire n20542;
wire n20543;
wire n20544;
wire n20545;
wire n20546;
wire n20547;
wire n20548;
wire n20549;
wire n20550;
wire n20551;
wire n20552;
wire n20553;
wire n20554;
wire n20555;
wire n20556;
wire n20557;
wire n20558;
wire n20559;
wire n20560;
wire n20561;
wire n20562;
wire n20563;
wire n20564;
wire n20565;
wire n20566;
wire n20567;
wire n20568;
wire n20569;
wire n20570;
wire n20571;
wire n20572;
wire n20573;
wire n20574;
wire n20575;
wire n20576;
wire n20577;
wire n20578;
wire n20579;
wire n20580;
wire n20581;
wire n20582;
wire n20583;
wire n20584;
wire n20585;
wire n20586;
wire n20587;
wire n20588;
wire n20589;
wire n20590;
wire n20591;
wire n20592;
wire n20593;
wire n20594;
wire n20595;
wire n20596;
wire n20597;
wire n20598;
wire n20599;
wire n20600;
wire n20601;
wire n20602;
wire n20603;
wire n20604;
wire n20605;
wire n20606;
wire n20607;
wire n20608;
wire n20609;
wire n20610;
wire n20611;
wire n20612;
wire n20613;
wire n20614;
wire n20615;
wire n20616;
wire n20617;
wire n20618;
wire n20619;
wire n20620;
wire n20621;
wire n20622;
wire n20623;
wire n20624;
wire n20625;
wire n20626;
wire n20627;
wire n20628;
wire n20629;
wire n20630;
wire n20631;
wire n20632;
wire n20633;
wire n20634;
wire n20635;
wire n20636;
wire n20637;
wire n20638;
wire n20639;
wire n20640;
wire n20641;
wire n20642;
wire n20643;
wire n20644;
wire n20645;
wire n20646;
wire n20647;
wire n20648;
wire n20649;
wire n20650;
wire n20651;
wire n20652;
wire n20653;
wire n20654;
wire n20655;
wire n20656;
wire n20657;
wire n20658;
wire n20659;
wire n20660;
wire n20661;
wire n20662;
wire n20663;
wire n20664;
wire n20665;
wire n20666;
wire n20667;
wire n20668;
wire n20669;
wire n20670;
wire n20671;
wire n20672;
wire n20673;
wire n20674;
wire n20675;
wire n20676;
wire n20677;
wire n20678;
wire n20679;
wire n20680;
wire n20681;
wire n20682;
wire n20683;
wire n20684;
wire n20685;
wire n20686;
wire n20687;
wire n20688;
wire n20689;
wire n20690;
wire n20691;
wire n20692;
wire n20693;
wire n20694;
wire n20695;
wire n20696;
wire n20697;
wire n20698;
wire n20699;
wire n20700;
wire n20701;
wire n20702;
wire n20703;
wire n20704;
wire n20705;
wire n20706;
wire n20707;
wire n20708;
wire n20709;
wire n20710;
wire n20711;
wire n20712;
wire n20713;
wire n20714;
wire n20715;
wire n20716;
wire n20717;
wire n20718;
wire n20719;
wire n20720;
wire n20721;
wire n20722;
wire n20723;
wire n20724;
wire n20725;
wire n20726;
wire n20727;
wire n20728;
wire n20729;
wire n20730;
wire n20731;
wire n20732;
wire n20733;
wire n20734;
wire n20735;
wire n20736;
wire n20737;
wire n20738;
wire n20739;
wire n20740;
wire n20741;
wire n20742;
wire n20743;
wire n20744;
wire n20745;
wire n20746;
wire n20747;
wire n20748;
wire n20749;
wire n20750;
wire n20751;
wire n20752;
wire n20753;
wire n20754;
wire n20755;
wire n20756;
wire n20757;
wire n20758;
wire n20759;
wire n20760;
wire n20761;
wire n20762;
wire n20763;
wire n20764;
wire n20765;
wire n20766;
wire n20767;
wire n20768;
wire n20769;
wire n20770;
wire n20771;
wire n20772;
wire n20773;
wire n20774;
wire n20775;
wire n20776;
wire n20777;
wire n20778;
wire n20779;
wire n20780;
wire n20781;
wire n20782;
wire n20783;
wire n20784;
wire n20785;
wire n20786;
wire n20787;
wire n20788;
wire n20789;
wire n20790;
wire n20791;
wire n20792;
wire n20793;
wire n20794;
wire n20795;
wire n20796;
wire n20797;
wire n20798;
wire n20799;
wire n20800;
wire n20801;
wire n20802;
wire n20803;
wire n20804;
wire n20805;
wire n20806;
wire n20807;
wire n20808;
wire n20809;
wire n20810;
wire n20811;
wire n20812;
wire n20813;
wire n20814;
wire n20815;
wire n20816;
wire n20817;
wire n20818;
wire n20819;
wire n20820;
wire n20821;
wire n20822;
wire n20823;
wire n20824;
wire n20825;
wire n20826;
wire n20827;
wire n20828;
wire n20829;
wire n20830;
wire n20831;
wire n20832;
wire n20833;
wire n20834;
wire n20835;
wire n20836;
wire n20837;
wire n20838;
wire n20839;
wire n20840;
wire n20841;
wire n20842;
wire n20843;
wire n20844;
wire n20845;
wire n20846;
wire n20847;
wire n20848;
wire n20849;
wire n20850;
wire n20851;
wire n20852;
wire n20853;
wire n20854;
wire n20855;
wire n20856;
wire n20857;
wire n20858;
wire n20859;
wire n20860;
wire n20861;
wire n20862;
wire n20863;
wire n20864;
wire n20865;
wire n20866;
wire n20867;
wire n20868;
wire n20869;
wire n20870;
wire n20871;
wire n20872;
wire n20873;
wire n20874;
wire n20875;
wire n20876;
wire n20877;
wire n20878;
wire n20879;
wire n20880;
wire n20881;
wire n20882;
wire n20883;
wire n20884;
wire n20885;
wire n20886;
wire n20887;
wire n20888;
wire n20889;
wire n20890;
wire n20891;
wire n20892;
wire n20893;
wire n20894;
wire n20895;
wire n20896;
wire n20897;
wire n20898;
wire n20899;
wire n20900;
wire n20901;
wire n20902;
wire n20903;
wire n20904;
wire n20905;
wire n20906;
wire n20907;
wire n20908;
wire n20909;
wire n20910;
wire n20911;
wire n20912;
wire n20913;
wire n20914;
wire n20915;
wire n20916;
wire n20917;
wire n20918;
wire n20919;
wire n20920;
wire n20921;
wire n20922;
wire n20923;
wire n20924;
wire n20925;
wire n20926;
wire n20927;
wire n20928;
wire n20929;
wire n20930;
wire n20931;
wire n20932;
wire n20933;
wire n20934;
wire n20935;
wire n20936;
wire n20937;
wire n20938;
wire n20939;
wire n20940;
wire n20941;
wire n20942;
wire n20943;
wire n20944;
wire n20945;
wire n20946;
wire n20947;
wire n20948;
wire n20949;
wire n20950;
wire n20951;
wire n20952;
wire n20953;
wire n20954;
wire n20955;
wire n20956;
wire n20957;
wire n20958;
wire n20959;
wire n20960;
wire n20961;
wire n20962;
wire n20963;
wire n20964;
wire n20965;
wire n20966;
wire n20967;
wire n20968;
wire n20969;
wire n20970;
wire n20971;
wire n20972;
wire n20973;
wire n20974;
wire n20975;
wire n20976;
wire n20977;
wire n20978;
wire n20979;
wire n20980;
wire n20981;
wire n20982;
wire n20983;
wire n20984;
wire n20985;
wire n20986;
wire n20987;
wire n20988;
wire n20989;
wire n20990;
wire n20991;
wire n20992;
wire n20993;
wire n20994;
wire n20995;
wire n20996;
wire n20997;
wire n20998;
wire n20999;
wire n21000;
wire n21001;
wire n21002;
wire n21003;
wire n21004;
wire n21005;
wire n21006;
wire n21007;
wire n21008;
wire n21009;
wire n21010;
wire n21011;
wire n21012;
wire n21013;
wire n21014;
wire n21015;
wire n21016;
wire n21017;
wire n21018;
wire n21019;
wire n21020;
wire n21021;
wire n21022;
wire n21023;
wire n21024;
wire n21025;
wire n21026;
wire n21027;
wire n21028;
wire n21029;
wire n21030;
wire n21031;
wire n21032;
wire n21033;
wire n21034;
wire n21035;
wire n21036;
wire n21037;
wire n21038;
wire n21039;
wire n21040;
wire n21041;
wire n21042;
wire n21043;
wire n21044;
wire n21045;
wire n21046;
wire n21047;
wire n21048;
wire n21049;
wire n21050;
wire n21051;
wire n21052;
wire n21053;
wire n21054;
wire n21055;
wire n21056;
wire n21057;
wire n21058;
wire n21059;
wire n21060;
wire n21061;
wire n21062;
wire n21063;
wire n21064;
wire n21065;
wire n21066;
wire n21067;
wire n21068;
wire n21069;
wire n21070;
wire n21071;
wire n21072;
wire n21073;
wire n21074;
wire n21075;
wire n21076;
wire n21077;
wire n21078;
wire n21079;
wire n21080;
wire n21081;
wire n21082;
wire n21083;
wire n21084;
wire n21085;
wire n21086;
wire n21087;
wire n21088;
wire n21089;
wire n21090;
wire n21091;
wire n21092;
wire n21093;
wire n21094;
wire n21095;
wire n21096;
wire n21097;
wire n21098;
wire n21099;
wire n21100;
wire n21101;
wire n21102;
wire n21103;
wire n21104;
wire n21105;
wire n21106;
wire n21107;
wire n21108;
wire n21109;
wire n21110;
wire n21111;
wire n21112;
wire n21113;
wire n21114;
wire n21115;
wire n21116;
wire n21117;
wire n21118;
wire n21119;
wire n21120;
wire n21121;
wire n21122;
wire n21123;
wire n21124;
wire n21125;
wire n21126;
wire n21127;
wire n21128;
wire n21129;
wire n21130;
wire n21131;
wire n21132;
wire n21133;
wire n21134;
wire n21135;
wire n21136;
wire n21137;
wire n21138;
wire n21139;
wire n21140;
wire n21141;
wire n21142;
wire n21143;
wire n21144;
wire n21145;
wire n21146;
wire n21147;
wire n21148;
wire n21149;
wire n21150;
wire n21151;
wire n21152;
wire n21153;
wire n21154;
wire n21155;
wire n21156;
wire n21157;
wire n21158;
wire n21159;
wire n21160;
wire n21161;
wire n21162;
wire n21163;
wire n21164;
wire n21165;
wire n21166;
wire n21167;
wire n21168;
wire n21169;
wire n21170;
wire n21171;
wire n21172;
wire n21173;
wire n21174;
wire n21175;
wire n21176;
wire n21177;
wire n21178;
wire n21179;
wire n21180;
wire n21181;
wire n21182;
wire n21183;
wire n21184;
wire n21185;
wire n21186;
wire n21187;
wire n21188;
wire n21189;
wire n21190;
wire n21191;
wire n21192;
wire n21193;
wire n21194;
wire n21195;
wire n21196;
wire n21197;
wire n21198;
wire n21199;
wire n21200;
wire n21201;
wire n21202;
wire n21203;
wire n21204;
wire n21205;
wire n21206;
wire n21207;
wire n21208;
wire n21209;
wire n21210;
wire n21211;
wire n21212;
wire n21213;
wire n21214;
wire n21215;
wire n21216;
wire n21217;
wire n21218;
wire n21219;
wire n21220;
wire n21221;
wire n21222;
wire n21223;
wire n21224;
wire n21225;
wire n21226;
wire n21227;
wire n21228;
wire n21229;
wire n21230;
wire n21231;
wire n21232;
wire n21233;
wire n21234;
wire n21235;
wire n21236;
wire n21237;
wire n21238;
wire n21239;
wire n21240;
wire n21241;
wire n21242;
wire n21243;
wire n21244;
wire n21245;
wire n21246;
wire n21247;
wire n21248;
wire n21249;
wire n21250;
wire n21251;
wire n21252;
wire n21253;
wire n21254;
wire n21255;
wire n21256;
wire n21257;
wire n21258;
wire n21259;
wire n21260;
wire n21261;
wire n21262;
wire n21263;
wire n21264;
wire n21265;
wire n21266;
wire n21267;
wire n21268;
wire n21269;
wire n21270;
wire n21271;
wire n21272;
wire n21273;
wire n21274;
wire n21275;
wire n21276;
wire n21277;
wire n21278;
wire n21279;
wire n21280;
wire n21281;
wire n21282;
wire n21283;
wire n21284;
wire n21285;
wire n21286;
wire n21287;
wire n21288;
wire n21289;
wire n21290;
wire n21291;
wire n21292;
wire n21293;
wire n21294;
wire n21295;
wire n21296;
wire n21297;
wire n21298;
wire n21299;
wire n21300;
wire n21301;
wire n21302;
wire n21303;
wire n21304;
wire n21305;
wire n21306;
wire n21307;
wire n21308;
wire n21309;
wire n21310;
wire n21311;
wire n21312;
wire n21313;
wire n21314;
wire n21315;
wire n21316;
wire n21317;
wire n21318;
wire n21319;
wire n21320;
wire n21321;
wire n21322;
wire n21323;
wire n21324;
wire n21325;
wire n21326;
wire n21327;
wire n21328;
wire n21329;
wire n21330;
wire n21331;
wire n21332;
wire n21333;
wire n21334;
wire n21335;
wire n21336;
wire n21337;
wire n21338;
wire n21339;
wire n21340;
wire n21341;
wire n21342;
wire n21343;
wire n21344;
wire n21345;
wire n21346;
wire n21347;
wire n21348;
wire n21349;
wire n21350;
wire n21351;
wire n21352;
wire n21353;
wire n21354;
wire n21355;
wire n21356;
wire n21357;
wire n21358;
wire n21359;
wire n21360;
wire n21361;
wire n21362;
wire n21363;
wire n21364;
wire n21365;
wire n21366;
wire n21367;
wire n21368;
wire n21369;
wire n21370;
wire n21371;
wire n21372;
wire n21373;
wire n21374;
wire n21375;
wire n21376;
wire n21377;
wire n21378;
wire n21379;
wire n21380;
wire n21381;
wire n21382;
wire n21383;
wire n21384;
wire n21385;
wire n21386;
wire n21387;
wire n21388;
wire n21389;
wire n21390;
wire n21391;
wire n21392;
wire n21393;
wire n21394;
wire n21395;
wire n21396;
wire n21397;
wire n21398;
wire n21399;
wire n21400;
wire n21401;
wire n21402;
wire n21403;
wire n21404;
wire n21405;
wire n21406;
wire n21407;
wire n21408;
wire n21409;
wire n21410;
wire n21411;
wire n21412;
wire n21413;
wire n21414;
wire n21415;
wire n21416;
wire n21417;
wire n21418;
wire n21419;
wire n21420;
wire n21421;
wire n21422;
wire n21423;
wire n21424;
wire n21425;
wire n21426;
wire n21427;
wire n21428;
wire n21429;
wire n21430;
wire n21431;
wire n21432;
wire n21433;
wire n21434;
wire n21435;
wire n21436;
wire n21437;
wire n21438;
wire n21439;
wire n21440;
wire n21441;
wire n21442;
wire n21443;
wire n21444;
wire n21445;
wire n21446;
wire n21447;
wire n21448;
wire n21449;
wire n21450;
wire n21451;
wire n21452;
wire n21453;
wire n21454;
wire n21455;
wire n21456;
wire n21457;
wire n21458;
wire n21459;
wire n21460;
wire n21461;
wire n21462;
wire n21463;
wire n21464;
wire n21465;
wire n21466;
wire n21467;
wire n21468;
wire n21469;
wire n21470;
wire n21471;
wire n21472;
wire n21473;
wire n21474;
wire n21475;
wire n21476;
wire n21477;
wire n21478;
wire n21479;
wire n21480;
wire n21481;
wire n21482;
wire n21483;
wire n21484;
wire n21485;
wire n21486;
wire n21487;
wire n21488;
wire n21489;
wire n21490;
wire n21491;
wire n21492;
wire n21493;
wire n21494;
wire n21495;
wire n21496;
wire n21497;
wire n21498;
wire n21499;
wire n21500;
wire n21501;
wire n21502;
wire n21503;
wire n21504;
wire n21505;
wire n21506;
wire n21507;
wire n21508;
wire n21509;
wire n21510;
wire n21511;
wire n21512;
wire n21513;
wire n21514;
wire n21515;
wire n21516;
wire n21517;
wire n21518;
wire n21519;
wire n21520;
wire n21521;
wire n21522;
wire n21523;
wire n21524;
wire n21525;
wire n21526;
wire n21527;
wire n21528;
wire n21529;
wire n21530;
wire n21531;
wire n21532;
wire n21533;
wire n21534;
wire n21535;
wire n21536;
wire n21537;
wire n21538;
wire n21539;
wire n21540;
wire n21541;
wire n21542;
wire n21543;
wire n21544;
wire n21545;
wire n21546;
wire n21547;
wire n21548;
wire n21549;
wire n21550;
wire n21551;
wire n21552;
wire n21553;
wire n21554;
wire n21555;
wire n21556;
wire n21557;
wire n21558;
wire n21559;
wire n21560;
wire n21561;
wire n21562;
wire n21563;
wire n21564;
wire n21565;
wire n21566;
wire n21567;
wire n21568;
wire n21569;
wire n21570;
wire n21571;
wire n21572;
wire n21573;
wire n21574;
wire n21575;
wire n21576;
wire n21577;
wire n21578;
wire n21579;
wire n21580;
wire n21581;
wire n21582;
wire n21583;
wire n21584;
wire n21585;
wire n21586;
wire n21587;
wire n21588;
wire n21589;
wire n21590;
wire n21591;
wire n21592;
wire n21593;
wire n21594;
wire n21595;
wire n21596;
wire n21597;
wire n21598;
wire n21599;
wire n21600;
wire n21601;
wire n21602;
wire n21603;
wire n21604;
wire n21605;
wire n21606;
wire n21607;
wire n21608;
wire n21609;
wire n21610;
wire n21611;
wire n21612;
wire n21613;
wire n21614;
wire n21615;
wire n21616;
wire n21617;
wire n21618;
wire n21619;
wire n21620;
wire n21621;
wire n21622;
wire n21623;
wire n21624;
wire n21625;
wire n21626;
wire n21627;
wire n21628;
wire n21629;
wire n21630;
wire n21631;
wire n21632;
wire n21633;
wire n21634;
wire n21635;
wire n21636;
wire n21637;
wire n21638;
wire n21639;
wire n21640;
wire n21641;
wire n21642;
wire n21643;
wire n21644;
wire n21645;
wire n21646;
wire n21647;
wire n21648;
wire n21649;
wire n21650;
wire n21651;
wire n21652;
wire n21653;
wire n21654;
wire n21655;
wire n21656;
wire n21657;
wire n21658;
wire n21659;
wire n21660;
wire n21661;
wire n21662;
wire n21663;
wire n21664;
wire n21665;
wire n21666;
wire n21667;
wire n21668;
wire n21669;
wire n21670;
wire n21671;
wire n21672;
wire n21673;
wire n21674;
wire n21675;
wire n21676;
wire n21677;
wire n21678;
wire n21679;
wire n21680;
wire n21681;
wire n21682;
wire n21683;
wire n21684;
wire n21685;
wire n21686;
wire n21687;
wire n21688;
wire n21689;
wire n21690;
wire n21691;
wire n21692;
wire n21693;
wire n21694;
wire n21695;
wire n21696;
wire n21697;
wire n21698;
wire n21699;
wire n21700;
wire n21701;
wire n21702;
wire n21703;
wire n21704;
wire n21705;
wire n21706;
wire n21707;
wire n21708;
wire n21709;
wire n21710;
wire n21711;
wire n21712;
wire n21713;
wire n21714;
wire n21715;
wire n21716;
wire n21717;
wire n21718;
wire n21719;
wire n21720;
wire n21721;
wire n21722;
wire n21723;
wire n21724;
wire n21725;
wire n21726;
wire n21727;
wire n21728;
wire n21729;
wire n21730;
wire n21731;
wire n21732;
wire n21733;
wire n21734;
wire n21735;
wire n21736;
wire n21737;
wire n21738;
wire n21739;
wire n21740;
wire n21741;
wire n21742;
wire n21743;
wire n21744;
wire n21745;
wire n21746;
wire n21747;
wire n21748;
wire n21749;
wire n21750;
wire n21751;
wire n21752;
wire n21753;
wire n21754;
wire n21755;
wire n21756;
wire n21757;
wire n21758;
wire n21759;
wire n21760;
wire n21761;
wire n21762;
wire n21763;
wire n21764;
wire n21765;
wire n21766;
wire n21767;
wire n21768;
wire n21769;
wire n21770;
wire n21771;
wire n21772;
wire n21773;
wire n21774;
wire n21775;
wire n21776;
wire n21777;
wire n21778;
wire n21779;
wire n21780;
wire n21781;
wire n21782;
wire n21783;
wire n21784;
wire n21785;
wire n21786;
wire n21787;
wire n21788;
wire n21789;
wire n21790;
wire n21791;
wire n21792;
wire n21793;
wire n21794;
wire n21795;
wire n21796;
wire n21797;
wire n21798;
wire n21799;
wire n21800;
wire n21801;
wire n21802;
wire n21803;
wire n21804;
wire n21805;
wire n21806;
wire n21807;
wire n21808;
wire n21809;
wire n21810;
wire n21811;
wire n21812;
wire n21813;
wire n21814;
wire n21815;
wire n21816;
wire n21817;
wire n21818;
wire n21819;
wire n21820;
wire n21821;
wire n21822;
wire n21823;
wire n21824;
wire n21825;
wire n21826;
wire n21827;
wire n21828;
wire n21829;
wire n21830;
wire n21831;
wire n21832;
wire n21833;
wire n21834;
wire n21835;
wire n21836;
wire n21837;
wire n21838;
wire n21839;
wire n21840;
wire n21841;
wire n21842;
wire n21843;
wire n21844;
wire n21845;
wire n21846;
wire n21847;
wire n21848;
wire n21849;
wire n21850;
wire n21851;
wire n21852;
wire n21853;
wire n21854;
wire n21855;
wire n21856;
wire n21857;
wire n21858;
wire n21859;
wire n21860;
wire n21861;
wire n21862;
wire n21863;
wire n21864;
wire n21865;
wire n21866;
wire n21867;
wire n21868;
wire n21869;
wire n21870;
wire n21871;
wire n21872;
wire n21873;
wire n21874;
wire n21875;
wire n21876;
wire n21877;
wire n21878;
wire n21879;
wire n21880;
wire n21881;
wire n21882;
wire n21883;
wire n21884;
wire n21885;
wire n21886;
wire n21887;
wire n21888;
wire n21889;
wire n21890;
wire n21891;
wire n21892;
wire n21893;
wire n21894;
wire n21895;
wire n21896;
wire n21897;
wire n21898;
wire n21899;
wire n21900;
wire n21901;
wire n21902;
wire n21903;
wire n21904;
wire n21905;
wire n21906;
wire n21907;
wire n21908;
wire n21909;
wire n21910;
wire n21911;
wire n21912;
wire n21913;
wire n21914;
wire n21915;
wire n21916;
wire n21917;
wire n21918;
wire n21919;
wire n21920;
wire n21921;
wire n21922;
wire n21923;
wire n21924;
wire n21925;
wire n21926;
wire n21927;
wire n21928;
wire n21929;
wire n21930;
wire n21931;
wire n21932;
wire n21933;
wire n21934;
wire n21935;
wire n21936;
wire n21937;
wire n21938;
wire n21939;
wire n21940;
wire n21941;
wire n21942;
wire n21943;
wire n21944;
wire n21945;
wire n21946;
wire n21947;
wire n21948;
wire n21949;
wire n21950;
wire n21951;
wire n21952;
wire n21953;
wire n21954;
wire n21955;
wire n21956;
wire n21957;
wire n21958;
wire n21959;
wire n21960;
wire n21961;
wire n21962;
wire n21963;
wire n21964;
wire n21965;
wire n21966;
wire n21967;
wire n21968;
wire n21969;
wire n21970;
wire n21971;
wire n21972;
wire n21973;
wire n21974;
wire n21975;
wire n21976;
wire n21977;
wire n21978;
wire n21979;
wire n21980;
wire n21981;
wire n21982;
wire n21983;
wire n21984;
wire n21985;
wire n21986;
wire n21987;
wire n21988;
wire n21989;
wire n21990;
wire n21991;
wire n21992;
wire n21993;
wire n21994;
wire n21995;
wire n21996;
wire n21997;
wire n21998;
wire n21999;
wire n22000;
wire n22001;
wire n22002;
wire n22003;
wire n22004;
wire n22005;
wire n22006;
wire n22007;
wire n22008;
wire n22009;
wire n22010;
wire n22011;
wire n22012;
wire n22013;
wire n22014;
wire n22015;
wire n22016;
wire n22017;
wire n22018;
wire n22019;
wire n22020;
wire n22021;
wire n22022;
wire n22023;
wire n22024;
wire n22025;
wire n22026;
wire n22027;
wire n22028;
wire n22029;
wire n22030;
wire n22031;
wire n22032;
wire n22033;
wire n22034;
wire n22035;
wire n22036;
wire n22037;
wire n22038;
wire n22039;
wire n22040;
wire n22041;
wire n22042;
wire n22043;
wire n22044;
wire n22045;
wire n22046;
wire n22047;
wire n22048;
wire n22049;
wire n22050;
wire n22051;
wire n22052;
wire n22053;
wire n22054;
wire n22055;
wire n22056;
wire n22057;
wire n22058;
wire n22059;
wire n22060;
wire n22061;
wire n22062;
wire n22063;
wire n22064;
wire n22065;
wire n22066;
wire n22067;
wire n22068;
wire n22069;
wire n22070;
wire n22071;
wire n22072;
wire n22073;
wire n22074;
wire n22075;
wire n22076;
wire n22077;
wire n22078;
wire n22079;
wire n22080;
wire n22081;
wire n22082;
wire n22083;
wire n22084;
wire n22085;
wire n22086;
wire n22087;
wire n22088;
wire n22089;
wire n22090;
wire n22091;
wire n22092;
wire n22093;
wire n22094;
wire n22095;
wire n22096;
wire n22097;
wire n22098;
wire n22099;
wire n22100;
wire n22101;
wire n22102;
wire n22103;
wire n22104;
wire n22105;
wire n22106;
wire n22107;
wire n22108;
wire n22109;
wire n22110;
wire n22111;
wire n22112;
wire n22113;
wire n22114;
wire n22115;
wire n22116;
wire n22117;
wire n22118;
wire n22119;
wire n22120;
wire n22121;
wire n22122;
wire n22123;
wire n22124;
wire n22125;
wire n22126;
wire n22127;
wire n22128;
wire n22129;
wire n22130;
wire n22131;
wire n22132;
wire n22133;
wire n22134;
wire n22135;
wire n22136;
wire n22137;
wire n22138;
wire n22139;
wire n22140;
wire n22141;
wire n22142;
wire n22143;
wire n22144;
wire n22145;
wire n22146;
wire n22147;
wire n22148;
wire n22149;
wire n22150;
wire n22151;
wire n22152;
wire n22153;
wire n22154;
wire n22155;
wire n22156;
wire n22157;
wire n22158;
wire n22159;
wire n22160;
wire n22161;
wire n22162;
wire n22163;
wire n22164;
wire n22165;
wire n22166;
wire n22167;
wire n22168;
wire n22169;
wire n22170;
wire n22171;
wire n22172;
wire n22173;
wire n22174;
wire n22175;
wire n22176;
wire n22177;
wire n22178;
wire n22179;
wire n22180;
wire n22181;
wire n22182;
wire n22183;
wire n22184;
wire n22185;
wire n22186;
wire n22187;
wire n22188;
wire n22189;
wire n22190;
wire n22191;
wire n22192;
wire n22193;
wire n22194;
wire n22195;
wire n22196;
wire n22197;
wire n22198;
wire n22199;
wire n22200;
wire n22201;
wire n22202;
wire n22203;
wire n22204;
wire n22205;
wire n22206;
wire n22207;
wire n22208;
wire n22209;
wire n22210;
wire n22211;
wire n22212;
wire n22213;
wire n22214;
wire n22215;
wire n22216;
wire n22217;
wire n22218;
wire n22219;
wire n22220;
wire n22221;
wire n22222;
wire n22223;
wire n22224;
wire n22225;
wire n22226;
wire n22227;
wire n22228;
wire n22229;
wire n22230;
wire n22231;
wire n22232;
wire n22233;
wire n22234;
wire n22235;
wire n22236;
wire n22237;
wire n22238;
wire n22239;
wire n22240;
wire n22241;
wire n22242;
wire n22243;
wire n22244;
wire n22245;
wire n22246;
wire n22247;
wire n22248;
wire n22249;
wire n22250;
wire n22251;
wire n22252;
wire n22253;
wire n22254;
wire n22255;
wire n22256;
wire n22257;
wire n22258;
wire n22259;
wire n22260;
wire n22261;
wire n22262;
wire n22263;
wire n22264;
wire n22265;
wire n22266;
wire n22267;
wire n22268;
wire n22269;
wire n22270;
wire n22271;
wire n22272;
wire n22273;
wire n22274;
wire n22275;
wire n22276;
wire n22277;
wire n22278;
wire n22279;
wire n22280;
wire n22281;
wire n22282;
wire n22283;
wire n22284;
wire n22285;
wire n22286;
wire n22287;
wire n22288;
wire n22289;
wire n22290;
wire n22291;
wire n22292;
wire n22293;
wire n22294;
wire n22295;
wire n22296;
wire n22297;
wire n22298;
wire n22299;
wire n22300;
wire n22301;
wire n22302;
wire n22303;
wire n22304;
wire n22305;
wire n22306;
wire n22307;
wire n22308;
wire n22309;
wire n22310;
wire n22311;
wire n22312;
wire n22313;
wire n22314;
wire n22315;
wire n22316;
wire n22317;
wire n22318;
wire n22319;
wire n22320;
wire n22321;
wire n22322;
wire n22323;
wire n22324;
wire n22325;
wire n22326;
wire n22327;
wire n22328;
wire n22329;
wire n22330;
wire n22331;
wire n22332;
wire n22333;
wire n22334;
wire n22335;
wire n22336;
wire n22337;
wire n22338;
wire n22339;
wire n22340;
wire n22341;
wire n22342;
wire n22343;
wire n22344;
wire n22345;
wire n22346;
wire n22347;
wire n22348;
wire n22349;
wire n22350;
wire n22351;
wire n22352;
wire n22353;
wire n22354;
wire n22355;
wire n22356;
wire n22357;
wire n22358;
wire n22359;
wire n22360;
wire n22361;
wire n22362;
wire n22363;
wire n22364;
wire n22365;
wire n22366;
wire n22367;
wire n22368;
wire n22369;
wire n22370;
wire n22371;
wire n22372;
wire n22373;
wire n22374;
wire n22375;
wire n22376;
wire n22377;
wire n22378;
wire n22379;
wire n22380;
wire n22381;
wire n22382;
wire n22383;
wire n22384;
wire n22385;
wire n22386;
wire n22387;
wire n22388;
wire n22389;
wire n22390;
wire n22391;
wire n22392;
wire n22393;
wire n22394;
wire n22395;
wire n22396;
wire n22397;
wire n22398;
wire n22399;
wire n22400;
wire n22401;
wire n22402;
wire n22403;
wire n22404;
wire n22405;
wire n22406;
wire n22407;
wire n22408;
wire n22409;
wire n22410;
wire n22411;
wire n22412;
wire n22413;
wire n22414;
wire n22415;
wire n22416;
wire n22417;
wire n22418;
wire n22419;
wire n22420;
wire n22421;
wire n22422;
wire n22423;
wire n22424;
wire n22425;
wire n22426;
wire n22427;
wire n22428;
wire n22429;
wire n22430;
wire n22431;
wire n22432;
wire n22433;
wire n22434;
wire n22435;
wire n22436;
wire n22437;
wire n22438;
wire n22439;
wire n22440;
wire n22441;
wire n22442;
wire n22443;
wire n22444;
wire n22445;
wire n22446;
wire n22447;
wire n22448;
wire n22449;
wire n22450;
wire n22451;
wire n22452;
wire n22453;
wire n22454;
wire n22455;
wire n22456;
wire n22457;
wire n22458;
wire n22459;
wire n22460;
wire n22461;
wire n22462;
wire n22463;
wire n22464;
wire n22465;
wire n22466;
wire n22467;
wire n22468;
wire n22469;
wire n22470;
wire n22471;
wire n22472;
wire n22473;
wire n22474;
wire n22475;
wire n22476;
wire n22477;
wire n22478;
wire n22479;
wire n22480;
wire n22481;
wire n22482;
wire n22483;
wire n22484;
wire n22485;
wire n22486;
wire n22487;
wire n22488;
wire n22489;
wire n22490;
wire n22491;
wire n22492;
wire n22493;
wire n22494;
wire n22495;
wire n22496;
wire n22497;
wire n22498;
wire n22499;
wire n22500;
wire n22501;
wire n22502;
wire n22503;
wire n22504;
wire n22505;
wire n22506;
wire n22507;
wire n22508;
wire n22509;
wire n22510;
wire n22511;
wire n22512;
wire n22513;
wire n22514;
wire n22515;
wire n22516;
wire n22517;
wire n22518;
wire n22519;
wire n22520;
wire n22521;
wire n22522;
wire n22523;
wire n22524;
wire n22525;
wire n22526;
wire n22527;
wire n22528;
wire n22529;
wire n22530;
wire n22531;
wire n22532;
wire n22533;
wire n22534;
wire n22535;
wire n22536;
wire n22537;
wire n22538;
wire n22539;
wire n22540;
wire n22541;
wire n22542;
wire n22543;
wire n22544;
wire n22545;
wire n22546;
wire n22547;
wire n22548;
wire n22549;
wire n22550;
wire n22551;
wire n22552;
wire n22553;
wire n22554;
wire n22555;
wire n22556;
wire n22557;
wire n22558;
wire n22559;
wire n22560;
wire n22561;
wire n22562;
wire n22563;
wire n22564;
wire n22565;
wire n22566;
wire n22567;
wire n22568;
wire n22569;
wire n22570;
wire n22571;
wire n22572;
wire n22573;
wire n22574;
wire n22575;
wire n22576;
wire n22577;
wire n22578;
wire n22579;
wire n22580;
wire n22581;
wire n22582;
wire n22583;
wire n22584;
wire n22585;
wire n22586;
wire n22587;
wire n22588;
wire n22589;
wire n22590;
wire n22591;
wire n22592;
wire n22593;
wire n22594;
wire n22595;
wire n22596;
wire n22597;
wire n22598;
wire n22599;
wire n22600;
wire n22601;
wire n22602;
wire n22603;
wire n22604;
wire n22605;
wire n22606;
wire n22607;
wire n22608;
wire n22609;
wire n22610;
wire n22611;
wire n22612;
wire n22613;
wire n22614;
wire n22615;
wire n22616;
wire n22617;
wire n22618;
wire n22619;
wire n22620;
wire n22621;
wire n22622;
wire n22623;
wire n22624;
wire n22625;
wire n22626;
wire n22627;
wire n22628;
wire n22629;
wire n22630;
wire n22631;
wire n22632;
wire n22633;
wire n22634;
wire n22635;
wire n22636;
wire n22637;
wire n22638;
wire n22639;
wire n22640;
wire n22641;
wire n22642;
wire n22643;
wire n22644;
wire n22645;
wire n22646;
wire n22647;
wire n22648;
wire n22649;
wire n22650;
wire n22651;
wire n22652;
wire n22653;
wire n22654;
wire n22655;
wire n22656;
wire n22657;
wire n22658;
wire n22659;
wire n22660;
wire n22661;
wire n22662;
wire n22663;
wire n22664;
wire n22665;
wire n22666;
wire n22667;
wire n22668;
wire n22669;
wire n22670;
wire n22671;
wire n22672;
wire n22673;
wire n22674;
wire n22675;
wire n22676;
wire n22677;
wire n22678;
wire n22679;
wire n22680;
wire n22681;
wire n22682;
wire n22683;
wire n22684;
wire n22685;
wire n22686;
wire n22687;
wire n22688;
wire n22689;
wire n22690;
wire n22691;
wire n22692;
wire n22693;
wire n22694;
wire n22695;
wire n22696;
wire n22697;
wire n22698;
wire n22699;
wire n22700;
wire n22701;
xor (out,n0,n10718);
nand (n0,n1,n10716);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
and (n5,n6,n10713);
nand (n6,n7,n10600);
not (n7,n8);
nor (n8,n9,n10463);
and (n9,n10,n10462);
nand (n10,n11,n3490,n7009);
not (n11,n12);
nor (n12,n13,n3483);
and (n13,n14,n3482);
nand (n14,n15,n2533,n3444,n3458);
nand (n15,n16,n1712);
nand (n16,n17,n1705);
or (n17,n18,n1395);
nor (n18,n19,n1394);
and (n19,n20,n1214);
not (n20,n21);
nor (n21,n22,n1201);
xor (n22,n23,n1035);
xor (n23,n24,n756);
xor (n24,n25,n616);
xor (n25,n26,n432);
or (n26,n27,n431);
and (n27,n28,n206);
xor (n28,n29,n110);
xor (n29,n30,n84);
xor (n30,n31,n56);
nand (n31,n32,n47);
or (n32,n33,n40);
not (n33,n34);
nand (n34,n35,n39);
or (n35,n36,n38);
not (n36,n37);
nand (n39,n36,n38);
not (n40,n41);
nand (n41,n42,n46);
or (n42,n43,n44);
not (n44,n45);
nand (n46,n44,n43);
nand (n47,n48,n51,n33);
nand (n48,n49,n50);
or (n49,n38,n44);
nand (n50,n44,n38);
nor (n51,n52,n54);
and (n52,n53,n45);
and (n54,n55,n44);
not (n55,n53);
nand (n56,n57,n78);
or (n57,n58,n65);
not (n58,n59);
nand (n59,n60,n64);
or (n60,n61,n63);
not (n61,n62);
nand (n64,n63,n61);
nand (n65,n66,n73);
or (n66,n67,n70);
not (n67,n68);
nand (n68,n61,n69);
not (n70,n71);
nand (n71,n72,n62);
not (n72,n69);
nor (n73,n74,n77);
and (n74,n75,n69);
not (n75,n76);
and (n77,n76,n72);
nand (n78,n79,n83);
nand (n79,n80,n82);
or (n80,n81,n61);
nand (n82,n81,n61);
not (n83,n73);
nand (n84,n85,n104);
or (n85,n86,n99);
nand (n86,n87,n94);
not (n87,n88);
nand (n88,n89,n93);
or (n89,n90,n92);
not (n90,n91);
nand (n93,n90,n92);
nand (n94,n95,n98);
or (n95,n96,n92);
not (n96,n97);
nand (n98,n96,n92);
nor (n99,n100,n103);
and (n100,n101,n96);
not (n101,n102);
and (n103,n102,n97);
or (n104,n105,n87);
nor (n105,n106,n109);
and (n106,n107,n96);
not (n107,n108);
and (n109,n108,n97);
xor (n110,n111,n166);
xor (n111,n112,n141);
nand (n112,n113,n133);
or (n113,n114,n128);
not (n114,n115);
nor (n115,n116,n123);
nor (n116,n117,n121);
and (n117,n118,n120);
not (n118,n119);
and (n121,n119,n122);
not (n122,n120);
nand (n123,n124,n127);
or (n124,n125,n120);
not (n125,n126);
nand (n127,n125,n120);
nor (n128,n129,n132);
and (n129,n118,n130);
not (n130,n131);
and (n132,n119,n131);
or (n133,n134,n135);
not (n134,n123);
not (n135,n136);
nor (n136,n137,n139);
and (n137,n118,n138);
and (n139,n119,n140);
not (n140,n138);
nand (n141,n142,n159);
or (n142,n143,n153);
not (n143,n144);
nor (n144,n145,n150);
nor (n145,n146,n148);
and (n146,n90,n147);
and (n148,n91,n149);
not (n149,n147);
nand (n150,n151,n152);
or (n151,n118,n147);
nand (n152,n118,n147);
not (n153,n154);
nand (n154,n155,n157);
or (n155,n91,n156);
not (n157,n158);
and (n158,n156,n91);
or (n159,n160,n165);
nor (n160,n161,n164);
and (n161,n162,n90);
not (n162,n163);
and (n164,n163,n91);
not (n165,n150);
xor (n166,n167,n194);
nand (n167,n168,n185);
or (n168,n169,n176);
not (n169,n170);
nand (n170,n171,n175);
or (n171,n172,n174);
not (n172,n173);
nand (n175,n174,n172);
not (n176,n177);
nand (n177,n178,n182);
nand (n178,n179,n180,n181);
not (n181,n174);
nand (n182,n183,n184,n174);
not (n183,n180);
not (n184,n179);
nand (n185,n186,n189);
nand (n186,n187,n188);
or (n187,n183,n179);
nand (n188,n183,n179);
nand (n189,n190,n193);
or (n190,n191,n174);
not (n191,n192);
nand (n193,n174,n191);
nand (n194,n195,n200);
or (n195,n196,n197);
not (n197,n198);
nand (n198,n179,n199);
not (n199,n196);
not (n200,n201);
nor (n201,n202,n204);
and (n202,n184,n203);
and (n204,n179,n205);
not (n205,n203);
or (n206,n207,n430);
and (n207,n208,n350);
xor (n208,n209,n270);
or (n209,n210,n269);
and (n210,n211,n243);
xor (n211,n212,n225);
nand (n212,n213,n220);
or (n213,n214,n219);
not (n214,n215);
nand (n215,n216,n218);
or (n216,n217,n44);
nand (n218,n44,n217);
nand (n219,n48,n33);
nand (n220,n221,n34);
nand (n221,n222,n224);
or (n222,n223,n44);
nand (n224,n44,n223);
nand (n225,n226,n237);
or (n226,n227,n231);
nand (n227,n228,n230);
not (n228,n229);
not (n231,n232);
nand (n232,n233,n235);
or (n233,n234,n230);
not (n235,n236);
and (n236,n234,n230);
nand (n237,n238,n229);
nand (n238,n239,n241);
or (n239,n240,n230);
not (n241,n242);
and (n242,n240,n230);
nand (n243,n244,n263);
or (n244,n245,n253);
not (n245,n246);
nor (n246,n247,n252);
and (n247,n248,n250);
not (n248,n249);
not (n250,n251);
and (n252,n249,n251);
not (n253,n254);
nor (n254,n255,n259);
nand (n255,n256,n258);
or (n256,n44,n257);
nand (n258,n44,n257);
nor (n259,n260,n261);
and (n260,n257,n250);
and (n261,n251,n262);
not (n262,n257);
nand (n263,n255,n264);
nand (n264,n265,n268);
or (n265,n266,n251);
not (n266,n267);
nand (n268,n251,n266);
and (n269,n212,n225);
or (n270,n271,n349);
and (n271,n272,n326);
xor (n272,n273,n300);
nand (n273,n274,n294);
or (n274,n275,n283);
not (n275,n276);
nor (n276,n277,n281);
and (n277,n278,n279);
not (n279,n280);
and (n281,n282,n280);
not (n282,n278);
nand (n283,n284,n290);
not (n284,n285);
nand (n285,n286,n289);
or (n286,n287,n288);
not (n287,n230);
nand (n289,n287,n288);
nand (n290,n291,n293);
or (n291,n292,n280);
not (n292,n288);
nand (n293,n280,n292);
nand (n294,n285,n295);
nand (n295,n296,n298);
or (n296,n297,n280);
not (n298,n299);
and (n299,n297,n280);
nand (n300,n301,n319);
or (n301,n302,n310);
not (n302,n303);
nor (n303,n304,n308);
and (n304,n305,n307);
not (n305,n306);
and (n308,n306,n309);
not (n309,n307);
nand (n310,n311,n316);
nor (n311,n312,n315);
and (n312,n313,n280);
not (n313,n314);
and (n315,n314,n279);
nand (n316,n317,n318);
or (n317,n314,n309);
nand (n318,n309,n314);
nand (n319,n320,n321);
not (n320,n311);
nand (n321,n322,n324);
or (n322,n323,n307);
not (n324,n325);
and (n325,n323,n307);
nand (n326,n327,n338);
or (n327,n328,n333);
not (n328,n329);
nand (n329,n330,n331);
or (n330,n43,n36);
or (n331,n37,n332);
not (n332,n43);
nor (n333,n334,n336);
and (n334,n181,n335);
and (n336,n174,n337);
not (n337,n335);
or (n338,n339,n345);
nand (n339,n340,n333);
or (n340,n341,n343);
not (n341,n342);
nand (n342,n36,n335);
not (n343,n344);
nand (n344,n337,n37);
not (n345,n346);
nand (n346,n347,n348);
or (n347,n37,n55);
nand (n348,n37,n55);
and (n349,n273,n300);
or (n350,n351,n429);
and (n351,n352,n406);
xor (n352,n353,n378);
nand (n353,n354,n373);
or (n354,n355,n363);
not (n355,n356);
nand (n356,n357,n361);
or (n357,n358,n359);
not (n359,n360);
or (n361,n362,n360);
not (n362,n358);
not (n363,n364);
nor (n364,n365,n370);
nor (n365,n366,n369);
and (n366,n360,n367);
not (n367,n368);
nor (n369,n367,n360);
nand (n370,n371,n372);
or (n371,n367,n251);
nand (n372,n367,n251);
nand (n373,n374,n370);
nand (n374,n375,n377);
or (n375,n376,n359);
nand (n377,n376,n359);
nand (n378,n379,n394);
or (n379,n380,n388);
not (n380,n381);
nor (n381,n382,n386);
and (n382,n383,n385);
not (n383,n384);
and (n386,n384,n387);
not (n387,n385);
not (n388,n389);
nand (n389,n390,n393);
or (n390,n391,n307);
not (n391,n392);
nand (n393,n391,n307);
or (n394,n395,n399);
nand (n395,n388,n396);
nand (n396,n397,n398);
or (n397,n392,n387);
nand (n398,n387,n392);
not (n399,n400);
nand (n400,n401,n404);
not (n401,n402);
and (n402,n403,n385);
nand (n404,n387,n405);
not (n405,n403);
nand (n406,n407,n424);
or (n407,n408,n412);
not (n408,n409);
nor (n409,n410,n411);
and (n410,n130,n126);
and (n411,n131,n125);
nand (n412,n413,n420);
or (n413,n414,n417);
not (n414,n415);
nand (n415,n125,n416);
not (n417,n418);
nand (n418,n419,n126);
not (n419,n416);
not (n420,n421);
nand (n421,n422,n423);
or (n422,n387,n416);
nand (n423,n387,n416);
nand (n424,n421,n425);
nand (n425,n426,n427);
or (n426,n126,n138);
not (n427,n428);
and (n428,n138,n126);
and (n429,n353,n378);
and (n430,n209,n270);
and (n431,n29,n110);
or (n432,n433,n615);
and (n433,n434,n580);
xor (n434,n435,n500);
or (n435,n436,n499);
and (n436,n437,n468);
xor (n437,n438,n445);
nand (n438,n439,n444);
or (n439,n114,n440);
not (n440,n441);
nor (n441,n442,n443);
and (n442,n162,n119);
and (n443,n163,n118);
or (n444,n134,n128);
xor (n445,n446,n462);
xor (n446,n447,n455);
nor (n447,n448,n61);
and (n448,n449,n453);
nand (n449,n450,n75);
not (n450,n451);
and (n451,n452,n69);
nand (n453,n454,n72);
not (n454,n452);
nor (n455,n456,n97);
and (n456,n457,n461);
nand (n457,n458,n91);
or (n458,n92,n459);
not (n459,n460);
nand (n461,n92,n459);
nand (n462,n463,n467);
or (n463,n198,n464);
nor (n464,n465,n466);
and (n465,n184,n192);
and (n466,n179,n191);
or (n467,n201,n199);
or (n468,n469,n498);
and (n469,n470,n485);
xor (n470,n471,n479);
nand (n471,n472,n477);
or (n472,n198,n473);
not (n473,n474);
nand (n474,n475,n476);
or (n475,n173,n184);
nand (n476,n184,n173);
nand (n477,n478,n196);
not (n478,n464);
nand (n479,n480,n484);
or (n480,n481,n483);
not (n481,n482);
nand (n482,n88,n460);
nand (n483,n83,n452);
nand (n484,n481,n483);
nand (n485,n486,n492);
nand (n486,n177,n487);
nand (n487,n488,n491);
or (n488,n489,n174);
not (n489,n490);
nand (n491,n174,n489);
nand (n492,n186,n493);
nand (n493,n494,n497);
or (n494,n495,n174);
not (n495,n496);
nand (n497,n174,n495);
and (n498,n471,n479);
and (n499,n438,n445);
or (n500,n501,n579);
and (n501,n502,n568);
xor (n502,n503,n540);
xor (n503,n504,n533);
xor (n504,n505,n511);
nand (n505,n506,n507);
or (n506,n380,n395);
nand (n507,n389,n508);
nor (n508,n509,n510);
and (n509,n305,n385);
and (n510,n306,n387);
nand (n511,n512,n522);
or (n512,n513,n519);
not (n513,n514);
nand (n514,n515,n518);
or (n515,n516,n360);
not (n516,n517);
nand (n518,n516,n360);
nor (n519,n520,n521);
and (n520,n362,n76);
and (n521,n358,n75);
nand (n522,n523,n528);
not (n523,n524);
nor (n524,n525,n526);
and (n525,n75,n81);
and (n526,n76,n527);
not (n527,n81);
not (n528,n529);
nand (n529,n513,n530);
nand (n530,n531,n532);
or (n531,n517,n75);
nand (n532,n75,n517);
nand (n533,n534,n536);
or (n534,n535,n412);
not (n535,n425);
nand (n536,n421,n537);
nor (n537,n538,n539);
and (n538,n405,n126);
and (n539,n403,n125);
xor (n540,n541,n559);
xor (n541,n542,n550);
nand (n542,n543,n545);
or (n543,n544,n253);
not (n544,n264);
nand (n545,n255,n546);
nand (n546,n547,n549);
or (n547,n548,n251);
not (n548,n217);
nand (n549,n251,n548);
nand (n550,n551,n553);
or (n551,n227,n552);
not (n552,n238);
nand (n553,n554,n229);
nand (n554,n555,n557);
or (n555,n556,n230);
not (n557,n558);
and (n558,n556,n230);
nand (n559,n560,n566);
or (n560,n561,n284);
not (n561,n562);
nor (n562,n563,n565);
and (n563,n564,n280);
not (n564,n234);
and (n565,n234,n279);
or (n566,n283,n567);
not (n567,n295);
xor (n568,n569,n578);
xor (n569,n570,n574);
nand (n570,n571,n573);
or (n571,n572,n176);
not (n572,n493);
nand (n573,n170,n186);
nand (n574,n575,n577);
or (n575,n219,n576);
not (n576,n221);
nand (n577,n34,n51);
nor (n578,n483,n482);
and (n579,n503,n540);
xor (n580,n581,n612);
xor (n581,n582,n585);
or (n582,n583,n584);
and (n583,n541,n559);
and (n584,n542,n550);
or (n585,n586,n611);
and (n586,n587,n602);
xor (n587,n588,n595);
nand (n588,n589,n590);
or (n589,n328,n339);
nand (n590,n591,n592);
not (n591,n333);
nand (n592,n593,n594);
or (n593,n489,n37);
nand (n594,n37,n489);
nand (n595,n596,n598);
or (n596,n597,n363);
not (n597,n374);
nand (n598,n599,n370);
nand (n599,n600,n601);
or (n600,n360,n248);
or (n601,n359,n249);
nand (n602,n603,n609);
or (n603,n604,n311);
not (n604,n605);
nand (n605,n606,n608);
not (n606,n607);
and (n607,n278,n307);
nand (n608,n309,n282);
or (n609,n310,n610);
not (n610,n321);
and (n611,n588,n595);
or (n612,n613,n614);
and (n613,n504,n533);
and (n614,n505,n511);
and (n615,n435,n500);
or (n616,n617,n755);
and (n617,n618,n683);
xor (n618,n619,n651);
xor (n619,n620,n648);
xor (n620,n621,n624);
or (n621,n622,n623);
and (n622,n446,n462);
and (n623,n447,n455);
or (n624,n625,n647);
and (n625,n626,n641);
xor (n626,n627,n633);
nand (n627,n628,n629);
or (n628,n73,n58);
or (n629,n65,n630);
nor (n630,n631,n632);
and (n631,n454,n62);
and (n632,n452,n61);
nand (n633,n634,n640);
or (n634,n143,n635);
not (n635,n636);
nand (n636,n637,n639);
not (n637,n638);
and (n638,n108,n91);
nand (n639,n90,n107);
nand (n640,n154,n150);
nand (n641,n642,n646);
or (n642,n86,n643);
nor (n643,n644,n645);
and (n644,n460,n97);
and (n645,n96,n459);
or (n646,n87,n99);
and (n647,n627,n633);
or (n648,n649,n650);
and (n649,n569,n578);
and (n650,n570,n574);
or (n651,n652,n682);
and (n652,n653,n681);
xor (n653,n654,n680);
or (n654,n655,n679);
and (n655,n656,n673);
xor (n656,n657,n665);
nand (n657,n658,n664);
or (n658,n659,n529);
not (n659,n660);
nor (n660,n661,n663);
and (n661,n75,n662);
not (n662,n63);
and (n663,n76,n63);
nand (n664,n523,n514);
nand (n665,n666,n672);
or (n666,n667,n114);
not (n667,n668);
nor (n668,n669,n670);
and (n669,n118,n156);
and (n670,n119,n671);
not (n671,n156);
nand (n672,n441,n123);
nand (n673,n674,n678);
or (n674,n143,n675);
nor (n675,n676,n677);
and (n676,n90,n101);
and (n677,n91,n102);
or (n678,n635,n165);
and (n679,n657,n665);
xor (n680,n626,n641);
xor (n681,n587,n602);
and (n682,n654,n680);
xor (n683,n684,n731);
xor (n684,n685,n710);
xor (n685,n686,n701);
xor (n686,n687,n694);
nand (n687,n688,n690);
or (n688,n689,n395);
not (n689,n508);
nand (n690,n389,n691);
nand (n691,n692,n693);
or (n692,n323,n385);
nand (n693,n385,n323);
nand (n694,n695,n697);
or (n695,n696,n412);
not (n696,n537);
nand (n697,n421,n698);
nor (n698,n699,n700);
and (n699,n383,n126);
and (n700,n384,n125);
nand (n701,n702,n708);
or (n702,n703,n513);
not (n703,n704);
nand (n704,n705,n707);
or (n705,n76,n706);
not (n706,n376);
nand (n707,n706,n76);
nand (n708,n709,n528);
not (n709,n519);
xor (n710,n711,n723);
xor (n711,n712,n715);
nand (n712,n713,n554);
or (n713,n229,n714);
not (n714,n227);
nand (n715,n716,n718);
or (n716,n717,n253);
not (n717,n546);
nand (n718,n255,n719);
nand (n719,n720,n721);
or (n720,n223,n250);
or (n721,n251,n722);
not (n722,n223);
nand (n723,n724,n730);
or (n724,n725,n284);
not (n725,n726);
nor (n726,n727,n728);
and (n727,n240,n279);
and (n728,n729,n280);
not (n729,n240);
or (n730,n283,n561);
xor (n731,n732,n746);
xor (n732,n733,n739);
nand (n733,n734,n735);
or (n734,n604,n310);
nand (n735,n320,n736);
nand (n736,n737,n738);
or (n737,n297,n307);
nand (n738,n307,n297);
nand (n739,n740,n742);
or (n740,n741,n339);
not (n741,n592);
nand (n742,n591,n743);
nand (n743,n744,n745);
or (n744,n495,n37);
nand (n745,n37,n495);
nand (n746,n747,n753);
or (n747,n748,n749);
not (n748,n370);
not (n749,n750);
nand (n750,n751,n752);
or (n751,n360,n266);
or (n752,n359,n267);
or (n753,n363,n754);
not (n754,n599);
and (n755,n619,n651);
or (n756,n757,n1034);
and (n757,n758,n773);
xor (n758,n759,n772);
or (n759,n760,n771);
and (n760,n761,n770);
xor (n761,n762,n763);
xor (n762,n437,n468);
or (n763,n764,n769);
and (n764,n765,n768);
xor (n765,n766,n767);
xor (n766,n656,n673);
xor (n767,n272,n326);
xor (n768,n211,n243);
and (n769,n766,n767);
xor (n770,n502,n568);
and (n771,n762,n763);
xor (n772,n434,n580);
or (n773,n774,n1033);
and (n774,n775,n930);
xor (n775,n776,n777);
xor (n776,n653,n681);
or (n777,n778,n929);
and (n778,n779,n894);
xor (n779,n780,n781);
xor (n780,n352,n406);
or (n781,n782,n893);
and (n782,n783,n857);
xor (n783,n784,n821);
or (n784,n785,n820);
and (n785,n786,n807);
xor (n786,n787,n797);
nand (n787,n788,n793);
or (n788,n789,n176);
not (n789,n790);
nand (n790,n791,n792);
or (n791,n55,n174);
nand (n792,n174,n55);
nand (n793,n794,n186);
nand (n794,n795,n796);
or (n795,n332,n174);
nand (n796,n174,n332);
nand (n797,n798,n803);
or (n798,n799,n219);
not (n799,n800);
nand (n800,n801,n802);
or (n801,n249,n44);
nand (n802,n44,n249);
nand (n803,n804,n34);
nand (n804,n805,n806);
or (n805,n266,n45);
nand (n806,n45,n266);
nand (n807,n808,n814);
or (n808,n228,n809);
not (n809,n810);
nand (n810,n811,n812);
or (n811,n297,n230);
not (n812,n813);
and (n813,n297,n230);
or (n814,n815,n227);
not (n815,n816);
nand (n816,n817,n818);
or (n817,n278,n230);
not (n818,n819);
and (n819,n278,n230);
and (n820,n787,n797);
or (n821,n822,n856);
and (n822,n823,n845);
xor (n823,n824,n835);
nand (n824,n825,n831);
or (n825,n284,n826);
not (n826,n827);
nand (n827,n828,n829);
or (n828,n323,n280);
not (n829,n830);
and (n830,n323,n280);
or (n831,n283,n832);
nor (n832,n833,n834);
and (n833,n279,n305);
and (n834,n280,n306);
nand (n835,n836,n841);
or (n836,n837,n253);
not (n837,n838);
nor (n838,n839,n840);
and (n839,n362,n250);
and (n840,n358,n251);
nand (n841,n255,n842);
nand (n842,n843,n844);
or (n843,n251,n706);
nand (n844,n251,n706);
nand (n845,n846,n852);
or (n846,n847,n311);
not (n847,n848);
nand (n848,n849,n851);
not (n849,n850);
and (n850,n384,n307);
nand (n851,n309,n383);
or (n852,n310,n853);
nor (n853,n854,n855);
and (n854,n309,n405);
and (n855,n307,n403);
and (n856,n824,n835);
or (n857,n858,n892);
and (n858,n859,n880);
xor (n859,n860,n870);
nand (n860,n861,n866);
or (n861,n862,n395);
not (n862,n863);
nor (n863,n864,n865);
and (n864,n130,n385);
and (n865,n131,n387);
nand (n866,n389,n867);
nor (n867,n868,n869);
and (n868,n138,n387);
and (n869,n140,n385);
nand (n870,n871,n876);
or (n871,n872,n363);
not (n872,n873);
nand (n873,n874,n875);
or (n874,n360,n662);
nand (n875,n662,n360);
nand (n876,n877,n370);
nor (n877,n878,n879);
and (n878,n359,n527);
and (n879,n360,n81);
nand (n880,n881,n887);
or (n881,n882,n412);
not (n882,n883);
nand (n883,n884,n885);
or (n884,n126,n156);
not (n885,n886);
and (n886,n156,n126);
nand (n887,n421,n888);
nand (n888,n889,n891);
not (n889,n890);
and (n890,n163,n126);
or (n891,n126,n163);
and (n892,n860,n870);
and (n893,n784,n821);
or (n894,n895,n928);
and (n895,n896,n909);
xor (n896,n897,n903);
nand (n897,n898,n902);
or (n898,n114,n899);
nor (n899,n900,n901);
and (n900,n118,n107);
and (n901,n119,n108);
or (n902,n134,n667);
nand (n903,n904,n908);
or (n904,n143,n905);
nor (n905,n906,n907);
and (n906,n459,n90);
and (n907,n460,n91);
or (n908,n675,n165);
xor (n909,n910,n922);
xor (n910,n911,n917);
nor (n911,n912,n75);
and (n912,n913,n916);
nand (n913,n914,n359);
not (n914,n915);
and (n915,n452,n517);
nand (n916,n454,n516);
nor (n917,n918,n91);
nor (n918,n919,n921);
nor (n919,n920,n118);
and (n920,n460,n149);
nor (n921,n460,n149);
nand (n922,n923,n927);
or (n923,n198,n924);
nor (n924,n925,n926);
and (n925,n496,n184);
and (n926,n495,n179);
or (n927,n473,n199);
and (n928,n897,n903);
and (n929,n780,n781);
or (n930,n931,n1032);
and (n931,n932,n1006);
xor (n932,n933,n972);
xor (n933,n934,n971);
xor (n934,n935,n953);
or (n935,n936,n952);
and (n936,n937,n948);
xor (n937,n938,n941);
nand (n938,n939,n940);
nand (n939,n848,n311,n316);
nand (n940,n320,n303);
nand (n941,n942,n947);
or (n942,n943,n339);
not (n943,n944);
nand (n944,n945,n946);
or (n945,n722,n37);
nand (n946,n37,n722);
nand (n947,n591,n346);
nand (n948,n949,n951);
or (n949,n950,n363);
not (n950,n877);
nand (n951,n370,n356);
and (n952,n938,n941);
or (n953,n954,n970);
and (n954,n955,n964);
xor (n955,n956,n960);
nand (n956,n957,n959);
or (n957,n958,n395);
not (n958,n867);
nand (n959,n400,n389);
nand (n960,n961,n963);
or (n961,n962,n412);
not (n962,n888);
nand (n963,n421,n409);
nand (n964,n965,n969);
or (n965,n529,n966);
nor (n966,n967,n968);
and (n967,n454,n76);
and (n968,n452,n75);
nand (n969,n660,n514);
and (n970,n956,n960);
xor (n971,n470,n485);
xor (n972,n973,n992);
xor (n973,n974,n977);
or (n974,n975,n976);
and (n975,n910,n922);
and (n976,n911,n917);
or (n977,n978,n991);
and (n978,n979,n988);
xor (n979,n980,n984);
nand (n980,n981,n983);
or (n981,n982,n176);
not (n982,n794);
nand (n983,n186,n487);
nand (n984,n985,n987);
or (n985,n986,n219);
not (n986,n804);
nand (n987,n34,n215);
nor (n988,n989,n990);
nand (n989,n452,n514);
nand (n990,n150,n460);
and (n991,n980,n984);
or (n992,n993,n1005);
and (n993,n994,n1002);
xor (n994,n995,n998);
nand (n995,n996,n997);
or (n996,n227,n809);
nand (n997,n232,n229);
nand (n998,n999,n1001);
or (n999,n1000,n253);
not (n1000,n842);
nand (n1001,n255,n246);
nand (n1002,n1003,n1004);
or (n1003,n275,n284);
or (n1004,n283,n826);
and (n1005,n995,n998);
or (n1006,n1007,n1031);
and (n1007,n1008,n1030);
xor (n1008,n1009,n1029);
or (n1009,n1010,n1028);
and (n1010,n1011,n1022);
xor (n1011,n1012,n1016);
nand (n1012,n1013,n1015);
or (n1013,n1014,n989);
not (n1014,n990);
nand (n1015,n1014,n989);
nand (n1016,n1017,n1021);
or (n1017,n114,n1018);
nor (n1018,n1019,n1020);
and (n1019,n118,n101);
and (n1020,n119,n102);
or (n1021,n134,n899);
nand (n1022,n1023,n1027);
or (n1023,n198,n1024);
nor (n1024,n1025,n1026);
and (n1025,n184,n490);
and (n1026,n179,n489);
or (n1027,n924,n199);
and (n1028,n1012,n1016);
xor (n1029,n979,n988);
xor (n1030,n955,n964);
and (n1031,n1009,n1029);
and (n1032,n933,n972);
and (n1033,n776,n777);
and (n1034,n759,n772);
xor (n1035,n1036,n1184);
xor (n1036,n1037,n1080);
xor (n1037,n1038,n1051);
xor (n1038,n1039,n1042);
or (n1039,n1040,n1041);
and (n1040,n620,n648);
and (n1041,n621,n624);
xor (n1042,n1043,n1048);
xor (n1043,n1044,n1045);
and (n1044,n167,n194);
or (n1045,n1046,n1047);
and (n1046,n30,n84);
and (n1047,n31,n56);
or (n1048,n1049,n1050);
and (n1049,n711,n723);
and (n1050,n712,n715);
xor (n1051,n1052,n1059);
xor (n1052,n1053,n1056);
or (n1053,n1054,n1055);
and (n1054,n732,n746);
and (n1055,n733,n739);
or (n1056,n1057,n1058);
and (n1057,n686,n701);
and (n1058,n687,n694);
xor (n1059,n1060,n1074);
xor (n1060,n1061,n1067);
nand (n1061,n1062,n1063);
or (n1062,n725,n283);
nand (n1063,n285,n1064);
nand (n1064,n1065,n1066);
or (n1065,n556,n280);
nand (n1066,n280,n556);
nand (n1067,n1068,n1070);
or (n1068,n1069,n310);
not (n1069,n736);
nand (n1070,n320,n1071);
nand (n1071,n1072,n1073);
or (n1072,n234,n307);
nand (n1073,n307,n234);
nand (n1074,n1075,n1076);
or (n1075,n749,n363);
nand (n1076,n1077,n370);
nor (n1077,n1078,n1079);
and (n1078,n548,n359);
and (n1079,n217,n360);
xor (n1080,n1081,n1150);
xor (n1081,n1082,n1085);
or (n1082,n1083,n1084);
and (n1083,n684,n731);
and (n1084,n685,n710);
xor (n1085,n1086,n1128);
xor (n1086,n1087,n1110);
xor (n1087,n1088,n1102);
xor (n1088,n1089,n1095);
nand (n1089,n1090,n1091);
or (n1090,n40,n219);
nand (n1091,n34,n1092);
nand (n1092,n1093,n1094);
or (n1093,n489,n45);
nand (n1094,n45,n489);
nand (n1095,n1096,n1097);
or (n1096,n105,n86);
nand (n1097,n1098,n88);
not (n1098,n1099);
nor (n1099,n1100,n1101);
and (n1100,n671,n96);
and (n1101,n156,n97);
nand (n1102,n1103,n1108);
or (n1103,n73,n1104);
not (n1104,n1105);
nor (n1105,n1106,n1107);
and (n1106,n61,n362);
and (n1107,n358,n62);
nand (n1108,n1109,n79);
not (n1109,n65);
nand (n1110,n1111,n1127);
or (n1111,n1112,n1119);
nor (n1112,n1113,n1115);
and (n1113,n1114,n743);
not (n1114,n339);
and (n1115,n591,n1116);
nand (n1116,n1117,n1118);
or (n1117,n172,n37);
nand (n1118,n37,n172);
not (n1119,n1120);
nand (n1120,n1121,n1123);
or (n1121,n1122,n253);
not (n1122,n719);
nand (n1123,n255,n1124);
nand (n1124,n1125,n1126);
or (n1125,n55,n251);
nand (n1126,n251,n55);
nand (n1127,n1119,n1112);
xor (n1128,n1129,n1142);
xor (n1129,n1130,n1136);
nand (n1130,n1131,n1132);
or (n1131,n703,n529);
nand (n1132,n514,n1133);
nand (n1133,n1134,n1135);
or (n1134,n76,n248);
nand (n1135,n76,n248);
nand (n1136,n1137,n1138);
or (n1137,n135,n114);
nand (n1138,n1139,n123);
nand (n1139,n1140,n1141);
or (n1140,n119,n403);
nand (n1141,n403,n119);
nand (n1142,n1143,n1144);
or (n1143,n143,n160);
or (n1144,n1145,n165);
not (n1145,n1146);
nand (n1146,n1147,n1149);
not (n1147,n1148);
and (n1148,n131,n91);
nand (n1149,n90,n130);
xor (n1150,n1151,n1181);
xor (n1151,n1152,n1178);
xor (n1152,n1153,n1169);
xor (n1153,n1154,n1162);
nand (n1154,n1155,n1157);
or (n1155,n1156,n395);
not (n1156,n691);
nand (n1157,n1158,n389);
nand (n1158,n1159,n1161);
not (n1159,n1160);
and (n1160,n278,n385);
nand (n1161,n387,n282);
nand (n1162,n1163,n1165);
or (n1163,n1164,n412);
not (n1164,n698);
nand (n1165,n421,n1166);
nor (n1166,n1167,n1168);
and (n1167,n305,n126);
and (n1168,n306,n125);
nand (n1169,n1170,n1172);
or (n1170,n176,n1171);
not (n1171,n189);
or (n1172,n1173,n1174);
not (n1173,n186);
not (n1174,n1175);
nand (n1175,n1176,n1177);
or (n1176,n203,n181);
nand (n1177,n181,n203);
or (n1178,n1179,n1180);
and (n1179,n111,n166);
and (n1180,n112,n141);
or (n1181,n1182,n1183);
and (n1182,n581,n612);
and (n1183,n582,n585);
or (n1184,n1185,n1200);
and (n1185,n1186,n1199);
xor (n1186,n1187,n1188);
xor (n1187,n28,n206);
or (n1188,n1189,n1198);
and (n1189,n1190,n1197);
xor (n1190,n1191,n1194);
or (n1191,n1192,n1193);
and (n1192,n973,n992);
and (n1193,n974,n977);
or (n1194,n1195,n1196);
and (n1195,n934,n971);
and (n1196,n935,n953);
xor (n1197,n208,n350);
and (n1198,n1191,n1194);
xor (n1199,n618,n683);
and (n1200,n1187,n1188);
or (n1201,n1202,n1213);
and (n1202,n1203,n1206);
xor (n1203,n1204,n1205);
xor (n1204,n1186,n1199);
xor (n1205,n758,n773);
or (n1206,n1207,n1212);
and (n1207,n1208,n1211);
xor (n1208,n1209,n1210);
xor (n1209,n761,n770);
xor (n1210,n1190,n1197);
xor (n1211,n775,n930);
and (n1212,n1209,n1210);
and (n1213,n1204,n1205);
not (n1214,n1215);
nand (n1215,n1216,n1217);
xor (n1216,n1203,n1206);
or (n1217,n1218,n1393);
and (n1218,n1219,n1392);
xor (n1219,n1220,n1373);
or (n1220,n1221,n1372);
and (n1221,n1222,n1231);
xor (n1222,n1223,n1224);
xor (n1223,n765,n768);
or (n1224,n1225,n1230);
and (n1225,n1226,n1229);
xor (n1226,n1227,n1228);
xor (n1227,n994,n1002);
xor (n1228,n937,n948);
xor (n1229,n896,n909);
and (n1230,n1227,n1228);
or (n1231,n1232,n1371);
and (n1232,n1233,n1370);
xor (n1233,n1234,n1299);
or (n1234,n1235,n1298);
and (n1235,n1236,n1272);
xor (n1236,n1237,n1244);
nand (n1237,n1238,n1243);
or (n1238,n339,n1239);
not (n1239,n1240);
nor (n1240,n1241,n1242);
and (n1241,n548,n36);
and (n1242,n217,n37);
or (n1243,n333,n943);
or (n1244,n1245,n1271);
and (n1245,n1246,n1262);
xor (n1246,n1247,n1254);
nand (n1247,n1248,n1253);
or (n1248,n1249,n219);
not (n1249,n1250);
nand (n1250,n1251,n1252);
or (n1251,n376,n44);
nand (n1252,n44,n376);
nand (n1253,n34,n800);
nand (n1254,n1255,n1261);
or (n1255,n227,n1256);
not (n1256,n1257);
nor (n1257,n1258,n1260);
and (n1258,n1259,n230);
not (n1259,n323);
and (n1260,n323,n287);
nand (n1261,n816,n229);
nand (n1262,n1263,n1269);
or (n1263,n283,n1264);
not (n1264,n1265);
nand (n1265,n1266,n1267);
or (n1266,n384,n280);
not (n1267,n1268);
and (n1268,n384,n280);
nand (n1269,n1270,n285);
not (n1270,n832);
and (n1271,n1247,n1254);
or (n1272,n1273,n1297);
and (n1273,n1274,n1289);
xor (n1274,n1275,n1282);
nand (n1275,n1276,n1281);
or (n1276,n1277,n253);
not (n1277,n1278);
nor (n1278,n1279,n1280);
and (n1279,n527,n250);
and (n1280,n81,n251);
nand (n1281,n255,n838);
nand (n1282,n1283,n1288);
or (n1283,n1284,n310);
not (n1284,n1285);
nor (n1285,n1286,n1287);
and (n1286,n140,n307);
and (n1287,n138,n309);
or (n1288,n311,n853);
nand (n1289,n1290,n1296);
or (n1290,n395,n1291);
not (n1291,n1292);
nand (n1292,n1293,n1295);
not (n1293,n1294);
and (n1294,n163,n385);
nand (n1295,n387,n162);
or (n1296,n388,n862);
and (n1297,n1275,n1282);
and (n1298,n1237,n1244);
or (n1299,n1300,n1369);
and (n1300,n1301,n1348);
xor (n1301,n1302,n1329);
or (n1302,n1303,n1328);
and (n1303,n1304,n1320);
xor (n1304,n1305,n1312);
nand (n1305,n1306,n1311);
or (n1306,n1307,n363);
not (n1307,n1308);
nor (n1308,n1309,n1310);
and (n1309,n359,n454);
and (n1310,n452,n360);
nand (n1311,n873,n370);
nand (n1312,n1313,n1319);
or (n1313,n1314,n412);
not (n1314,n1315);
nand (n1315,n1316,n1317);
or (n1316,n126,n108);
not (n1317,n1318);
and (n1318,n108,n126);
nand (n1319,n883,n421);
nand (n1320,n1321,n1327);
or (n1321,n1322,n114);
not (n1322,n1323);
nand (n1323,n1324,n1325);
or (n1324,n460,n119);
not (n1325,n1326);
and (n1326,n460,n119);
or (n1327,n1018,n134);
and (n1328,n1305,n1312);
or (n1329,n1330,n1347);
and (n1330,n1331,n1344);
xor (n1331,n1332,n1338);
nand (n1332,n1333,n1337);
or (n1333,n198,n1334);
nor (n1334,n1335,n1336);
and (n1335,n184,n43);
and (n1336,n179,n332);
or (n1337,n1024,n199);
nand (n1338,n1339,n1343);
or (n1339,n339,n1340);
nor (n1340,n1341,n1342);
and (n1341,n266,n37);
and (n1342,n267,n36);
nand (n1343,n1240,n591);
and (n1344,n1345,n1346);
and (n1345,n123,n460);
and (n1346,n370,n452);
and (n1347,n1332,n1338);
or (n1348,n1349,n1368);
and (n1349,n1350,n1361);
xor (n1350,n1351,n1356);
nor (n1351,n1352,n359);
nor (n1352,n1353,n1354);
and (n1353,n454,n367);
and (n1354,n1355,n250);
nand (n1355,n452,n368);
and (n1356,n1357,n118);
nand (n1357,n1358,n1360);
nand (n1358,n1359,n126);
or (n1359,n120,n459);
nand (n1360,n459,n120);
nand (n1361,n1362,n1367);
or (n1362,n1363,n176);
not (n1363,n1364);
nor (n1364,n1365,n1366);
and (n1365,n722,n181);
and (n1366,n223,n174);
nand (n1367,n186,n790);
and (n1368,n1351,n1356);
and (n1369,n1302,n1329);
xor (n1370,n783,n857);
and (n1371,n1234,n1299);
and (n1372,n1223,n1224);
or (n1373,n1374,n1391);
and (n1374,n1375,n1378);
xor (n1375,n1376,n1377);
xor (n1376,n779,n894);
xor (n1377,n932,n1006);
or (n1378,n1379,n1390);
and (n1379,n1380,n1389);
xor (n1380,n1381,n1388);
or (n1381,n1382,n1387);
and (n1382,n1383,n1386);
xor (n1383,n1384,n1385);
xor (n1384,n859,n880);
xor (n1385,n1011,n1022);
xor (n1386,n786,n807);
and (n1387,n1384,n1385);
xor (n1388,n1008,n1030);
xor (n1389,n1226,n1229);
and (n1390,n1381,n1388);
and (n1391,n1376,n1377);
xor (n1392,n1208,n1211);
and (n1393,n1220,n1373);
and (n1394,n22,n1201);
not (n1395,n1396);
nor (n1396,n1397,n1700);
nor (n1397,n1398,n1689);
xor (n1398,n1399,n1680);
xor (n1399,n1400,n1490);
or (n1400,n1401,n1489);
and (n1401,n1402,n1473);
xor (n1402,n1403,n1470);
xor (n1403,n1404,n1450);
xor (n1404,n1405,n1425);
xor (n1405,n1406,n1416);
xor (n1406,n1407,n1409);
nand (n1407,n1408,n1175);
or (n1408,n186,n177);
nand (n1409,n1410,n1412);
or (n1410,n1411,n529);
not (n1411,n1133);
nand (n1412,n1413,n514);
nand (n1413,n1414,n1415);
or (n1414,n267,n75);
or (n1415,n266,n76);
nand (n1416,n1417,n1419);
or (n1417,n114,n1418);
not (n1418,n1139);
or (n1419,n134,n1420);
not (n1420,n1421);
nand (n1421,n1422,n1424);
not (n1422,n1423);
and (n1423,n384,n119);
nand (n1424,n118,n383);
xor (n1425,n1426,n1442);
xor (n1426,n1427,n1434);
nand (n1427,n1428,n1430);
or (n1428,n1429,n363);
not (n1429,n1077);
nand (n1430,n1431,n370);
nor (n1431,n1432,n1433);
and (n1432,n722,n359);
and (n1433,n223,n360);
nand (n1434,n1435,n1437);
or (n1435,n1436,n395);
not (n1436,n1158);
nand (n1437,n389,n1438);
nor (n1438,n1439,n1441);
and (n1439,n1440,n385);
not (n1440,n297);
and (n1441,n297,n387);
nand (n1442,n1443,n1445);
or (n1443,n412,n1444);
not (n1444,n1166);
or (n1445,n420,n1446);
not (n1446,n1447);
nor (n1447,n1448,n1449);
and (n1448,n1259,n126);
and (n1449,n323,n125);
xor (n1450,n1451,n1467);
xor (n1451,n1452,n1458);
nand (n1452,n1453,n1454);
or (n1453,n1104,n65);
or (n1454,n1455,n73);
or (n1455,n1456,n1457);
and (n1456,n706,n61);
and (n1457,n376,n62);
not (n1458,n1459);
nand (n1459,n1460,n1462);
or (n1460,n339,n1461);
not (n1461,n1116);
or (n1462,n333,n1463);
not (n1463,n1464);
nand (n1464,n1465,n1466);
or (n1465,n192,n36);
nand (n1466,n36,n192);
or (n1467,n1468,n1469);
and (n1468,n1129,n1142);
and (n1469,n1130,n1136);
or (n1470,n1471,n1472);
and (n1471,n1038,n1051);
and (n1472,n1039,n1042);
xor (n1473,n1474,n1486);
xor (n1474,n1475,n1478);
or (n1475,n1476,n1477);
and (n1476,n1043,n1048);
and (n1477,n1044,n1045);
xor (n1478,n1479,n1483);
xor (n1479,n1127,n1480);
or (n1480,n1481,n1482);
and (n1481,n1060,n1074);
and (n1482,n1061,n1067);
or (n1483,n1484,n1485);
and (n1484,n1153,n1169);
and (n1485,n1154,n1162);
or (n1486,n1487,n1488);
and (n1487,n1052,n1059);
and (n1488,n1053,n1056);
and (n1489,n1403,n1470);
xor (n1490,n1491,n1656);
xor (n1491,n1492,n1645);
xor (n1492,n1493,n1576);
xor (n1493,n1494,n1547);
xor (n1494,n1495,n1520);
xor (n1495,n1496,n1517);
or (n1496,n1497,n1516);
and (n1497,n1498,n1509);
xor (n1498,n1499,n1506);
nand (n1499,n1500,n1502);
or (n1500,n1501,n253);
not (n1501,n1124);
nand (n1502,n255,n1503);
nand (n1503,n1504,n1505);
or (n1504,n332,n251);
nand (n1505,n251,n332);
nand (n1506,n1507,n1064);
or (n1507,n285,n1508);
not (n1508,n283);
nand (n1509,n1510,n1512);
or (n1510,n310,n1511);
not (n1511,n1071);
or (n1512,n311,n1513);
nor (n1513,n1514,n1515);
and (n1514,n240,n307);
and (n1515,n729,n309);
and (n1516,n1499,n1506);
or (n1517,n1518,n1519);
and (n1518,n1426,n1442);
and (n1519,n1427,n1434);
xor (n1520,n1521,n1539);
xor (n1521,n1522,n1528);
nand (n1522,n1523,n1524);
or (n1523,n1455,n65);
nand (n1524,n1525,n83);
nand (n1525,n1526,n1527);
or (n1526,n249,n61);
nand (n1527,n249,n61);
nand (n1528,n1529,n1535);
or (n1529,n1530,n86);
not (n1530,n1531);
nand (n1531,n1532,n1533);
or (n1532,n97,n163);
not (n1533,n1534);
and (n1534,n163,n97);
or (n1535,n1536,n87);
nor (n1536,n1537,n1538);
and (n1537,n96,n130);
and (n1538,n131,n97);
nand (n1539,n1540,n1546);
or (n1540,n1541,n311);
not (n1541,n1542);
nor (n1542,n1543,n1545);
and (n1543,n1544,n307);
not (n1544,n556);
and (n1545,n556,n309);
or (n1546,n310,n1513);
or (n1547,n1548,n1575);
and (n1548,n1549,n1574);
xor (n1549,n1550,n1553);
or (n1550,n1551,n1552);
and (n1551,n1088,n1102);
and (n1552,n1089,n1095);
xor (n1553,n1554,n1570);
xor (n1554,n1555,n1563);
nand (n1555,n1556,n1562);
or (n1556,n165,n1557);
not (n1557,n1558);
nand (n1558,n1559,n1561);
not (n1559,n1560);
and (n1560,n138,n91);
or (n1561,n91,n138);
nand (n1562,n144,n1146);
nand (n1563,n1564,n1566);
or (n1564,n1565,n219);
not (n1565,n1092);
nand (n1566,n34,n1567);
nand (n1567,n1568,n1569);
or (n1568,n495,n45);
nand (n1569,n45,n495);
nand (n1570,n1571,n1572);
or (n1571,n1530,n87);
nand (n1572,n1098,n1573);
not (n1573,n86);
xor (n1574,n1498,n1509);
and (n1575,n1550,n1553);
xor (n1576,n1577,n1622);
xor (n1577,n1578,n1600);
xor (n1578,n1579,n1593);
xor (n1579,n1580,n1586);
nand (n1580,n1581,n1582);
or (n1581,n1463,n339);
nand (n1582,n1583,n591);
nand (n1583,n1584,n1585);
or (n1584,n203,n36);
nand (n1585,n36,n203);
nand (n1586,n1587,n1589);
or (n1587,n1588,n219);
not (n1588,n1567);
nand (n1589,n34,n1590);
nand (n1590,n1591,n1592);
or (n1591,n172,n45);
nand (n1592,n45,n172);
nand (n1593,n1594,n1596);
or (n1594,n1595,n363);
not (n1595,n1431);
nand (n1596,n1597,n370);
nand (n1597,n1598,n1599);
or (n1598,n55,n360);
nand (n1599,n55,n360);
xor (n1600,n1601,n1615);
xor (n1601,n1602,n1609);
nand (n1602,n1603,n1604);
or (n1603,n1420,n114);
nand (n1604,n1605,n123);
nand (n1605,n1606,n1608);
not (n1606,n1607);
and (n1607,n306,n119);
nand (n1608,n118,n305);
nand (n1609,n1610,n1611);
or (n1610,n1557,n143);
nand (n1611,n1612,n150);
nand (n1612,n1613,n1614);
or (n1613,n403,n91);
nand (n1614,n91,n403);
nand (n1615,n1616,n1618);
or (n1616,n1617,n253);
not (n1617,n1503);
nand (n1618,n255,n1619);
nor (n1619,n1620,n1621);
and (n1620,n489,n250);
and (n1621,n490,n251);
xor (n1622,n1623,n1637);
xor (n1623,n1624,n1631);
nand (n1624,n1625,n1627);
or (n1625,n1626,n395);
not (n1626,n1438);
nand (n1627,n389,n1628);
nand (n1628,n1629,n1630);
or (n1629,n234,n385);
nand (n1630,n385,n234);
nand (n1631,n1632,n1633);
or (n1632,n1446,n412);
nand (n1633,n421,n1634);
nor (n1634,n1635,n1636);
and (n1635,n282,n126);
and (n1636,n278,n125);
nand (n1637,n1638,n1643);
or (n1638,n1639,n513);
not (n1639,n1640);
nand (n1640,n1641,n1642);
or (n1641,n217,n75);
nand (n1642,n75,n217);
or (n1643,n529,n1644);
not (n1644,n1413);
or (n1645,n1646,n1655);
and (n1646,n1647,n1652);
xor (n1647,n1648,n1651);
or (n1648,n1649,n1650);
and (n1649,n1086,n1128);
and (n1650,n1087,n1110);
xor (n1651,n1549,n1574);
or (n1652,n1653,n1654);
and (n1653,n1151,n1181);
and (n1654,n1152,n1178);
and (n1655,n1648,n1651);
xor (n1656,n1657,n1664);
xor (n1657,n1658,n1661);
or (n1658,n1659,n1660);
and (n1659,n1404,n1450);
and (n1660,n1405,n1425);
or (n1661,n1662,n1663);
and (n1662,n1474,n1486);
and (n1663,n1475,n1478);
xor (n1664,n1665,n1672);
xor (n1665,n1666,n1669);
or (n1666,n1667,n1668);
and (n1667,n1451,n1467);
and (n1668,n1452,n1458);
or (n1669,n1670,n1671);
and (n1670,n1479,n1483);
and (n1671,n1127,n1480);
xor (n1672,n1673,n1677);
xor (n1673,n1459,n1674);
or (n1674,n1675,n1676);
and (n1675,n1406,n1416);
and (n1676,n1407,n1409);
or (n1677,n1678,n1679);
and (n1678,n1554,n1570);
and (n1679,n1555,n1563);
or (n1680,n1681,n1688);
and (n1681,n1682,n1687);
xor (n1682,n1683,n1684);
xor (n1683,n1647,n1652);
or (n1684,n1685,n1686);
and (n1685,n1081,n1150);
and (n1686,n1082,n1085);
xor (n1687,n1402,n1473);
and (n1688,n1683,n1684);
or (n1689,n1690,n1699);
and (n1690,n1691,n1696);
xor (n1691,n1692,n1695);
or (n1692,n1693,n1694);
and (n1693,n25,n616);
and (n1694,n26,n432);
xor (n1695,n1682,n1687);
or (n1696,n1697,n1698);
and (n1697,n1036,n1184);
and (n1698,n1037,n1080);
and (n1699,n1692,n1695);
nor (n1700,n1701,n1702);
xor (n1701,n1691,n1696);
or (n1702,n1703,n1704);
and (n1703,n23,n1035);
and (n1704,n24,n756);
or (n1705,n1706,n1397);
not (n1706,n1707);
nand (n1707,n1708,n1711);
or (n1708,n1709,n1710);
not (n1709,n1398);
not (n1710,n1689);
nand (n1711,n1701,n1702);
and (n1712,n1713,n1971);
nor (n1713,n1714,n1852);
and (n1714,n1715,n1848);
not (n1715,n1716);
xor (n1716,n1717,n1845);
xor (n1717,n1718,n1818);
xor (n1718,n1719,n1815);
xor (n1719,n1720,n1765);
xor (n1720,n1721,n1744);
xor (n1721,n1722,n1725);
or (n1722,n1723,n1724);
and (n1723,n1623,n1637);
and (n1724,n1624,n1631);
xor (n1725,n1726,n1736);
xor (n1726,n1727,n1729);
nand (n1727,n1728,n1583);
or (n1728,n591,n1114);
nand (n1729,n1730,n1732);
or (n1730,n1731,n253);
not (n1731,n1619);
nand (n1732,n255,n1733);
nor (n1733,n1734,n1735);
and (n1734,n495,n250);
and (n1735,n496,n251);
nand (n1736,n1737,n1742);
or (n1737,n1738,n87);
not (n1738,n1739);
nor (n1739,n1740,n1741);
and (n1740,n138,n96);
and (n1741,n140,n97);
nand (n1742,n1743,n1573);
not (n1743,n1536);
xor (n1744,n1745,n1758);
xor (n1745,n1746,n1753);
nand (n1746,n1747,n1749);
or (n1747,n1748,n363);
not (n1748,n1597);
nand (n1749,n1750,n370);
nand (n1750,n1751,n1752);
or (n1751,n43,n359);
nand (n1752,n359,n43);
nand (n1753,n1754,n1756);
or (n1754,n1755,n395);
not (n1755,n1628);
nand (n1756,n389,n1757);
xor (n1757,n729,n385);
nand (n1758,n1759,n1761);
or (n1759,n412,n1760);
not (n1760,n1634);
or (n1761,n420,n1762);
nor (n1762,n1763,n1764);
and (n1763,n125,n1440);
and (n1764,n297,n126);
xor (n1765,n1766,n1812);
xor (n1766,n1767,n1790);
xor (n1767,n1768,n1782);
xor (n1768,n1769,n1775);
nand (n1769,n1770,n1771);
or (n1770,n1639,n529);
nand (n1771,n1772,n514);
nor (n1772,n1773,n1774);
and (n1773,n722,n75);
and (n1774,n223,n76);
nand (n1775,n1776,n1778);
or (n1776,n1777,n114);
not (n1777,n1605);
nand (n1778,n123,n1779);
nand (n1779,n1780,n1781);
or (n1780,n119,n323);
nand (n1781,n119,n323);
nand (n1782,n1783,n1788);
or (n1783,n165,n1784);
not (n1784,n1785);
nor (n1785,n1786,n1787);
and (n1786,n383,n91);
and (n1787,n384,n90);
or (n1788,n143,n1789);
not (n1789,n1612);
xor (n1790,n1791,n1803);
xor (n1791,n1792,n1800);
nand (n1792,n1793,n1798);
or (n1793,n73,n1794);
not (n1794,n1795);
nor (n1795,n1796,n1797);
and (n1796,n61,n266);
and (n1797,n267,n62);
or (n1798,n65,n1799);
not (n1799,n1525);
nand (n1800,n1801,n1542);
or (n1801,n320,n1802);
not (n1802,n310);
not (n1803,n1804);
nand (n1804,n1805,n1807);
or (n1805,n219,n1806);
not (n1806,n1590);
or (n1807,n33,n1808);
not (n1808,n1809);
nor (n1809,n1810,n1811);
and (n1810,n191,n44);
and (n1811,n192,n45);
or (n1812,n1813,n1814);
and (n1813,n1673,n1677);
and (n1814,n1459,n1674);
or (n1815,n1816,n1817);
and (n1816,n1665,n1672);
and (n1817,n1666,n1669);
xor (n1818,n1819,n1842);
xor (n1819,n1820,n1839);
xor (n1820,n1821,n1828);
xor (n1821,n1822,n1825);
or (n1822,n1823,n1824);
and (n1823,n1577,n1622);
and (n1824,n1578,n1600);
or (n1825,n1826,n1827);
and (n1826,n1495,n1520);
and (n1827,n1496,n1517);
xor (n1828,n1829,n1836);
xor (n1829,n1830,n1833);
or (n1830,n1831,n1832);
and (n1831,n1601,n1615);
and (n1832,n1602,n1609);
or (n1833,n1834,n1835);
and (n1834,n1521,n1539);
and (n1835,n1522,n1528);
or (n1836,n1837,n1838);
and (n1837,n1579,n1593);
and (n1838,n1580,n1586);
or (n1839,n1840,n1841);
and (n1840,n1493,n1576);
and (n1841,n1494,n1547);
or (n1842,n1843,n1844);
and (n1843,n1657,n1664);
and (n1844,n1658,n1661);
or (n1845,n1846,n1847);
and (n1846,n1491,n1656);
and (n1847,n1492,n1645);
not (n1848,n1849);
or (n1849,n1850,n1851);
and (n1850,n1399,n1680);
and (n1851,n1400,n1490);
nor (n1852,n1853,n1856);
or (n1853,n1854,n1855);
and (n1854,n1717,n1845);
and (n1855,n1718,n1818);
xor (n1856,n1857,n1968);
xor (n1857,n1858,n1861);
or (n1858,n1859,n1860);
and (n1859,n1719,n1815);
and (n1860,n1720,n1765);
xor (n1861,n1862,n1885);
xor (n1862,n1863,n1882);
xor (n1863,n1864,n1879);
xor (n1864,n1865,n1868);
or (n1865,n1866,n1867);
and (n1866,n1829,n1836);
and (n1867,n1830,n1833);
xor (n1868,n1869,n1876);
xor (n1869,n1870,n1804);
nand (n1870,n1871,n1872);
or (n1871,n412,n1762);
or (n1872,n420,n1873);
nor (n1873,n1874,n1875);
and (n1874,n125,n564);
and (n1875,n234,n126);
or (n1876,n1877,n1878);
and (n1877,n1745,n1758);
and (n1878,n1746,n1753);
or (n1879,n1880,n1881);
and (n1880,n1721,n1744);
and (n1881,n1722,n1725);
or (n1882,n1883,n1884);
and (n1883,n1821,n1828);
and (n1884,n1822,n1825);
xor (n1885,n1886,n1965);
xor (n1886,n1887,n1916);
xor (n1887,n1888,n1895);
xor (n1888,n1889,n1892);
or (n1889,n1890,n1891);
and (n1890,n1768,n1782);
and (n1891,n1769,n1775);
or (n1892,n1893,n1894);
and (n1893,n1726,n1736);
and (n1894,n1727,n1729);
xor (n1895,n1896,n1910);
xor (n1896,n1897,n1904);
nand (n1897,n1898,n1900);
or (n1898,n1899,n114);
not (n1899,n1779);
nand (n1900,n1901,n123);
nand (n1901,n1902,n1903);
or (n1902,n278,n119);
nand (n1903,n119,n278);
nand (n1904,n1905,n1906);
or (n1905,n1784,n143);
nand (n1906,n1907,n150);
nor (n1907,n1908,n1909);
and (n1908,n305,n91);
and (n1909,n306,n90);
nand (n1910,n1911,n1912);
or (n1911,n1794,n65);
or (n1912,n1913,n73);
nor (n1913,n1914,n1915);
and (n1914,n61,n217);
and (n1915,n62,n548);
xor (n1916,n1917,n1962);
xor (n1917,n1918,n1940);
xor (n1918,n1919,n1933);
xor (n1919,n1920,n1926);
nand (n1920,n1921,n1922);
or (n1921,n1738,n86);
nand (n1922,n1923,n88);
nor (n1923,n1924,n1925);
and (n1924,n96,n403);
and (n1925,n97,n405);
nand (n1926,n1927,n1929);
or (n1927,n1928,n363);
not (n1928,n1750);
nand (n1929,n1930,n370);
nor (n1930,n1931,n1932);
and (n1931,n489,n359);
and (n1932,n490,n360);
nand (n1933,n1934,n1936);
or (n1934,n1935,n395);
not (n1935,n1757);
nand (n1936,n389,n1937);
nor (n1937,n1938,n1939);
and (n1938,n1544,n385);
and (n1939,n556,n387);
xor (n1940,n1941,n1955);
xor (n1941,n1942,n1948);
nand (n1942,n1943,n1944);
or (n1943,n1808,n219);
nand (n1944,n34,n1945);
nor (n1945,n1946,n1947);
and (n1946,n205,n44);
and (n1947,n203,n45);
nand (n1948,n1949,n1951);
or (n1949,n1950,n253);
not (n1950,n1733);
nand (n1951,n255,n1952);
nor (n1952,n1953,n1954);
and (n1953,n173,n251);
and (n1954,n172,n250);
nand (n1955,n1956,n1961);
or (n1956,n1957,n513);
not (n1957,n1958);
nand (n1958,n1959,n1960);
or (n1959,n76,n55);
nand (n1960,n76,n55);
nand (n1961,n1772,n528);
or (n1962,n1963,n1964);
and (n1963,n1791,n1803);
and (n1964,n1792,n1800);
or (n1965,n1966,n1967);
and (n1966,n1766,n1812);
and (n1967,n1767,n1790);
or (n1968,n1969,n1970);
and (n1969,n1819,n1842);
and (n1970,n1820,n1839);
nor (n1971,n1972,n2184);
nand (n1972,n1973,n2084);
nand (n1973,n1974,n1978);
not (n1974,n1975);
or (n1975,n1976,n1977);
and (n1976,n1857,n1968);
and (n1977,n1858,n1861);
not (n1978,n1979);
xor (n1979,n1980,n2081);
xor (n1980,n1981,n2047);
xor (n1981,n1982,n1997);
xor (n1982,n1983,n1994);
xor (n1983,n1984,n1991);
xor (n1984,n1985,n1988);
nor (n1985,n1986,n1987);
and (n1986,n219,n33);
not (n1987,n1945);
or (n1988,n1989,n1990);
and (n1989,n1941,n1955);
and (n1990,n1942,n1948);
or (n1991,n1992,n1993);
and (n1992,n1896,n1910);
and (n1993,n1897,n1904);
or (n1994,n1995,n1996);
and (n1995,n1917,n1962);
and (n1996,n1918,n1940);
xor (n1997,n1998,n2024);
xor (n1998,n1999,n2002);
or (n1999,n2000,n2001);
and (n2000,n1919,n1933);
and (n2001,n1920,n1926);
xor (n2002,n2003,n2017);
xor (n2003,n2004,n2010);
nand (n2004,n2005,n2006);
or (n2005,n1957,n529);
nand (n2006,n2007,n514);
nor (n2007,n2008,n2009);
and (n2008,n332,n75);
and (n2009,n43,n76);
nand (n2010,n2011,n2013);
or (n2011,n2012,n114);
not (n2012,n1901);
nand (n2013,n2014,n123);
nor (n2014,n2015,n2016);
and (n2015,n1440,n119);
and (n2016,n297,n118);
nand (n2017,n2018,n2020);
or (n2018,n143,n2019);
not (n2019,n1907);
or (n2020,n2021,n165);
nor (n2021,n2022,n2023);
and (n2022,n90,n1259);
and (n2023,n323,n91);
xor (n2024,n2025,n2041);
xor (n2025,n2026,n2033);
nand (n2026,n2027,n2029);
or (n2027,n2028,n253);
not (n2028,n1952);
nand (n2029,n255,n2030);
nor (n2030,n2031,n2032);
and (n2031,n191,n250);
and (n2032,n192,n251);
nand (n2033,n2034,n2036);
or (n2034,n2035,n86);
not (n2035,n1923);
nand (n2036,n2037,n88);
nand (n2037,n2038,n2039);
or (n2038,n384,n97);
not (n2039,n2040);
and (n2040,n384,n97);
nand (n2041,n2042,n2043);
or (n2042,n65,n1913);
or (n2043,n2044,n73);
nor (n2044,n2045,n2046);
and (n2045,n61,n223);
and (n2046,n62,n722);
xor (n2047,n2048,n2078);
xor (n2048,n2049,n2075);
xor (n2049,n2050,n2072);
xor (n2050,n2051,n2069);
xor (n2051,n2052,n2063);
xor (n2052,n2053,n2060);
nand (n2053,n2054,n2056);
or (n2054,n363,n2055);
not (n2055,n1930);
or (n2056,n748,n2057);
nor (n2057,n2058,n2059);
and (n2058,n496,n359);
and (n2059,n495,n360);
nand (n2060,n2061,n1937);
or (n2061,n389,n2062);
not (n2062,n395);
nand (n2063,n2064,n2065);
or (n2064,n412,n1873);
or (n2065,n420,n2066);
nor (n2066,n2067,n2068);
and (n2067,n125,n729);
and (n2068,n240,n126);
or (n2069,n2070,n2071);
and (n2070,n1869,n1876);
and (n2071,n1870,n1804);
or (n2072,n2073,n2074);
and (n2073,n1888,n1895);
and (n2074,n1889,n1892);
or (n2075,n2076,n2077);
and (n2076,n1864,n1879);
and (n2077,n1865,n1868);
or (n2078,n2079,n2080);
and (n2079,n1886,n1965);
and (n2080,n1887,n1916);
or (n2081,n2082,n2083);
and (n2082,n1862,n1885);
and (n2083,n1863,n1882);
nand (n2084,n2085,n2180);
not (n2085,n2086);
xor (n2086,n2087,n2177);
xor (n2087,n2088,n2107);
xor (n2088,n2089,n2096);
xor (n2089,n2090,n2093);
or (n2090,n2091,n2092);
and (n2091,n1984,n1991);
and (n2092,n1985,n1988);
or (n2093,n2094,n2095);
and (n2094,n1998,n2024);
and (n2095,n1999,n2002);
xor (n2096,n2097,n2104);
xor (n2097,n2098,n2101);
or (n2098,n2099,n2100);
and (n2099,n2003,n2017);
and (n2100,n2004,n2010);
or (n2101,n2102,n2103);
and (n2102,n2025,n2041);
and (n2103,n2026,n2033);
or (n2104,n2105,n2106);
and (n2105,n2052,n2063);
and (n2106,n2053,n2060);
xor (n2107,n2108,n2174);
xor (n2108,n2109,n2171);
xor (n2109,n2110,n2155);
xor (n2110,n2111,n2133);
xor (n2111,n2112,n2127);
xor (n2112,n2113,n2120);
nand (n2113,n2114,n2116);
or (n2114,n2115,n253);
not (n2115,n2030);
nand (n2116,n255,n2117);
nor (n2117,n2118,n2119);
and (n2118,n205,n250);
and (n2119,n203,n251);
nand (n2120,n2121,n2126);
or (n2121,n2122,n748);
not (n2122,n2123);
nor (n2123,n2124,n2125);
and (n2124,n172,n359);
and (n2125,n173,n360);
or (n2126,n363,n2057);
nand (n2127,n2128,n2129);
or (n2128,n65,n2044);
or (n2129,n2130,n73);
nor (n2130,n2131,n2132);
and (n2131,n61,n53);
and (n2132,n62,n55);
xor (n2133,n2134,n2148);
xor (n2134,n2135,n2142);
nand (n2135,n2136,n2138);
or (n2136,n2137,n86);
not (n2137,n2037);
nand (n2138,n2139,n88);
nor (n2139,n2140,n2141);
and (n2140,n306,n96);
and (n2141,n305,n97);
nand (n2142,n2143,n2144);
or (n2143,n2066,n412);
nand (n2144,n421,n2145);
nor (n2145,n2146,n2147);
and (n2146,n1544,n126);
and (n2147,n556,n125);
nand (n2148,n2149,n2151);
or (n2149,n529,n2150);
not (n2150,n2007);
or (n2151,n513,n2152);
nor (n2152,n2153,n2154);
and (n2153,n75,n490);
and (n2154,n76,n489);
xor (n2155,n2156,n2170);
xor (n2156,n2157,n2164);
nand (n2157,n2158,n2160);
or (n2158,n114,n2159);
not (n2159,n2014);
or (n2160,n134,n2161);
nor (n2161,n2162,n2163);
and (n2162,n118,n564);
and (n2163,n234,n119);
nand (n2164,n2165,n2166);
or (n2165,n143,n2021);
or (n2166,n2167,n165);
nor (n2167,n2168,n2169);
and (n2168,n90,n282);
and (n2169,n278,n91);
not (n2170,n1985);
or (n2171,n2172,n2173);
and (n2172,n2050,n2072);
and (n2173,n2051,n2069);
or (n2174,n2175,n2176);
and (n2175,n1982,n1997);
and (n2176,n1983,n1994);
or (n2177,n2178,n2179);
and (n2178,n2048,n2078);
and (n2179,n2049,n2075);
not (n2180,n2181);
or (n2181,n2182,n2183);
and (n2182,n1980,n2081);
and (n2183,n1981,n2047);
nand (n2184,n2185,n2270,n2514);
nand (n2185,n2186,n2190);
not (n2186,n2187);
or (n2187,n2188,n2189);
and (n2188,n2087,n2177);
and (n2189,n2088,n2107);
not (n2190,n2191);
xor (n2191,n2192,n2267);
xor (n2192,n2193,n2196);
or (n2193,n2194,n2195);
and (n2194,n2089,n2096);
and (n2195,n2090,n2093);
xor (n2196,n2197,n2245);
xor (n2197,n2198,n2242);
xor (n2198,n2199,n2225);
xor (n2199,n2200,n2203);
or (n2200,n2201,n2202);
and (n2201,n2134,n2148);
and (n2202,n2135,n2142);
xor (n2203,n2204,n2219);
xor (n2204,n2205,n2212);
nand (n2205,n2206,n2207);
or (n2206,n2122,n363);
nand (n2207,n2208,n370);
not (n2208,n2209);
nor (n2209,n2210,n2211);
and (n2210,n191,n360);
and (n2211,n192,n359);
nand (n2212,n2213,n2215);
or (n2213,n2214,n86);
not (n2214,n2139);
or (n2215,n87,n2216);
nor (n2216,n2217,n2218);
and (n2217,n96,n1259);
and (n2218,n323,n97);
nand (n2219,n2220,n2221);
or (n2220,n65,n2130);
or (n2221,n2222,n73);
nor (n2222,n2223,n2224);
and (n2223,n61,n43);
and (n2224,n62,n332);
xor (n2225,n2226,n2236);
xor (n2226,n2227,n2230);
nand (n2227,n2228,n2145);
or (n2228,n421,n2229);
not (n2229,n412);
nand (n2230,n2231,n2232);
or (n2231,n529,n2152);
or (n2232,n513,n2233);
nor (n2233,n2234,n2235);
and (n2234,n75,n496);
and (n2235,n76,n495);
nand (n2236,n2237,n2238);
or (n2237,n114,n2161);
or (n2238,n134,n2239);
nor (n2239,n2240,n2241);
and (n2240,n118,n729);
and (n2241,n240,n119);
or (n2242,n2243,n2244);
and (n2243,n2110,n2155);
and (n2244,n2111,n2133);
xor (n2245,n2246,n2264);
xor (n2246,n2247,n2250);
or (n2247,n2248,n2249);
and (n2248,n2156,n2170);
and (n2249,n2157,n2164);
xor (n2250,n2251,n2261);
xor (n2251,n2252,n2258);
nand (n2252,n2253,n2254);
or (n2253,n143,n2167);
or (n2254,n2255,n165);
nor (n2255,n2256,n2257);
and (n2256,n297,n91);
and (n2257,n1440,n90);
and (n2258,n2259,n2117);
nand (n2259,n2260,n253);
not (n2260,n255);
or (n2261,n2262,n2263);
and (n2262,n2112,n2127);
and (n2263,n2113,n2120);
or (n2264,n2265,n2266);
and (n2265,n2097,n2104);
and (n2266,n2098,n2101);
or (n2267,n2268,n2269);
and (n2268,n2108,n2174);
and (n2269,n2109,n2171);
nor (n2270,n2271,n2343);
nor (n2271,n2272,n2340);
xor (n2272,n2273,n2337);
xor (n2273,n2274,n2320);
xor (n2274,n2275,n2317);
xor (n2275,n2276,n2296);
xor (n2276,n2277,n2290);
xor (n2277,n2278,n2284);
nand (n2278,n2279,n2280);
or (n2279,n143,n2255);
or (n2280,n2281,n165);
nor (n2281,n2282,n2283);
and (n2282,n564,n90);
and (n2283,n234,n91);
nand (n2284,n2285,n2286);
or (n2285,n65,n2222);
or (n2286,n2287,n73);
nor (n2287,n2288,n2289);
and (n2288,n61,n490);
and (n2289,n62,n489);
nand (n2290,n2291,n2292);
or (n2291,n86,n2216);
or (n2292,n87,n2293);
nor (n2293,n2294,n2295);
and (n2294,n96,n282);
and (n2295,n278,n97);
xor (n2296,n2297,n2311);
xor (n2297,n2298,n2305);
nand (n2298,n2299,n2304);
or (n2299,n2300,n748);
not (n2300,n2301);
nand (n2301,n2302,n2303);
or (n2302,n360,n205);
or (n2303,n359,n203);
or (n2304,n363,n2209);
nand (n2305,n2306,n2307);
or (n2306,n529,n2233);
or (n2307,n513,n2308);
nor (n2308,n2309,n2310);
and (n2309,n75,n173);
and (n2310,n76,n172);
nand (n2311,n2312,n2313);
or (n2312,n114,n2239);
or (n2313,n134,n2314);
nor (n2314,n2315,n2316);
and (n2315,n118,n1544);
and (n2316,n556,n119);
or (n2317,n2318,n2319);
and (n2318,n2251,n2261);
and (n2319,n2252,n2258);
xor (n2320,n2321,n2334);
xor (n2321,n2322,n2331);
xor (n2322,n2323,n2328);
xor (n2323,n2324,n2325);
not (n2324,n2258);
or (n2325,n2326,n2327);
and (n2326,n2204,n2219);
and (n2327,n2205,n2212);
or (n2328,n2329,n2330);
and (n2329,n2226,n2236);
and (n2330,n2227,n2230);
or (n2331,n2332,n2333);
and (n2332,n2199,n2225);
and (n2333,n2200,n2203);
or (n2334,n2335,n2336);
and (n2335,n2246,n2264);
and (n2336,n2247,n2250);
or (n2337,n2338,n2339);
and (n2338,n2197,n2245);
and (n2339,n2198,n2242);
or (n2340,n2341,n2342);
and (n2341,n2192,n2267);
and (n2342,n2193,n2196);
nand (n2343,n2344,n2470);
or (n2344,n2345,n2438);
or (n2345,n2346,n2437);
and (n2346,n2347,n2428);
xor (n2347,n2348,n2371);
or (n2348,n2349,n2370);
and (n2349,n2350,n2357);
xor (n2350,n2351,n2354);
or (n2351,n2352,n2353);
and (n2352,n2277,n2290);
and (n2353,n2278,n2284);
or (n2354,n2355,n2356);
and (n2355,n2297,n2311);
and (n2356,n2298,n2305);
xor (n2357,n2358,n2368);
xor (n2358,n2359,n2362);
nand (n2359,n2360,n2361);
or (n2360,n123,n115);
not (n2361,n2314);
nand (n2362,n2363,n2364);
or (n2363,n143,n2281);
or (n2364,n2365,n165);
nor (n2365,n2366,n2367);
and (n2366,n90,n729);
and (n2367,n240,n91);
nand (n2368,n2369,n2301);
or (n2369,n364,n370);
and (n2370,n2351,n2354);
xor (n2371,n2372,n2417);
xor (n2372,n2373,n2402);
xor (n2373,n2374,n2393);
xor (n2374,n2375,n2384);
nand (n2375,n2376,n2380);
or (n2376,n529,n2377);
nor (n2377,n2378,n2379);
and (n2378,n75,n192);
and (n2379,n76,n191);
or (n2380,n513,n2381);
nor (n2381,n2382,n2383);
and (n2382,n75,n203);
and (n2383,n76,n205);
nand (n2384,n2385,n2389);
or (n2385,n65,n2386);
nor (n2386,n2387,n2388);
and (n2387,n61,n496);
and (n2388,n62,n495);
or (n2389,n2390,n73);
nor (n2390,n2391,n2392);
and (n2391,n61,n173);
and (n2392,n62,n172);
nand (n2393,n2394,n2398);
or (n2394,n86,n2395);
nor (n2395,n2396,n2397);
and (n2396,n96,n1440);
and (n2397,n297,n97);
or (n2398,n87,n2399);
nor (n2399,n2400,n2401);
and (n2400,n96,n564);
and (n2401,n234,n97);
or (n2402,n2403,n2416);
and (n2403,n2404,n2411);
xor (n2404,n2405,n2408);
nand (n2405,n2406,n2407);
or (n2406,n86,n2293);
or (n2407,n87,n2395);
nand (n2408,n2409,n2410);
or (n2409,n65,n2287);
or (n2410,n2386,n73);
not (n2411,n2412);
nand (n2412,n2413,n2414);
or (n2413,n2308,n529);
nand (n2414,n2415,n514);
not (n2415,n2377);
and (n2416,n2405,n2408);
xor (n2417,n2418,n2425);
xor (n2418,n2419,n2412);
nand (n2419,n2420,n2421);
or (n2420,n143,n2365);
or (n2421,n2422,n165);
nor (n2422,n2423,n2424);
and (n2423,n90,n1544);
and (n2424,n556,n91);
or (n2425,n2426,n2427);
and (n2426,n2358,n2368);
and (n2427,n2359,n2362);
or (n2428,n2429,n2436);
and (n2429,n2430,n2435);
xor (n2430,n2431,n2432);
xor (n2431,n2404,n2411);
or (n2432,n2433,n2434);
and (n2433,n2323,n2328);
and (n2434,n2324,n2325);
xor (n2435,n2350,n2357);
and (n2436,n2431,n2432);
and (n2437,n2348,n2371);
xor (n2438,n2439,n2467);
xor (n2439,n2440,n2443);
or (n2440,n2441,n2442);
and (n2441,n2418,n2425);
and (n2442,n2419,n2412);
xor (n2443,n2444,n2450);
xor (n2444,n2445,n2447);
nor (n2445,n2446,n2381);
and (n2446,n529,n513);
or (n2447,n2448,n2449);
and (n2448,n2374,n2393);
and (n2449,n2375,n2384);
xor (n2450,n2451,n2464);
xor (n2451,n2452,n2458);
nand (n2452,n2453,n2454);
or (n2453,n86,n2399);
or (n2454,n87,n2455);
nor (n2455,n2456,n2457);
and (n2456,n96,n729);
and (n2457,n240,n97);
nand (n2458,n2459,n2460);
or (n2459,n65,n2390);
or (n2460,n2461,n73);
nor (n2461,n2462,n2463);
and (n2462,n61,n192);
and (n2463,n62,n191);
nand (n2464,n2465,n2466);
or (n2465,n150,n144);
not (n2466,n2422);
or (n2467,n2468,n2469);
and (n2468,n2372,n2417);
and (n2469,n2373,n2402);
nor (n2470,n2471,n2499);
nor (n2471,n2472,n2475);
or (n2472,n2473,n2474);
and (n2473,n2439,n2467);
and (n2474,n2440,n2443);
xor (n2475,n2476,n2496);
xor (n2476,n2477,n2480);
or (n2477,n2478,n2479);
and (n2478,n2451,n2464);
and (n2479,n2452,n2458);
xor (n2480,n2481,n2495);
xor (n2481,n2482,n2489);
nand (n2482,n2483,n2488);
or (n2483,n73,n2484);
not (n2484,n2485);
nand (n2485,n2486,n2487);
or (n2486,n62,n205);
or (n2487,n61,n203);
or (n2488,n65,n2461);
nand (n2489,n2490,n2491);
or (n2490,n86,n2455);
or (n2491,n87,n2492);
nor (n2492,n2493,n2494);
and (n2493,n96,n1544);
and (n2494,n556,n97);
not (n2495,n2445);
or (n2496,n2497,n2498);
and (n2497,n2444,n2450);
and (n2498,n2445,n2447);
and (n2499,n2500,n2504);
not (n2500,n2501);
or (n2501,n2502,n2503);
and (n2502,n2476,n2496);
and (n2503,n2477,n2480);
not (n2504,n2505);
xor (n2505,n2506,n2511);
xor (n2506,n2507,n2509);
nand (n2507,n2508,n2485);
or (n2508,n1109,n83);
nor (n2509,n2510,n2492);
and (n2510,n86,n87);
or (n2511,n2512,n2513);
and (n2512,n2481,n2495);
and (n2513,n2482,n2489);
nor (n2514,n2515,n2528);
nor (n2515,n2516,n2519);
or (n2516,n2517,n2518);
and (n2517,n2273,n2337);
and (n2518,n2274,n2320);
xor (n2519,n2520,n2525);
xor (n2520,n2521,n2524);
or (n2521,n2522,n2523);
and (n2522,n2275,n2317);
and (n2523,n2276,n2296);
xor (n2524,n2430,n2435);
or (n2525,n2526,n2527);
and (n2526,n2321,n2334);
and (n2527,n2322,n2331);
nor (n2528,n2529,n2532);
or (n2529,n2530,n2531);
and (n2530,n2520,n2525);
and (n2531,n2521,n2524);
xor (n2532,n2347,n2428);
nand (n2533,n1712,n2534,n2539);
nor (n2534,n1395,n2535);
nand (n2535,n20,n2536);
nand (n2536,n2537,n2538);
not (n2537,n1216);
not (n2538,n1217);
nand (n2539,n2540,n3431);
or (n2540,n2541,n2792);
not (n2541,n2542);
nor (n2542,n2543,n2648);
nor (n2543,n2544,n2545);
xor (n2544,n1219,n1392);
or (n2545,n2546,n2647);
and (n2546,n2547,n2646);
xor (n2547,n2548,n2549);
xor (n2548,n1222,n1231);
or (n2549,n2550,n2645);
and (n2550,n2551,n2638);
xor (n2551,n2552,n2553);
xor (n2552,n1233,n1370);
or (n2553,n2554,n2637);
and (n2554,n2555,n2607);
xor (n2555,n2556,n2557);
xor (n2556,n823,n845);
or (n2557,n2558,n2606);
and (n2558,n2559,n2580);
xor (n2559,n2560,n2561);
xor (n2560,n1350,n1361);
or (n2561,n2562,n2579);
and (n2562,n2563,n2572);
xor (n2563,n2564,n2571);
nand (n2564,n2565,n2570);
or (n2565,n2566,n176);
not (n2566,n2567);
nor (n2567,n2568,n2569);
and (n2568,n548,n181);
and (n2569,n217,n174);
nand (n2570,n186,n1364);
xor (n2571,n1345,n1346);
nand (n2572,n2573,n2578);
or (n2573,n219,n2574);
not (n2574,n2575);
nor (n2575,n2576,n2577);
and (n2576,n362,n44);
and (n2577,n358,n45);
or (n2578,n33,n1249);
and (n2579,n2564,n2571);
or (n2580,n2581,n2605);
and (n2581,n2582,n2598);
xor (n2582,n2583,n2591);
nand (n2583,n2584,n2590);
or (n2584,n2585,n283);
not (n2585,n2586);
nand (n2586,n2587,n2588);
or (n2587,n403,n280);
not (n2588,n2589);
and (n2589,n403,n280);
nand (n2590,n285,n1265);
nand (n2591,n2592,n2597);
or (n2592,n2593,n310);
not (n2593,n2594);
nor (n2594,n2595,n2596);
and (n2595,n130,n307);
and (n2596,n131,n309);
nand (n2597,n320,n1285);
nand (n2598,n2599,n2604);
or (n2599,n2600,n253);
not (n2600,n2601);
nand (n2601,n2602,n2603);
or (n2602,n251,n662);
nand (n2603,n251,n662);
nand (n2604,n255,n1278);
and (n2605,n2583,n2591);
and (n2606,n2560,n2561);
or (n2607,n2608,n2636);
and (n2608,n2609,n2635);
xor (n2609,n2610,n2634);
or (n2610,n2611,n2633);
and (n2611,n2612,n2627);
xor (n2612,n2613,n2621);
nand (n2613,n2614,n2620);
or (n2614,n2615,n395);
not (n2615,n2616);
nand (n2616,n2617,n2619);
not (n2617,n2618);
and (n2618,n156,n385);
nand (n2619,n671,n387);
nand (n2620,n1292,n389);
nand (n2621,n2622,n2626);
or (n2622,n2623,n412);
nor (n2623,n2624,n2625);
and (n2624,n125,n101);
and (n2625,n126,n102);
nand (n2626,n1315,n421);
nand (n2627,n2628,n2632);
or (n2628,n198,n2629);
nor (n2629,n2630,n2631);
and (n2630,n179,n55);
nor (n2631,n55,n179);
or (n2632,n1334,n199);
and (n2633,n2613,n2621);
xor (n2634,n1331,n1344);
xor (n2635,n1246,n1262);
and (n2636,n2610,n2634);
and (n2637,n2556,n2557);
or (n2638,n2639,n2644);
and (n2639,n2640,n2643);
xor (n2640,n2641,n2642);
xor (n2641,n1301,n1348);
xor (n2642,n1236,n1272);
xor (n2643,n1383,n1386);
and (n2644,n2641,n2642);
and (n2645,n2552,n2553);
xor (n2646,n1375,n1378);
and (n2647,n2548,n2549);
nor (n2648,n2649,n2650);
xor (n2649,n2547,n2646);
or (n2650,n2651,n2791);
and (n2651,n2652,n2790);
xor (n2652,n2653,n2654);
xor (n2653,n1380,n1389);
or (n2654,n2655,n2789);
and (n2655,n2656,n2788);
xor (n2656,n2657,n2701);
or (n2657,n2658,n2700);
and (n2658,n2659,n2662);
xor (n2659,n2660,n2661);
xor (n2660,n1274,n1289);
xor (n2661,n1304,n1320);
or (n2662,n2663,n2699);
and (n2663,n2664,n2679);
xor (n2664,n2665,n2672);
nand (n2665,n2666,n2671);
or (n2666,n339,n2667);
not (n2667,n2668);
nor (n2668,n2669,n2670);
and (n2669,n36,n248);
and (n2670,n37,n249);
or (n2671,n333,n1340);
nand (n2672,n2673,n2674);
or (n2673,n228,n1256);
nand (n2674,n2675,n714);
not (n2675,n2676);
nor (n2676,n2677,n2678);
and (n2677,n287,n305);
and (n2678,n230,n306);
or (n2679,n2680,n2698);
and (n2680,n2681,n2695);
xor (n2681,n2682,n2689);
nand (n2682,n2683,n2688);
or (n2683,n198,n2684);
not (n2684,n2685);
nand (n2685,n2686,n2687);
or (n2686,n722,n179);
nand (n2687,n179,n722);
or (n2688,n2629,n199);
nand (n2689,n2690,n2691);
or (n2690,n2667,n333);
nand (n2691,n2692,n1114);
nor (n2692,n2693,n2694);
and (n2693,n706,n36);
and (n2694,n376,n37);
nor (n2695,n2696,n2697);
nand (n2696,n255,n452);
nand (n2697,n421,n460);
and (n2698,n2682,n2689);
and (n2699,n2665,n2672);
and (n2700,n2660,n2661);
or (n2701,n2702,n2787);
and (n2702,n2703,n2786);
xor (n2703,n2704,n2779);
or (n2704,n2705,n2778);
and (n2705,n2706,n2753);
xor (n2706,n2707,n2732);
or (n2707,n2708,n2731);
and (n2708,n2709,n2725);
xor (n2709,n2710,n2717);
nand (n2710,n2711,n2712);
or (n2711,n2260,n2600);
nand (n2712,n2260,n2713,n2716);
nand (n2713,n2714,n2715);
or (n2714,n251,n454);
nand (n2715,n454,n251);
not (n2716,n259);
nand (n2717,n2718,n2724);
or (n2718,n2719,n395);
not (n2719,n2720);
nand (n2720,n2721,n2722);
or (n2721,n385,n108);
not (n2722,n2723);
and (n2723,n108,n385);
nand (n2724,n389,n2616);
nand (n2725,n2726,n2730);
or (n2726,n412,n2727);
nor (n2727,n2728,n2729);
and (n2728,n459,n125);
and (n2729,n460,n126);
or (n2730,n420,n2623);
and (n2731,n2710,n2717);
or (n2732,n2733,n2752);
and (n2733,n2734,n2746);
xor (n2734,n2735,n2741);
nor (n2735,n2736,n250);
and (n2736,n2737,n2740);
nand (n2737,n2738,n44);
not (n2738,n2739);
and (n2739,n452,n257);
nand (n2740,n454,n262);
nor (n2741,n2742,n126);
nor (n2742,n2743,n2745);
and (n2743,n2744,n385);
nand (n2744,n460,n419);
and (n2745,n459,n416);
nand (n2746,n2747,n2751);
or (n2747,n2748,n176);
nor (n2748,n2749,n2750);
and (n2749,n267,n181);
and (n2750,n266,n174);
nand (n2751,n2567,n186);
and (n2752,n2735,n2741);
or (n2753,n2754,n2777);
and (n2754,n2755,n2770);
xor (n2755,n2756,n2763);
nand (n2756,n2757,n2762);
or (n2757,n2758,n219);
not (n2758,n2759);
nand (n2759,n2760,n2761);
or (n2760,n81,n44);
nand (n2761,n44,n81);
nand (n2762,n34,n2575);
nand (n2763,n2764,n2769);
or (n2764,n283,n2765);
not (n2765,n2766);
nor (n2766,n2767,n2768);
and (n2767,n140,n280);
and (n2768,n138,n279);
nand (n2769,n285,n2586);
nand (n2770,n2771,n2776);
or (n2771,n2772,n310);
not (n2772,n2773);
nor (n2773,n2774,n2775);
and (n2774,n162,n307);
and (n2775,n163,n309);
nand (n2776,n320,n2594);
and (n2777,n2756,n2763);
and (n2778,n2707,n2732);
or (n2779,n2780,n2785);
and (n2780,n2781,n2784);
xor (n2781,n2782,n2783);
xor (n2782,n2612,n2627);
xor (n2783,n2582,n2598);
xor (n2784,n2563,n2572);
and (n2785,n2782,n2783);
xor (n2786,n2559,n2580);
and (n2787,n2704,n2779);
xor (n2788,n2555,n2607);
and (n2789,n2657,n2701);
xor (n2790,n2551,n2638);
and (n2791,n2653,n2654);
not (n2792,n2793);
nor (n2793,n2794,n3412);
nor (n2794,n2795,n3411);
and (n2795,n2796,n3394);
nand (n2796,n2797,n3393);
or (n2797,n2798,n3070);
not (n2798,n2799);
or (n2799,n2800,n2990);
xor (n2800,n2801,n2905);
xor (n2801,n2802,n2898);
or (n2802,n2803,n2897);
and (n2803,n2804,n2890);
xor (n2804,n2805,n2860);
xor (n2805,n2806,n2836);
xor (n2806,n2807,n2814);
nand (n2807,n2808,n2813);
or (n2808,n227,n2809);
not (n2809,n2810);
nor (n2810,n2811,n2812);
and (n2811,n383,n230);
and (n2812,n384,n287);
or (n2813,n2676,n228);
or (n2814,n2815,n2835);
and (n2815,n2816,n2828);
xor (n2816,n2817,n2821);
nand (n2817,n2818,n2820);
or (n2818,n2819,n2697);
not (n2819,n2696);
nand (n2820,n2819,n2697);
nand (n2821,n2822,n2827);
or (n2822,n198,n2823);
not (n2823,n2824);
nor (n2824,n2825,n2826);
and (n2825,n217,n179);
and (n2826,n548,n184);
nand (n2827,n2685,n196);
nand (n2828,n2829,n2834);
or (n2829,n176,n2830);
not (n2830,n2831);
nor (n2831,n2832,n2833);
and (n2832,n248,n181);
and (n2833,n249,n174);
or (n2834,n1173,n2748);
and (n2835,n2817,n2821);
or (n2836,n2837,n2859);
and (n2837,n2838,n2852);
xor (n2838,n2839,n2845);
nand (n2839,n2840,n2844);
nand (n2840,n1114,n2841);
nand (n2841,n2842,n2843);
or (n2842,n358,n36);
nand (n2843,n36,n358);
nand (n2844,n2692,n591);
nand (n2845,n2846,n2847);
or (n2846,n228,n2809);
nand (n2847,n2848,n714);
nand (n2848,n2849,n2851);
not (n2849,n2850);
and (n2850,n403,n230);
nand (n2851,n287,n405);
nand (n2852,n2853,n2858);
or (n2853,n2854,n283);
not (n2854,n2855);
nor (n2855,n2856,n2857);
and (n2856,n130,n280);
and (n2857,n131,n279);
nand (n2858,n285,n2766);
and (n2859,n2839,n2845);
or (n2860,n2861,n2889);
and (n2861,n2862,n2888);
xor (n2862,n2863,n2864);
xor (n2863,n2838,n2852);
xor (n2864,n2865,n2880);
xor (n2865,n2866,n2873);
nand (n2866,n2867,n2872);
or (n2867,n2868,n219);
not (n2868,n2869);
nand (n2869,n2870,n2871);
or (n2870,n63,n44);
nand (n2871,n44,n63);
nand (n2872,n2759,n34);
nand (n2873,n2874,n2879);
or (n2874,n2875,n310);
not (n2875,n2876);
nor (n2876,n2877,n2878);
and (n2877,n671,n307);
and (n2878,n156,n309);
nand (n2879,n320,n2773);
nand (n2880,n2881,n2887);
or (n2881,n2882,n395);
not (n2882,n2883);
nand (n2883,n2884,n2885);
or (n2884,n385,n102);
not (n2885,n2886);
and (n2886,n102,n385);
nand (n2887,n389,n2720);
xor (n2888,n2816,n2828);
and (n2889,n2863,n2864);
xor (n2890,n2891,n2896);
xor (n2891,n2892,n2893);
xor (n2892,n2734,n2746);
or (n2893,n2894,n2895);
and (n2894,n2865,n2880);
and (n2895,n2866,n2873);
xor (n2896,n2755,n2770);
and (n2897,n2805,n2860);
xor (n2898,n2899,n2904);
xor (n2899,n2900,n2903);
or (n2900,n2901,n2902);
and (n2901,n2806,n2836);
and (n2902,n2807,n2814);
xor (n2903,n2664,n2679);
xor (n2904,n2706,n2753);
xor (n2905,n2906,n2911);
xor (n2906,n2907,n2910);
or (n2907,n2908,n2909);
and (n2908,n2891,n2896);
and (n2909,n2892,n2893);
xor (n2910,n2781,n2784);
or (n2911,n2912,n2989);
and (n2912,n2913,n2916);
xor (n2913,n2914,n2915);
xor (n2914,n2681,n2695);
xor (n2915,n2709,n2725);
or (n2916,n2917,n2988);
and (n2917,n2918,n2963);
xor (n2918,n2919,n2940);
or (n2919,n2920,n2939);
and (n2920,n2921,n2932);
xor (n2921,n2922,n2929);
nand (n2922,n2923,n2928);
or (n2923,n2924,n176);
not (n2924,n2925);
nand (n2925,n2926,n2927);
or (n2926,n706,n174);
nand (n2927,n174,n706);
nand (n2928,n2831,n186);
nor (n2929,n2930,n2931);
nand (n2930,n34,n452);
nand (n2931,n389,n460);
nand (n2932,n2933,n2938);
or (n2933,n2934,n339);
not (n2934,n2935);
nand (n2935,n2936,n2937);
or (n2936,n81,n36);
or (n2937,n37,n527);
nand (n2938,n591,n2841);
and (n2939,n2922,n2929);
or (n2940,n2941,n2962);
and (n2941,n2942,n2955);
xor (n2942,n2943,n2950);
nor (n2943,n2944,n44);
and (n2944,n2945,n2948);
nand (n2945,n2946,n36);
not (n2946,n2947);
and (n2947,n452,n38);
nand (n2948,n2949,n454);
not (n2949,n38);
nor (n2950,n2951,n385);
nor (n2951,n2952,n2954);
and (n2952,n2953,n307);
nand (n2953,n460,n391);
and (n2954,n459,n392);
nand (n2955,n2956,n2961);
or (n2956,n2957,n219);
not (n2957,n2958);
nor (n2958,n2959,n2960);
and (n2959,n44,n454);
and (n2960,n452,n45);
nand (n2961,n2869,n34);
and (n2962,n2943,n2950);
or (n2963,n2964,n2987);
and (n2964,n2965,n2980);
xor (n2965,n2966,n2973);
nand (n2966,n2967,n2972);
or (n2967,n2968,n310);
not (n2968,n2969);
nor (n2969,n2970,n2971);
and (n2970,n107,n307);
and (n2971,n108,n309);
nand (n2972,n320,n2876);
nand (n2973,n2974,n2975);
or (n2974,n388,n2882);
nand (n2975,n2976,n2062);
not (n2976,n2977);
nor (n2977,n2978,n2979);
and (n2978,n459,n387);
and (n2979,n460,n385);
nand (n2980,n2981,n2986);
or (n2981,n198,n2982);
not (n2982,n2983);
nand (n2983,n2984,n2985);
or (n2984,n267,n184);
nand (n2985,n184,n267);
or (n2986,n2823,n199);
and (n2987,n2966,n2973);
and (n2988,n2919,n2940);
and (n2989,n2914,n2915);
or (n2990,n2991,n3069);
and (n2991,n2992,n3068);
xor (n2992,n2993,n2994);
xor (n2993,n2913,n2916);
or (n2994,n2995,n3067);
and (n2995,n2996,n3066);
xor (n2996,n2997,n3037);
or (n2997,n2998,n3036);
and (n2998,n2999,n3014);
xor (n2999,n3000,n3007);
nand (n3000,n3001,n3005);
or (n3001,n3002,n227);
nor (n3002,n3003,n3004);
and (n3003,n287,n140);
and (n3004,n230,n138);
or (n3005,n3006,n228);
not (n3006,n2848);
nand (n3007,n3008,n3013);
or (n3008,n3009,n283);
not (n3009,n3010);
nor (n3010,n3011,n3012);
and (n3011,n162,n280);
and (n3012,n163,n279);
nand (n3013,n285,n2855);
or (n3014,n3015,n3035);
and (n3015,n3016,n3028);
xor (n3016,n3017,n3024);
nand (n3017,n3018,n3023);
or (n3018,n3019,n198);
not (n3019,n3020);
nor (n3020,n3021,n3022);
and (n3021,n249,n179);
and (n3022,n248,n184);
nand (n3023,n2983,n196);
nand (n3024,n3025,n3027);
or (n3025,n3026,n2931);
not (n3026,n2930);
nand (n3027,n3026,n2931);
nand (n3028,n3029,n3034);
or (n3029,n176,n3030);
not (n3030,n3031);
nand (n3031,n3032,n3033);
or (n3032,n362,n174);
nand (n3033,n174,n362);
or (n3034,n1173,n2924);
and (n3035,n3017,n3024);
and (n3036,n3000,n3007);
or (n3037,n3038,n3065);
and (n3038,n3039,n3064);
xor (n3039,n3040,n3041);
xor (n3040,n2942,n2955);
or (n3041,n3042,n3063);
and (n3042,n3043,n3057);
xor (n3043,n3044,n3050);
nand (n3044,n3045,n3049);
or (n3045,n3046,n227);
nor (n3046,n3047,n3048);
and (n3047,n287,n130);
and (n3048,n230,n131);
or (n3049,n3002,n228);
nand (n3050,n3051,n3056);
or (n3051,n3052,n339);
not (n3052,n3053);
nor (n3053,n3054,n3055);
and (n3054,n662,n36);
and (n3055,n63,n37);
nand (n3056,n2935,n591);
nand (n3057,n3058,n3062);
or (n3058,n283,n3059);
nor (n3059,n3060,n3061);
and (n3060,n279,n671);
and (n3061,n280,n156);
nand (n3062,n285,n3010);
and (n3063,n3044,n3050);
xor (n3064,n2965,n2980);
and (n3065,n3040,n3041);
xor (n3066,n2918,n2963);
and (n3067,n2997,n3037);
xor (n3068,n2804,n2890);
and (n3069,n2993,n2994);
not (n3070,n3071);
nand (n3071,n3072,n3389,n3392);
nand (n3072,n3073,n3143,n3384);
nand (n3073,n3074,n3076);
not (n3074,n3075);
xor (n3075,n2992,n3068);
not (n3076,n3077);
or (n3077,n3078,n3142);
and (n3078,n3079,n3141);
xor (n3079,n3080,n3081);
xor (n3080,n2862,n2888);
or (n3081,n3082,n3140);
and (n3082,n3083,n3139);
xor (n3083,n3084,n3085);
xor (n3084,n2921,n2932);
or (n3085,n3086,n3138);
and (n3086,n3087,n3117);
xor (n3087,n3088,n3096);
nand (n3088,n3089,n3095);
or (n3089,n3090,n310);
not (n3090,n3091);
nand (n3091,n3092,n3093);
or (n3092,n307,n102);
not (n3093,n3094);
and (n3094,n102,n307);
nand (n3095,n320,n2969);
or (n3096,n3097,n3116);
and (n3097,n3098,n3109);
xor (n3098,n3099,n3106);
nand (n3099,n3100,n3105);
or (n3100,n3101,n176);
not (n3101,n3102);
nand (n3102,n3103,n3104);
or (n3103,n81,n181);
nand (n3104,n181,n81);
nand (n3105,n3031,n186);
nor (n3106,n3107,n3108);
nand (n3107,n320,n460);
nand (n3108,n591,n452);
nand (n3109,n3110,n3115);
or (n3110,n227,n3111);
not (n3111,n3112);
nor (n3112,n3113,n3114);
and (n3113,n163,n287);
and (n3114,n162,n230);
or (n3115,n3046,n228);
and (n3116,n3099,n3106);
or (n3117,n3118,n3137);
and (n3118,n3119,n3131);
xor (n3119,n3120,n3126);
nor (n3120,n3121,n36);
and (n3121,n3122,n3125);
nand (n3122,n3123,n181);
not (n3123,n3124);
and (n3124,n452,n335);
nand (n3125,n454,n337);
and (n3126,n3127,n309);
nand (n3127,n3128,n3129);
or (n3128,n313,n460);
nand (n3129,n3130,n280);
or (n3130,n314,n459);
nand (n3131,n3132,n3133);
or (n3132,n199,n3019);
nand (n3133,n3134,n197);
nand (n3134,n3135,n3136);
or (n3135,n376,n184);
nand (n3136,n184,n376);
and (n3137,n3120,n3126);
and (n3138,n3088,n3096);
xor (n3139,n2999,n3014);
and (n3140,n3084,n3085);
xor (n3141,n2996,n3066);
and (n3142,n3080,n3081);
nand (n3143,n3144,n3383);
or (n3144,n3145,n3369);
not (n3145,n3146);
nand (n3146,n3147,n3368);
or (n3147,n3148,n3351);
nor (n3148,n3149,n3350);
and (n3149,n3150,n3263);
nand (n3150,n3151,n3232);
not (n3151,n3152);
xor (n3152,n3153,n3206);
xor (n3153,n3154,n3176);
xor (n3154,n3155,n3170);
xor (n3155,n3156,n3163);
nand (n3156,n3157,n3162);
or (n3157,n3158,n339);
not (n3158,n3159);
nand (n3159,n3160,n3161);
or (n3160,n452,n36);
or (n3161,n454,n37);
nand (n3162,n3053,n591);
nand (n3163,n3164,n3169);
or (n3164,n3165,n283);
not (n3165,n3166);
nor (n3166,n3167,n3168);
and (n3167,n108,n279);
and (n3168,n107,n280);
or (n3169,n284,n3059);
nand (n3170,n3171,n3172);
or (n3171,n311,n3090);
or (n3172,n310,n3173);
nor (n3173,n3174,n3175);
and (n3174,n459,n309);
and (n3175,n460,n307);
or (n3176,n3177,n3205);
and (n3177,n3178,n3193);
xor (n3178,n3179,n3185);
nand (n3179,n3180,n3184);
or (n3180,n3181,n283);
nor (n3181,n3182,n3183);
and (n3182,n102,n280);
and (n3183,n101,n279);
nand (n3184,n3166,n285);
nand (n3185,n3186,n3191);
or (n3186,n198,n3187);
not (n3187,n3188);
nor (n3188,n3189,n3190);
and (n3189,n358,n179);
and (n3190,n362,n184);
or (n3191,n3192,n199);
not (n3192,n3134);
and (n3193,n3194,n3200);
nor (n3194,n3195,n181);
and (n3195,n3196,n3199);
nand (n3196,n3197,n184);
not (n3197,n3198);
and (n3198,n452,n180);
nand (n3199,n183,n454);
nor (n3200,n3201,n280);
and (n3201,n3202,n3204);
nand (n3202,n3203,n230);
or (n3203,n459,n288);
nand (n3204,n459,n288);
and (n3205,n3179,n3185);
xor (n3206,n3207,n3231);
xor (n3207,n3208,n3230);
or (n3208,n3209,n3229);
and (n3209,n3210,n3225);
xor (n3210,n3211,n3218);
nand (n3211,n3212,n3217);
or (n3212,n3213,n176);
not (n3213,n3214);
nand (n3214,n3215,n3216);
or (n3215,n63,n181);
nand (n3216,n181,n63);
nand (n3217,n3102,n186);
nand (n3218,n3219,n3220);
or (n3219,n228,n3111);
nand (n3220,n3221,n714);
nand (n3221,n3222,n3224);
not (n3222,n3223);
and (n3223,n156,n230);
nand (n3224,n287,n671);
nand (n3225,n3226,n3228);
or (n3226,n3227,n3107);
not (n3227,n3108);
nand (n3228,n3227,n3107);
and (n3229,n3211,n3218);
xor (n3230,n3119,n3131);
xor (n3231,n3098,n3109);
not (n3232,n3233);
or (n3233,n3234,n3262);
and (n3234,n3235,n3261);
xor (n3235,n3236,n3260);
or (n3236,n3237,n3259);
and (n3237,n3238,n3253);
xor (n3238,n3239,n3246);
nand (n3239,n3240,n3245);
or (n3240,n3241,n176);
not (n3241,n3242);
nor (n3242,n3243,n3244);
and (n3243,n454,n181);
and (n3244,n452,n174);
nand (n3245,n3214,n186);
nand (n3246,n3247,n3252);
or (n3247,n227,n3248);
not (n3248,n3249);
nor (n3249,n3250,n3251);
and (n3250,n108,n287);
and (n3251,n107,n230);
nand (n3252,n3221,n229);
nand (n3253,n3254,n3258);
or (n3254,n283,n3255);
nor (n3255,n3256,n3257);
and (n3256,n279,n459);
and (n3257,n460,n280);
or (n3258,n284,n3181);
and (n3259,n3239,n3246);
xor (n3260,n3210,n3225);
xor (n3261,n3178,n3193);
and (n3262,n3236,n3260);
nand (n3263,n3264,n3349);
or (n3264,n3265,n3308);
not (n3265,n3266);
nand (n3266,n3267,n3269);
not (n3267,n3268);
xor (n3268,n3235,n3261);
not (n3269,n3270);
or (n3270,n3271,n3307);
and (n3271,n3272,n3285);
xor (n3272,n3273,n3280);
nand (n3273,n3274,n3275);
or (n3274,n199,n3187);
or (n3275,n198,n3276);
not (n3276,n3277);
nor (n3277,n3278,n3279);
and (n3278,n81,n179);
and (n3279,n527,n184);
xor (n3280,n3281,n3282);
xor (n3281,n3194,n3200);
nor (n3282,n3283,n3284);
nand (n3283,n285,n460);
nand (n3284,n186,n452);
or (n3285,n3286,n3306);
and (n3286,n3287,n3299);
xor (n3287,n3288,n3295);
nand (n3288,n3289,n3294);
or (n3289,n198,n3290);
not (n3290,n3291);
nor (n3291,n3292,n3293);
and (n3292,n662,n184);
and (n3293,n63,n179);
nand (n3294,n3277,n196);
nand (n3295,n3296,n3298);
or (n3296,n3284,n3297);
not (n3297,n3283);
nand (n3298,n3297,n3284);
nand (n3299,n3300,n3305);
or (n3300,n227,n3301);
not (n3301,n3302);
nor (n3302,n3303,n3304);
and (n3303,n102,n287);
and (n3304,n101,n230);
nand (n3305,n3249,n229);
and (n3306,n3288,n3295);
and (n3307,n3273,n3280);
not (n3308,n3309);
nand (n3309,n3310,n3348);
or (n3310,n3311,n3314);
nor (n3311,n3312,n3313);
xor (n3312,n3272,n3285);
xor (n3313,n3238,n3253);
nor (n3314,n3315,n3346);
and (n3315,n3316,n3333);
nand (n3316,n3317,n3319);
not (n3317,n3318);
xor (n3318,n3287,n3299);
not (n3319,n3320);
or (n3320,n3321,n3332);
and (n3321,n3322,n3326);
xor (n3322,n3323,n3325);
nor (n3323,n3324,n184);
and (n3324,n452,n196);
and (n3325,n287,n459,n229);
nand (n3326,n3327,n3328);
or (n3327,n228,n3301);
or (n3328,n3329,n227);
nor (n3329,n3330,n3331);
and (n3330,n287,n459);
and (n3331,n460,n230);
and (n3332,n3323,n3325);
or (n3333,n3334,n3345);
and (n3334,n3335,n3344);
xor (n3335,n3336,n3338);
and (n3336,n3324,n3337);
and (n3337,n460,n229);
nand (n3338,n3339,n3340);
or (n3339,n199,n3290);
nand (n3340,n3341,n197);
nand (n3341,n3342,n3343);
or (n3342,n184,n452);
or (n3343,n454,n179);
xor (n3344,n3322,n3326);
and (n3345,n3336,n3338);
not (n3346,n3347);
nand (n3347,n3318,n3320);
nand (n3348,n3312,n3313);
nand (n3349,n3268,n3270);
and (n3350,n3152,n3233);
nor (n3351,n3352,n3365);
xor (n3352,n3353,n3358);
xor (n3353,n3354,n3355);
xor (n3354,n3087,n3117);
or (n3355,n3356,n3357);
and (n3356,n3207,n3231);
and (n3357,n3208,n3230);
xor (n3358,n3359,n3364);
xor (n3359,n3360,n3363);
or (n3360,n3361,n3362);
and (n3361,n3155,n3170);
and (n3362,n3156,n3163);
xor (n3363,n3043,n3057);
xor (n3364,n3016,n3028);
or (n3365,n3366,n3367);
and (n3366,n3153,n3206);
and (n3367,n3154,n3176);
nand (n3368,n3352,n3365);
not (n3369,n3370);
nand (n3370,n3371,n3379);
not (n3371,n3372);
xor (n3372,n3373,n3378);
xor (n3373,n3374,n3377);
or (n3374,n3375,n3376);
and (n3375,n3359,n3364);
and (n3376,n3360,n3363);
xor (n3377,n3039,n3064);
xor (n3378,n3083,n3139);
not (n3379,n3380);
or (n3380,n3381,n3382);
and (n3381,n3353,n3358);
and (n3382,n3354,n3355);
nand (n3383,n3372,n3380);
or (n3384,n3385,n3386);
xor (n3385,n3079,n3141);
or (n3386,n3387,n3388);
and (n3387,n3373,n3378);
and (n3388,n3374,n3377);
nand (n3389,n3073,n3390);
not (n3390,n3391);
nand (n3391,n3385,n3386);
nand (n3392,n3075,n3077);
nand (n3393,n2800,n2990);
or (n3394,n3395,n3408);
xor (n3395,n3396,n3401);
xor (n3396,n3397,n3398);
xor (n3397,n2703,n2786);
or (n3398,n3399,n3400);
and (n3399,n2906,n2911);
and (n3400,n2907,n2910);
xor (n3401,n3402,n3405);
xor (n3402,n3403,n3404);
xor (n3403,n2609,n2635);
xor (n3404,n2659,n2662);
or (n3405,n3406,n3407);
and (n3406,n2899,n2904);
and (n3407,n2900,n2903);
or (n3408,n3409,n3410);
and (n3409,n2801,n2905);
and (n3410,n2802,n2898);
and (n3411,n3395,n3408);
nand (n3412,n3413,n3426);
nand (n3413,n3414,n3416);
not (n3414,n3415);
xor (n3415,n2652,n2790);
not (n3416,n3417);
or (n3417,n3418,n3425);
and (n3418,n3419,n3424);
xor (n3419,n3420,n3421);
xor (n3420,n2640,n2643);
or (n3421,n3422,n3423);
and (n3422,n3402,n3405);
and (n3423,n3403,n3404);
xor (n3424,n2656,n2788);
and (n3425,n3420,n3421);
or (n3426,n3427,n3428);
xor (n3427,n3419,n3424);
or (n3428,n3429,n3430);
and (n3429,n3396,n3401);
and (n3430,n3397,n3398);
nand (n3431,n3432,n3443);
or (n3432,n3433,n3436);
nand (n3433,n3434,n3435);
nand (n3434,n2544,n2545);
nand (n3435,n2649,n2650);
nor (n3436,n3437,n2648);
nand (n3437,n3438,n3413);
or (n3438,n3439,n3441);
not (n3439,n3440);
nand (n3440,n3427,n3428);
not (n3441,n3442);
nand (n3442,n3415,n3417);
not (n3443,n2543);
nor (n3444,n3445,n3448);
and (n3445,n1971,n3446);
nor (n3446,n1852,n3447);
nand (n3447,n1716,n1849);
nand (n3448,n3449,n3453);
or (n3449,n3450,n3452);
not (n3450,n3451);
and (n3451,n1853,n1856);
not (n3452,n1971);
nand (n3453,n3454,n3455,n2084);
not (n3454,n2184);
nand (n3455,n3456,n3457);
or (n3456,n1974,n1978);
or (n3457,n2085,n2180);
nor (n3458,n3459,n3475);
and (n3459,n3460,n3474);
nand (n3460,n3461,n3470);
or (n3461,n3462,n3463);
not (n3462,n2514);
not (n3463,n3464);
nand (n3464,n3465,n3468);
or (n3465,n3466,n3467);
not (n3466,n2272);
not (n3467,n2340);
or (n3468,n3469,n2271);
nand (n3469,n2187,n2191);
nor (n3470,n3471,n3473);
and (n3471,n2516,n3472,n2519);
not (n3472,n2528);
and (n3473,n2529,n2532);
not (n3474,n2343);
nand (n3475,n3476,n3481);
or (n3476,n3477,n2499);
nor (n3477,n3478,n3480);
and (n3478,n2345,n3479,n2438);
not (n3479,n2471);
and (n3480,n2472,n2475);
or (n3481,n2500,n2504);
nor (n3482,n3483,n3488);
and (n3483,n3484,n3487);
or (n3484,n3485,n3486);
and (n3485,n2506,n2511);
and (n3486,n2507,n2509);
not (n3487,n2509);
and (n3488,n3489,n2509);
not (n3489,n3484);
not (n3490,n3491);
nor (n3491,n3492,n7002);
and (n3492,n3493,n7001);
nand (n3493,n3494,n6943,n6960,n6979);
nand (n3494,n3495,n5322,n6019);
not (n3495,n3496);
nand (n3496,n3497,n5073);
and (n3497,n3498,n4721);
nor (n3498,n3499,n4620);
and (n3499,n3500,n4510);
not (n3500,n3501);
or (n3501,n3502,n4509);
and (n3502,n3503,n4316);
xor (n3503,n3504,n4100);
or (n3504,n3505,n4099);
and (n3505,n3506,n3940);
xor (n3506,n3507,n3714);
xor (n3507,n3508,n3672);
xor (n3508,n3509,n3595);
or (n3509,n3510,n3594);
and (n3510,n3511,n3568);
xor (n3511,n3512,n3539);
nand (n3512,n3513,n3534);
or (n3513,n3514,n3523);
not (n3514,n3515);
nand (n3515,n3516,n3520);
not (n3516,n3517);
and (n3517,n3518,n3519);
nand (n3520,n3521,n3522);
not (n3521,n3519);
not (n3522,n3518);
nand (n3523,n3524,n3531);
not (n3524,n3525);
nand (n3525,n3526,n3530);
or (n3526,n3527,n3529);
not (n3527,n3528);
nand (n3530,n3527,n3529);
nand (n3531,n3532,n3533);
or (n3532,n3529,n3521);
nand (n3533,n3521,n3529);
nand (n3534,n3525,n3535);
nand (n3535,n3536,n3538);
or (n3536,n3537,n3519);
nand (n3538,n3519,n3537);
nand (n3539,n3540,n3561);
or (n3540,n3541,n3549);
not (n3541,n3542);
nor (n3542,n3543,n3547);
and (n3543,n3544,n3546);
not (n3544,n3545);
and (n3547,n3545,n3548);
not (n3548,n3546);
nand (n3549,n3550,n3557);
or (n3550,n3551,n3555);
not (n3551,n3552);
nand (n3552,n3553,n3546);
not (n3553,n3554);
not (n3555,n3556);
nand (n3556,n3548,n3554);
not (n3557,n3558);
nand (n3558,n3559,n3560);
or (n3559,n3521,n3554);
nand (n3560,n3521,n3554);
nand (n3561,n3562,n3558);
not (n3562,n3563);
nor (n3563,n3564,n3567);
and (n3564,n3548,n3565);
not (n3565,n3566);
and (n3567,n3566,n3546);
nand (n3568,n3569,n3588);
or (n3569,n3570,n3583);
nand (n3570,n3571,n3578);
nor (n3571,n3572,n3576);
and (n3572,n3573,n3574);
not (n3574,n3575);
and (n3576,n3577,n3575);
not (n3577,n3573);
nand (n3578,n3579,n3582);
or (n3579,n3575,n3580);
not (n3580,n3581);
nand (n3582,n3580,n3575);
not (n3583,n3584);
nand (n3584,n3585,n3587);
or (n3585,n3586,n3580);
nand (n3587,n3580,n3586);
or (n3588,n3589,n3571);
not (n3589,n3590);
nand (n3590,n3591,n3593);
or (n3591,n3592,n3580);
nand (n3593,n3580,n3592);
and (n3594,n3512,n3539);
xor (n3595,n3596,n3644);
xor (n3596,n3597,n3617);
nand (n3597,n3598,n3613);
or (n3598,n3599,n3605);
nand (n3599,n3600,n3604);
or (n3600,n3601,n3603);
not (n3601,n3602);
nand (n3604,n3601,n3603);
not (n3605,n3606);
nand (n3606,n3607,n3608);
not (n3607,n3599);
nand (n3608,n3609,n3612);
or (n3609,n3602,n3610);
not (n3610,n3611);
nand (n3612,n3610,n3602);
nand (n3613,n3614,n3616);
or (n3614,n3615,n3610);
nand (n3616,n3610,n3615);
nand (n3617,n3618,n3638);
or (n3618,n3619,n3627);
not (n3619,n3620);
nand (n3620,n3621,n3625);
or (n3621,n3622,n3623);
not (n3623,n3624);
or (n3625,n3624,n3626);
not (n3626,n3622);
nand (n3627,n3628,n3635);
not (n3628,n3629);
nand (n3629,n3630,n3634);
or (n3630,n3631,n3633);
not (n3631,n3632);
nand (n3634,n3631,n3633);
nand (n3635,n3636,n3637);
or (n3636,n3633,n3623);
nand (n3637,n3623,n3633);
nand (n3638,n3629,n3639);
nor (n3639,n3640,n3642);
and (n3640,n3641,n3624);
and (n3642,n3643,n3623);
not (n3643,n3641);
nand (n3644,n3645,n3661);
or (n3645,n3646,n3654);
not (n3646,n3647);
nor (n3647,n3648,n3652);
and (n3648,n3649,n3651);
not (n3649,n3650);
and (n3652,n3650,n3653);
not (n3653,n3651);
not (n3654,n3655);
nand (n3655,n3656,n3660);
or (n3656,n3657,n3658);
not (n3658,n3659);
nand (n3660,n3658,n3657);
nand (n3661,n3662,n3667);
not (n3662,n3663);
nand (n3663,n3654,n3664);
nand (n3664,n3665,n3666);
or (n3665,n3649,n3657);
nand (n3666,n3649,n3657);
nand (n3667,n3668,n3671);
not (n3668,n3669);
and (n3669,n3670,n3650);
or (n3671,n3650,n3670);
xor (n3672,n3673,n3706);
xor (n3673,n3674,n3697);
nand (n3674,n3675,n3692);
or (n3675,n3676,n3682);
not (n3676,n3677);
nand (n3677,n3678,n3681);
or (n3678,n3679,n3573);
not (n3679,n3680);
nand (n3681,n3679,n3573);
not (n3682,n3683);
nor (n3683,n3684,n3689);
nor (n3684,n3685,n3688);
and (n3685,n3573,n3686);
not (n3686,n3687);
nor (n3688,n3686,n3573);
nand (n3689,n3690,n3691);
or (n3690,n3686,n3624);
nand (n3691,n3686,n3624);
nand (n3692,n3689,n3693);
nand (n3693,n3694,n3696);
or (n3694,n3695,n3577);
nand (n3696,n3577,n3695);
nand (n3697,n3698,n3700);
or (n3698,n3699,n3523);
not (n3699,n3535);
nand (n3700,n3525,n3701);
nor (n3701,n3702,n3705);
and (n3702,n3703,n3519);
not (n3703,n3704);
and (n3705,n3704,n3521);
nand (n3706,n3707,n3713);
or (n3707,n3557,n3708);
not (n3708,n3709);
nand (n3709,n3710,n3711);
or (n3710,n3546,n3518);
not (n3711,n3712);
and (n3712,n3518,n3546);
or (n3713,n3549,n3563);
xor (n3714,n3715,n3845);
xor (n3715,n3716,n3776);
xor (n3716,n3717,n3752);
xor (n3717,n3718,n3726);
nand (n3718,n3719,n3720);
or (n3719,n3589,n3570);
nand (n3720,n3721,n3725);
nand (n3721,n3722,n3724);
or (n3722,n3723,n3580);
nand (n3724,n3580,n3723);
not (n3725,n3571);
nand (n3726,n3727,n3747);
or (n3727,n3728,n3737);
not (n3728,n3729);
nand (n3729,n3730,n3734);
not (n3730,n3731);
and (n3731,n3732,n3733);
nand (n3734,n3735,n3736);
not (n3735,n3733);
not (n3736,n3732);
not (n3737,n3738);
nor (n3738,n3739,n3743);
nand (n3739,n3740,n3742);
or (n3740,n3548,n3741);
nand (n3742,n3548,n3741);
nor (n3743,n3744,n3745);
and (n3744,n3735,n3741);
and (n3745,n3733,n3746);
not (n3746,n3741);
nand (n3747,n3739,n3748);
nand (n3748,n3749,n3751);
not (n3749,n3750);
and (n3750,n3545,n3733);
nand (n3751,n3735,n3544);
nand (n3752,n3753,n3765);
or (n3753,n3754,n3759);
nor (n3754,n3755,n3757);
and (n3755,n3735,n3756);
and (n3757,n3733,n3758);
not (n3758,n3756);
not (n3759,n3760);
nor (n3760,n3761,n3764);
and (n3761,n3762,n3659);
not (n3762,n3763);
and (n3764,n3763,n3658);
or (n3765,n3766,n3771);
not (n3766,n3767);
and (n3767,n3768,n3754);
nor (n3768,n3769,n3770);
and (n3769,n3658,n3758);
and (n3770,n3659,n3756);
not (n3771,n3772);
nand (n3772,n3773,n3775);
or (n3773,n3774,n3659);
nand (n3775,n3659,n3774);
xor (n3776,n3777,n3822);
xor (n3777,n3778,n3802);
nand (n3778,n3779,n3793);
or (n3779,n3780,n3786);
not (n3780,n3781);
nand (n3781,n3782,n3784);
nand (n3782,n3580,n3783);
nand (n3784,n3785,n3581);
not (n3785,n3783);
not (n3786,n3787);
nor (n3787,n3788,n3792);
and (n3788,n3789,n3791);
not (n3789,n3790);
not (n3791,n3586);
and (n3792,n3586,n3790);
nand (n3793,n3794,n3798);
nor (n3794,n3781,n3795);
nor (n3795,n3796,n3797);
and (n3796,n3789,n3783);
and (n3797,n3790,n3785);
nand (n3798,n3799,n3801);
or (n3799,n3800,n3789);
nand (n3801,n3800,n3789);
nand (n3802,n3803,n3817);
or (n3803,n3804,n3810);
nand (n3804,n3805,n3809);
or (n3805,n3806,n3807);
not (n3807,n3808);
nand (n3809,n3807,n3806);
not (n3810,n3811);
nand (n3811,n3812,n3813);
not (n3812,n3804);
nand (n3813,n3814,n3816);
or (n3814,n3815,n3528);
not (n3815,n3806);
nand (n3816,n3528,n3815);
nand (n3817,n3818,n3821);
not (n3818,n3819);
and (n3819,n3820,n3528);
or (n3821,n3528,n3820);
nor (n3822,n3823,n3839);
and (n3823,n3824,n3834);
not (n3824,n3825);
nand (n3825,n3826,n3830);
nand (n3826,n3827,n3829);
or (n3827,n3828,n3631);
nand (n3829,n3631,n3828);
not (n3830,n3831);
nand (n3831,n3832,n3833);
or (n3832,n3610,n3828);
nand (n3833,n3610,n3828);
nand (n3834,n3835,n3838);
or (n3835,n3836,n3632);
not (n3836,n3837);
nand (n3838,n3632,n3836);
and (n3839,n3831,n3840);
nand (n3840,n3841,n3844);
or (n3841,n3842,n3632);
not (n3842,n3843);
nand (n3844,n3632,n3842);
or (n3845,n3846,n3939);
and (n3846,n3847,n3899);
xor (n3847,n3848,n3858);
nand (n3848,n3849,n3854);
or (n3849,n3850,n3606);
not (n3850,n3851);
nor (n3851,n3852,n3853);
and (n3852,n3837,n3611);
and (n3853,n3836,n3610);
nand (n3854,n3599,n3855);
nand (n3855,n3856,n3857);
or (n3856,n3843,n3610);
nand (n3857,n3610,n3843);
or (n3858,n3859,n3898);
and (n3859,n3860,n3885);
xor (n3860,n3861,n3877);
nand (n3861,n3862,n3874);
or (n3862,n3863,n3869);
nand (n3863,n3864,n3868);
or (n3864,n3865,n3867);
not (n3865,n3866);
nand (n3868,n3865,n3867);
nand (n3869,n3870,n3872);
nand (n3870,n3866,n3867,n3871);
not (n3871,n3603);
nand (n3872,n3865,n3873,n3603);
not (n3873,n3867);
nand (n3874,n3875,n3876);
or (n3875,n3615,n3871);
nand (n3876,n3871,n3615);
nand (n3877,n3878,n3884);
or (n3878,n3570,n3879);
not (n3879,n3880);
nand (n3880,n3881,n3883);
or (n3881,n3581,n3882);
not (n3882,n3800);
nand (n3883,n3581,n3882);
nand (n3884,n3725,n3584);
nand (n3885,n3886,n3893);
or (n3886,n3887,n3892);
not (n3887,n3888);
nand (n3888,n3889,n3891);
not (n3889,n3890);
and (n3890,n3763,n3733);
nand (n3891,n3735,n3762);
not (n3892,n3739);
or (n3893,n3737,n3894);
not (n3894,n3895);
nand (n3895,n3896,n3897);
or (n3896,n3733,n3774);
nand (n3897,n3774,n3733);
and (n3898,n3861,n3877);
or (n3899,n3900,n3938);
and (n3900,n3901,n3924);
xor (n3901,n3902,n3914);
nand (n3902,n3903,n3908);
or (n3903,n3754,n3904);
not (n3904,n3905);
nand (n3905,n3906,n3907);
or (n3906,n3651,n3659);
nand (n3907,n3659,n3651);
nand (n3908,n3767,n3909);
nand (n3909,n3910,n3912);
not (n3910,n3911);
and (n3911,n3670,n3659);
nand (n3912,n3658,n3913);
not (n3913,n3670);
nand (n3914,n3915,n3920);
or (n3915,n3916,n3825);
not (n3916,n3917);
nand (n3917,n3918,n3919);
or (n3918,n3626,n3632);
nand (n3919,n3632,n3626);
nand (n3920,n3831,n3921);
nand (n3921,n3922,n3923);
or (n3922,n3643,n3632);
nand (n3923,n3632,n3643);
nand (n3924,n3925,n3931);
or (n3925,n3926,n3654);
not (n3926,n3927);
nand (n3927,n3928,n3930);
or (n3928,n3650,n3929);
nand (n3930,n3929,n3650);
nand (n3931,n3932,n3662);
nand (n3932,n3933,n3936);
not (n3933,n3934);
and (n3934,n3935,n3650);
nand (n3936,n3937,n3649);
not (n3937,n3935);
and (n3938,n3902,n3914);
and (n3939,n3848,n3858);
or (n3940,n3941,n4098);
and (n3941,n3942,n4097);
xor (n3942,n3943,n3990);
or (n3943,n3944,n3989);
and (n3944,n3945,n3962);
xor (n3945,n3946,n3961);
nand (n3946,n3947,n3955);
or (n3947,n3948,n3954);
not (n3948,n3949);
nor (n3949,n3950,n3953);
and (n3950,n3789,n3951);
not (n3951,n3952);
and (n3953,n3952,n3790);
not (n3954,n3794);
or (n3955,n3956,n3780);
not (n3956,n3957);
nand (n3957,n3958,n3960);
or (n3958,n3959,n3789);
nand (n3960,n3959,n3789);
not (n3961,n3848);
or (n3962,n3963,n3988);
and (n3963,n3964,n3980);
xor (n3964,n3965,n3973);
nand (n3965,n3966,n3972);
or (n3966,n3967,n3570);
not (n3967,n3968);
nand (n3968,n3969,n3971);
or (n3969,n3581,n3970);
not (n3970,n3959);
nand (n3971,n3970,n3581);
nand (n3972,n3880,n3725);
nand (n3973,n3974,n3979);
or (n3974,n3975,n3737);
not (n3975,n3976);
nor (n3976,n3977,n3978);
and (n3977,n3735,n3651);
and (n3978,n3733,n3653);
nand (n3979,n3895,n3739);
nand (n3980,n3981,n3986);
or (n3981,n3766,n3982);
nor (n3982,n3983,n3985);
and (n3983,n3984,n3658);
not (n3984,n3929);
and (n3985,n3929,n3659);
or (n3986,n3987,n3754);
not (n3987,n3909);
and (n3988,n3965,n3973);
and (n3989,n3946,n3961);
or (n3990,n3991,n4096);
and (n3991,n3992,n4061);
xor (n3992,n3993,n4012);
or (n3993,n3994,n4005);
nand (n3994,n3995,n4001);
or (n3995,n3996,n3627);
not (n3996,n3997);
nor (n3997,n3998,n4000);
and (n3998,n3999,n3623);
not (n3999,n3723);
and (n4000,n3723,n3624);
nand (n4001,n3629,n4002);
nand (n4002,n4003,n4004);
or (n4003,n3679,n3624);
nand (n4004,n3624,n3679);
nand (n4005,n4006,n4011);
or (n4006,n4007,n3606);
not (n4007,n4008);
nor (n4008,n4009,n4010);
and (n4009,n3643,n3610);
and (n4010,n3641,n3611);
nand (n4011,n3599,n3851);
or (n4012,n4013,n4060);
and (n4013,n4014,n4049);
xor (n4014,n4015,n4039);
nand (n4015,n4016,n4034);
or (n4016,n4017,n4021);
not (n4017,n4018);
nor (n4018,n4019,n4020);
and (n4019,n3704,n3807);
and (n4020,n3703,n3808);
nand (n4021,n4022,n4029);
or (n4022,n4023,n4026);
not (n4023,n4024);
nand (n4024,n3807,n4025);
not (n4026,n4027);
nand (n4027,n3808,n4028);
not (n4028,n4025);
nor (n4029,n4030,n4033);
and (n4030,n4031,n4025);
not (n4031,n4032);
and (n4033,n4032,n4028);
nand (n4034,n4035,n4036);
not (n4035,n4029);
nand (n4036,n4037,n4038);
or (n4037,n3820,n3808);
nand (n4038,n3808,n3820);
nand (n4039,n4040,n4045);
or (n4040,n4041,n3811);
not (n4041,n4042);
nand (n4042,n4043,n4044);
or (n4043,n3518,n3528);
nand (n4044,n3528,n3518);
nand (n4045,n3804,n4046);
nand (n4046,n4047,n4048);
or (n4047,n3537,n3528);
nand (n4048,n3528,n3537);
nand (n4049,n4050,n4055);
or (n4050,n4051,n3682);
not (n4051,n4052);
nand (n4052,n4053,n4054);
or (n4053,n3573,n3791);
or (n4054,n3577,n3586);
nand (n4055,n4056,n3689);
nor (n4056,n4057,n4059);
and (n4057,n4058,n3577);
not (n4058,n3592);
and (n4059,n3592,n3573);
and (n4060,n4015,n4039);
or (n4061,n4062,n4095);
and (n4062,n4063,n4085);
xor (n4063,n4064,n4075);
nand (n4064,n4065,n4070);
or (n4065,n4066,n3523);
not (n4066,n4067);
nand (n4067,n4068,n4069);
or (n4068,n3545,n3519);
nand (n4069,n3519,n3545);
nand (n4070,n4071,n3525);
nand (n4071,n4072,n4074);
not (n4072,n4073);
and (n4073,n3566,n3519);
nand (n4074,n3521,n3565);
nand (n4075,n4076,n4081);
or (n4076,n4077,n3549);
not (n4077,n4078);
nor (n4078,n4079,n4080);
and (n4079,n3762,n3546);
and (n4080,n3763,n3548);
nand (n4081,n3558,n4082);
nor (n4082,n4083,n4084);
and (n4083,n3736,n3546);
and (n4084,n3732,n3548);
nand (n4085,n4086,n4092);
or (n4086,n4087,n4088);
not (n4087,n3869);
not (n4088,n4089);
nand (n4089,n4090,n4091);
or (n4090,n3842,n3603);
nand (n4091,n3603,n3842);
or (n4092,n4093,n4094);
not (n4093,n3863);
not (n4094,n3874);
and (n4095,n4064,n4075);
and (n4096,n3993,n4012);
xor (n4097,n3847,n3899);
and (n4098,n3943,n3990);
and (n4099,n3507,n3714);
xor (n4100,n4101,n4228);
xor (n4101,n4102,n4180);
xor (n4102,n4103,n4177);
xor (n4103,n4104,n4163);
or (n4104,n4105,n4162);
and (n4105,n4106,n4143);
xor (n4106,n4107,n4126);
or (n4107,n4108,n4125);
and (n4108,n4109,n4117);
xor (n4109,n4110,n4113);
nand (n4110,n4111,n4112);
or (n4111,n3887,n3737);
nand (n4112,n3729,n3739);
nand (n4113,n4114,n4115);
or (n4114,n3904,n3766);
nand (n4115,n3772,n4116);
not (n4116,n3754);
nand (n4117,n4118,n4124);
or (n4118,n4119,n3627);
not (n4119,n4120);
nand (n4120,n4121,n4123);
or (n4121,n4122,n3624);
not (n4122,n3695);
nand (n4123,n3624,n4122);
nand (n4124,n3629,n3620);
and (n4125,n4110,n4113);
or (n4126,n4127,n4142);
and (n4127,n4128,n4135);
xor (n4128,n4129,n4132);
nand (n4129,n4130,n4131);
or (n4130,n3956,n3954);
nand (n4131,n3798,n3781);
nand (n4132,n4133,n4134);
or (n4133,n3926,n3663);
nand (n4134,n3667,n3655);
nand (n4135,n4136,n4138);
or (n4136,n4137,n3812);
not (n4137,n3817);
or (n4138,n3811,n4139);
nor (n4139,n4140,n4141);
and (n4140,n3527,n3703);
and (n4141,n3704,n3528);
and (n4142,n4129,n4132);
or (n4143,n4144,n4161);
and (n4144,n4145,n4154);
xor (n4145,n4146,n4150);
nand (n4146,n4147,n4149);
or (n4147,n4148,n3606);
not (n4148,n3855);
nand (n4149,n3613,n3599);
nand (n4150,n4151,n4153);
or (n4151,n4152,n3825);
not (n4152,n3921);
nand (n4153,n3831,n3834);
nand (n4154,n4155,n4160);
or (n4155,n4156,n3682);
not (n4156,n4157);
nand (n4157,n4158,n4159);
or (n4158,n3723,n3577);
nand (n4159,n3577,n3723);
nand (n4160,n3689,n3677);
and (n4161,n4146,n4150);
and (n4162,n4107,n4126);
xor (n4163,n4164,n4174);
xor (n4164,n4165,n4173);
nand (n4165,n4166,n4167);
or (n4166,n3708,n3549);
nand (n4167,n4168,n3558);
not (n4168,n4169);
nor (n4169,n4170,n4172);
and (n4170,n4171,n3548);
not (n4171,n3537);
and (n4172,n3537,n3546);
not (n4173,n3822);
or (n4174,n4175,n4176);
and (n4175,n3673,n3706);
and (n4176,n3674,n3697);
or (n4177,n4178,n4179);
and (n4178,n3508,n3672);
and (n4179,n3509,n3595);
or (n4180,n4181,n4227);
and (n4181,n4182,n4226);
xor (n4182,n4183,n4190);
or (n4183,n4184,n4189);
and (n4184,n4185,n4188);
xor (n4185,n4186,n4187);
xor (n4186,n4145,n4154);
xor (n4187,n4109,n4117);
xor (n4188,n3511,n3568);
and (n4189,n4186,n4187);
or (n4190,n4191,n4225);
and (n4191,n4192,n4224);
xor (n4192,n4193,n4208);
or (n4193,n4194,n4207);
and (n4194,n4195,n4203);
xor (n4195,n4196,n4200);
nand (n4196,n4197,n4199);
or (n4197,n4198,n3627);
not (n4198,n4002);
nand (n4199,n3629,n4120);
nand (n4200,n4201,n4036);
or (n4201,n4035,n4202);
not (n4202,n4021);
nand (n4203,n4204,n4205);
or (n4204,n4139,n3812);
or (n4205,n3811,n4206);
not (n4206,n4046);
and (n4207,n4196,n4200);
or (n4208,n4209,n4223);
and (n4209,n4210,n4219);
xor (n4210,n4211,n4215);
nand (n4211,n4212,n4214);
or (n4212,n4213,n3682);
not (n4213,n4056);
nand (n4214,n4157,n3689);
nand (n4215,n4216,n4218);
or (n4216,n4217,n3523);
not (n4217,n4071);
nand (n4218,n3525,n3515);
nand (n4219,n4220,n4221);
or (n4220,n3541,n3557);
or (n4221,n3549,n4222);
not (n4222,n4082);
and (n4223,n4211,n4215);
xor (n4224,n4128,n4135);
and (n4225,n4193,n4208);
xor (n4226,n4106,n4143);
and (n4227,n4183,n4190);
xor (n4228,n4229,n4313);
xor (n4229,n4230,n4260);
xor (n4230,n4231,n4238);
xor (n4231,n4232,n4235);
or (n4232,n4233,n4234);
and (n4233,n3717,n3752);
and (n4234,n3718,n3726);
or (n4235,n4236,n4237);
and (n4236,n3596,n3644);
and (n4237,n3597,n3617);
xor (n4238,n4239,n4254);
xor (n4239,n4240,n4247);
nand (n4240,n4241,n4242);
nand (n4241,n3738,n3748);
nand (n4242,n3739,n4243);
nand (n4243,n4244,n4246);
not (n4244,n4245);
and (n4245,n3566,n3733);
nand (n4246,n3735,n3565);
nand (n4247,n4248,n4253);
not (n4248,n4249);
nor (n4249,n4250,n3754);
nor (n4250,n4251,n4252);
and (n4251,n3658,n3736);
and (n4252,n3732,n3659);
nand (n4253,n3767,n3760);
nand (n4254,n4255,n4256);
or (n4255,n3786,n3954);
nand (n4256,n4257,n3781);
nor (n4257,n4258,n4259);
and (n4258,n4058,n3789);
and (n4259,n3592,n3790);
xor (n4260,n4261,n4310);
xor (n4261,n4262,n4286);
xor (n4262,n4263,n4279);
xor (n4263,n4264,n4272);
nand (n4264,n4265,n4266);
or (n4265,n3646,n3663);
nand (n4266,n4267,n3655);
nand (n4267,n4268,n4270);
not (n4268,n4269);
and (n4269,n3774,n3650);
nand (n4270,n4271,n3649);
not (n4271,n3774);
nand (n4272,n4273,n4275);
or (n4273,n4274,n3682);
not (n4274,n3693);
nand (n4275,n4276,n3689);
nor (n4276,n4277,n4278);
and (n4277,n3626,n3577);
and (n4278,n3622,n3573);
nand (n4279,n4280,n4282);
or (n4280,n4281,n3523);
not (n4281,n3701);
nand (n4282,n3525,n4283);
nand (n4283,n4284,n4285);
or (n4284,n3820,n3519);
nand (n4285,n3519,n3820);
xor (n4286,n4287,n4303);
xor (n4287,n4288,n4296);
nand (n4288,n4289,n4291);
or (n4289,n4290,n3825);
not (n4290,n3840);
nand (n4291,n3831,n4292);
nand (n4292,n4293,n4295);
or (n4293,n4294,n3632);
not (n4294,n3615);
nand (n4295,n3632,n4294);
nand (n4296,n4297,n4299);
or (n4297,n4298,n3627);
not (n4298,n3639);
nand (n4299,n3629,n4300);
nand (n4300,n4301,n4302);
or (n4301,n3836,n3624);
nand (n4302,n3624,n3836);
nand (n4303,n4304,n4306);
or (n4304,n4305,n3570);
not (n4305,n3721);
nand (n4306,n3725,n4307);
nand (n4307,n4308,n4309);
or (n4308,n3581,n3679);
nand (n4309,n3679,n3581);
or (n4310,n4311,n4312);
and (n4311,n3777,n3822);
and (n4312,n3778,n3802);
or (n4313,n4314,n4315);
and (n4314,n3715,n3845);
and (n4315,n3716,n3776);
or (n4316,n4317,n4508);
and (n4317,n4318,n4358);
xor (n4318,n4319,n4320);
xor (n4319,n4182,n4226);
or (n4320,n4321,n4357);
and (n4321,n4322,n4356);
xor (n4322,n4323,n4324);
xor (n4323,n4192,n4224);
or (n4324,n4325,n4355);
and (n4325,n4326,n4354);
xor (n4326,n4327,n4353);
or (n4327,n4328,n4352);
and (n4328,n4329,n4345);
xor (n4329,n4330,n4337);
nand (n4330,n4331,n4336);
or (n4331,n4332,n3825);
not (n4332,n4333);
nand (n4333,n4334,n4335);
or (n4334,n3695,n3631);
nand (n4335,n3631,n3695);
nand (n4336,n3831,n3917);
nand (n4337,n4338,n4344);
or (n4338,n4339,n3663);
nor (n4339,n4340,n4343);
and (n4340,n4341,n3649);
not (n4341,n4342);
and (n4343,n4342,n3650);
nand (n4344,n3932,n3655);
nand (n4345,n4346,n4347);
or (n4346,n3780,n3948);
nand (n4347,n3794,n4348);
nand (n4348,n4349,n4351);
or (n4349,n4350,n3789);
nand (n4351,n4350,n3789);
and (n4352,n4330,n4337);
xor (n4353,n3901,n3924);
xor (n4354,n4195,n4203);
and (n4355,n4327,n4353);
xor (n4356,n4185,n4188);
and (n4357,n4323,n4324);
or (n4358,n4359,n4507);
and (n4359,n4360,n4506);
xor (n4360,n4361,n4368);
or (n4361,n4362,n4367);
and (n4362,n4363,n4366);
xor (n4363,n4364,n4365);
xor (n4364,n3860,n3885);
xor (n4365,n4210,n4219);
xor (n4366,n3945,n3962);
and (n4367,n4364,n4365);
or (n4368,n4369,n4505);
and (n4369,n4370,n4448);
xor (n4370,n4371,n4447);
or (n4371,n4372,n4446);
and (n4372,n4373,n4418);
xor (n4373,n4374,n4392);
and (n4374,n4375,n4382);
nand (n4375,n4376,n4381);
or (n4376,n4377,n4087);
not (n4377,n4378);
nand (n4378,n4379,n4380);
or (n4379,n3836,n3603);
nand (n4380,n3603,n3836);
nand (n4381,n3863,n4089);
nand (n4382,n4383,n4388);
or (n4383,n4384,n4385);
not (n4385,n4386);
nand (n4386,n4387,n3867);
not (n4387,n4384);
not (n4388,n4389);
nor (n4389,n4390,n4391);
and (n4390,n3873,n3615);
and (n4391,n3867,n4294);
or (n4392,n4393,n4417);
and (n4393,n4394,n4409);
xor (n4394,n4395,n4401);
nand (n4395,n4396,n4397);
or (n4396,n3830,n4332);
nand (n4397,n3830,n4398,n3826);
nor (n4398,n4399,n4400);
and (n4399,n3680,n3632);
and (n4400,n3679,n3631);
nand (n4401,n4402,n4408);
or (n4402,n4403,n3954);
not (n4403,n4404);
nand (n4404,n4405,n4407);
or (n4405,n3789,n4406);
nand (n4407,n4406,n3789);
nand (n4408,n4348,n3781);
nand (n4409,n4410,n4416);
or (n4410,n3663,n4411);
nor (n4411,n4412,n4414);
and (n4412,n3650,n4413);
and (n4414,n3649,n4415);
not (n4415,n4413);
or (n4416,n4339,n3654);
and (n4417,n4395,n4401);
or (n4418,n4419,n4445);
and (n4419,n4420,n4438);
xor (n4420,n4421,n4431);
nand (n4421,n4422,n4427);
or (n4422,n4423,n4424);
not (n4424,n4425);
nand (n4425,n4426,n4032);
not (n4426,n4423);
nand (n4427,n4428,n4429);
or (n4428,n3820,n4032);
not (n4429,n4430);
and (n4430,n3820,n4032);
nand (n4431,n4432,n4437);
or (n4432,n4433,n3627);
not (n4433,n4434);
nand (n4434,n4435,n4436);
or (n4435,n4058,n3624);
nand (n4436,n3624,n4058);
nand (n4437,n3629,n3997);
nand (n4438,n4439,n4440);
or (n4439,n4017,n4029);
or (n4440,n4021,n4441);
not (n4441,n4442);
nor (n4442,n4443,n4444);
and (n4443,n4171,n3808);
and (n4444,n3537,n3807);
and (n4445,n4421,n4431);
and (n4446,n4374,n4392);
xor (n4447,n3992,n4061);
or (n4448,n4449,n4504);
and (n4449,n4450,n4503);
xor (n4450,n4451,n4478);
or (n4451,n4452,n4477);
and (n4452,n4453,n4469);
xor (n4453,n4454,n4462);
nand (n4454,n4455,n4461);
or (n4455,n4456,n3811);
not (n4456,n4457);
nand (n4457,n4458,n4460);
not (n4458,n4459);
and (n4459,n3566,n3528);
nand (n4460,n3527,n3565);
nand (n4461,n3804,n4042);
nand (n4462,n4463,n4468);
or (n4463,n4464,n3606);
not (n4464,n4465);
nand (n4465,n4466,n4467);
or (n4466,n3626,n3611);
nand (n4467,n3611,n3626);
nand (n4468,n3599,n4008);
nand (n4469,n4470,n4472);
or (n4470,n4471,n4051);
not (n4471,n3689);
or (n4472,n3682,n4473);
not (n4473,n4474);
nand (n4474,n4475,n4476);
or (n4475,n3573,n3882);
or (n4476,n3577,n3800);
and (n4477,n4454,n4462);
or (n4478,n4479,n4502);
and (n4479,n4480,n4495);
xor (n4480,n4481,n4488);
nand (n4481,n4482,n4487);
or (n4482,n4483,n3523);
not (n4483,n4484);
nor (n4484,n4485,n4486);
and (n4485,n3736,n3519);
and (n4486,n3732,n3521);
nand (n4487,n3525,n4067);
nand (n4488,n4489,n4494);
or (n4489,n4490,n3549);
not (n4490,n4491);
nor (n4491,n4492,n4493);
and (n4492,n4271,n3546);
and (n4493,n3774,n3548);
nand (n4494,n3558,n4078);
nand (n4495,n4496,n4497);
or (n4496,n3967,n3571);
nand (n4497,n4498,n4499);
not (n4498,n3570);
nor (n4499,n4500,n4501);
and (n4500,n3951,n3580);
and (n4501,n3952,n3581);
and (n4502,n4481,n4488);
xor (n4503,n4014,n4049);
and (n4504,n4451,n4478);
and (n4505,n4371,n4447);
xor (n4506,n3942,n4097);
and (n4507,n4361,n4368);
and (n4508,n4319,n4320);
and (n4509,n3504,n4100);
not (n4510,n4511);
xor (n4511,n4512,n4617);
xor (n4512,n4513,n4581);
xor (n4513,n4514,n4529);
xor (n4514,n4515,n4526);
xor (n4515,n4516,n4523);
xor (n4516,n4517,n4520);
nor (n4517,n4518,n4519);
and (n4518,n3825,n3830);
not (n4519,n4292);
or (n4520,n4521,n4522);
and (n4521,n4287,n4303);
and (n4522,n4288,n4296);
or (n4523,n4524,n4525);
and (n4524,n4239,n4254);
and (n4525,n4240,n4247);
or (n4526,n4527,n4528);
and (n4527,n4261,n4310);
and (n4528,n4262,n4286);
xor (n4529,n4530,n4557);
xor (n4530,n4531,n4534);
or (n4531,n4532,n4533);
and (n4532,n4263,n4279);
and (n4533,n4264,n4272);
xor (n4534,n4535,n4551);
xor (n4535,n4536,n4543);
nand (n4536,n4537,n4539);
or (n4537,n4538,n3570);
not (n4538,n4307);
nand (n4539,n4540,n3725);
nor (n4540,n4541,n4542);
and (n4541,n4122,n3580);
and (n4542,n3695,n3581);
nand (n4543,n4544,n4546);
or (n4544,n4545,n3737);
not (n4545,n4243);
nand (n4546,n3739,n4547);
nand (n4547,n4548,n4550);
not (n4548,n4549);
and (n4549,n3518,n3733);
nand (n4550,n3735,n3522);
nand (n4551,n4552,n4556);
or (n4552,n3754,n4553);
nor (n4553,n4554,n4555);
and (n4554,n3658,n3544);
and (n4555,n3545,n3659);
or (n4556,n3766,n4250);
xor (n4557,n4558,n4574);
xor (n4558,n4559,n4566);
nand (n4559,n4560,n4562);
or (n4560,n4561,n3627);
not (n4561,n4300);
nand (n4562,n3629,n4563);
nand (n4563,n4564,n4565);
or (n4564,n3842,n3624);
nand (n4565,n3624,n3842);
nand (n4566,n4567,n4569);
or (n4567,n4568,n3663);
not (n4568,n4267);
nand (n4569,n4570,n3655);
nand (n4570,n4571,n4573);
not (n4571,n4572);
and (n4572,n3763,n3650);
or (n4573,n3763,n3650);
nand (n4574,n4575,n4577);
or (n4575,n3954,n4576);
not (n4576,n4257);
or (n4577,n4578,n3780);
nor (n4578,n4579,n4580);
and (n4579,n3789,n3723);
and (n4580,n3790,n3999);
xor (n4581,n4582,n4614);
xor (n4582,n4583,n4611);
xor (n4583,n4584,n4608);
xor (n4584,n4585,n4605);
xor (n4585,n4586,n4597);
xor (n4586,n4587,n4594);
nand (n4587,n4588,n4590);
or (n4588,n4589,n3682);
not (n4589,n4276);
nand (n4590,n3689,n4591);
nor (n4591,n4592,n4593);
and (n4592,n3643,n3577);
and (n4593,n3641,n3573);
nand (n4594,n4595,n4283);
or (n4595,n3525,n4596);
not (n4596,n3523);
nand (n4597,n4598,n4604);
or (n4598,n4599,n3557);
not (n4599,n4600);
nand (n4600,n4601,n4602);
or (n4601,n3546,n3704);
not (n4602,n4603);
and (n4603,n3704,n3546);
or (n4604,n3549,n4169);
or (n4605,n4606,n4607);
and (n4606,n4164,n4174);
and (n4607,n4165,n4173);
or (n4608,n4609,n4610);
and (n4609,n4231,n4238);
and (n4610,n4232,n4235);
or (n4611,n4612,n4613);
and (n4612,n4103,n4177);
and (n4613,n4104,n4163);
or (n4614,n4615,n4616);
and (n4615,n4229,n4313);
and (n4616,n4230,n4260);
or (n4617,n4618,n4619);
and (n4618,n4101,n4228);
and (n4619,n4102,n4180);
nor (n4620,n4621,n4718);
xor (n4621,n4622,n4715);
xor (n4622,n4623,n4642);
xor (n4623,n4624,n4631);
xor (n4624,n4625,n4628);
or (n4625,n4626,n4627);
and (n4626,n4516,n4523);
and (n4627,n4517,n4520);
or (n4628,n4629,n4630);
and (n4629,n4530,n4557);
and (n4630,n4531,n4534);
xor (n4631,n4632,n4639);
xor (n4632,n4633,n4636);
or (n4633,n4634,n4635);
and (n4634,n4535,n4551);
and (n4635,n4536,n4543);
or (n4636,n4637,n4638);
and (n4637,n4558,n4574);
and (n4638,n4559,n4566);
or (n4639,n4640,n4641);
and (n4640,n4586,n4597);
and (n4641,n4587,n4594);
xor (n4642,n4643,n4712);
xor (n4643,n4644,n4709);
xor (n4644,n4645,n4692);
xor (n4645,n4646,n4668);
xor (n4646,n4647,n4662);
xor (n4647,n4648,n4655);
nand (n4648,n4649,n4651);
or (n4649,n4650,n3627);
not (n4650,n4563);
nand (n4651,n3629,n4652);
nand (n4652,n4653,n4654);
or (n4653,n4294,n3624);
nand (n4654,n3624,n4294);
nand (n4655,n4656,n4658);
or (n4656,n4657,n3682);
not (n4657,n4591);
nand (n4658,n3689,n4659);
nor (n4659,n4660,n4661);
and (n4660,n3836,n3577);
and (n4661,n3837,n3573);
nand (n4662,n4663,n4664);
or (n4663,n3954,n4578);
or (n4664,n4665,n3780);
nor (n4665,n4666,n4667);
and (n4666,n3679,n3790);
and (n4667,n3789,n3680);
xor (n4668,n4669,n4684);
xor (n4669,n4670,n4677);
nand (n4670,n4671,n4673);
or (n4671,n4672,n3663);
not (n4672,n4570);
nand (n4673,n4674,n3655);
nand (n4674,n4675,n4676);
or (n4675,n3650,n3732);
nand (n4676,n3732,n3650);
nand (n4677,n4678,n4679);
or (n4678,n4599,n3549);
nand (n4679,n3558,n4680);
nor (n4680,n4681,n4683);
and (n4681,n4682,n3546);
not (n4682,n3820);
and (n4683,n3820,n3548);
nand (n4684,n4685,n4690);
or (n4685,n4686,n3571);
not (n4686,n4687);
nand (n4687,n4688,n4689);
or (n4688,n3581,n3626);
or (n4689,n3580,n3622);
or (n4690,n3570,n4691);
not (n4691,n4540);
xor (n4692,n4693,n4708);
xor (n4693,n4694,n4702);
nand (n4694,n4695,n4697);
or (n4695,n4696,n3737);
not (n4696,n4547);
nand (n4697,n4698,n3739);
not (n4698,n4699);
nor (n4699,n4700,n4701);
and (n4700,n3735,n4171);
and (n4701,n3537,n3733);
nand (n4702,n4703,n4704);
or (n4703,n3766,n4553);
or (n4704,n4705,n3754);
nor (n4705,n4706,n4707);
and (n4706,n3658,n3565);
and (n4707,n3566,n3659);
not (n4708,n4517);
or (n4709,n4710,n4711);
and (n4710,n4584,n4608);
and (n4711,n4585,n4605);
or (n4712,n4713,n4714);
and (n4713,n4514,n4529);
and (n4714,n4515,n4526);
or (n4715,n4716,n4717);
and (n4716,n4582,n4614);
and (n4717,n4583,n4611);
or (n4718,n4719,n4720);
and (n4719,n4512,n4617);
and (n4720,n4513,n4581);
nor (n4721,n4722,n4984);
nand (n4722,n4723,n4808);
or (n4723,n4724,n4727);
or (n4724,n4725,n4726);
and (n4725,n4622,n4715);
and (n4726,n4623,n4642);
xor (n4727,n4728,n4805);
xor (n4728,n4729,n4732);
or (n4729,n4730,n4731);
and (n4730,n4624,n4631);
and (n4731,n4625,n4628);
xor (n4732,n4733,n4784);
xor (n4733,n4734,n4781);
xor (n4734,n4735,n4763);
xor (n4735,n4736,n4739);
or (n4736,n4737,n4738);
and (n4737,n4669,n4684);
and (n4738,n4670,n4677);
xor (n4739,n4740,n4757);
xor (n4740,n4741,n4749);
nand (n4741,n4742,n4744);
or (n4742,n4743,n3682);
not (n4743,n4659);
nand (n4744,n4745,n3689);
not (n4745,n4746);
nor (n4746,n4747,n4748);
and (n4747,n3842,n3573);
and (n4748,n3843,n3577);
nand (n4749,n4750,n4752);
or (n4750,n4751,n3663);
not (n4751,n4674);
nand (n4752,n4753,n3655);
not (n4753,n4754);
nor (n4754,n4755,n4756);
and (n4755,n3649,n3544);
and (n4756,n3545,n3650);
nand (n4757,n4758,n4759);
or (n4758,n3954,n4665);
or (n4759,n4760,n3780);
nor (n4760,n4761,n4762);
and (n4761,n3789,n3695);
and (n4762,n3790,n4122);
xor (n4763,n4764,n4775);
xor (n4764,n4765,n4768);
nand (n4765,n4766,n4680);
or (n4766,n3558,n4767);
not (n4767,n3549);
nand (n4768,n4769,n4770);
or (n4769,n4686,n3570);
nand (n4770,n4771,n3725);
not (n4771,n4772);
nor (n4772,n4773,n4774);
and (n4773,n3580,n3641);
and (n4774,n3581,n3643);
nand (n4775,n4776,n4777);
or (n4776,n3737,n4699);
or (n4777,n3892,n4778);
nor (n4778,n4779,n4780);
and (n4779,n3735,n3703);
and (n4780,n3704,n3733);
or (n4781,n4782,n4783);
and (n4782,n4645,n4692);
and (n4783,n4646,n4668);
xor (n4784,n4785,n4802);
xor (n4785,n4786,n4789);
or (n4786,n4787,n4788);
and (n4787,n4693,n4708);
and (n4788,n4694,n4702);
xor (n4789,n4790,n4799);
xor (n4790,n4791,n4797);
nand (n4791,n4792,n4793);
or (n4792,n3766,n4705);
or (n4793,n4794,n3754);
nor (n4794,n4795,n4796);
and (n4795,n3658,n3522);
and (n4796,n3518,n3659);
and (n4797,n4798,n4652);
nand (n4798,n3627,n3628);
or (n4799,n4800,n4801);
and (n4800,n4647,n4662);
and (n4801,n4648,n4655);
or (n4802,n4803,n4804);
and (n4803,n4632,n4639);
and (n4804,n4633,n4636);
or (n4805,n4806,n4807);
and (n4806,n4643,n4712);
and (n4807,n4644,n4709);
nor (n4808,n4809,n4936);
nor (n4809,n4810,n4880);
or (n4810,n4811,n4879);
and (n4811,n4812,n4876);
xor (n4812,n4813,n4859);
xor (n4813,n4814,n4856);
xor (n4814,n4815,n4835);
xor (n4815,n4816,n4829);
xor (n4816,n4817,n4823);
nand (n4817,n4818,n4819);
or (n4818,n4794,n3766);
nand (n4819,n4820,n4116);
nor (n4820,n4821,n4822);
and (n4821,n3537,n3658);
and (n4822,n4171,n3659);
nand (n4823,n4824,n4825);
or (n4824,n3954,n4760);
or (n4825,n4826,n3780);
nor (n4826,n4827,n4828);
and (n4827,n3789,n3622);
and (n4828,n3790,n3626);
nand (n4829,n4830,n4831);
or (n4830,n3663,n4754);
or (n4831,n3654,n4832);
nor (n4832,n4833,n4834);
and (n4833,n3649,n3565);
and (n4834,n3566,n3650);
xor (n4835,n4836,n4850);
xor (n4836,n4837,n4844);
nand (n4837,n4838,n4843);
or (n4838,n4839,n4471);
not (n4839,n4840);
nand (n4840,n4841,n4842);
or (n4841,n3573,n4294);
or (n4842,n3577,n3615);
nand (n4843,n4745,n3683);
nand (n4844,n4845,n4846);
or (n4845,n3570,n4772);
or (n4846,n3571,n4847);
nor (n4847,n4848,n4849);
and (n4848,n3580,n3837);
and (n4849,n3581,n3836);
nand (n4850,n4851,n4852);
or (n4851,n3737,n4778);
or (n4852,n3892,n4853);
nor (n4853,n4854,n4855);
and (n4854,n3735,n4682);
and (n4855,n3820,n3733);
or (n4856,n4857,n4858);
and (n4857,n4790,n4799);
and (n4858,n4791,n4797);
xor (n4859,n4860,n4873);
xor (n4860,n4861,n4870);
xor (n4861,n4862,n4867);
xor (n4862,n4863,n4864);
not (n4863,n4797);
or (n4864,n4865,n4866);
and (n4865,n4740,n4757);
and (n4866,n4741,n4749);
or (n4867,n4868,n4869);
and (n4868,n4764,n4775);
and (n4869,n4765,n4768);
or (n4870,n4871,n4872);
and (n4871,n4735,n4763);
and (n4872,n4736,n4739);
or (n4873,n4874,n4875);
and (n4874,n4785,n4802);
and (n4875,n4786,n4789);
or (n4876,n4877,n4878);
and (n4877,n4733,n4784);
and (n4878,n4734,n4781);
and (n4879,n4813,n4859);
xor (n4880,n4881,n4933);
xor (n4881,n4882,n4885);
or (n4882,n4883,n4884);
and (n4883,n4814,n4856);
and (n4884,n4815,n4835);
xor (n4885,n4886,n4911);
xor (n4886,n4887,n4908);
xor (n4887,n4888,n4901);
xor (n4888,n4889,n4895);
nand (n4889,n4890,n4891);
or (n4890,n3663,n4832);
or (n4891,n3654,n4892);
nor (n4892,n4893,n4894);
and (n4893,n3649,n3522);
and (n4894,n3518,n3650);
nand (n4895,n4896,n4897);
or (n4896,n3954,n4826);
or (n4897,n4898,n3780);
nor (n4898,n4899,n4900);
and (n4899,n3789,n3641);
and (n4900,n3790,n3643);
not (n4901,n4902);
nand (n4902,n4903,n4904);
or (n4903,n3570,n4847);
or (n4904,n3571,n4905);
nor (n4905,n4906,n4907);
and (n4906,n3580,n3843);
and (n4907,n3581,n3842);
or (n4908,n4909,n4910);
and (n4909,n4862,n4867);
and (n4910,n4863,n4864);
xor (n4911,n4912,n4919);
xor (n4912,n4913,n4916);
or (n4913,n4914,n4915);
and (n4914,n4816,n4829);
and (n4915,n4817,n4823);
or (n4916,n4917,n4918);
and (n4917,n4836,n4850);
and (n4918,n4837,n4844);
xor (n4919,n4920,n4931);
xor (n4920,n4921,n4924);
nand (n4921,n4922,n4923);
or (n4922,n3739,n3738);
not (n4923,n4853);
nand (n4924,n4925,n4927);
or (n4925,n3766,n4926);
not (n4926,n4820);
or (n4927,n4928,n3754);
nor (n4928,n4929,n4930);
and (n4929,n3658,n3703);
and (n4930,n3704,n3659);
nand (n4931,n4932,n4840);
or (n4932,n3683,n3689);
or (n4933,n4934,n4935);
and (n4934,n4860,n4873);
and (n4935,n4861,n4870);
nor (n4936,n4937,n4940);
or (n4937,n4938,n4939);
and (n4938,n4881,n4933);
and (n4939,n4882,n4885);
xor (n4940,n4941,n4981);
xor (n4941,n4942,n4945);
or (n4942,n4943,n4944);
and (n4943,n4912,n4919);
and (n4944,n4913,n4916);
xor (n4945,n4946,n4970);
xor (n4946,n4947,n4967);
xor (n4947,n4948,n4961);
xor (n4948,n4949,n4955);
nand (n4949,n4950,n4951);
or (n4950,n3570,n4905);
or (n4951,n3571,n4952);
nor (n4952,n4953,n4954);
and (n4953,n3580,n3615);
and (n4954,n3581,n4294);
nand (n4955,n4956,n4957);
or (n4956,n3954,n4898);
or (n4957,n4958,n3780);
nor (n4958,n4959,n4960);
and (n4959,n3837,n3789);
and (n4960,n3836,n3790);
nand (n4961,n4962,n4963);
or (n4962,n3663,n4892);
or (n4963,n3654,n4964);
nor (n4964,n4965,n4966);
and (n4965,n3649,n4171);
and (n4966,n3537,n3650);
or (n4967,n4968,n4969);
and (n4968,n4888,n4901);
and (n4969,n4889,n4895);
xor (n4970,n4971,n4978);
xor (n4971,n4972,n4902);
nand (n4972,n4973,n4974);
or (n4973,n3766,n4928);
or (n4974,n4975,n3754);
nor (n4975,n4976,n4977);
and (n4976,n3658,n4682);
and (n4977,n3820,n3659);
or (n4978,n4979,n4980);
and (n4979,n4920,n4931);
and (n4980,n4921,n4924);
or (n4981,n4982,n4983);
and (n4982,n4886,n4911);
and (n4983,n4887,n4908);
nand (n4984,n4985,n4992);
nand (n4985,n4986,n4988);
not (n4986,n4987);
xor (n4987,n4812,n4876);
not (n4988,n4989);
or (n4989,n4990,n4991);
and (n4990,n4728,n4805);
and (n4991,n4729,n4732);
nor (n4992,n4993,n5029);
nor (n4993,n4994,n4997);
or (n4994,n4995,n4996);
and (n4995,n4941,n4981);
and (n4996,n4942,n4945);
xor (n4997,n4998,n5026);
xor (n4998,n4999,n5002);
or (n4999,n5000,n5001);
and (n5000,n4971,n4978);
and (n5001,n4972,n4902);
xor (n5002,n5003,n5009);
xor (n5003,n5004,n5006);
nor (n5004,n5005,n4952);
and (n5005,n3570,n3571);
or (n5006,n5007,n5008);
and (n5007,n4948,n4961);
and (n5008,n4949,n4955);
xor (n5009,n5010,n5023);
xor (n5010,n5011,n5017);
nand (n5011,n5012,n5013);
or (n5012,n3663,n4964);
or (n5013,n3654,n5014);
nor (n5014,n5015,n5016);
and (n5015,n3649,n3703);
and (n5016,n3704,n3650);
nand (n5017,n5018,n5019);
or (n5018,n3954,n4958);
or (n5019,n5020,n3780);
nor (n5020,n5021,n5022);
and (n5021,n3789,n3843);
and (n5022,n3790,n3842);
nand (n5023,n5024,n5025);
or (n5024,n4116,n3767);
not (n5025,n4975);
or (n5026,n5027,n5028);
and (n5027,n4946,n4970);
and (n5028,n4947,n4967);
nand (n5029,n5030,n5058);
or (n5030,n5031,n5055);
xor (n5031,n5032,n5052);
xor (n5032,n5033,n5036);
or (n5033,n5034,n5035);
and (n5034,n5010,n5023);
and (n5035,n5011,n5017);
xor (n5036,n5037,n5051);
xor (n5037,n5038,n5045);
nand (n5038,n5039,n5044);
or (n5039,n3780,n5040);
not (n5040,n5041);
nand (n5041,n5042,n5043);
or (n5042,n3790,n4294);
or (n5043,n3789,n3615);
or (n5044,n3954,n5020);
nand (n5045,n5046,n5047);
or (n5046,n3663,n5014);
or (n5047,n3654,n5048);
nor (n5048,n5049,n5050);
and (n5049,n3649,n4682);
and (n5050,n3820,n3650);
not (n5051,n5004);
or (n5052,n5053,n5054);
and (n5053,n5003,n5009);
and (n5054,n5004,n5006);
or (n5055,n5056,n5057);
and (n5056,n4998,n5026);
and (n5057,n4999,n5002);
nand (n5058,n5059,n5063);
not (n5059,n5060);
or (n5060,n5061,n5062);
and (n5061,n5032,n5052);
and (n5062,n5033,n5036);
not (n5063,n5064);
xor (n5064,n5065,n5070);
xor (n5065,n5066,n5068);
nand (n5066,n5067,n5041);
or (n5067,n3794,n3781);
nor (n5068,n5069,n5048);
and (n5069,n3663,n3654);
or (n5070,n5071,n5072);
and (n5071,n5037,n5051);
and (n5072,n5038,n5045);
nor (n5073,n5074,n5210);
nor (n5074,n5075,n5209);
or (n5075,n5076,n5208);
and (n5076,n5077,n5080);
xor (n5077,n5078,n5079);
xor (n5078,n3506,n3940);
xor (n5079,n4318,n4358);
or (n5080,n5081,n5207);
and (n5081,n5082,n5206);
xor (n5082,n5083,n5084);
xor (n5083,n4322,n4356);
or (n5084,n5085,n5205);
and (n5085,n5086,n5098);
xor (n5086,n5087,n5097);
or (n5087,n5088,n5096);
and (n5088,n5089,n5095);
xor (n5089,n5090,n5091);
xor (n5090,n4329,n4345);
nand (n5091,n5092,n3993);
or (n5092,n5093,n5094);
not (n5093,n4005);
not (n5094,n3994);
xor (n5095,n3964,n3980);
and (n5096,n5090,n5091);
xor (n5097,n4326,n4354);
or (n5098,n5099,n5204);
and (n5099,n5100,n5124);
xor (n5100,n5101,n5102);
xor (n5101,n4063,n4085);
or (n5102,n5103,n5123);
and (n5103,n5104,n5119);
xor (n5104,n5105,n5111);
nand (n5105,n5106,n5110);
or (n5106,n3737,n5107);
nor (n5107,n5108,n5109);
and (n5108,n3735,n3913);
and (n5109,n3733,n3670);
or (n5110,n3892,n3975);
nand (n5111,n5112,n5118);
or (n5112,n3766,n5113);
not (n5113,n5114);
nand (n5114,n5115,n5116);
or (n5115,n3659,n3935);
not (n5116,n5117);
and (n5117,n3935,n3659);
or (n5118,n3982,n3754);
nand (n5119,n5120,n5122);
or (n5120,n4382,n5121);
not (n5121,n4375);
nand (n5122,n5121,n4382);
and (n5123,n5105,n5111);
or (n5124,n5125,n5203);
and (n5125,n5126,n5178);
xor (n5126,n5127,n5154);
or (n5127,n5128,n5153);
and (n5128,n5129,n5145);
xor (n5129,n5130,n5137);
nand (n5130,n5131,n5136);
or (n5131,n5132,n3627);
not (n5132,n5133);
nand (n5133,n5134,n5135);
or (n5134,n3791,n3624);
nand (n5135,n3624,n3791);
nand (n5136,n3629,n4434);
nand (n5137,n5138,n5144);
or (n5138,n4425,n5139);
not (n5139,n5140);
nand (n5140,n5141,n5142);
or (n5141,n3704,n4032);
not (n5142,n5143);
and (n5143,n3704,n4032);
nand (n5144,n4427,n4423);
nand (n5145,n5146,n5147);
or (n5146,n4441,n4029);
or (n5147,n4021,n5148);
not (n5148,n5149);
nand (n5149,n5150,n5151);
or (n5150,n3518,n3808);
not (n5151,n5152);
and (n5152,n3518,n3808);
and (n5153,n5130,n5137);
or (n5154,n5155,n5177);
and (n5155,n5156,n5171);
xor (n5156,n5157,n5164);
nand (n5157,n5158,n5163);
or (n5158,n5159,n3606);
not (n5159,n5160);
nand (n5160,n5161,n5162);
or (n5161,n3695,n3610);
or (n5162,n3611,n4122);
nand (n5163,n3599,n4465);
nand (n5164,n5165,n5170);
or (n5165,n5166,n3682);
not (n5166,n5167);
nor (n5167,n5168,n5169);
and (n5168,n3577,n3970);
and (n5169,n3573,n3959);
nand (n5170,n4474,n3689);
nand (n5171,n5172,n5173);
or (n5172,n4456,n3812);
or (n5173,n3811,n5174);
nor (n5174,n5175,n5176);
and (n5175,n3527,n3544);
and (n5176,n3528,n3545);
and (n5177,n5157,n5164);
or (n5178,n5179,n5202);
and (n5179,n5180,n5196);
xor (n5180,n5181,n5188);
nand (n5181,n5182,n5187);
or (n5182,n5183,n3523);
not (n5183,n5184);
nor (n5184,n5185,n5186);
and (n5185,n3763,n3521);
and (n5186,n3762,n3519);
nand (n5187,n3525,n4484);
nand (n5188,n5189,n5195);
or (n5189,n5190,n3570);
not (n5190,n5191);
nand (n5191,n5192,n5194);
or (n5192,n3581,n5193);
not (n5193,n4350);
nand (n5194,n5193,n3581);
nand (n5195,n4499,n3725);
nand (n5196,n5197,n5201);
or (n5197,n5198,n3549);
nor (n5198,n5199,n5200);
and (n5199,n3548,n3653);
and (n5200,n3546,n3651);
nand (n5201,n3558,n4491);
and (n5202,n5181,n5188);
and (n5203,n5127,n5154);
and (n5204,n5101,n5102);
and (n5205,n5087,n5097);
xor (n5206,n4360,n4506);
and (n5207,n5083,n5084);
and (n5208,n5078,n5079);
xor (n5209,n3503,n4316);
nor (n5210,n5211,n5212);
xor (n5211,n5077,n5080);
or (n5212,n5213,n5321);
and (n5213,n5214,n5302);
xor (n5214,n5215,n5301);
or (n5215,n5216,n5300);
and (n5216,n5217,n5299);
xor (n5217,n5218,n5219);
xor (n5218,n4363,n4366);
or (n5219,n5220,n5298);
and (n5220,n5221,n5297);
xor (n5221,n5222,n5296);
or (n5222,n5223,n5295);
and (n5223,n5224,n5274);
xor (n5224,n5225,n5250);
or (n5225,n5226,n5249);
and (n5226,n5227,n5243);
xor (n5227,n5228,n5236);
nor (n5228,n5229,n3789);
and (n5229,n5230,n5234);
nand (n5230,n5231,n3580);
not (n5231,n5232);
and (n5232,n5233,n3783);
nand (n5234,n5235,n3785);
not (n5235,n5233);
nor (n5236,n5237,n3650);
and (n5237,n5238,n5242);
nand (n5238,n5239,n3659);
or (n5239,n3657,n5240);
not (n5240,n5241);
nand (n5242,n3657,n5240);
nand (n5243,n5244,n5248);
or (n5244,n4386,n5245);
nor (n5245,n5246,n5247);
and (n5246,n3873,n3843);
and (n5247,n3867,n3842);
or (n5248,n4389,n4387);
and (n5249,n5228,n5236);
or (n5250,n5251,n5273);
and (n5251,n5252,n5267);
xor (n5252,n5253,n5259);
nand (n5253,n5254,n5255);
or (n5254,n3780,n4403);
or (n5255,n3954,n5256);
nor (n5256,n5257,n5258);
and (n5257,n5235,n3790);
and (n5258,n5233,n3789);
nand (n5259,n5260,n5266);
or (n5260,n3766,n5261);
not (n5261,n5262);
nand (n5262,n5263,n5265);
not (n5263,n5264);
and (n5264,n4342,n3659);
nand (n5265,n3658,n4341);
nand (n5266,n5114,n4116);
nand (n5267,n5268,n5272);
or (n5268,n3663,n5269);
nor (n5269,n5270,n5271);
and (n5270,n5241,n3650);
and (n5271,n3649,n5240);
or (n5272,n3654,n4411);
and (n5273,n5253,n5259);
or (n5274,n5275,n5294);
and (n5275,n5276,n5291);
xor (n5276,n5277,n5284);
nand (n5277,n5278,n5283);
or (n5278,n5279,n4087);
not (n5279,n5280);
nand (n5280,n5281,n5282);
or (n5281,n3643,n3603);
nand (n5282,n3603,n3643);
nand (n5283,n4378,n3863);
nand (n5284,n5285,n5290);
or (n5285,n3825,n5286);
not (n5286,n5287);
nand (n5287,n5288,n5289);
or (n5288,n3723,n3631);
nand (n5289,n3631,n3723);
nand (n5290,n3831,n4398);
nor (n5291,n5292,n5293);
nand (n5292,n3781,n5233);
nand (n5293,n3655,n5241);
and (n5294,n5277,n5284);
and (n5295,n5225,n5250);
xor (n5296,n4373,n4418);
xor (n5297,n4450,n4503);
and (n5298,n5222,n5296);
xor (n5299,n4370,n4448);
and (n5300,n5218,n5219);
xor (n5301,n5082,n5206);
or (n5302,n5303,n5320);
and (n5303,n5304,n5319);
xor (n5304,n5305,n5306);
xor (n5305,n5086,n5098);
or (n5306,n5307,n5318);
and (n5307,n5308,n5317);
xor (n5308,n5309,n5316);
or (n5309,n5310,n5315);
and (n5310,n5311,n5314);
xor (n5311,n5312,n5313);
xor (n5312,n4480,n4495);
xor (n5313,n4420,n4438);
xor (n5314,n4453,n4469);
and (n5315,n5312,n5313);
xor (n5316,n5089,n5095);
xor (n5317,n5100,n5124);
and (n5318,n5309,n5316);
xor (n5319,n5217,n5299);
and (n5320,n5305,n5306);
and (n5321,n5215,n5301);
nor (n5322,n5323,n5820);
not (n5323,n5324);
nor (n5324,n5325,n5651);
nor (n5325,n5326,n5327);
xor (n5326,n5214,n5302);
or (n5327,n5328,n5650);
and (n5328,n5329,n5506);
xor (n5329,n5330,n5505);
or (n5330,n5331,n5504);
and (n5331,n5332,n5467);
xor (n5332,n5333,n5421);
or (n5333,n5334,n5420);
and (n5334,n5335,n5338);
xor (n5335,n5336,n5337);
xor (n5336,n4394,n4409);
xor (n5337,n5104,n5119);
or (n5338,n5339,n5419);
and (n5339,n5340,n5393);
xor (n5340,n5341,n5367);
or (n5341,n5342,n5366);
and (n5342,n5343,n5359);
xor (n5343,n5344,n5351);
nand (n5344,n5345,n5350);
or (n5345,n5346,n3825);
not (n5346,n5347);
nand (n5347,n5348,n5349);
or (n5348,n3592,n3631);
nand (n5349,n3631,n3592);
nand (n5350,n5287,n3831);
nand (n5351,n5352,n5358);
or (n5352,n4425,n5353);
not (n5353,n5354);
nand (n5354,n5355,n5356);
or (n5355,n3537,n4032);
not (n5356,n5357);
and (n5357,n3537,n4032);
nand (n5358,n5140,n4423);
nand (n5359,n5360,n5365);
or (n5360,n5361,n3627);
not (n5361,n5362);
nor (n5362,n5363,n5364);
and (n5363,n3882,n3623);
and (n5364,n3800,n3624);
nand (n5365,n3629,n5133);
and (n5366,n5344,n5351);
or (n5367,n5368,n5392);
and (n5368,n5369,n5385);
xor (n5369,n5370,n5377);
nand (n5370,n5371,n5376);
or (n5371,n5372,n4021);
not (n5372,n5373);
nor (n5373,n5374,n5375);
and (n5374,n3566,n3807);
and (n5375,n3565,n3808);
nand (n5376,n4035,n5149);
nand (n5377,n5378,n5383);
or (n5378,n5379,n3811);
not (n5379,n5380);
nor (n5380,n5381,n5382);
and (n5381,n3736,n3528);
and (n5382,n3732,n3527);
nand (n5383,n5384,n3804);
not (n5384,n5174);
nand (n5385,n5386,n5387);
or (n5386,n5159,n3607);
or (n5387,n3606,n5388);
not (n5388,n5389);
nand (n5389,n5390,n5391);
or (n5390,n3611,n3679);
nand (n5391,n3611,n3679);
and (n5392,n5370,n5377);
or (n5393,n5394,n5418);
and (n5394,n5395,n5410);
xor (n5395,n5396,n5403);
nand (n5396,n5397,n5402);
or (n5397,n5398,n3682);
not (n5398,n5399);
nor (n5399,n5400,n5401);
and (n5400,n3951,n3577);
and (n5401,n3952,n3573);
nand (n5402,n5167,n3689);
nand (n5403,n5404,n5405);
or (n5404,n5183,n3524);
nand (n5405,n5406,n4596);
nand (n5406,n5407,n5409);
not (n5407,n5408);
and (n5408,n3774,n3519);
nand (n5409,n3521,n4271);
nand (n5410,n5411,n5417);
or (n5411,n3549,n5412);
not (n5412,n5413);
nand (n5413,n5414,n5416);
not (n5414,n5415);
and (n5415,n3670,n3546);
nand (n5416,n3548,n3913);
or (n5417,n3557,n5198);
and (n5418,n5396,n5403);
and (n5419,n5341,n5367);
and (n5420,n5336,n5337);
or (n5421,n5422,n5466);
and (n5422,n5423,n5465);
xor (n5423,n5424,n5458);
or (n5424,n5425,n5457);
and (n5425,n5426,n5435);
xor (n5426,n5427,n5434);
nand (n5427,n5428,n5433);
or (n5428,n3737,n5429);
not (n5429,n5430);
nor (n5430,n5431,n5432);
and (n5431,n3984,n3733);
and (n5432,n3929,n3735);
or (n5433,n3892,n5107);
xor (n5434,n5227,n5243);
or (n5435,n5436,n5456);
and (n5436,n5437,n5450);
xor (n5437,n5438,n5446);
nand (n5438,n5439,n5444);
or (n5439,n4386,n5440);
not (n5440,n5441);
nand (n5441,n5442,n5443);
or (n5442,n3837,n3873);
nand (n5443,n3873,n3837);
nand (n5444,n5445,n4384);
not (n5445,n5245);
nand (n5446,n5447,n5449);
or (n5447,n5448,n5292);
not (n5448,n5293);
nand (n5449,n5448,n5292);
nand (n5450,n5451,n5455);
nand (n5451,n3869,n5452);
nand (n5452,n5453,n5454);
or (n5453,n3626,n3603);
nand (n5454,n3603,n3626);
nand (n5455,n3863,n5280);
and (n5456,n5438,n5446);
and (n5457,n5427,n5434);
or (n5458,n5459,n5464);
and (n5459,n5460,n5463);
xor (n5460,n5461,n5462);
xor (n5461,n5180,n5196);
xor (n5462,n5129,n5145);
xor (n5463,n5276,n5291);
and (n5464,n5461,n5462);
xor (n5465,n5126,n5178);
and (n5466,n5424,n5458);
or (n5467,n5468,n5503);
and (n5468,n5469,n5502);
xor (n5469,n5470,n5471);
xor (n5470,n5224,n5274);
or (n5471,n5472,n5501);
and (n5472,n5473,n5500);
xor (n5473,n5474,n5499);
or (n5474,n5475,n5498);
and (n5475,n5476,n5492);
xor (n5476,n5477,n5485);
nand (n5477,n5478,n5484);
or (n5478,n5479,n3570);
not (n5479,n5480);
nor (n5480,n5481,n5483);
and (n5481,n3580,n5482);
not (n5482,n4406);
and (n5483,n3581,n4406);
nand (n5484,n5191,n3725);
nand (n5485,n5486,n5491);
or (n5486,n5487,n3737);
not (n5487,n5488);
nor (n5488,n5489,n5490);
and (n5489,n3735,n3935);
and (n5490,n3733,n3937);
nand (n5491,n5430,n3739);
nand (n5492,n5493,n5494);
or (n5493,n5261,n3754);
or (n5494,n3766,n5495);
nor (n5495,n5496,n5497);
and (n5496,n3658,n4415);
and (n5497,n3659,n4413);
and (n5498,n5477,n5485);
xor (n5499,n5252,n5267);
xor (n5500,n5156,n5171);
and (n5501,n5474,n5499);
xor (n5502,n5311,n5314);
and (n5503,n5470,n5471);
and (n5504,n5333,n5421);
xor (n5505,n5304,n5319);
or (n5506,n5507,n5649);
and (n5507,n5508,n5511);
xor (n5508,n5509,n5510);
xor (n5509,n5221,n5297);
xor (n5510,n5308,n5317);
or (n5511,n5512,n5648);
and (n5512,n5513,n5647);
xor (n5513,n5514,n5515);
xor (n5514,n5335,n5338);
or (n5515,n5516,n5646);
and (n5516,n5517,n5645);
xor (n5517,n5518,n5589);
or (n5518,n5519,n5588);
and (n5519,n5520,n5561);
xor (n5520,n5521,n5540);
or (n5521,n5522,n5539);
and (n5522,n5523,n5535);
xor (n5523,n5524,n5530);
nor (n5524,n5525,n3580);
and (n5525,n5526,n5529);
nand (n5526,n5527,n3577);
not (n5527,n5528);
and (n5528,n5233,n3575);
nand (n5529,n3574,n5235);
nor (n5530,n5531,n3659);
and (n5531,n5532,n5534);
nand (n5532,n5533,n3733);
or (n5533,n3756,n5240);
nand (n5534,n5240,n3756);
nand (n5535,n5536,n5538);
or (n5536,n4386,n5537);
xnor (n5537,n3641,n3867);
or (n5538,n5440,n4387);
and (n5539,n5524,n5530);
or (n5540,n5541,n5560);
and (n5541,n5542,n5557);
xor (n5542,n5543,n5550);
nand (n5543,n5544,n5549);
or (n5544,n5545,n4087);
not (n5545,n5546);
nand (n5546,n5547,n5548);
or (n5547,n4122,n3603);
nand (n5548,n3603,n4122);
nand (n5549,n3863,n5452);
nand (n5550,n5551,n5556);
or (n5551,n5552,n3825);
not (n5552,n5553);
nand (n5553,n5554,n5555);
or (n5554,n3791,n3632);
nand (n5555,n3632,n3791);
nand (n5556,n3831,n5347);
nor (n5557,n5558,n5559);
nand (n5558,n3725,n5233);
nand (n5559,n5241,n4116);
and (n5560,n5543,n5550);
or (n5561,n5562,n5587);
and (n5562,n5563,n5579);
xor (n5563,n5564,n5572);
nand (n5564,n5565,n5571);
or (n5565,n4425,n5566);
not (n5566,n5567);
nand (n5567,n5568,n5569);
or (n5568,n3518,n4032);
not (n5569,n5570);
and (n5570,n3518,n4032);
nand (n5571,n5354,n4423);
nand (n5572,n5573,n5578);
or (n5573,n5574,n3627);
not (n5574,n5575);
nand (n5575,n5576,n5577);
or (n5576,n3624,n3970);
nand (n5577,n3624,n3970);
nand (n5578,n3629,n5362);
nand (n5579,n5580,n5581);
or (n5580,n5372,n4029);
or (n5581,n4021,n5582);
not (n5582,n5583);
nand (n5583,n5584,n5585);
or (n5584,n3545,n3808);
not (n5585,n5586);
and (n5586,n3545,n3808);
and (n5587,n5564,n5572);
and (n5588,n5521,n5540);
or (n5589,n5590,n5644);
and (n5590,n5591,n5643);
xor (n5591,n5592,n5617);
or (n5592,n5593,n5616);
and (n5593,n5594,n5609);
xor (n5594,n5595,n5602);
nand (n5595,n5596,n5601);
nand (n5596,n3812,n5597,n3813);
nand (n5597,n5598,n5600);
not (n5598,n5599);
and (n5599,n3763,n3528);
nand (n5600,n3527,n3762);
nand (n5601,n3804,n5380);
nand (n5602,n5603,n5608);
or (n5603,n5604,n3606);
not (n5604,n5605);
nand (n5605,n5606,n5607);
or (n5606,n3999,n3611);
nand (n5607,n3611,n3999);
nand (n5608,n3599,n5389);
nand (n5609,n5610,n5615);
or (n5610,n5611,n3682);
not (n5611,n5612);
nor (n5612,n5613,n5614);
and (n5613,n3577,n5193);
and (n5614,n3573,n4350);
nand (n5615,n3689,n5399);
and (n5616,n5595,n5602);
or (n5617,n5618,n5642);
and (n5618,n5619,n5636);
xor (n5619,n5620,n5628);
nand (n5620,n5621,n5627);
or (n5621,n5622,n3523);
not (n5622,n5623);
nand (n5623,n5624,n5626);
not (n5624,n5625);
and (n5625,n3651,n3519);
nand (n5626,n3521,n3653);
nand (n5627,n5406,n3525);
nand (n5628,n5629,n5635);
or (n5629,n5630,n3549);
not (n5630,n5631);
nand (n5631,n5632,n5633);
or (n5632,n3546,n3929);
not (n5633,n5634);
and (n5634,n3929,n3546);
nand (n5635,n3558,n5413);
nand (n5636,n5637,n5641);
or (n5637,n3570,n5638);
nor (n5638,n5639,n5640);
and (n5639,n3580,n5233);
and (n5640,n3581,n5235);
nand (n5641,n3725,n5480);
and (n5642,n5620,n5628);
xor (n5643,n5437,n5450);
and (n5644,n5592,n5617);
xor (n5645,n5340,n5393);
and (n5646,n5518,n5589);
xor (n5647,n5469,n5502);
and (n5648,n5514,n5515);
and (n5649,n5509,n5510);
and (n5650,n5330,n5505);
nor (n5651,n5652,n5653);
xor (n5652,n5329,n5506);
or (n5653,n5654,n5819);
and (n5654,n5655,n5818);
xor (n5655,n5656,n5657);
xor (n5656,n5332,n5467);
or (n5657,n5658,n5817);
and (n5658,n5659,n5674);
xor (n5659,n5660,n5673);
or (n5660,n5661,n5672);
and (n5661,n5662,n5671);
xor (n5662,n5663,n5664);
xor (n5663,n5426,n5435);
or (n5664,n5665,n5670);
and (n5665,n5666,n5669);
xor (n5666,n5667,n5668);
xor (n5667,n5476,n5492);
xor (n5668,n5369,n5385);
xor (n5669,n5343,n5359);
and (n5670,n5667,n5668);
xor (n5671,n5460,n5463);
and (n5672,n5663,n5664);
xor (n5673,n5423,n5465);
or (n5674,n5675,n5816);
and (n5675,n5676,n5782);
xor (n5676,n5677,n5678);
xor (n5677,n5473,n5500);
or (n5678,n5679,n5781);
and (n5679,n5680,n5764);
xor (n5680,n5681,n5682);
xor (n5681,n5395,n5410);
or (n5682,n5683,n5763);
and (n5683,n5684,n5737);
xor (n5684,n5685,n5711);
or (n5685,n5686,n5710);
and (n5686,n5687,n5702);
xor (n5687,n5688,n5695);
nand (n5688,n5689,n5694);
or (n5689,n5690,n4087);
not (n5690,n5691);
nand (n5691,n5692,n5693);
or (n5692,n3679,n3603);
nand (n5693,n3603,n3679);
nand (n5694,n5546,n3863);
nand (n5695,n5696,n5701);
or (n5696,n5697,n3825);
not (n5697,n5698);
nand (n5698,n5699,n5700);
or (n5699,n3800,n3631);
nand (n5700,n3631,n3800);
nand (n5701,n5553,n3831);
nand (n5702,n5703,n5704);
or (n5703,n4426,n5566);
or (n5704,n5705,n4425);
not (n5705,n5706);
nand (n5706,n5707,n5708);
or (n5707,n3566,n4032);
not (n5708,n5709);
and (n5709,n3566,n4032);
and (n5710,n5688,n5695);
or (n5711,n5712,n5736);
and (n5712,n5713,n5729);
xor (n5713,n5714,n5722);
nand (n5714,n5715,n5721);
or (n5715,n5716,n4021);
not (n5716,n5717);
nand (n5717,n5718,n5719);
or (n5718,n3732,n3808);
not (n5719,n5720);
and (n5720,n3732,n3808);
nand (n5721,n4035,n5583);
nand (n5722,n5723,n5728);
or (n5723,n5724,n3627);
not (n5724,n5725);
nand (n5725,n5726,n5727);
or (n5726,n3952,n3623);
nand (n5727,n3623,n3952);
nand (n5728,n3629,n5575);
nand (n5729,n5730,n5732);
or (n5730,n5731,n3812);
not (n5731,n5597);
or (n5732,n3811,n5733);
nor (n5733,n5734,n5735);
and (n5734,n3527,n4271);
and (n5735,n3528,n3774);
and (n5736,n5714,n5722);
or (n5737,n5738,n5762);
and (n5738,n5739,n5754);
xor (n5739,n5740,n5747);
nand (n5740,n5741,n5746);
or (n5741,n5742,n3523);
not (n5742,n5743);
nor (n5743,n5744,n5745);
and (n5744,n3670,n3521);
and (n5745,n3913,n3519);
nand (n5746,n3525,n5623);
nand (n5747,n5748,n5753);
or (n5748,n5749,n3682);
not (n5749,n5750);
nand (n5750,n5751,n5752);
or (n5751,n3573,n5482);
nand (n5752,n5482,n3573);
nand (n5753,n5612,n3689);
nand (n5754,n5755,n5761);
or (n5755,n5756,n3549);
not (n5756,n5757);
nand (n5757,n5758,n5759);
or (n5758,n3546,n3935);
not (n5759,n5760);
and (n5760,n3935,n3546);
nand (n5761,n3558,n5631);
and (n5762,n5740,n5747);
and (n5763,n5685,n5711);
or (n5764,n5765,n5780);
and (n5765,n5766,n5779);
xor (n5766,n5767,n5773);
nand (n5767,n5768,n5772);
or (n5768,n3737,n5769);
nor (n5769,n5770,n5771);
and (n5770,n3735,n4341);
and (n5771,n3733,n4342);
or (n5772,n3892,n5487);
nand (n5773,n5774,n5778);
or (n5774,n3766,n5775);
nor (n5775,n5776,n5777);
and (n5776,n5240,n3658);
and (n5777,n5241,n3659);
or (n5778,n5495,n3754);
xor (n5779,n5523,n5535);
and (n5780,n5767,n5773);
and (n5781,n5681,n5682);
or (n5782,n5783,n5815);
and (n5783,n5784,n5787);
xor (n5784,n5785,n5786);
xor (n5785,n5591,n5643);
xor (n5786,n5520,n5561);
or (n5787,n5788,n5814);
and (n5788,n5789,n5813);
xor (n5789,n5790,n5812);
or (n5790,n5791,n5811);
and (n5791,n5792,n5805);
xor (n5792,n5793,n5797);
nand (n5793,n5794,n5796);
or (n5794,n5795,n5558);
not (n5795,n5559);
nand (n5796,n5795,n5558);
nand (n5797,n5798,n5804);
or (n5798,n3737,n5799);
not (n5799,n5800);
nand (n5800,n5801,n5802);
or (n5801,n4413,n3733);
not (n5802,n5803);
and (n5803,n4413,n3733);
or (n5804,n3892,n5769);
nand (n5805,n5806,n5810);
or (n5806,n4386,n5807);
nor (n5807,n5808,n5809);
and (n5808,n3873,n3622);
and (n5809,n3867,n3626);
or (n5810,n5537,n4387);
and (n5811,n5793,n5797);
xor (n5812,n5542,n5557);
xor (n5813,n5619,n5636);
and (n5814,n5790,n5812);
and (n5815,n5785,n5786);
and (n5816,n5677,n5678);
and (n5817,n5660,n5673);
xor (n5818,n5508,n5511);
and (n5819,n5656,n5657);
nand (n5820,n5821,n5837);
not (n5821,n5822);
nor (n5822,n5823,n5824);
xor (n5823,n5655,n5818);
or (n5824,n5825,n5836);
and (n5825,n5826,n5829);
xor (n5826,n5827,n5828);
xor (n5827,n5513,n5647);
xor (n5828,n5659,n5674);
or (n5829,n5830,n5835);
and (n5830,n5831,n5834);
xor (n5831,n5832,n5833);
xor (n5832,n5662,n5671);
xor (n5833,n5517,n5645);
xor (n5834,n5676,n5782);
and (n5835,n5832,n5833);
and (n5836,n5827,n5828);
nand (n5837,n5838,n5840);
not (n5838,n5839);
xor (n5839,n5826,n5829);
not (n5840,n5841);
or (n5841,n5842,n6018);
and (n5842,n5843,n6017);
xor (n5843,n5844,n5998);
or (n5844,n5845,n5997);
and (n5845,n5846,n5855);
xor (n5846,n5847,n5848);
xor (n5847,n5666,n5669);
or (n5848,n5849,n5854);
and (n5849,n5850,n5853);
xor (n5850,n5851,n5852);
xor (n5851,n5563,n5579);
xor (n5852,n5594,n5609);
xor (n5853,n5766,n5779);
and (n5854,n5851,n5852);
or (n5855,n5856,n5996);
and (n5856,n5857,n5995);
xor (n5857,n5858,n5924);
or (n5858,n5859,n5923);
and (n5859,n5860,n5895);
xor (n5860,n5861,n5868);
nand (n5861,n5862,n5867);
or (n5862,n3606,n5863);
not (n5863,n5864);
nand (n5864,n5865,n5866);
or (n5865,n3592,n3610);
nand (n5866,n3610,n3592);
or (n5867,n3607,n5604);
or (n5868,n5869,n5894);
and (n5869,n5870,n5886);
xor (n5870,n5871,n5878);
nand (n5871,n5872,n5877);
or (n5872,n5873,n3825);
not (n5873,n5874);
nand (n5874,n5875,n5876);
or (n5875,n3959,n3631);
nand (n5876,n3631,n3959);
nand (n5877,n3831,n5698);
nand (n5878,n5879,n5885);
or (n5879,n4425,n5880);
not (n5880,n5881);
nand (n5881,n5882,n5883);
or (n5882,n3545,n4032);
not (n5883,n5884);
and (n5884,n3545,n4032);
nand (n5885,n5706,n4423);
nand (n5886,n5887,n5888);
or (n5887,n5716,n4029);
or (n5888,n4021,n5889);
not (n5889,n5890);
nand (n5890,n5891,n5892);
or (n5891,n3763,n3808);
not (n5892,n5893);
and (n5893,n3763,n3808);
and (n5894,n5871,n5878);
or (n5895,n5896,n5922);
and (n5896,n5897,n5914);
xor (n5897,n5898,n5905);
nand (n5898,n5899,n5904);
or (n5899,n5900,n3627);
not (n5900,n5901);
nand (n5901,n5902,n5903);
or (n5902,n4350,n3623);
or (n5903,n5193,n3624);
nand (n5904,n3629,n5725);
nand (n5905,n5906,n5912);
or (n5906,n5907,n3811);
not (n5907,n5908);
nand (n5908,n5909,n5910);
or (n5909,n3651,n3528);
not (n5910,n5911);
and (n5911,n3651,n3528);
nand (n5912,n5913,n3804);
not (n5913,n5733);
nand (n5914,n5915,n5921);
or (n5915,n3523,n5916);
not (n5916,n5917);
nand (n5917,n5918,n5920);
not (n5918,n5919);
and (n5919,n3929,n3519);
nand (n5920,n3521,n3984);
or (n5921,n3524,n5742);
and (n5922,n5898,n5905);
and (n5923,n5861,n5868);
or (n5924,n5925,n5994);
and (n5925,n5926,n5973);
xor (n5926,n5927,n5953);
or (n5927,n5928,n5952);
and (n5928,n5929,n5945);
xor (n5929,n5930,n5937);
nand (n5930,n5931,n5936);
or (n5931,n5932,n3682);
not (n5932,n5933);
nor (n5933,n5934,n5935);
and (n5934,n3577,n5235);
and (n5935,n5233,n3573);
nand (n5936,n5750,n3689);
nand (n5937,n5938,n5944);
or (n5938,n5939,n3549);
not (n5939,n5940);
nand (n5940,n5941,n5943);
not (n5941,n5942);
and (n5942,n4342,n3546);
nand (n5943,n3548,n4341);
nand (n5944,n5757,n3558);
nand (n5945,n5946,n5951);
or (n5946,n5947,n3737);
not (n5947,n5948);
nor (n5948,n5949,n5950);
and (n5949,n3735,n5241);
and (n5950,n3733,n5240);
nand (n5951,n5800,n3739);
and (n5952,n5930,n5937);
or (n5953,n5954,n5972);
and (n5954,n5955,n5968);
xor (n5955,n5956,n5962);
nand (n5956,n5957,n5961);
or (n5957,n4386,n5958);
nor (n5958,n5959,n5960);
and (n5959,n3873,n3695);
and (n5960,n3867,n4122);
or (n5961,n5807,n4387);
nand (n5962,n5963,n5967);
or (n5963,n3606,n5964);
nor (n5964,n5965,n5966);
and (n5965,n3791,n3611);
and (n5966,n3586,n3610);
nand (n5967,n5864,n3599);
nor (n5968,n5969,n5971);
not (n5969,n5970);
and (n5970,n3689,n5233);
nand (n5971,n3739,n5241);
and (n5972,n5956,n5962);
or (n5973,n5974,n5993);
and (n5974,n5975,n5986);
xor (n5975,n5976,n5981);
nor (n5976,n5977,n3577);
nor (n5977,n5978,n5980);
nor (n5978,n5979,n3624);
and (n5979,n5233,n3687);
nor (n5980,n5233,n3687);
and (n5981,n5982,n3735);
nand (n5982,n5983,n5984);
or (n5983,n3746,n5241);
nand (n5984,n5985,n3546);
or (n5985,n5240,n3741);
nand (n5986,n5987,n5992);
or (n5987,n5988,n4087);
not (n5988,n5989);
nand (n5989,n5990,n5991);
or (n5990,n3723,n3871);
or (n5991,n3603,n3999);
nand (n5992,n3863,n5691);
and (n5993,n5976,n5981);
and (n5994,n5927,n5953);
xor (n5995,n5684,n5737);
and (n5996,n5858,n5924);
and (n5997,n5847,n5848);
or (n5998,n5999,n6016);
and (n5999,n6000,n6003);
xor (n6000,n6001,n6002);
xor (n6001,n5680,n5764);
xor (n6002,n5784,n5787);
or (n6003,n6004,n6015);
and (n6004,n6005,n6014);
xor (n6005,n6006,n6013);
or (n6006,n6007,n6012);
and (n6007,n6008,n6011);
xor (n6008,n6009,n6010);
xor (n6009,n5739,n5754);
xor (n6010,n5792,n5805);
xor (n6011,n5687,n5702);
and (n6012,n6009,n6010);
xor (n6013,n5789,n5813);
xor (n6014,n5850,n5853);
and (n6015,n6006,n6013);
and (n6016,n6001,n6002);
xor (n6017,n5831,n5834);
and (n6018,n5844,n5998);
nand (n6019,n6020,n6930);
or (n6020,n6021,n6278);
not (n6021,n6022);
nor (n6022,n6023,n6134);
nor (n6023,n6024,n6025);
xor (n6024,n5843,n6017);
or (n6025,n6026,n6133);
and (n6026,n6027,n6132);
xor (n6027,n6028,n6029);
xor (n6028,n5846,n5855);
or (n6029,n6030,n6131);
and (n6030,n6031,n6124);
xor (n6031,n6032,n6033);
xor (n6032,n5857,n5995);
or (n6033,n6034,n6123);
and (n6034,n6035,n6089);
xor (n6035,n6036,n6037);
xor (n6036,n5713,n5729);
or (n6037,n6038,n6088);
and (n6038,n6039,n6062);
xor (n6039,n6040,n6041);
xor (n6040,n5975,n5986);
or (n6041,n6042,n6061);
and (n6042,n6043,n6054);
xor (n6043,n6044,n6051);
nand (n6044,n6045,n6050);
or (n6045,n6046,n4087);
not (n6046,n6047);
nor (n6047,n6048,n6049);
and (n6048,n4058,n3871);
and (n6049,n3592,n3603);
nand (n6050,n3863,n5989);
nand (n6051,n6052,n6053);
or (n6052,n5970,n5971);
nand (n6053,n5971,n5970);
nand (n6054,n6055,n6060);
or (n6055,n3825,n6056);
not (n6056,n6057);
nand (n6057,n6058,n6059);
or (n6058,n3951,n3632);
nand (n6059,n3632,n3951);
or (n6060,n3830,n5873);
and (n6061,n6044,n6051);
or (n6062,n6063,n6087);
and (n6063,n6064,n6080);
xor (n6064,n6065,n6073);
nand (n6065,n6066,n6072);
or (n6066,n6067,n4021);
not (n6067,n6068);
nand (n6068,n6069,n6070);
or (n6069,n3774,n3808);
not (n6070,n6071);
and (n6071,n3774,n3808);
nand (n6072,n4035,n5890);
nand (n6073,n6074,n6079);
or (n6074,n6075,n3811);
not (n6075,n6076);
nor (n6076,n6077,n6078);
and (n6077,n3670,n3527);
and (n6078,n3913,n3528);
nand (n6079,n3804,n5908);
nand (n6080,n6081,n6086);
or (n6081,n6082,n3627);
not (n6082,n6083);
nand (n6083,n6084,n6085);
or (n6084,n3624,n5482);
nand (n6085,n3624,n5482);
nand (n6086,n3629,n5901);
and (n6087,n6065,n6073);
and (n6088,n6040,n6041);
or (n6089,n6090,n6122);
and (n6090,n6091,n6121);
xor (n6091,n6092,n6120);
or (n6092,n6093,n6119);
and (n6093,n6094,n6111);
xor (n6094,n6095,n6103);
nand (n6095,n6096,n6102);
or (n6096,n6097,n3523);
not (n6097,n6098);
nand (n6098,n6099,n6101);
not (n6099,n6100);
and (n6100,n3935,n3519);
nand (n6101,n3937,n3521);
nand (n6102,n5917,n3525);
nand (n6103,n6104,n6110);
or (n6104,n6105,n3549);
not (n6105,n6106);
nand (n6106,n6107,n6108);
or (n6107,n4413,n3546);
not (n6108,n6109);
and (n6109,n4413,n3546);
nand (n6110,n5940,n3558);
nand (n6111,n6112,n6117);
or (n6112,n6113,n4386);
not (n6113,n6114);
nor (n6114,n6115,n6116);
and (n6115,n3679,n3873);
and (n6116,n3680,n3867);
nand (n6117,n6118,n4384);
not (n6118,n5958);
and (n6119,n6095,n6103);
xor (n6120,n5955,n5968);
xor (n6121,n5870,n5886);
and (n6122,n6092,n6120);
and (n6123,n6036,n6037);
or (n6124,n6125,n6130);
and (n6125,n6126,n6129);
xor (n6126,n6127,n6128);
xor (n6127,n5926,n5973);
xor (n6128,n5860,n5895);
xor (n6129,n6008,n6011);
and (n6130,n6127,n6128);
and (n6131,n6032,n6033);
xor (n6132,n6000,n6003);
and (n6133,n6028,n6029);
nor (n6134,n6135,n6136);
xor (n6135,n6027,n6132);
or (n6136,n6137,n6277);
and (n6137,n6138,n6276);
xor (n6138,n6139,n6140);
xor (n6139,n6005,n6014);
or (n6140,n6141,n6275);
and (n6141,n6142,n6274);
xor (n6142,n6143,n6187);
or (n6143,n6144,n6186);
and (n6144,n6145,n6148);
xor (n6145,n6146,n6147);
xor (n6146,n5897,n5914);
xor (n6147,n5929,n5945);
or (n6148,n6149,n6185);
and (n6149,n6150,n6164);
xor (n6150,n6151,n6157);
nand (n6151,n6152,n6156);
or (n6152,n3606,n6153);
nor (n6153,n6154,n6155);
and (n6154,n3610,n3800);
and (n6155,n3611,n3882);
or (n6156,n3607,n5964);
nand (n6157,n6158,n6159);
or (n6158,n4426,n5880);
nand (n6159,n6160,n4424);
not (n6160,n6161);
nor (n6161,n6162,n6163);
and (n6162,n4031,n3736);
and (n6163,n4032,n3732);
or (n6164,n6165,n6184);
and (n6165,n6166,n6181);
xor (n6166,n6167,n6173);
nand (n6167,n6168,n6169);
or (n6168,n4387,n6113);
nand (n6169,n6170,n4385);
nor (n6170,n6171,n6172);
and (n6171,n3723,n3867);
and (n6172,n3999,n3873);
nand (n6173,n6174,n6179);
or (n6174,n6175,n3606);
not (n6175,n6176);
nand (n6176,n6177,n6178);
or (n6177,n3959,n3610);
nand (n6178,n3610,n3959);
nand (n6179,n6180,n3599);
not (n6180,n6153);
nor (n6181,n6182,n6183);
nand (n6182,n3629,n5233);
nand (n6183,n3558,n5241);
and (n6184,n6167,n6173);
and (n6185,n6151,n6157);
and (n6186,n6146,n6147);
or (n6187,n6188,n6273);
and (n6188,n6189,n6272);
xor (n6189,n6190,n6265);
or (n6190,n6191,n6264);
and (n6191,n6192,n6239);
xor (n6192,n6193,n6217);
or (n6193,n6194,n6216);
and (n6194,n6195,n6210);
xor (n6195,n6196,n6202);
nand (n6196,n6197,n6198);
or (n6197,n3628,n6082);
nand (n6198,n3628,n6199,n3635);
nand (n6199,n6200,n6201);
or (n6200,n3624,n5235);
nand (n6201,n5235,n3624);
nand (n6202,n6203,n6209);
or (n6203,n6204,n3523);
not (n6204,n6205);
nand (n6205,n6206,n6207);
or (n6206,n3519,n4342);
not (n6207,n6208);
and (n6208,n4342,n3519);
nand (n6209,n3525,n6098);
nand (n6210,n6211,n6212);
or (n6211,n6105,n3557);
or (n6212,n3549,n6213);
nor (n6213,n6214,n6215);
and (n6214,n3548,n5240);
and (n6215,n5241,n3546);
and (n6216,n6196,n6202);
or (n6217,n6218,n6238);
and (n6218,n6219,n6232);
xor (n6219,n6220,n6227);
nor (n6220,n6221,n3623);
and (n6221,n6222,n6225);
nand (n6222,n6223,n3631);
not (n6223,n6224);
and (n6224,n5233,n3633);
nand (n6225,n5235,n6226);
not (n6226,n3633);
nor (n6227,n6228,n3546);
nor (n6228,n6229,n6231);
and (n6229,n6230,n3519);
nand (n6230,n5241,n3553);
and (n6231,n5240,n3554);
nand (n6232,n6233,n6237);
or (n6233,n6234,n4087);
nor (n6234,n6235,n6236);
and (n6235,n3791,n3603);
and (n6236,n3586,n3871);
nand (n6237,n6047,n3863);
and (n6238,n6220,n6227);
or (n6239,n6240,n6263);
and (n6240,n6241,n6256);
xor (n6241,n6242,n6249);
nand (n6242,n6243,n6248);
or (n6243,n6244,n3825);
not (n6244,n6245);
nand (n6245,n6246,n6247);
or (n6246,n4350,n3631);
nand (n6247,n3631,n4350);
nand (n6248,n3831,n6057);
nand (n6249,n6250,n6255);
or (n6250,n4021,n6251);
not (n6251,n6252);
nor (n6252,n6253,n6254);
and (n6253,n3653,n3808);
and (n6254,n3651,n3807);
nand (n6255,n4035,n6068);
nand (n6256,n6257,n6262);
or (n6257,n6258,n3811);
not (n6258,n6259);
nor (n6259,n6260,n6261);
and (n6260,n3984,n3528);
and (n6261,n3929,n3527);
nand (n6262,n3804,n6076);
and (n6263,n6242,n6249);
and (n6264,n6193,n6217);
or (n6265,n6266,n6271);
and (n6266,n6267,n6270);
xor (n6267,n6268,n6269);
xor (n6268,n6094,n6111);
xor (n6269,n6064,n6080);
xor (n6270,n6043,n6054);
and (n6271,n6268,n6269);
xor (n6272,n6039,n6062);
and (n6273,n6190,n6265);
xor (n6274,n6035,n6089);
and (n6275,n6143,n6187);
xor (n6276,n6031,n6124);
and (n6277,n6139,n6140);
not (n6278,n6279);
nor (n6279,n6280,n6911);
nor (n6280,n6281,n6910);
and (n6281,n6282,n6893);
nand (n6282,n6283,n6892);
or (n6283,n6284,n6558);
not (n6284,n6285);
or (n6285,n6286,n6476);
xor (n6286,n6287,n6390);
xor (n6287,n6288,n6383);
or (n6288,n6289,n6382);
and (n6289,n6290,n6375);
xor (n6290,n6291,n6346);
xor (n6291,n6292,n6321);
xor (n6292,n6293,n6300);
nand (n6293,n6294,n6299);
or (n6294,n4425,n6295);
not (n6295,n6296);
nor (n6296,n6297,n6298);
and (n6297,n3763,n4031);
and (n6298,n3762,n4032);
or (n6299,n6161,n4426);
or (n6300,n6301,n6320);
and (n6301,n6302,n6313);
xor (n6302,n6303,n6307);
nand (n6303,n6304,n6306);
or (n6304,n6305,n6183);
not (n6305,n6182);
nand (n6306,n6305,n6183);
nand (n6307,n6308,n6312);
or (n6308,n4386,n6309);
nor (n6309,n6310,n6311);
and (n6310,n3592,n3873);
and (n6311,n4058,n3867);
nand (n6312,n6170,n4384);
nand (n6313,n6314,n6319);
or (n6314,n4087,n6315);
not (n6315,n6316);
nor (n6316,n6317,n6318);
and (n6317,n3882,n3871);
and (n6318,n3800,n3603);
or (n6319,n4093,n6234);
and (n6320,n6303,n6307);
or (n6321,n6322,n6345);
and (n6322,n6323,n6338);
xor (n6323,n6324,n6331);
nand (n6324,n6325,n6330);
or (n6325,n6326,n3606);
not (n6326,n6327);
nand (n6327,n6328,n6329);
or (n6328,n3952,n3610);
nand (n6329,n3610,n3952);
nand (n6330,n3599,n6176);
nand (n6331,n6332,n6333);
or (n6332,n4426,n6295);
nand (n6333,n6334,n4424);
nand (n6334,n6335,n6337);
not (n6335,n6336);
and (n6336,n3774,n4032);
nand (n6337,n4271,n4031);
nand (n6338,n6339,n6344);
or (n6339,n6340,n4021);
not (n6340,n6341);
nor (n6341,n6342,n6343);
and (n6342,n3913,n3808);
and (n6343,n3670,n3807);
nand (n6344,n4035,n6252);
and (n6345,n6324,n6331);
or (n6346,n6347,n6374);
and (n6347,n6348,n6373);
xor (n6348,n6349,n6350);
xor (n6349,n6323,n6338);
xor (n6350,n6351,n6366);
xor (n6351,n6352,n6359);
nand (n6352,n6353,n6358);
or (n6353,n6354,n3825);
not (n6354,n6355);
nand (n6355,n6356,n6357);
or (n6356,n4406,n3631);
nand (n6357,n3631,n4406);
nand (n6358,n6245,n3831);
nand (n6359,n6360,n6365);
or (n6360,n6361,n3811);
not (n6361,n6362);
nor (n6362,n6363,n6364);
and (n6363,n3937,n3528);
and (n6364,n3935,n3527);
nand (n6365,n3804,n6259);
nand (n6366,n6367,n6372);
or (n6367,n6368,n3523);
not (n6368,n6369);
nor (n6369,n6370,n6371);
and (n6370,n4415,n3519);
and (n6371,n4413,n3521);
nand (n6372,n3525,n6205);
xor (n6373,n6302,n6313);
and (n6374,n6349,n6350);
xor (n6375,n6376,n6381);
xor (n6376,n6377,n6378);
xor (n6377,n6219,n6232);
or (n6378,n6379,n6380);
and (n6379,n6351,n6366);
and (n6380,n6352,n6359);
xor (n6381,n6241,n6256);
and (n6382,n6291,n6346);
xor (n6383,n6384,n6389);
xor (n6384,n6385,n6388);
or (n6385,n6386,n6387);
and (n6386,n6292,n6321);
and (n6387,n6293,n6300);
xor (n6388,n6150,n6164);
xor (n6389,n6192,n6239);
xor (n6390,n6391,n6396);
xor (n6391,n6392,n6395);
or (n6392,n6393,n6394);
and (n6393,n6376,n6381);
and (n6394,n6377,n6378);
xor (n6395,n6267,n6270);
or (n6396,n6397,n6475);
and (n6397,n6398,n6401);
xor (n6398,n6399,n6400);
xor (n6399,n6166,n6181);
xor (n6400,n6195,n6210);
or (n6401,n6402,n6474);
and (n6402,n6403,n6449);
xor (n6403,n6404,n6425);
or (n6404,n6405,n6424);
and (n6405,n6406,n6417);
xor (n6406,n6407,n6414);
nand (n6407,n6408,n6413);
or (n6408,n6409,n4087);
not (n6409,n6410);
nand (n6410,n6411,n6412);
or (n6411,n3970,n3603);
nand (n6412,n3603,n3970);
nand (n6413,n6316,n3863);
nor (n6414,n6415,n6416);
nand (n6415,n3831,n5233);
nand (n6416,n3525,n5241);
nand (n6417,n6418,n6423);
or (n6418,n6419,n3606);
not (n6419,n6420);
nand (n6420,n6421,n6422);
or (n6421,n4350,n3610);
nand (n6422,n4350,n3610);
nand (n6423,n3599,n6327);
and (n6424,n6407,n6414);
or (n6425,n6426,n6448);
and (n6426,n6427,n6441);
xor (n6427,n6428,n6435);
nor (n6428,n6429,n3631);
and (n6429,n6430,n6433);
nand (n6430,n6431,n3610);
not (n6431,n6432);
and (n6432,n5233,n3828);
nand (n6433,n5235,n6434);
not (n6434,n3828);
nor (n6435,n6436,n3519);
nor (n6436,n6437,n6440);
and (n6437,n6438,n3528);
nand (n6438,n5241,n6439);
not (n6439,n3529);
nor (n6440,n5241,n6439);
nand (n6441,n6442,n6447);
or (n6442,n6443,n3825);
not (n6443,n6444);
nor (n6444,n6445,n6446);
and (n6445,n3631,n5235);
and (n6446,n5233,n3632);
nand (n6447,n6355,n3831);
and (n6448,n6428,n6435);
or (n6449,n6450,n6473);
and (n6450,n6451,n6466);
xor (n6451,n6452,n6459);
nand (n6452,n6453,n6458);
or (n6453,n6454,n3811);
not (n6454,n6455);
nor (n6455,n6456,n6457);
and (n6456,n4341,n3528);
and (n6457,n4342,n3527);
nand (n6458,n3804,n6362);
nand (n6459,n6460,n6461);
or (n6460,n3524,n6368);
nand (n6461,n6462,n4596);
not (n6462,n6463);
nor (n6463,n6464,n6465);
and (n6464,n5240,n3521);
and (n6465,n5241,n3519);
nand (n6466,n6467,n6472);
or (n6467,n4386,n6468);
not (n6468,n6469);
nand (n6469,n6470,n6471);
or (n6470,n3586,n3873);
nand (n6471,n3873,n3586);
or (n6472,n6309,n4387);
and (n6473,n6452,n6459);
and (n6474,n6404,n6425);
and (n6475,n6399,n6400);
or (n6476,n6477,n6557);
and (n6477,n6478,n6556);
xor (n6478,n6479,n6480);
xor (n6479,n6398,n6401);
or (n6480,n6481,n6555);
and (n6481,n6482,n6554);
xor (n6482,n6483,n6523);
or (n6483,n6484,n6522);
and (n6484,n6485,n6500);
xor (n6485,n6486,n6493);
nand (n6486,n6487,n6491);
or (n6487,n6488,n4425);
nor (n6488,n6489,n6490);
and (n6489,n4031,n3653);
and (n6490,n4032,n3651);
or (n6491,n6492,n4426);
not (n6492,n6334);
nand (n6493,n6494,n6499);
or (n6494,n6495,n4021);
not (n6495,n6496);
nor (n6496,n6497,n6498);
and (n6497,n3984,n3808);
and (n6498,n3929,n3807);
nand (n6499,n4035,n6341);
or (n6500,n6501,n6521);
and (n6501,n6502,n6514);
xor (n6502,n6503,n6510);
nand (n6503,n6504,n6509);
or (n6504,n6505,n4386);
not (n6505,n6506);
nor (n6506,n6507,n6508);
and (n6507,n3800,n3867);
and (n6508,n3882,n3873);
nand (n6509,n6469,n4384);
nand (n6510,n6511,n6513);
or (n6511,n6512,n6416);
not (n6512,n6415);
nand (n6513,n6512,n6416);
nand (n6514,n6515,n6520);
or (n6515,n6516,n4087);
not (n6516,n6517);
nor (n6517,n6518,n6519);
and (n6518,n3951,n3871);
and (n6519,n3952,n3603);
or (n6520,n4093,n6409);
and (n6521,n6503,n6510);
and (n6522,n6486,n6493);
or (n6523,n6524,n6553);
and (n6524,n6525,n6552);
xor (n6525,n6526,n6527);
xor (n6526,n6427,n6441);
or (n6527,n6528,n6551);
and (n6528,n6529,n6543);
xor (n6529,n6530,n6536);
nand (n6530,n6531,n6535);
or (n6531,n6532,n4425);
or (n6532,n6533,n6534);
and (n6533,n3670,n4031);
and (n6534,n3913,n4032);
or (n6535,n6488,n4426);
nand (n6536,n6537,n6542);
or (n6537,n6538,n3606);
not (n6538,n6539);
nor (n6539,n6540,n6541);
and (n6540,n5482,n3610);
and (n6541,n4406,n3611);
nand (n6542,n6420,n3599);
nand (n6543,n6544,n6550);
or (n6544,n6545,n4021);
not (n6545,n6546);
nand (n6546,n6547,n6548);
or (n6547,n3935,n3808);
not (n6548,n6549);
and (n6549,n3935,n3808);
nand (n6550,n4035,n6496);
and (n6551,n6530,n6536);
xor (n6552,n6451,n6466);
and (n6553,n6526,n6527);
xor (n6554,n6403,n6449);
and (n6555,n6483,n6523);
xor (n6556,n6290,n6375);
and (n6557,n6479,n6480);
not (n6558,n6559);
nand (n6559,n6560,n6889,n6891);
nand (n6560,n6561,n6633,n6882);
nand (n6561,n6562,n6564);
not (n6562,n6563);
xor (n6563,n6478,n6556);
not (n6564,n6565);
or (n6565,n6566,n6632);
and (n6566,n6567,n6631);
xor (n6567,n6568,n6569);
xor (n6568,n6348,n6373);
or (n6569,n6570,n6630);
and (n6570,n6571,n6629);
xor (n6571,n6572,n6573);
xor (n6572,n6406,n6417);
or (n6573,n6574,n6628);
and (n6574,n6575,n6607);
xor (n6575,n6576,n6583);
nand (n6576,n6577,n6582);
or (n6577,n6578,n3811);
not (n6578,n6579);
nor (n6579,n6580,n6581);
and (n6580,n4415,n3528);
and (n6581,n4413,n3527);
nand (n6582,n3804,n6455);
or (n6583,n6584,n6606);
and (n6584,n6585,n6597);
xor (n6585,n6586,n6593);
nand (n6586,n6587,n6592);
or (n6587,n6588,n4087);
not (n6588,n6589);
nand (n6589,n6590,n6591);
or (n6590,n4350,n3871);
nand (n6591,n3871,n4350);
nand (n6592,n6517,n3863);
nor (n6593,n6594,n6596);
not (n6594,n6595);
and (n6595,n3804,n5241);
nand (n6596,n5233,n3599);
nand (n6597,n6598,n6604);
or (n6598,n4425,n6599);
not (n6599,n6600);
nand (n6600,n6601,n6603);
not (n6601,n6602);
and (n6602,n3929,n4032);
nand (n6603,n4031,n3984);
nand (n6604,n6605,n4423);
not (n6605,n6532);
and (n6606,n6586,n6593);
or (n6607,n6608,n6627);
and (n6608,n6609,n6621);
xor (n6609,n6610,n6616);
nor (n6610,n6611,n3610);
and (n6611,n6612,n6615);
nand (n6612,n6613,n3871);
not (n6613,n6614);
and (n6614,n5233,n3602);
nand (n6615,n5235,n3601);
nor (n6616,n6617,n3528);
nor (n6617,n6618,n6620);
and (n6618,n6619,n3808);
nand (n6619,n5241,n3815);
and (n6620,n5240,n3806);
nand (n6621,n6622,n6623);
or (n6622,n4387,n6505);
nand (n6623,n6624,n4385);
nor (n6624,n6625,n6626);
and (n6625,n3959,n3867);
and (n6626,n3970,n3873);
and (n6627,n6610,n6616);
and (n6628,n6576,n6583);
xor (n6629,n6485,n6500);
and (n6630,n6572,n6573);
xor (n6631,n6482,n6554);
and (n6632,n6568,n6569);
nand (n6633,n6634,n6881);
or (n6634,n6635,n6867);
not (n6635,n6636);
nand (n6636,n6637,n6866);
or (n6637,n6638,n6738);
not (n6638,n6639);
nand (n6639,n6640,n6702);
not (n6640,n6641);
xor (n6641,n6642,n6672);
xor (n6642,n6643,n6644);
xor (n6643,n6575,n6607);
or (n6644,n6645,n6671);
and (n6645,n6646,n6670);
xor (n6646,n6647,n6669);
or (n6647,n6648,n6668);
and (n6648,n6649,n6664);
xor (n6649,n6650,n6657);
nand (n6650,n6651,n6656);
or (n6651,n6652,n4087);
not (n6652,n6653);
nand (n6653,n6654,n6655);
or (n6654,n4406,n3871);
nand (n6655,n3871,n4406);
nand (n6656,n6589,n3863);
nand (n6657,n6658,n6659);
or (n6658,n4426,n6599);
nand (n6659,n6660,n4424);
nand (n6660,n6661,n6663);
not (n6661,n6662);
and (n6662,n3935,n4032);
nand (n6663,n4031,n3937);
nand (n6664,n6665,n6667);
or (n6665,n6666,n6594);
not (n6666,n6596);
or (n6667,n6595,n6596);
and (n6668,n6650,n6657);
xor (n6669,n6609,n6621);
xor (n6670,n6585,n6597);
and (n6671,n6647,n6669);
xor (n6672,n6673,n6701);
xor (n6673,n6674,n6700);
or (n6674,n6675,n6699);
and (n6675,n6676,n6691);
xor (n6676,n6677,n6684);
nand (n6677,n6678,n6683);
or (n6678,n6679,n3606);
not (n6679,n6680);
nor (n6680,n6681,n6682);
and (n6681,n3610,n5235);
and (n6682,n5233,n3611);
nand (n6683,n6539,n3599);
nand (n6684,n6685,n6690);
or (n6685,n6686,n4021);
not (n6686,n6687);
nor (n6687,n6688,n6689);
and (n6688,n4342,n3807);
and (n6689,n4341,n3808);
nand (n6690,n4035,n6546);
nand (n6691,n6692,n6698);
or (n6692,n6693,n3811);
not (n6693,n6694);
nand (n6694,n6695,n6696);
or (n6695,n5241,n3528);
not (n6696,n6697);
and (n6697,n5241,n3528);
nand (n6698,n3804,n6579);
and (n6699,n6677,n6684);
xor (n6700,n6529,n6543);
xor (n6701,n6502,n6514);
not (n6702,n6703);
or (n6703,n6704,n6737);
and (n6704,n6705,n6736);
xor (n6705,n6706,n6707);
xor (n6706,n6676,n6691);
or (n6707,n6708,n6735);
and (n6708,n6709,n6723);
xor (n6709,n6710,n6716);
nand (n6710,n6711,n6715);
or (n6711,n6712,n4021);
nor (n6712,n6713,n6714);
and (n6713,n4415,n3807);
and (n6714,n4413,n3808);
nand (n6715,n6687,n4035);
nand (n6716,n6717,n6722);
or (n6717,n4386,n6718);
not (n6718,n6719);
nor (n6719,n6720,n6721);
and (n6720,n3952,n3867);
and (n6721,n3951,n3873);
nand (n6722,n6624,n4384);
and (n6723,n6724,n6730);
nor (n6724,n6725,n3871);
and (n6725,n6726,n6729);
nand (n6726,n6727,n3873);
not (n6727,n6728);
and (n6728,n5233,n3866);
nand (n6729,n3865,n5235);
nor (n6730,n6731,n3808);
and (n6731,n6732,n6734);
nand (n6732,n6733,n4032);
or (n6733,n5240,n4025);
nand (n6734,n5240,n4025);
and (n6735,n6710,n6716);
xor (n6736,n6646,n6670);
and (n6737,n6706,n6707);
not (n6738,n6739);
nand (n6739,n6740,n6865);
or (n6740,n6741,n6857);
not (n6741,n6742);
nand (n6742,n6743,n6856);
or (n6743,n6744,n6815);
not (n6744,n6745);
nand (n6745,n6746,n6776);
not (n6746,n6747);
xor (n6747,n6748,n6775);
xor (n6748,n6749,n6774);
or (n6749,n6750,n6773);
and (n6750,n6751,n6767);
xor (n6751,n6752,n6759);
nand (n6752,n6753,n6758);
or (n6753,n6754,n4087);
not (n6754,n6755);
nand (n6755,n6756,n6757);
or (n6756,n5233,n3871);
nand (n6757,n3871,n5233);
nand (n6758,n6653,n3863);
nand (n6759,n6760,n6766);
or (n6760,n6761,n4425);
not (n6761,n6762);
nand (n6762,n6763,n6765);
not (n6763,n6764);
and (n6764,n4342,n4032);
nand (n6765,n4031,n4341);
nand (n6766,n6660,n4423);
nand (n6767,n6768,n6772);
or (n6768,n4021,n6769);
nor (n6769,n6770,n6771);
and (n6770,n3807,n5240);
and (n6771,n5241,n3808);
or (n6772,n4029,n6712);
and (n6773,n6752,n6759);
xor (n6774,n6649,n6664);
xor (n6775,n6709,n6723);
not (n6776,n6777);
or (n6777,n6778,n6814);
and (n6778,n6779,n6792);
xor (n6779,n6780,n6787);
nand (n6780,n6781,n6782);
or (n6781,n4387,n6718);
or (n6782,n4386,n6783);
not (n6783,n6784);
nor (n6784,n6785,n6786);
and (n6785,n4350,n3867);
and (n6786,n5193,n3873);
xor (n6787,n6788,n6789);
xor (n6788,n6724,n6730);
nor (n6789,n6790,n6791);
nand (n6790,n4035,n5241);
nand (n6791,n3863,n5233);
or (n6792,n6793,n6813);
and (n6793,n6794,n6806);
xor (n6794,n6795,n6802);
nand (n6795,n6796,n6801);
or (n6796,n4386,n6797);
not (n6797,n6798);
nor (n6798,n6799,n6800);
and (n6799,n5482,n3873);
and (n6800,n4406,n3867);
nand (n6801,n6784,n4384);
nand (n6802,n6803,n6805);
or (n6803,n6791,n6804);
not (n6804,n6790);
nand (n6805,n6804,n6791);
nand (n6806,n6807,n6812);
or (n6807,n4425,n6808);
not (n6808,n6809);
nor (n6809,n6810,n6811);
and (n6810,n4415,n4032);
and (n6811,n4413,n4031);
nand (n6812,n6762,n4423);
and (n6813,n6795,n6802);
and (n6814,n6780,n6787);
not (n6815,n6816);
nand (n6816,n6817,n6855);
or (n6817,n6818,n6821);
nor (n6818,n6819,n6820);
xor (n6819,n6779,n6792);
xor (n6820,n6751,n6767);
nor (n6821,n6822,n6853);
and (n6822,n6823,n6840);
nand (n6823,n6824,n6826);
not (n6824,n6825);
xor (n6825,n6794,n6806);
not (n6826,n6827);
or (n6827,n6828,n6839);
and (n6828,n6829,n6833);
xor (n6829,n6830,n6832);
nor (n6830,n6831,n3873);
and (n6831,n5233,n4384);
and (n6832,n4031,n5240,n4423);
nand (n6833,n6834,n6835);
or (n6834,n4426,n6808);
nand (n6835,n6836,n4424);
nor (n6836,n6837,n6838);
and (n6837,n5240,n4032);
and (n6838,n5241,n4031);
and (n6839,n6830,n6832);
or (n6840,n6841,n6852);
and (n6841,n6842,n6851);
xor (n6842,n6843,n6845);
and (n6843,n6831,n6844);
and (n6844,n5241,n4423);
nand (n6845,n6846,n6847);
or (n6846,n4387,n6797);
nand (n6847,n6848,n4385);
nand (n6848,n6849,n6850);
or (n6849,n3873,n5233);
or (n6850,n5235,n3867);
xor (n6851,n6829,n6833);
and (n6852,n6843,n6845);
not (n6853,n6854);
nand (n6854,n6825,n6827);
nand (n6855,n6819,n6820);
nand (n6856,n6747,n6777);
not (n6857,n6858);
nand (n6858,n6859,n6861);
not (n6859,n6860);
xor (n6860,n6705,n6736);
not (n6861,n6862);
or (n6862,n6863,n6864);
and (n6863,n6748,n6775);
and (n6864,n6749,n6774);
nand (n6865,n6860,n6862);
nand (n6866,n6641,n6703);
not (n6867,n6868);
nand (n6868,n6869,n6877);
not (n6869,n6870);
xor (n6870,n6871,n6876);
xor (n6871,n6872,n6875);
or (n6872,n6873,n6874);
and (n6873,n6673,n6701);
and (n6874,n6674,n6700);
xor (n6875,n6525,n6552);
xor (n6876,n6571,n6629);
not (n6877,n6878);
or (n6878,n6879,n6880);
and (n6879,n6642,n6672);
and (n6880,n6643,n6644);
nand (n6881,n6870,n6878);
nand (n6882,n6883,n6885);
not (n6883,n6884);
xor (n6884,n6567,n6631);
not (n6885,n6886);
or (n6886,n6887,n6888);
and (n6887,n6871,n6876);
and (n6888,n6872,n6875);
nand (n6889,n6561,n6890);
nor (n6890,n6883,n6885);
nand (n6891,n6563,n6565);
nand (n6892,n6286,n6476);
or (n6893,n6894,n6907);
xor (n6894,n6895,n6900);
xor (n6895,n6896,n6897);
xor (n6896,n6189,n6272);
or (n6897,n6898,n6899);
and (n6898,n6391,n6396);
and (n6899,n6392,n6395);
xor (n6900,n6901,n6904);
xor (n6901,n6902,n6903);
xor (n6902,n6091,n6121);
xor (n6903,n6145,n6148);
or (n6904,n6905,n6906);
and (n6905,n6384,n6389);
and (n6906,n6385,n6388);
or (n6907,n6908,n6909);
and (n6908,n6287,n6390);
and (n6909,n6288,n6383);
and (n6910,n6894,n6907);
nand (n6911,n6912,n6925);
nand (n6912,n6913,n6915);
not (n6913,n6914);
xor (n6914,n6138,n6276);
not (n6915,n6916);
or (n6916,n6917,n6924);
and (n6917,n6918,n6923);
xor (n6918,n6919,n6920);
xor (n6919,n6126,n6129);
or (n6920,n6921,n6922);
and (n6921,n6901,n6904);
and (n6922,n6902,n6903);
xor (n6923,n6142,n6274);
and (n6924,n6919,n6920);
or (n6925,n6926,n6927);
xor (n6926,n6918,n6923);
or (n6927,n6928,n6929);
and (n6928,n6895,n6900);
and (n6929,n6896,n6897);
nand (n6930,n6931,n6942);
or (n6931,n6932,n6935);
nand (n6932,n6933,n6934);
nand (n6933,n6024,n6025);
nand (n6934,n6135,n6136);
nor (n6935,n6936,n6134);
nand (n6936,n6937,n6912);
or (n6937,n6938,n6940);
not (n6938,n6939);
nand (n6939,n6926,n6927);
not (n6940,n6941);
nand (n6941,n6914,n6916);
not (n6942,n6023);
nand (n6943,n6944,n3495);
nand (n6944,n6945,n6953);
or (n6945,n6946,n5323);
not (n6946,n6947);
nand (n6947,n6948,n6951);
or (n6948,n6949,n6950);
not (n6949,n5823);
not (n6950,n5824);
or (n6951,n5822,n6952);
nand (n6952,n5839,n5841);
nand (n6953,n6954,n6955);
not (n6954,n5325);
nand (n6955,n6956,n6959);
or (n6956,n6957,n6958);
not (n6957,n5327);
not (n6958,n5326);
nand (n6959,n5652,n5653);
nor (n6960,n6961,n6973);
nand (n6961,n6962,n6968);
or (n6962,n6963,n6967);
not (n6963,n6964);
nor (n6964,n6965,n6966);
not (n6965,n5075);
not (n6966,n5209);
not (n6967,n3497);
nand (n6968,n6969,n4721,n6970);
not (n6969,n4620);
nand (n6970,n6971,n6972);
or (n6971,n3500,n4510);
nand (n6972,n4621,n4718);
nor (n6973,n6967,n6974);
nand (n6974,n6975,n6976);
not (n6975,n5074);
nor (n6976,n6977,n6978);
not (n6977,n5211);
not (n6978,n5212);
nor (n6979,n6980,n6994);
and (n6980,n6981,n4992);
nand (n6981,n6982,n6990);
or (n6982,n6983,n6984);
not (n6983,n4808);
not (n6984,n6985);
nand (n6985,n6986,n6987);
or (n6986,n4986,n4988);
or (n6987,n6988,n6989);
nand (n6988,n4724,n4727);
not (n6989,n4985);
nor (n6990,n6991,n6993);
and (n6991,n4810,n6992,n4880);
not (n6992,n4936);
and (n6993,n4937,n4940);
nand (n6994,n6995,n7000);
or (n6995,n6996,n6999);
nor (n6996,n6997,n6998);
and (n6997,n4994,n5030,n4997);
and (n6998,n5055,n5031);
not (n6999,n5058);
or (n7000,n5059,n5063);
nor (n7001,n7002,n7007);
and (n7002,n7003,n7006);
or (n7003,n7004,n7005);
and (n7004,n5065,n5070);
and (n7005,n5066,n5068);
not (n7006,n5068);
and (n7007,n7008,n5068);
not (n7008,n7003);
not (n7009,n7010);
nor (n7010,n7011,n10455);
and (n7011,n7012,n10454);
nand (n7012,n7013,n10403,n10420,n10432);
nand (n7013,n7014,n8918,n9580);
nand (n7014,n7015,n8913);
or (n7015,n7016,n8284);
not (n7016,n7017);
nor (n7017,n7018,n8143);
nor (n7018,n7019,n8038);
xor (n7019,n7020,n7830);
xor (n7020,n7021,n7671);
or (n7021,n7022,n7670);
and (n7022,n7023,n7396);
xor (n7023,n7024,n7272);
xor (n7024,n7025,n7196);
xor (n7025,n7026,n7112);
xor (n7026,n7027,n7086);
xor (n7027,n7028,n7058);
nand (n7028,n7029,n7051);
or (n7029,n7030,n7038);
not (n7030,n7031);
nor (n7031,n7032,n7037);
and (n7032,n7033,n7035);
not (n7033,n7034);
not (n7035,n7036);
and (n7037,n7034,n7036);
nand (n7038,n7039,n7046);
or (n7039,n7040,n7043);
not (n7040,n7041);
nand (n7041,n7035,n7042);
not (n7043,n7044);
nand (n7044,n7045,n7036);
not (n7045,n7042);
nor (n7046,n7047,n7050);
and (n7047,n7048,n7042);
not (n7048,n7049);
and (n7050,n7049,n7045);
nand (n7051,n7052,n7057);
nor (n7052,n7053,n7056);
and (n7053,n7054,n7035);
not (n7054,n7055);
and (n7056,n7055,n7036);
not (n7057,n7046);
nand (n7058,n7059,n7080);
or (n7059,n7060,n7068);
not (n7060,n7061);
nor (n7061,n7062,n7066);
and (n7062,n7063,n7065);
not (n7063,n7064);
and (n7066,n7064,n7067);
not (n7067,n7065);
not (n7068,n7069);
nor (n7069,n7070,n7075);
nor (n7070,n7071,n7073);
and (n7071,n7067,n7072);
and (n7073,n7065,n7074);
not (n7074,n7072);
nand (n7075,n7076,n7079);
or (n7076,n7077,n7072);
not (n7077,n7078);
nand (n7079,n7077,n7072);
nand (n7080,n7081,n7075);
nor (n7081,n7082,n7085);
and (n7082,n7083,n7065);
not (n7083,n7084);
and (n7085,n7084,n7067);
nand (n7086,n7087,n7104);
or (n7087,n7088,n7099);
nand (n7088,n7089,n7095);
nand (n7089,n7090,n7094);
or (n7090,n7091,n7092);
not (n7092,n7093);
nand (n7094,n7092,n7091);
nor (n7095,n7096,n7097);
and (n7096,n7067,n7091);
and (n7097,n7065,n7098);
not (n7098,n7091);
nor (n7099,n7100,n7103);
and (n7100,n7092,n7101);
not (n7101,n7102);
and (n7103,n7102,n7093);
or (n7104,n7105,n7095);
not (n7105,n7106);
nand (n7106,n7107,n7110);
not (n7107,n7108);
and (n7108,n7109,n7093);
nand (n7110,n7092,n7111);
not (n7111,n7109);
xor (n7112,n7113,n7167);
xor (n7113,n7114,n7140);
nand (n7114,n7115,n7131);
or (n7115,n7116,n7126);
not (n7116,n7117);
nand (n7117,n7118,n7125);
or (n7118,n7119,n7121);
not (n7119,n7120);
not (n7121,n7122);
nor (n7122,n7123,n7124);
nand (n7125,n7119,n7124,n7123);
not (n7126,n7127);
nand (n7127,n7128,n7130);
or (n7128,n7129,n7120);
nand (n7130,n7120,n7129);
nand (n7131,n7132,n7136);
nand (n7132,n7133,n7135);
or (n7133,n7134,n7120);
nand (n7135,n7120,n7134);
nand (n7136,n7137,n7139);
or (n7137,n7124,n7138);
not (n7138,n7123);
nand (n7139,n7138,n7124);
nand (n7140,n7141,n7160);
or (n7141,n7142,n7150);
not (n7142,n7143);
nor (n7143,n7144,n7148);
and (n7144,n7145,n7147);
not (n7145,n7146);
and (n7148,n7146,n7149);
not (n7149,n7147);
not (n7150,n7151);
nor (n7151,n7152,n7157);
nor (n7152,n7153,n7155);
and (n7153,n7149,n7154);
and (n7155,n7147,n7156);
not (n7156,n7154);
nand (n7157,n7158,n7159);
or (n7158,n7119,n7154);
nand (n7159,n7119,n7154);
nand (n7160,n7161,n7157);
not (n7161,n7162);
nor (n7162,n7163,n7166);
and (n7163,n7149,n7164);
not (n7164,n7165);
and (n7166,n7165,n7147);
nand (n7167,n7168,n7183);
or (n7168,n7169,n7176);
not (n7169,n7170);
nand (n7170,n7171,n7175);
or (n7171,n7172,n7174);
not (n7172,n7173);
nand (n7175,n7174,n7172);
not (n7176,n7177);
nand (n7177,n7178,n7182);
or (n7178,n7179,n7181);
not (n7179,n7180);
nand (n7182,n7179,n7181);
or (n7183,n7184,n7191);
not (n7184,n7185);
nor (n7185,n7186,n7177);
nor (n7186,n7187,n7189);
and (n7187,n7181,n7188);
not (n7188,n7174);
and (n7189,n7174,n7190);
not (n7190,n7181);
not (n7191,n7192);
nand (n7192,n7193,n7195);
or (n7193,n7194,n7188);
nand (n7195,n7188,n7194);
xor (n7196,n7197,n7245);
xor (n7197,n7198,n7227);
nand (n7198,n7199,n7219);
or (n7199,n7200,n7207);
not (n7200,n7201);
nand (n7201,n7202,n7206);
or (n7202,n7203,n7205);
not (n7203,n7204);
nand (n7206,n7205,n7203);
not (n7207,n7208);
and (n7208,n7209,n7214,n7216);
nand (n7209,n7210,n7213);
or (n7210,n7211,n7212);
not (n7211,n7205);
nand (n7213,n7211,n7212);
not (n7214,n7215);
and (n7215,n7212,n7188);
not (n7216,n7217);
and (n7217,n7218,n7174);
not (n7218,n7212);
nand (n7219,n7220,n7225);
nor (n7220,n7221,n7224);
and (n7221,n7222,n7211);
not (n7222,n7223);
and (n7224,n7223,n7205);
not (n7225,n7226);
nor (n7226,n7217,n7215);
nand (n7227,n7228,n7238);
or (n7228,n7229,n7235);
not (n7229,n7230);
nor (n7230,n7231,n7233);
and (n7231,n7232,n7138);
and (n7233,n7234,n7123);
not (n7234,n7232);
nand (n7235,n7123,n7236);
not (n7236,n7237);
nand (n7238,n7239,n7237);
nand (n7239,n7240,n7243);
not (n7240,n7241);
and (n7241,n7242,n7123);
nand (n7243,n7138,n7244);
not (n7244,n7242);
nand (n7245,n7246,n7263);
or (n7246,n7247,n7255);
not (n7247,n7248);
nor (n7248,n7249,n7254);
and (n7249,n7250,n7252);
not (n7250,n7251);
not (n7252,n7253);
and (n7254,n7251,n7253);
not (n7255,n7256);
nand (n7256,n7257,n7262);
or (n7257,n7211,n7258);
not (n7258,n7259);
nor (n7259,n7260,n7253);
not (n7260,n7261);
nand (n7262,n7253,n7211,n7260);
nand (n7263,n7264,n7267);
nand (n7264,n7265,n7266);
or (n7265,n7211,n7261);
nand (n7266,n7211,n7261);
nand (n7267,n7268,n7271);
or (n7268,n7269,n7253);
not (n7269,n7270);
nand (n7271,n7253,n7269);
or (n7272,n7273,n7395);
and (n7273,n7274,n7341);
xor (n7274,n7275,n7300);
xor (n7275,n7276,n7292);
xor (n7276,n7277,n7283);
nand (n7277,n7278,n7279);
or (n7278,n7236,n7229);
or (n7279,n7280,n7235);
nor (n7280,n7281,n7282);
and (n7281,n7134,n7123);
nor (n7282,n7123,n7134);
nand (n7283,n7284,n7291);
or (n7284,n7285,n7255);
not (n7285,n7286);
nor (n7286,n7287,n7290);
and (n7287,n7288,n7252);
not (n7288,n7289);
and (n7290,n7289,n7253);
nand (n7291,n7248,n7264);
nand (n7292,n7293,n7298);
or (n7293,n7116,n7294);
not (n7294,n7295);
nand (n7295,n7296,n7297);
or (n7296,n7165,n7120);
nand (n7297,n7120,n7165);
or (n7298,n7299,n7126);
not (n7299,n7136);
xor (n7300,n7301,n7319);
xor (n7301,n7302,n7312);
nand (n7302,n7303,n7311);
or (n7303,n7304,n7150);
not (n7304,n7305);
nand (n7305,n7306,n7309);
not (n7306,n7307);
and (n7307,n7308,n7147);
nand (n7309,n7149,n7310);
not (n7310,n7308);
nand (n7311,n7143,n7157);
nand (n7312,n7313,n7318);
or (n7313,n7314,n7184);
not (n7314,n7315);
nand (n7315,n7316,n7317);
or (n7316,n7222,n7174);
nand (n7317,n7174,n7222);
nand (n7318,n7192,n7177);
nand (n7319,n7320,n7335);
or (n7320,n7321,n7325);
not (n7321,n7322);
nor (n7322,n7323,n7324);
and (n7323,n7054,n7048);
and (n7324,n7055,n7049);
nand (n7325,n7326,n7332);
not (n7326,n7327);
nand (n7327,n7328,n7331);
or (n7328,n7329,n7253);
not (n7329,n7330);
nand (n7331,n7329,n7253);
nand (n7332,n7333,n7334);
or (n7333,n7329,n7049);
nand (n7334,n7049,n7329);
nand (n7335,n7336,n7327);
nand (n7336,n7337,n7340);
or (n7337,n7049,n7338);
not (n7338,n7339);
nand (n7340,n7049,n7338);
xor (n7341,n7342,n7359);
xor (n7342,n7343,n7350);
nand (n7343,n7344,n7348);
or (n7344,n7068,n7345);
nor (n7345,n7346,n7347);
and (n7346,n7067,n7111);
and (n7347,n7109,n7065);
or (n7348,n7349,n7060);
not (n7349,n7075);
nand (n7350,n7351,n7358);
or (n7351,n7352,n7088);
not (n7352,n7353);
nand (n7353,n7354,n7356);
or (n7354,n7093,n7355);
not (n7356,n7357);
and (n7357,n7355,n7093);
or (n7358,n7099,n7095);
xor (n7359,n7360,n7375);
xor (n7360,n7361,n7369);
nor (n7361,n7362,n7035);
and (n7362,n7363,n7367);
nand (n7363,n7364,n7048);
not (n7364,n7365);
and (n7365,n7366,n7042);
nand (n7367,n7368,n7045);
not (n7368,n7366);
nor (n7369,n7370,n7093);
nor (n7370,n7371,n7373);
and (n7371,n7065,n7372);
nand (n7372,n7098,n7355);
and (n7373,n7374,n7091);
not (n7374,n7355);
nand (n7375,n7376,n7387);
or (n7376,n7377,n7379);
not (n7377,n7378);
not (n7379,n7380);
nor (n7380,n7381,n7386);
and (n7381,n7382,n7384);
not (n7382,n7383);
not (n7384,n7385);
and (n7386,n7383,n7385);
nand (n7387,n7388,n7393);
nor (n7388,n7389,n7392);
and (n7389,n7390,n7384);
not (n7390,n7391);
and (n7392,n7391,n7385);
not (n7393,n7394);
nand (n7394,n7385,n7377);
and (n7395,n7275,n7300);
or (n7396,n7397,n7669);
and (n7397,n7398,n7609);
xor (n7398,n7399,n7501);
or (n7399,n7400,n7500);
and (n7400,n7401,n7444);
xor (n7401,n7402,n7409);
nand (n7402,n7403,n7408);
or (n7403,n7184,n7404);
not (n7404,n7405);
nand (n7405,n7406,n7407);
or (n7406,n7204,n7188);
or (n7407,n7174,n7203);
or (n7408,n7176,n7314);
or (n7409,n7410,n7443);
and (n7410,n7411,n7431);
xor (n7411,n7412,n7422);
nand (n7412,n7413,n7418);
or (n7413,n7414,n7207);
not (n7414,n7415);
nor (n7415,n7416,n7417);
and (n7416,n7288,n7211);
and (n7417,n7289,n7205);
nand (n7418,n7225,n7419);
nand (n7419,n7420,n7421);
or (n7420,n7251,n7211);
nand (n7421,n7211,n7251);
nand (n7422,n7423,n7427);
or (n7423,n7235,n7424);
or (n7424,n7425,n7426);
and (n7425,n7165,n7138);
and (n7426,n7164,n7123);
or (n7427,n7428,n7236);
nor (n7428,n7429,n7430);
and (n7429,n7129,n7123);
nor (n7430,n7123,n7129);
nand (n7431,n7432,n7437);
or (n7432,n7433,n7299);
not (n7433,n7434);
nand (n7434,n7435,n7436);
or (n7435,n7146,n7120);
nand (n7436,n7120,n7146);
or (n7437,n7116,n7438);
not (n7438,n7439);
nand (n7439,n7440,n7442);
not (n7440,n7441);
and (n7441,n7308,n7120);
nand (n7442,n7119,n7310);
and (n7443,n7412,n7422);
or (n7444,n7445,n7499);
and (n7445,n7446,n7473);
xor (n7446,n7447,n7457);
nand (n7447,n7448,n7453);
or (n7448,n7449,n7255);
not (n7449,n7450);
nor (n7450,n7451,n7452);
and (n7451,n7054,n7252);
and (n7452,n7055,n7253);
nand (n7453,n7264,n7454);
nor (n7454,n7455,n7456);
and (n7455,n7338,n7252);
and (n7456,n7339,n7253);
nand (n7457,n7458,n7466);
or (n7458,n7150,n7459);
not (n7459,n7460);
nand (n7460,n7461,n7464);
not (n7461,n7462);
and (n7462,n7463,n7147);
nand (n7464,n7149,n7465);
not (n7465,n7463);
or (n7466,n7467,n7468);
not (n7467,n7157);
nor (n7468,n7469,n7472);
and (n7469,n7149,n7470);
not (n7470,n7471);
and (n7472,n7471,n7147);
nand (n7473,n7474,n7492);
or (n7474,n7475,n7487);
nand (n7475,n7476,n7481);
not (n7476,n7477);
nand (n7477,n7478,n7480);
or (n7478,n7149,n7479);
nand (n7480,n7149,n7479);
nand (n7481,n7482,n7485);
nand (n7482,n7483,n7484);
not (n7484,n7479);
nand (n7485,n7486,n7479);
not (n7486,n7483);
not (n7487,n7488);
nand (n7488,n7489,n7491);
not (n7489,n7490);
and (n7490,n7084,n7483);
nand (n7491,n7486,n7083);
or (n7492,n7476,n7493);
not (n7493,n7494);
nor (n7494,n7495,n7498);
and (n7495,n7496,n7483);
not (n7496,n7497);
and (n7498,n7497,n7486);
and (n7499,n7447,n7457);
and (n7500,n7402,n7409);
or (n7501,n7502,n7608);
and (n7502,n7503,n7570);
xor (n7503,n7504,n7545);
or (n7504,n7505,n7544);
and (n7505,n7506,n7536);
xor (n7506,n7507,n7517);
nand (n7507,n7508,n7513);
or (n7508,n7509,n7325);
not (n7509,n7510);
nand (n7510,n7511,n7512);
or (n7511,n7049,n7368);
nand (n7512,n7368,n7049);
nand (n7513,n7514,n7327);
nand (n7514,n7515,n7516);
or (n7515,n7034,n7048);
nand (n7516,n7034,n7048);
nand (n7517,n7518,n7532);
or (n7518,n7519,n7523);
not (n7519,n7520);
nor (n7520,n7521,n7522);
and (n7521,n7111,n7078);
and (n7522,n7109,n7077);
nand (n7523,n7524,n7529);
not (n7524,n7525);
nand (n7525,n7526,n7528);
or (n7526,n7486,n7527);
nand (n7528,n7486,n7527);
nand (n7529,n7530,n7531);
or (n7530,n7527,n7077);
nand (n7531,n7077,n7527);
nand (n7532,n7525,n7533);
nand (n7533,n7534,n7535);
or (n7534,n7064,n7078);
nand (n7535,n7078,n7064);
nand (n7536,n7537,n7540);
or (n7537,n7349,n7538);
not (n7538,n7539);
xor (n7539,n7101,n7065);
or (n7540,n7068,n7541);
nor (n7541,n7542,n7543);
and (n7542,n7067,n7374);
and (n7543,n7355,n7065);
and (n7544,n7507,n7517);
or (n7545,n7546,n7569);
and (n7546,n7547,n7566);
xor (n7547,n7548,n7560);
nand (n7548,n7549,n7554);
or (n7549,n7550,n7394);
not (n7550,n7551);
nand (n7551,n7552,n7553);
or (n7552,n7173,n7384);
nand (n7553,n7384,n7173);
nand (n7554,n7555,n7378);
nor (n7555,n7556,n7559);
and (n7556,n7557,n7384);
not (n7557,n7558);
and (n7559,n7558,n7385);
nand (n7560,n7561,n7565);
or (n7561,n7184,n7562);
nor (n7562,n7563,n7564);
and (n7563,n7270,n7188);
and (n7564,n7269,n7174);
nand (n7565,n7177,n7405);
and (n7566,n7567,n7568);
and (n7567,n7075,n7355);
and (n7568,n7327,n7366);
and (n7569,n7548,n7560);
or (n7570,n7571,n7607);
and (n7571,n7572,n7585);
xor (n7572,n7573,n7580);
nor (n7573,n7574,n7048);
and (n7574,n7575,n7578);
not (n7575,n7576);
nor (n7576,n7577,n7253);
and (n7577,n7366,n7330);
not (n7578,n7579);
nor (n7579,n7366,n7330);
and (n7580,n7581,n7067);
nand (n7581,n7582,n7583);
or (n7582,n7074,n7355);
nand (n7583,n7584,n7078);
or (n7584,n7072,n7374);
nand (n7585,n7586,n7602);
or (n7586,n7587,n7591);
not (n7587,n7588);
nor (n7588,n7589,n7590);
and (n7589,n7222,n7179);
and (n7590,n7223,n7180);
nand (n7591,n7592,n7599);
or (n7592,n7593,n7596);
not (n7593,n7594);
nand (n7594,n7179,n7595);
not (n7596,n7597);
nand (n7597,n7598,n7180);
not (n7598,n7595);
nor (n7599,n7600,n7601);
and (n7600,n7598,n7385);
and (n7601,n7384,n7595);
nand (n7602,n7603,n7604);
not (n7603,n7599);
nand (n7604,n7605,n7606);
or (n7605,n7194,n7179);
nand (n7606,n7179,n7194);
and (n7607,n7573,n7580);
and (n7608,n7504,n7545);
xor (n7609,n7610,n7646);
xor (n7610,n7611,n7632);
or (n7611,n7612,n7631);
and (n7612,n7613,n7628);
xor (n7613,n7614,n7621);
nand (n7614,n7615,n7617);
or (n7615,n7616,n7591);
not (n7616,n7604);
nand (n7617,n7618,n7603);
nand (n7618,n7619,n7620);
or (n7619,n7173,n7179);
nand (n7620,n7179,n7173);
nand (n7621,n7622,n7624);
or (n7622,n7207,n7623);
not (n7623,n7419);
nand (n7624,n7625,n7225);
nand (n7625,n7626,n7627);
or (n7626,n7269,n7205);
nand (n7627,n7205,n7269);
nand (n7628,n7629,n7630);
or (n7629,n7428,n7235);
or (n7630,n7280,n7236);
and (n7631,n7614,n7621);
or (n7632,n7633,n7645);
and (n7633,n7634,n7642);
xor (n7634,n7635,n7638);
nand (n7635,n7636,n7637);
or (n7636,n7116,n7433);
nand (n7637,n7295,n7136);
nand (n7638,n7639,n7641);
or (n7639,n7640,n7255);
not (n7640,n7454);
nand (n7641,n7286,n7264);
nand (n7642,n7643,n7644);
or (n7643,n7304,n7467);
or (n7644,n7150,n7468);
and (n7645,n7635,n7638);
or (n7646,n7647,n7668);
and (n7647,n7648,n7660);
xor (n7648,n7649,n7656);
nand (n7649,n7650,n7651);
or (n7650,n7493,n7475);
nand (n7651,n7477,n7652);
nand (n7652,n7653,n7655);
not (n7653,n7654);
and (n7654,n7463,n7483);
nand (n7655,n7486,n7465);
nand (n7656,n7657,n7659);
or (n7657,n7325,n7658);
not (n7658,n7514);
nand (n7659,n7322,n7327);
nand (n7660,n7661,n7666);
or (n7661,n7662,n7524);
not (n7662,n7663);
nor (n7663,n7664,n7665);
and (n7664,n7083,n7078);
and (n7665,n7084,n7077);
or (n7666,n7523,n7667);
not (n7667,n7533);
and (n7668,n7649,n7656);
and (n7669,n7399,n7501);
and (n7670,n7024,n7272);
or (n7671,n7672,n7829);
and (n7672,n7673,n7816);
xor (n7673,n7674,n7712);
xor (n7674,n7675,n7709);
xor (n7675,n7676,n7706);
xor (n7676,n7677,n7696);
xor (n7677,n7678,n7685);
nand (n7678,n7679,n7681);
or (n7679,n7325,n7680);
not (n7680,n7336);
nand (n7681,n7682,n7327);
nand (n7682,n7683,n7684);
or (n7683,n7049,n7288);
or (n7684,n7048,n7289);
nand (n7685,n7686,n7692);
or (n7686,n7475,n7687);
not (n7687,n7688);
nand (n7688,n7689,n7691);
not (n7689,n7690);
and (n7690,n7471,n7483);
nand (n7691,n7486,n7470);
nand (n7692,n7477,n7693);
nor (n7693,n7694,n7695);
and (n7694,n7310,n7483);
and (n7695,n7308,n7486);
nand (n7696,n7697,n7702);
or (n7697,n7523,n7698);
not (n7698,n7699);
nor (n7699,n7700,n7701);
and (n7700,n7497,n7077);
and (n7701,n7496,n7078);
or (n7702,n7524,n7703);
nor (n7703,n7704,n7705);
and (n7704,n7465,n7077);
and (n7705,n7463,n7078);
or (n7706,n7707,n7708);
and (n7707,n7610,n7646);
and (n7708,n7611,n7632);
or (n7709,n7710,n7711);
and (n7710,n7342,n7359);
and (n7711,n7343,n7350);
xor (n7712,n7713,n7794);
xor (n7713,n7714,n7770);
xor (n7714,n7715,n7737);
xor (n7715,n7716,n7719);
or (n7716,n7717,n7718);
and (n7717,n7301,n7319);
and (n7718,n7302,n7312);
or (n7719,n7720,n7736);
and (n7720,n7721,n7729);
xor (n7721,n7722,n7726);
nand (n7722,n7723,n7725);
or (n7723,n7724,n7475);
not (n7724,n7652);
nand (n7725,n7688,n7477);
nand (n7726,n7727,n7728);
or (n7727,n7662,n7523);
nand (n7728,n7699,n7525);
nand (n7729,n7730,n7735);
or (n7730,n7731,n7038);
not (n7731,n7732);
nand (n7732,n7733,n7734);
or (n7733,n7035,n7366);
or (n7734,n7368,n7036);
nand (n7735,n7057,n7031);
and (n7736,n7722,n7726);
xor (n7737,n7738,n7760);
xor (n7738,n7739,n7747);
nand (n7739,n7740,n7741);
or (n7740,n7394,n7379);
nand (n7741,n7742,n7378);
nand (n7742,n7743,n7746);
or (n7743,n7744,n7385);
not (n7744,n7745);
nand (n7746,n7385,n7744);
xor (n7747,n7748,n7755);
and (n7748,n7749,n7355);
not (n7749,n7750);
nor (n7750,n7751,n7754);
and (n7751,n7093,n7752);
not (n7752,n7753);
and (n7754,n7092,n7753);
and (n7755,n7756,n7366);
nand (n7756,n7757,n7759);
or (n7757,n7758,n7035);
nand (n7759,n7035,n7758);
nand (n7760,n7761,n7766);
or (n7761,n7762,n7591);
not (n7762,n7763);
nand (n7763,n7764,n7765);
or (n7764,n7557,n7180);
nand (n7765,n7180,n7557);
nand (n7766,n7603,n7767);
nor (n7767,n7768,n7769);
and (n7768,n7390,n7179);
and (n7769,n7391,n7180);
xor (n7770,n7771,n7791);
xor (n7771,n7772,n7775);
or (n7772,n7773,n7774);
and (n7773,n7360,n7375);
and (n7774,n7361,n7369);
or (n7775,n7776,n7790);
and (n7776,n7777,n7786);
xor (n7777,n7778,n7782);
nand (n7778,n7779,n7780);
or (n7779,n7599,n7762);
or (n7780,n7591,n7781);
not (n7781,n7618);
nand (n7782,n7783,n7785);
or (n7783,n7784,n7207);
not (n7784,n7625);
nand (n7785,n7225,n7201);
nor (n7786,n7787,n7789);
nand (n7787,n7788,n7355);
not (n7788,n7095);
nand (n7789,n7057,n7366);
and (n7790,n7778,n7782);
or (n7791,n7792,n7793);
and (n7792,n7276,n7292);
and (n7793,n7277,n7283);
or (n7794,n7795,n7815);
and (n7795,n7796,n7814);
xor (n7796,n7797,n7813);
or (n7797,n7798,n7812);
and (n7798,n7799,n7807);
xor (n7799,n7800,n7804);
nand (n7800,n7801,n7803);
or (n7801,n7802,n7787);
not (n7802,n7789);
nand (n7803,n7802,n7787);
nand (n7804,n7805,n7806);
or (n7805,n7538,n7068);
or (n7806,n7345,n7349);
nand (n7807,n7808,n7810);
or (n7808,n7394,n7809);
not (n7809,n7555);
or (n7810,n7811,n7377);
not (n7811,n7388);
and (n7812,n7800,n7804);
xor (n7813,n7777,n7786);
xor (n7814,n7721,n7729);
and (n7815,n7797,n7813);
or (n7816,n7817,n7828);
and (n7817,n7818,n7827);
xor (n7818,n7819,n7826);
or (n7819,n7820,n7825);
and (n7820,n7821,n7824);
xor (n7821,n7822,n7823);
xor (n7822,n7648,n7660);
xor (n7823,n7799,n7807);
xor (n7824,n7613,n7628);
and (n7825,n7822,n7823);
xor (n7826,n7796,n7814);
xor (n7827,n7274,n7341);
and (n7828,n7819,n7826);
and (n7829,n7674,n7712);
xor (n7830,n7831,n7963);
xor (n7831,n7832,n7944);
xor (n7832,n7833,n7875);
xor (n7833,n7834,n7872);
xor (n7834,n7835,n7869);
xor (n7835,n7836,n7843);
nand (n7836,n7837,n7839);
or (n7837,n7068,n7838);
not (n7838,n7081);
or (n7839,n7349,n7840);
nor (n7840,n7841,n7842);
and (n7841,n7067,n7496);
and (n7842,n7497,n7065);
xor (n7843,n7844,n7860);
xor (n7844,n7845,n7854);
nor (n7845,n7846,n7852);
and (n7846,n7847,n7850);
nand (n7847,n7848,n7035);
not (n7848,n7849);
and (n7849,n7366,n7758);
nand (n7850,n7368,n7851);
not (n7851,n7758);
not (n7852,n7853);
nor (n7854,n7855,n7859);
and (n7855,n7856,n7858);
nand (n7856,n7857,n7093);
or (n7857,n7753,n7374);
nand (n7858,n7374,n7753);
nand (n7860,n7861,n7863);
or (n7861,n7394,n7862);
not (n7862,n7742);
nand (n7863,n7864,n7378);
nand (n7864,n7865,n7868);
or (n7865,n7866,n7385);
not (n7866,n7867);
nand (n7868,n7385,n7866);
or (n7869,n7870,n7871);
and (n7870,n7738,n7760);
and (n7871,n7739,n7747);
or (n7872,n7873,n7874);
and (n7873,n7025,n7196);
and (n7874,n7026,n7112);
xor (n7875,n7876,n7927);
xor (n7876,n7877,n7902);
xor (n7877,n7878,n7893);
xor (n7878,n7879,n7886);
nand (n7879,n7880,n7882);
or (n7880,n7881,n7475);
not (n7881,n7693);
nand (n7882,n7477,n7883);
nand (n7883,n7884,n7885);
or (n7884,n7146,n7483);
nand (n7885,n7483,n7146);
nand (n7886,n7887,n7889);
or (n7887,n7888,n7038);
not (n7888,n7052);
nand (n7889,n7890,n7057);
nor (n7890,n7891,n7892);
and (n7891,n7338,n7035);
and (n7892,n7339,n7036);
nand (n7893,n7894,n7899);
or (n7894,n7895,n7524);
not (n7895,n7896);
nor (n7896,n7897,n7898);
and (n7897,n7470,n7078);
and (n7898,n7471,n7077);
nand (n7899,n7900,n7901);
not (n7900,n7703);
not (n7901,n7523);
xor (n7902,n7903,n7920);
xor (n7903,n7904,n7911);
nand (n7904,n7905,n7907);
or (n7905,n7906,n7255);
not (n7906,n7267);
nand (n7907,n7908,n7264);
nand (n7908,n7909,n7910);
or (n7909,n7203,n7253);
nand (n7910,n7253,n7203);
nand (n7911,n7912,n7914);
or (n7912,n7235,n7913);
not (n7913,n7239);
or (n7914,n7915,n7236);
nor (n7915,n7916,n7918);
and (n7916,n7917,n7123);
and (n7918,n7919,n7138);
not (n7919,n7917);
nand (n7920,n7921,n7923);
or (n7921,n7116,n7922);
not (n7922,n7132);
or (n7923,n7299,n7924);
nor (n7924,n7925,n7926);
and (n7925,n7234,n7119);
and (n7926,n7232,n7120);
xor (n7927,n7928,n7943);
xor (n7928,n7929,n7936);
nand (n7929,n7930,n7932);
or (n7930,n7931,n7591);
not (n7931,n7767);
nand (n7932,n7933,n7603);
nand (n7933,n7934,n7935);
or (n7934,n7383,n7179);
nand (n7935,n7179,n7383);
nand (n7936,n7937,n7939);
or (n7937,n7938,n7207);
not (n7938,n7220);
nand (n7939,n7225,n7940);
nand (n7940,n7941,n7942);
or (n7941,n7194,n7211);
nand (n7942,n7211,n7194);
and (n7943,n7748,n7755);
xor (n7944,n7945,n7952);
xor (n7945,n7946,n7949);
or (n7946,n7947,n7948);
and (n7947,n7771,n7791);
and (n7948,n7772,n7775);
or (n7949,n7950,n7951);
and (n7950,n7715,n7737);
and (n7951,n7716,n7719);
xor (n7952,n7953,n7960);
xor (n7953,n7954,n7957);
or (n7954,n7955,n7956);
and (n7955,n7197,n7245);
and (n7956,n7198,n7227);
or (n7957,n7958,n7959);
and (n7958,n7113,n7167);
and (n7959,n7114,n7140);
or (n7960,n7961,n7962);
and (n7961,n7677,n7696);
and (n7962,n7678,n7685);
xor (n7963,n7964,n8035);
xor (n7964,n7965,n8032);
xor (n7965,n7966,n8010);
xor (n7966,n7967,n7970);
or (n7967,n7968,n7969);
and (n7968,n7027,n7086);
and (n7969,n7028,n7058);
xor (n7970,n7971,n7996);
xor (n7971,n7972,n7988);
nand (n7972,n7973,n7984);
or (n7973,n7974,n7978);
not (n7974,n7975);
nor (n7975,n7976,n7977);
and (n7976,n7368,n7852);
and (n7977,n7366,n7853);
not (n7978,n7979);
nor (n7979,n7980,n7982);
and (n7980,n7035,n7981);
nand (n7981,n7851,n7853);
and (n7982,n7036,n7983);
nand (n7983,n7758,n7852);
nand (n7984,n7756,n7985);
nand (n7985,n7986,n7987);
or (n7986,n7034,n7852);
nand (n7987,n7852,n7034);
nand (n7988,n7989,n7995);
or (n7989,n7095,n7990);
not (n7990,n7991);
nand (n7991,n7992,n7994);
not (n7992,n7993);
and (n7993,n7064,n7093);
nand (n7994,n7092,n7063);
nand (n7995,n7106,n7089,n7095);
nand (n7996,n7997,n8006);
or (n7997,n7998,n8003);
nand (n7998,n7750,n7999);
nor (n7999,n8000,n8001);
and (n8000,n7859,n7753);
and (n8001,n8002,n7752);
not (n8002,n7859);
nor (n8003,n8004,n8005);
and (n8004,n7374,n8002);
and (n8005,n7355,n7859);
or (n8006,n8007,n7750);
nor (n8007,n8008,n8009);
and (n8008,n7102,n7859);
and (n8009,n7101,n8002);
xor (n8010,n8011,n8025);
xor (n8011,n8012,n8018);
nand (n8012,n8013,n8014);
or (n8013,n7169,n7184);
nand (n8014,n8015,n7177);
nand (n8015,n8016,n8017);
or (n8016,n7557,n7174);
nand (n8017,n7174,n7557);
nand (n8018,n8019,n8021);
or (n8019,n8020,n7325);
not (n8020,n7682);
nand (n8021,n7327,n8022);
nand (n8022,n8023,n8024);
or (n8023,n7251,n7048);
nand (n8024,n7251,n7048);
nand (n8025,n8026,n8031);
or (n8026,n8027,n7467);
not (n8027,n8028);
nand (n8028,n8029,n8030);
or (n8029,n7129,n7147);
nand (n8030,n7147,n7129);
or (n8031,n7150,n7162);
or (n8032,n8033,n8034);
and (n8033,n7675,n7709);
and (n8034,n7676,n7706);
or (n8035,n8036,n8037);
and (n8036,n7713,n7794);
and (n8037,n7714,n7770);
or (n8038,n8039,n8142);
and (n8039,n8040,n8141);
xor (n8040,n8041,n8042);
xor (n8041,n7023,n7396);
or (n8042,n8043,n8140);
and (n8043,n8044,n8133);
xor (n8044,n8045,n8046);
xor (n8045,n7398,n7609);
or (n8046,n8047,n8132);
and (n8047,n8048,n8099);
xor (n8048,n8049,n8050);
xor (n8049,n7634,n7642);
or (n8050,n8051,n8098);
and (n8051,n8052,n8073);
xor (n8052,n8053,n8054);
xor (n8053,n7572,n7585);
or (n8054,n8055,n8072);
and (n8055,n8056,n8065);
xor (n8056,n8057,n8064);
nand (n8057,n8058,n8063);
or (n8058,n8059,n7591);
not (n8059,n8060);
nor (n8060,n8061,n8062);
and (n8061,n7203,n7179);
and (n8062,n7204,n7180);
nand (n8063,n7603,n7588);
xor (n8064,n7567,n7568);
nand (n8065,n8066,n8071);
or (n8066,n7207,n8067);
not (n8067,n8068);
nand (n8068,n8069,n8070);
or (n8069,n7338,n7205);
nand (n8070,n7205,n7338);
or (n8071,n7226,n7414);
and (n8072,n8057,n8064);
or (n8073,n8074,n8097);
and (n8074,n8075,n8090);
xor (n8075,n8076,n8083);
nand (n8076,n8077,n8082);
or (n8077,n8078,n7116);
not (n8078,n8079);
nand (n8079,n8080,n8081);
or (n8080,n7471,n7120);
nand (n8081,n7120,n7471);
nand (n8082,n7439,n7136);
nand (n8083,n8084,n8089);
or (n8084,n8085,n7150);
not (n8085,n8086);
nor (n8086,n8087,n8088);
and (n8087,n7496,n7147);
and (n8088,n7497,n7149);
nand (n8089,n7460,n7157);
nand (n8090,n8091,n8096);
or (n8091,n8092,n7255);
not (n8092,n8093);
nand (n8093,n8094,n8095);
or (n8094,n7034,n7252);
nand (n8095,n7034,n7252);
nand (n8096,n7264,n7450);
and (n8097,n8076,n8083);
and (n8098,n8053,n8054);
or (n8099,n8100,n8131);
and (n8100,n8101,n8130);
xor (n8101,n8102,n8129);
or (n8102,n8103,n8128);
and (n8103,n8104,n8120);
xor (n8104,n8105,n8113);
nand (n8105,n8106,n8112);
or (n8106,n8107,n7475);
not (n8107,n8108);
nand (n8108,n8109,n8111);
not (n8109,n8110);
and (n8110,n7064,n7483);
nand (n8111,n7486,n7063);
nand (n8112,n7477,n7488);
nand (n8113,n8114,n8119);
or (n8114,n8115,n7523);
not (n8115,n8116);
nor (n8116,n8117,n8118);
and (n8117,n7102,n7077);
and (n8118,n7101,n7078);
nand (n8119,n7525,n7520);
nand (n8120,n8121,n8127);
or (n8121,n8122,n7394);
not (n8122,n8123);
nor (n8123,n8124,n8126);
and (n8124,n8125,n7384);
not (n8125,n7194);
and (n8126,n7194,n7385);
nand (n8127,n7551,n7378);
and (n8128,n8105,n8113);
xor (n8129,n7547,n7566);
xor (n8130,n7411,n7431);
and (n8131,n8102,n8129);
and (n8132,n8049,n8050);
or (n8133,n8134,n8139);
and (n8134,n8135,n8138);
xor (n8135,n8136,n8137);
xor (n8136,n7503,n7570);
xor (n8137,n7401,n7444);
xor (n8138,n7821,n7824);
and (n8139,n8136,n8137);
and (n8140,n8045,n8046);
xor (n8141,n7673,n7816);
and (n8142,n8041,n8042);
nor (n8143,n8144,n8145);
xor (n8144,n8040,n8141);
or (n8145,n8146,n8283);
and (n8146,n8147,n8282);
xor (n8147,n8148,n8149);
xor (n8148,n7818,n7827);
or (n8149,n8150,n8281);
and (n8150,n8151,n8280);
xor (n8151,n8152,n8195);
or (n8152,n8153,n8194);
and (n8153,n8154,n8157);
xor (n8154,n8155,n8156);
xor (n8155,n7446,n7473);
xor (n8156,n7506,n7536);
or (n8157,n8158,n8193);
and (n8158,n8159,n8173);
xor (n8159,n8160,n8167);
nand (n8160,n8161,n8166);
or (n8161,n8162,n7184);
not (n8162,n8163);
nor (n8163,n8164,n8165);
and (n8164,n7250,n7188);
and (n8165,n7251,n7174);
or (n8166,n7176,n7562);
nand (n8167,n8168,n8172);
or (n8168,n7235,n8169);
nor (n8169,n8170,n8171);
and (n8170,n7138,n7145);
and (n8171,n7146,n7123);
or (n8172,n7424,n7236);
or (n8173,n8174,n8192);
and (n8174,n8175,n8189);
xor (n8175,n8176,n8182);
nand (n8176,n8177,n8178);
or (n8177,n7377,n8122);
nand (n8178,n8179,n7393);
nor (n8179,n8180,n8181);
and (n8180,n7384,n7222);
and (n8181,n7223,n7385);
nand (n8182,n8183,n8188);
or (n8183,n8184,n7184);
not (n8184,n8185);
nor (n8185,n8186,n8187);
and (n8186,n7288,n7188);
and (n8187,n7289,n7174);
nand (n8188,n8163,n7177);
and (n8189,n8190,n8191);
and (n8190,n7525,n7355);
and (n8191,n7264,n7366);
and (n8192,n8176,n8182);
and (n8193,n8160,n8167);
and (n8194,n8155,n8156);
or (n8195,n8196,n8279);
and (n8196,n8197,n8278);
xor (n8197,n8198,n8271);
or (n8198,n8199,n8270);
and (n8199,n8200,n8247);
xor (n8200,n8201,n8225);
or (n8201,n8202,n8224);
and (n8202,n8203,n8218);
xor (n8203,n8204,n8211);
nand (n8204,n8205,n8210);
or (n8205,n8206,n7255);
not (n8206,n8207);
nor (n8207,n8208,n8209);
and (n8208,n7368,n7252);
and (n8209,n7366,n7253);
nand (n8210,n7264,n8093);
nand (n8211,n8212,n8217);
or (n8212,n8213,n7475);
not (n8213,n8214);
nand (n8214,n8215,n8216);
or (n8215,n7109,n7483);
nand (n8216,n7483,n7109);
nand (n8217,n7477,n8108);
nand (n8218,n8219,n8223);
or (n8219,n7523,n8220);
nor (n8220,n8221,n8222);
and (n8221,n7077,n7374);
and (n8222,n7355,n7078);
nand (n8223,n7525,n8116);
and (n8224,n8204,n8211);
or (n8225,n8226,n8246);
and (n8226,n8227,n8239);
xor (n8227,n8228,n8233);
nor (n8228,n8229,n7252);
nor (n8229,n8230,n8231);
and (n8230,n7368,n7260);
nor (n8231,n8232,n7205);
and (n8232,n7366,n7261);
and (n8233,n8234,n7077);
nand (n8234,n8235,n8237);
or (n8235,n7355,n8236);
not (n8236,n7527);
nand (n8237,n8238,n7483);
or (n8238,n7527,n7374);
nand (n8239,n8240,n8245);
or (n8240,n8241,n7591);
not (n8241,n8242);
nor (n8242,n8243,n8244);
and (n8243,n7269,n7179);
and (n8244,n7270,n7180);
nand (n8245,n8060,n7603);
and (n8246,n8228,n8233);
or (n8247,n8248,n8269);
and (n8248,n8249,n8263);
xor (n8249,n8250,n8257);
nand (n8250,n8251,n8256);
or (n8251,n7207,n8252);
not (n8252,n8253);
nand (n8253,n8254,n8255);
or (n8254,n7055,n7211);
nand (n8255,n7211,n7055);
nand (n8256,n7225,n8068);
nand (n8257,n8258,n8259);
or (n8258,n8078,n7299);
or (n8259,n7116,n8260);
nor (n8260,n8261,n8262);
and (n8261,n7119,n7465);
and (n8262,n7463,n7120);
nand (n8263,n8264,n8268);
or (n8264,n7150,n8265);
nor (n8265,n8266,n8267);
and (n8266,n7149,n7083);
and (n8267,n7084,n7147);
or (n8268,n7467,n8085);
and (n8269,n8250,n8257);
and (n8270,n8201,n8225);
or (n8271,n8272,n8277);
and (n8272,n8273,n8276);
xor (n8273,n8274,n8275);
xor (n8274,n8104,n8120);
xor (n8275,n8075,n8090);
xor (n8276,n8056,n8065);
and (n8277,n8274,n8275);
xor (n8278,n8052,n8073);
and (n8279,n8198,n8271);
xor (n8280,n8048,n8099);
and (n8281,n8152,n8195);
xor (n8282,n8044,n8133);
and (n8283,n8148,n8149);
not (n8284,n8285);
nand (n8285,n8286,n8907);
or (n8286,n8287,n8487);
not (n8287,n8288);
nor (n8288,n8289,n8363);
nor (n8289,n8290,n8291);
xor (n8290,n8147,n8282);
or (n8291,n8292,n8362);
and (n8292,n8293,n8361);
xor (n8293,n8294,n8295);
xor (n8294,n8135,n8138);
or (n8295,n8296,n8360);
and (n8296,n8297,n8300);
xor (n8297,n8298,n8299);
xor (n8298,n8101,n8130);
xor (n8299,n8154,n8157);
or (n8300,n8301,n8359);
and (n8301,n8302,n8358);
xor (n8302,n8303,n8357);
or (n8303,n8304,n8356);
and (n8304,n8305,n8332);
xor (n8305,n8306,n8313);
nand (n8306,n8307,n8312);
or (n8307,n7235,n8308);
not (n8308,n8309);
nor (n8309,n8310,n8311);
and (n8310,n7310,n7123);
and (n8311,n7308,n7138);
or (n8312,n8169,n7236);
or (n8313,n8314,n8331);
and (n8314,n8315,n8324);
xor (n8315,n8316,n8317);
xor (n8316,n8190,n8191);
nand (n8317,n8318,n8320);
or (n8318,n7377,n8319);
not (n8319,n8179);
nand (n8320,n8321,n7393);
nor (n8321,n8322,n8323);
and (n8322,n7203,n7384);
and (n8323,n7204,n7385);
nand (n8324,n8325,n8330);
or (n8325,n7591,n8326);
not (n8326,n8327);
nand (n8327,n8328,n8329);
or (n8328,n7251,n7179);
nand (n8329,n7179,n7251);
nand (n8330,n7603,n8242);
and (n8331,n8316,n8317);
or (n8332,n8333,n8355);
and (n8333,n8334,n8349);
xor (n8334,n8335,n8342);
nand (n8335,n8336,n8341);
or (n8336,n8337,n7184);
not (n8337,n8338);
nor (n8338,n8339,n8340);
and (n8339,n7338,n7188);
and (n8340,n7339,n7174);
nand (n8341,n8185,n7177);
nand (n8342,n8343,n8348);
or (n8343,n8344,n7235);
not (n8344,n8345);
nor (n8345,n8346,n8347);
and (n8346,n7470,n7123);
and (n8347,n7471,n7138);
nand (n8348,n8309,n7237);
nand (n8349,n8350,n8354);
or (n8350,n7116,n8351);
nor (n8351,n8352,n8353);
and (n8352,n7496,n7119);
and (n8353,n7497,n7120);
or (n8354,n7299,n8260);
and (n8355,n8335,n8342);
and (n8356,n8306,n8313);
xor (n8357,n8159,n8173);
xor (n8358,n8200,n8247);
and (n8359,n8303,n8357);
and (n8360,n8298,n8299);
xor (n8361,n8151,n8280);
and (n8362,n8294,n8295);
nor (n8363,n8364,n8365);
xor (n8364,n8293,n8361);
or (n8365,n8366,n8486);
and (n8366,n8367,n8485);
xor (n8367,n8368,n8369);
xor (n8368,n8197,n8278);
or (n8369,n8370,n8484);
and (n8370,n8371,n8403);
xor (n8371,n8372,n8402);
or (n8372,n8373,n8401);
and (n8373,n8374,n8400);
xor (n8374,n8375,n8376);
xor (n8375,n8227,n8239);
or (n8376,n8377,n8399);
and (n8377,n8378,n8393);
xor (n8378,n8379,n8386);
nand (n8379,n8380,n8385);
or (n8380,n8381,n7207);
not (n8381,n8382);
nor (n8382,n8383,n8384);
and (n8383,n7034,n7205);
and (n8384,n7033,n7211);
nand (n8385,n7225,n8253);
nand (n8386,n8387,n8392);
or (n8387,n8388,n7150);
not (n8388,n8389);
nor (n8389,n8390,n8391);
and (n8390,n7063,n7147);
and (n8391,n7064,n7149);
or (n8392,n7467,n8265);
nand (n8393,n8394,n8398);
or (n8394,n7475,n8395);
nor (n8395,n8396,n8397);
and (n8396,n7101,n7486);
and (n8397,n7102,n7483);
or (n8398,n7476,n8213);
and (n8399,n8379,n8386);
xor (n8400,n8249,n8263);
and (n8401,n8375,n8376);
xor (n8402,n8273,n8276);
or (n8403,n8404,n8483);
and (n8404,n8405,n8408);
xor (n8405,n8406,n8407);
xor (n8406,n8175,n8189);
xor (n8407,n8203,n8218);
or (n8408,n8409,n8482);
and (n8409,n8410,n8455);
xor (n8410,n8411,n8432);
or (n8411,n8412,n8431);
and (n8412,n8413,n8425);
xor (n8413,n8414,n8421);
nand (n8414,n8415,n8420);
or (n8415,n8416,n7591);
not (n8416,n8417);
nor (n8417,n8418,n8419);
and (n8418,n7288,n7179);
and (n8419,n7289,n7180);
nand (n8420,n8327,n7603);
nor (n8421,n8422,n8423);
nand (n8422,n7225,n7366);
not (n8423,n8424);
and (n8424,n7477,n7355);
nand (n8425,n8426,n8427);
or (n8426,n8337,n7176);
or (n8427,n7184,n8428);
nor (n8428,n8429,n8430);
and (n8429,n7188,n7055);
and (n8430,n7174,n7054);
and (n8431,n8414,n8421);
or (n8432,n8433,n8454);
and (n8433,n8434,n8447);
xor (n8434,n8435,n8442);
nor (n8435,n8436,n7211);
and (n8436,n8437,n8440);
not (n8437,n8438);
nor (n8438,n8439,n7174);
and (n8439,n7366,n7212);
not (n8440,n8441);
nor (n8441,n7366,n7212);
and (n8442,n8443,n7486);
nand (n8443,n8444,n8445);
or (n8444,n7484,n7355);
nand (n8445,n8446,n7147);
or (n8446,n7479,n7374);
nand (n8447,n8448,n8453);
or (n8448,n8449,n7207);
not (n8449,n8450);
nand (n8450,n8451,n8452);
or (n8451,n7211,n7366);
or (n8452,n7368,n7205);
nand (n8453,n7225,n8382);
and (n8454,n8435,n8442);
or (n8455,n8456,n8481);
and (n8456,n8457,n8473);
xor (n8457,n8458,n8464);
nand (n8458,n8459,n8463);
or (n8459,n8460,n7150);
nor (n8460,n8461,n8462);
and (n8461,n7109,n7147);
and (n8462,n7111,n7149);
nand (n8463,n7157,n8389);
nand (n8464,n8465,n8471);
or (n8465,n8466,n7475);
not (n8466,n8467);
nand (n8467,n8468,n8469);
or (n8468,n7483,n7355);
not (n8469,n8470);
and (n8470,n7355,n7483);
nand (n8471,n8472,n7477);
not (n8472,n8395);
nand (n8473,n8474,n8479);
or (n8474,n7394,n8475);
not (n8475,n8476);
nand (n8476,n8477,n8478);
or (n8477,n7270,n7384);
nand (n8478,n7384,n7270);
or (n8479,n8480,n7377);
not (n8480,n8321);
and (n8481,n8458,n8464);
and (n8482,n8411,n8432);
and (n8483,n8406,n8407);
and (n8484,n8372,n8402);
xor (n8485,n8297,n8300);
and (n8486,n8368,n8369);
not (n8487,n8488);
nand (n8488,n8489,n8894,n8901);
nand (n8489,n8490,n8590);
nor (n8490,n8491,n8513);
not (n8491,n8492);
or (n8492,n8493,n8494);
xor (n8493,n8367,n8485);
or (n8494,n8495,n8512);
and (n8495,n8496,n8511);
xor (n8496,n8497,n8510);
or (n8497,n8498,n8509);
and (n8498,n8499,n8508);
xor (n8499,n8500,n8501);
xor (n8500,n8305,n8332);
or (n8501,n8502,n8507);
and (n8502,n8503,n8506);
xor (n8503,n8504,n8505);
xor (n8504,n8334,n8349);
xor (n8505,n8378,n8393);
xor (n8506,n8315,n8324);
and (n8507,n8504,n8505);
xor (n8508,n8374,n8400);
and (n8509,n8500,n8501);
xor (n8510,n8302,n8358);
xor (n8511,n8371,n8403);
and (n8512,n8497,n8510);
nor (n8513,n8514,n8515);
xor (n8514,n8496,n8511);
or (n8515,n8516,n8589);
and (n8516,n8517,n8588);
xor (n8517,n8518,n8519);
xor (n8518,n8405,n8408);
or (n8519,n8520,n8587);
and (n8520,n8521,n8586);
xor (n8521,n8522,n8559);
or (n8522,n8523,n8558);
and (n8523,n8524,n8537);
xor (n8524,n8525,n8531);
nand (n8525,n8526,n8530);
or (n8526,n7235,n8527);
nor (n8527,n8528,n8529);
and (n8528,n7138,n7465);
and (n8529,n7463,n7123);
or (n8530,n8344,n7236);
nand (n8531,n8532,n8536);
or (n8532,n7116,n8533);
nor (n8533,n8534,n8535);
and (n8534,n7119,n7083);
and (n8535,n7084,n7120);
or (n8536,n7299,n8351);
or (n8537,n8538,n8557);
and (n8538,n8539,n8550);
xor (n8539,n8540,n8547);
nand (n8540,n8541,n8546);
or (n8541,n8542,n7394);
not (n8542,n8543);
nand (n8543,n8544,n8545);
or (n8544,n7251,n7384);
or (n8545,n7250,n7385);
nand (n8546,n8476,n7378);
nand (n8547,n8548,n8549);
or (n8548,n8424,n8422);
nand (n8549,n8422,n8424);
nand (n8550,n8551,n8556);
or (n8551,n7591,n8552);
not (n8552,n8553);
nor (n8553,n8554,n8555);
and (n8554,n7338,n7179);
and (n8555,n7339,n7180);
or (n8556,n7599,n8416);
and (n8557,n8540,n8547);
and (n8558,n8525,n8531);
or (n8559,n8560,n8585);
and (n8560,n8561,n8584);
xor (n8561,n8562,n8563);
xor (n8562,n8434,n8447);
or (n8563,n8564,n8583);
and (n8564,n8565,n8577);
xor (n8565,n8566,n8570);
nand (n8566,n8567,n8569);
or (n8567,n7235,n8568);
xor (n8568,n7496,n7138);
or (n8569,n8527,n7236);
nand (n8570,n8571,n8576);
or (n8571,n7184,n8572);
not (n8572,n8573);
nand (n8573,n8574,n8575);
or (n8574,n7034,n7188);
nand (n8575,n7188,n7034);
or (n8576,n8428,n7176);
nand (n8577,n8578,n8582);
or (n8578,n7116,n8579);
nor (n8579,n8580,n8581);
and (n8580,n7119,n7063);
and (n8581,n7064,n7120);
or (n8582,n7299,n8533);
and (n8583,n8566,n8570);
xor (n8584,n8457,n8473);
and (n8585,n8562,n8563);
xor (n8586,n8410,n8455);
and (n8587,n8522,n8559);
xor (n8588,n8499,n8508);
and (n8589,n8518,n8519);
nor (n8590,n8591,n8876);
and (n8591,n8592,n8868);
nor (n8592,n8593,n8864);
and (n8593,n8594,n8756);
nor (n8594,n8595,n8719);
nor (n8595,n8596,n8686);
xor (n8596,n8597,n8634);
xor (n8597,n8598,n8633);
or (n8598,n8599,n8632);
and (n8599,n8600,n8631);
xor (n8600,n8601,n8630);
or (n8601,n8602,n8629);
and (n8602,n8603,n8620);
xor (n8603,n8604,n8611);
nand (n8604,n8605,n8610);
or (n8605,n8606,n7184);
not (n8606,n8607);
nand (n8607,n8608,n8609);
or (n8608,n7188,n7366);
or (n8609,n7368,n7174);
nand (n8610,n8573,n7177);
nand (n8611,n8612,n8618);
or (n8612,n8613,n7116);
not (n8613,n8614);
nand (n8614,n8615,n8616);
or (n8615,n7120,n7109);
not (n8616,n8617);
and (n8617,n7109,n7120);
nand (n8618,n8619,n7136);
not (n8619,n8579);
nand (n8620,n8621,n8625);
or (n8621,n7150,n8622);
nor (n8622,n8623,n8624);
and (n8623,n7149,n7374);
and (n8624,n7355,n7147);
or (n8625,n7467,n8626);
nor (n8626,n8627,n8628);
and (n8627,n7149,n7101);
and (n8628,n7102,n7147);
and (n8629,n8604,n8611);
xor (n8630,n8565,n8577);
xor (n8631,n8539,n8550);
and (n8632,n8601,n8630);
xor (n8633,n8561,n8584);
xor (n8634,n8635,n8685);
xor (n8635,n8636,n8637);
xor (n8636,n8413,n8425);
or (n8637,n8638,n8684);
and (n8638,n8639,n8663);
xor (n8639,n8640,n8643);
nand (n8640,n8641,n8642);
or (n8641,n7150,n8626);
or (n8642,n7467,n8460);
or (n8643,n8644,n8662);
and (n8644,n8645,n8656);
xor (n8645,n8646,n8653);
nand (n8646,n8647,n8652);
or (n8647,n8648,n7591);
not (n8648,n8649);
nand (n8649,n8650,n8651);
or (n8650,n7054,n7180);
nand (n8651,n7180,n7054);
nand (n8652,n8553,n7603);
nor (n8653,n8654,n8655);
nand (n8654,n7177,n7366);
nand (n8655,n7157,n7355);
nand (n8656,n8657,n8661);
or (n8657,n7235,n8658);
nor (n8658,n8659,n8660);
and (n8659,n7083,n7138);
and (n8660,n7084,n7123);
or (n8661,n8568,n7236);
and (n8662,n8646,n8653);
or (n8663,n8664,n8683);
and (n8664,n8665,n8677);
xor (n8665,n8666,n8672);
nor (n8666,n8667,n7188);
and (n8667,n8668,n8671);
nand (n8668,n8669,n7179);
not (n8669,n8670);
and (n8670,n7366,n7181);
nand (n8671,n7368,n7190);
nor (n8672,n8673,n7147);
and (n8673,n8674,n8676);
nand (n8674,n8675,n7120);
or (n8675,n7154,n7374);
nand (n8676,n7374,n7154);
nand (n8677,n8678,n8679);
or (n8678,n7377,n8542);
or (n8679,n7394,n8680);
nor (n8680,n8681,n8682);
and (n8681,n7384,n7289);
and (n8682,n7385,n7288);
and (n8683,n8666,n8672);
and (n8684,n8640,n8643);
xor (n8685,n8524,n8537);
or (n8686,n8687,n8718);
and (n8687,n8688,n8717);
xor (n8688,n8689,n8690);
xor (n8689,n8639,n8663);
or (n8690,n8691,n8716);
and (n8691,n8692,n8715);
xor (n8692,n8693,n8714);
or (n8693,n8694,n8713);
and (n8694,n8695,n8708);
xor (n8695,n8696,n8702);
nand (n8696,n8697,n8701);
or (n8697,n8698,n7591);
nor (n8698,n8699,n8700);
and (n8699,n7034,n7179);
and (n8700,n7033,n7180);
nand (n8701,n7603,n8649);
nand (n8702,n8703,n8707);
or (n8703,n7235,n8704);
nor (n8704,n8705,n8706);
and (n8705,n7138,n7063);
and (n8706,n7064,n7123);
or (n8707,n8658,n7236);
nand (n8708,n8709,n8711);
or (n8709,n8710,n8655);
not (n8710,n8654);
or (n8711,n8712,n8654);
not (n8712,n8655);
and (n8713,n8696,n8702);
xor (n8714,n8665,n8677);
xor (n8715,n8645,n8656);
and (n8716,n8693,n8714);
xor (n8717,n8600,n8631);
and (n8718,n8689,n8690);
nor (n8719,n8720,n8721);
xor (n8720,n8688,n8717);
or (n8721,n8722,n8755);
and (n8722,n8723,n8754);
xor (n8723,n8724,n8725);
xor (n8724,n8603,n8620);
or (n8725,n8726,n8753);
and (n8726,n8727,n8740);
xor (n8727,n8728,n8734);
nand (n8728,n8729,n8730);
or (n8729,n8613,n7299);
or (n8730,n7116,n8731);
nor (n8731,n8732,n8733);
and (n8732,n7119,n7101);
and (n8733,n7102,n7120);
nand (n8734,n8735,n8739);
or (n8735,n7394,n8736);
nor (n8736,n8737,n8738);
and (n8737,n7384,n7339);
and (n8738,n7385,n7338);
or (n8739,n8680,n7377);
and (n8740,n8741,n8747);
nor (n8741,n8742,n7179);
and (n8742,n8743,n8746);
nand (n8743,n8744,n7384);
not (n8744,n8745);
and (n8745,n7366,n7595);
nand (n8746,n7368,n7598);
nor (n8747,n8748,n7120);
nor (n8748,n8749,n8752);
and (n8749,n8750,n7123);
nand (n8750,n7355,n8751);
not (n8751,n7124);
and (n8752,n7374,n7124);
and (n8753,n8728,n8734);
xor (n8754,n8692,n8715);
and (n8755,n8724,n8725);
nor (n8756,n8757,n8787);
nor (n8757,n8758,n8759);
xor (n8758,n8723,n8754);
or (n8759,n8760,n8786);
and (n8760,n8761,n8785);
xor (n8761,n8762,n8784);
or (n8762,n8763,n8783);
and (n8763,n8764,n8777);
xor (n8764,n8765,n8771);
nand (n8765,n8766,n8770);
or (n8766,n7591,n8767);
nor (n8767,n8768,n8769);
and (n8768,n7368,n7180);
and (n8769,n7179,n7366);
or (n8770,n7599,n8698);
nand (n8771,n8772,n8776);
or (n8772,n7235,n8773);
nor (n8773,n8774,n8775);
and (n8774,n7138,n7111);
and (n8775,n7109,n7123);
or (n8776,n8704,n7236);
nand (n8777,n8778,n8779);
or (n8778,n8731,n7299);
or (n8779,n7116,n8780);
nor (n8780,n8781,n8782);
and (n8781,n7355,n7120);
and (n8782,n7119,n7374);
and (n8783,n8765,n8771);
xor (n8784,n8695,n8708);
xor (n8785,n8727,n8740);
and (n8786,n8762,n8784);
nand (n8787,n8788,n8859);
or (n8788,n8789,n8846);
nand (n8789,n8790,n8843);
or (n8790,n8791,n8826);
nor (n8791,n8792,n8793);
xor (n8792,n8764,n8777);
xor (n8793,n8794,n8806);
xor (n8794,n8795,n8801);
nand (n8795,n8796,n8800);
or (n8796,n7394,n8797);
nor (n8797,n8798,n8799);
and (n8798,n7384,n7055);
and (n8799,n7385,n7054);
or (n8800,n8736,n7377);
xor (n8801,n8802,n8803);
xor (n8802,n8741,n8747);
nor (n8803,n8804,n8805);
nand (n8804,n7136,n7355);
nand (n8805,n7603,n7366);
or (n8806,n8807,n8825);
and (n8807,n8808,n8819);
xor (n8808,n8809,n8815);
nand (n8809,n8810,n8814);
or (n8810,n7394,n8811);
nor (n8811,n8812,n8813);
and (n8812,n7384,n7034);
and (n8813,n7385,n7033);
or (n8814,n8797,n7377);
nand (n8815,n8816,n8818);
or (n8816,n8817,n8805);
not (n8817,n8804);
nand (n8818,n8817,n8805);
nand (n8819,n8820,n8824);
or (n8820,n7235,n8821);
nor (n8821,n8822,n8823);
and (n8822,n7138,n7101);
and (n8823,n7102,n7123);
or (n8824,n8773,n7236);
and (n8825,n8809,n8815);
nand (n8826,n8827,n8828);
xor (n8827,n8808,n8819);
or (n8828,n8829,n8842);
and (n8829,n8830,n8834);
xor (n8830,n8831,n8833);
nor (n8831,n8832,n7384);
and (n8832,n7366,n7378);
nor (n8833,n7123,n7355,n7236);
nand (n8834,n8835,n8841);
or (n8835,n8836,n7235);
not (n8836,n8837);
nand (n8837,n8838,n8839);
or (n8838,n7123,n7355);
not (n8839,n8840);
and (n8840,n7355,n7123);
or (n8841,n8821,n7236);
and (n8842,n8831,n8833);
or (n8843,n8844,n8845);
not (n8844,n8793);
not (n8845,n8792);
nor (n8846,n8791,n8847);
nand (n8847,n8848,n8849,n8852);
or (n8848,n8827,n8828);
or (n8849,n8850,n8851);
and (n8850,n8832,n7355,n7237);
xor (n8851,n8830,n8834);
nand (n8852,n8853,n8857,n8858);
or (n8853,n8854,n7394);
nor (n8854,n8855,n8856);
and (n8855,n7368,n7385);
and (n8856,n7384,n7366);
or (n8857,n7377,n8811);
nand (n8858,n8851,n8850);
or (n8859,n8860,n8861);
xor (n8860,n8761,n8785);
or (n8861,n8862,n8863);
and (n8862,n8794,n8806);
and (n8863,n8795,n8801);
nand (n8864,n8865,n8867);
or (n8865,n8595,n8866);
nand (n8866,n8720,n8721);
nand (n8867,n8596,n8686);
nand (n8868,n8869,n8594);
or (n8869,n8870,n8872);
not (n8870,n8871);
nand (n8871,n8758,n8759);
not (n8872,n8873);
nand (n8873,n8874,n8875);
not (n8874,n8757);
and (n8875,n8860,n8861);
not (n8876,n8877);
nor (n8877,n8878,n8889);
nor (n8878,n8879,n8880);
xor (n8879,n8517,n8588);
or (n8880,n8881,n8888);
and (n8881,n8882,n8887);
xor (n8882,n8883,n8884);
xor (n8883,n8503,n8506);
or (n8884,n8885,n8886);
and (n8885,n8635,n8685);
and (n8886,n8636,n8637);
xor (n8887,n8521,n8586);
and (n8888,n8883,n8884);
nor (n8889,n8890,n8891);
xor (n8890,n8882,n8887);
or (n8891,n8892,n8893);
and (n8892,n8597,n8634);
and (n8893,n8598,n8633);
nand (n8894,n8490,n8895);
nand (n8895,n8896,n8899);
or (n8896,n8897,n8898);
not (n8897,n8880);
not (n8898,n8879);
or (n8899,n8878,n8900);
nand (n8900,n8890,n8891);
nand (n8901,n8492,n8902);
nand (n8902,n8903,n8906);
or (n8903,n8904,n8905);
not (n8904,n8494);
not (n8905,n8493);
nand (n8906,n8514,n8515);
nor (n8907,n8908,n8912);
and (n8908,n8909,n8910);
not (n8909,n8289);
not (n8910,n8911);
nand (n8911,n8364,n8365);
and (n8912,n8290,n8291);
nor (n8913,n8914,n8917);
and (n8914,n8915,n8916);
not (n8915,n7018);
and (n8916,n8144,n8145);
and (n8917,n7019,n8038);
nor (n8918,n8919,n9560);
not (n8919,n8920);
nor (n8920,n8921,n9541);
nor (n8921,n8922,n9488);
xor (n8922,n8923,n9469);
xor (n8923,n8924,n9228);
or (n8924,n8925,n9227);
and (n8925,n8926,n9187);
xor (n8926,n8927,n9042);
xor (n8927,n8928,n8991);
xor (n8928,n8929,n8957);
xor (n8929,n8930,n8947);
xor (n8930,n8931,n8937);
nand (n8931,n8932,n8934);
or (n8932,n7603,n8933);
not (n8933,n7591);
nor (n8934,n8935,n8936);
and (n8935,n7866,n7179);
and (n8936,n7867,n7180);
nand (n8937,n8938,n8943);
or (n8938,n8939,n7038);
not (n8939,n8940);
nand (n8940,n8941,n8942);
or (n8941,n7251,n7035);
nand (n8942,n7035,n7251);
nand (n8943,n8944,n7057);
nor (n8944,n8945,n8946);
and (n8945,n7269,n7035);
and (n8946,n7270,n7036);
nand (n8947,n8948,n8953);
or (n8948,n8949,n7068);
not (n8949,n8950);
nor (n8950,n8951,n8952);
and (n8951,n7470,n7065);
and (n8952,n7471,n7067);
nand (n8953,n7075,n8954);
nand (n8954,n8955,n8956);
or (n8955,n7308,n7065);
nand (n8956,n7065,n7308);
xor (n8957,n8958,n8979);
xor (n8958,n8959,n8969);
nand (n8959,n8960,n8965);
or (n8960,n8961,n7325);
not (n8961,n8962);
nand (n8962,n8963,n8964);
or (n8963,n7204,n7048);
nand (n8964,n7204,n7048);
nand (n8965,n8966,n7327);
nand (n8966,n8967,n8968);
or (n8967,n7223,n7048);
nand (n8968,n7048,n7223);
nand (n8969,n8970,n8974);
or (n8970,n8971,n7475);
nor (n8971,n8972,n8973);
and (n8972,n7129,n7483);
nor (n8973,n7483,n7129);
nand (n8974,n8975,n7477);
nor (n8975,n8976,n8978);
and (n8976,n8977,n7483);
not (n8977,n7134);
and (n8978,n7134,n7486);
nand (n8979,n8980,n8986);
or (n8980,n8981,n7524);
not (n8981,n8982);
nand (n8982,n8983,n8984);
or (n8983,n7078,n7165);
not (n8984,n8985);
and (n8985,n7165,n7078);
or (n8986,n7523,n8987);
not (n8987,n8988);
nand (n8988,n8989,n8990);
or (n8989,n7146,n7078);
nand (n8990,n7078,n7146);
xor (n8991,n8992,n9015);
xor (n8992,n8993,n9005);
nand (n8993,n8994,n8999);
or (n8994,n7978,n8995);
not (n8995,n8996);
nand (n8996,n8997,n8998);
or (n8997,n7339,n7852);
nand (n8998,n7339,n7852);
or (n8999,n9000,n9001);
not (n9000,n7756);
not (n9001,n9002);
nor (n9002,n9003,n9004);
and (n9003,n7288,n7852);
and (n9004,n7289,n7853);
not (n9005,n9006);
nand (n9006,n9007,n9011);
or (n9007,n9008,n7184);
nor (n9008,n9009,n9010);
and (n9009,n7383,n7188);
and (n9010,n7382,n7174);
nand (n9011,n7177,n9012);
nor (n9012,n9013,n9014);
and (n9013,n7744,n7188);
and (n9014,n7745,n7174);
or (n9015,n9016,n9041);
and (n9016,n9017,n9032);
xor (n9017,n9018,n9025);
nand (n9018,n9019,n9024);
or (n9019,n9020,n7038);
not (n9020,n9021);
nand (n9021,n9022,n9023);
or (n9022,n7289,n7035);
nand (n9023,n7035,n7289);
nand (n9024,n8940,n7057);
nand (n9025,n9026,n9031);
or (n9026,n9027,n7068);
not (n9027,n9028);
nor (n9028,n9029,n9030);
and (n9029,n7465,n7065);
and (n9030,n7463,n7067);
nand (n9031,n8950,n7075);
nand (n9032,n9033,n9037);
or (n9033,n7088,n9034);
nor (n9034,n9035,n9036);
and (n9035,n7084,n7093);
and (n9036,n7083,n7092);
or (n9037,n9038,n7095);
nor (n9038,n9039,n9040);
and (n9039,n7092,n7496);
and (n9040,n7497,n7093);
and (n9041,n9018,n9025);
or (n9042,n9043,n9186);
and (n9043,n9044,n9117);
xor (n9044,n9045,n9058);
or (n9045,n9046,n9057);
and (n9046,n9047,n9054);
xor (n9047,n9048,n9051);
or (n9048,n9049,n9050);
and (n9049,n7844,n7860);
and (n9050,n7845,n7854);
or (n9051,n9052,n9053);
and (n9052,n7971,n7996);
and (n9053,n7972,n7988);
or (n9054,n9055,n9056);
and (n9055,n7928,n7943);
and (n9056,n7929,n7936);
and (n9057,n9048,n9051);
xor (n9058,n9059,n9094);
xor (n9059,n9060,n9070);
and (n9060,n9061,n9068);
nand (n9061,n9062,n9064);
or (n9062,n9063,n7591);
not (n9063,n7933);
nand (n9064,n7603,n9065);
nor (n9065,n9066,n9067);
and (n9066,n7744,n7179);
and (n9067,n7745,n7180);
nand (n9068,n9069,n7864);
or (n9069,n7378,n7393);
or (n9070,n9071,n9093);
and (n9071,n9072,n9087);
xor (n9072,n9073,n9080);
nand (n9073,n9074,n9076);
or (n9074,n9075,n7207);
not (n9075,n7940);
nand (n9076,n7225,n9077);
nand (n9077,n9078,n9079);
or (n9078,n7173,n7211);
nand (n9079,n7211,n7173);
nand (n9080,n9081,n9083);
or (n9081,n9082,n7978);
not (n9082,n7985);
nand (n9083,n7756,n9084);
nand (n9084,n9085,n9086);
or (n9085,n7055,n7852);
nand (n9086,n7852,n7055);
nand (n9087,n9088,n9089);
or (n9088,n7998,n8007);
or (n9089,n9090,n7750);
nor (n9090,n9091,n9092);
and (n9091,n8002,n7111);
and (n9092,n7109,n7859);
and (n9093,n9073,n9080);
or (n9094,n9095,n9116);
and (n9095,n9096,n9108);
xor (n9096,n9097,n9101);
nand (n9097,n9098,n9100);
or (n9098,n7237,n9099);
not (n9099,n7235);
not (n9100,n7915);
nand (n9101,n9102,n9104);
or (n9102,n9103,n7255);
not (n9103,n7908);
nand (n9104,n9105,n7264);
nand (n9105,n9106,n9107);
or (n9106,n7223,n7252);
nand (n9107,n7252,n7223);
nand (n9108,n9109,n9115);
or (n9109,n9110,n7299);
not (n9110,n9111);
nand (n9111,n9112,n9114);
not (n9112,n9113);
and (n9113,n7242,n7120);
nand (n9114,n7119,n7244);
or (n9115,n7116,n7924);
and (n9116,n9097,n9101);
xor (n9117,n9118,n9168);
xor (n9118,n9119,n9145);
or (n9119,n9120,n9144);
and (n9120,n9121,n9136);
xor (n9121,n9122,n9129);
nand (n9122,n9123,n9124);
or (n9123,n8027,n7150);
nand (n9124,n9125,n7157);
nand (n9125,n9126,n9128);
not (n9126,n9127);
and (n9127,n7134,n7147);
nand (n9128,n7149,n8977);
nand (n9129,n9130,n9132);
or (n9130,n9131,n7184);
not (n9131,n8015);
nand (n9132,n9133,n7177);
nand (n9133,n9134,n9135);
or (n9134,n7390,n7174);
nand (n9135,n7174,n7390);
nand (n9136,n9137,n9142);
or (n9137,n7326,n9138);
not (n9138,n9139);
nor (n9139,n9140,n9141);
and (n9140,n7269,n7048);
and (n9141,n7270,n7049);
or (n9142,n7325,n9143);
not (n9143,n8022);
and (n9144,n9122,n9129);
or (n9145,n9146,n9167);
and (n9146,n9147,n9163);
xor (n9147,n9148,n9156);
nand (n9148,n9149,n9151);
or (n9149,n9150,n7475);
not (n9150,n7883);
nand (n9151,n9152,n7477);
not (n9152,n9153);
nor (n9153,n9154,n9155);
and (n9154,n7486,n7164);
and (n9155,n7165,n7483);
nand (n9156,n9157,n9158);
or (n9157,n7895,n7523);
nand (n9158,n7525,n9159);
nand (n9159,n9160,n9162);
not (n9160,n9161);
and (n9161,n7308,n7078);
nand (n9162,n7077,n7310);
nand (n9163,n9164,n9166);
or (n9164,n9165,n7038);
not (n9165,n7890);
nand (n9166,n7057,n9021);
and (n9167,n9148,n9156);
xor (n9168,n9169,n9183);
xor (n9169,n9170,n9176);
nand (n9170,n9171,n9172);
or (n9171,n7116,n9110);
nand (n9172,n9173,n7136);
nor (n9173,n9174,n9175);
and (n9174,n7919,n7120);
and (n9175,n7917,n7119);
nand (n9176,n9177,n9179);
or (n9177,n9178,n7150);
not (n9178,n9125);
nand (n9179,n9180,n7157);
nor (n9180,n9181,n9182);
and (n9181,n7234,n7147);
and (n9182,n7232,n7149);
nand (n9183,n9184,n9185);
or (n9184,n9138,n7325);
nand (n9185,n8962,n7327);
and (n9186,n9045,n9058);
xor (n9187,n9188,n9224);
xor (n9188,n9189,n9192);
or (n9189,n9190,n9191);
and (n9190,n9059,n9094);
and (n9191,n9060,n9070);
xor (n9192,n9193,n9209);
xor (n9193,n9194,n9206);
nand (n9194,n9195,n9198);
nor (n9195,n9196,n9197);
and (n9196,n7185,n9133);
nor (n9197,n7176,n9008);
nor (n9198,n9199,n9200);
and (n9199,n7256,n9105);
nor (n9200,n9201,n9205);
not (n9201,n9202);
nand (n9202,n9203,n9204);
or (n9203,n7194,n7252);
nand (n9204,n7252,n7194);
not (n9205,n7264);
or (n9206,n9207,n9208);
and (n9207,n9169,n9183);
and (n9208,n9170,n9176);
or (n9209,n9210,n9223);
and (n9210,n9211,n9219);
xor (n9211,n9212,n9215);
nand (n9212,n9213,n9214);
or (n9213,n7475,n9153);
or (n9214,n7476,n8971);
nand (n9215,n9216,n9218);
or (n9216,n9217,n7523);
not (n9217,n9159);
nand (n9218,n8988,n7525);
nand (n9219,n9220,n9222);
or (n9220,n9221,n7591);
not (n9221,n9065);
nand (n9222,n7603,n8934);
and (n9223,n9212,n9215);
or (n9224,n9225,n9226);
and (n9225,n9118,n9168);
and (n9226,n9119,n9145);
and (n9227,n8927,n9042);
xor (n9228,n9229,n9445);
xor (n9229,n9230,n9401);
xor (n9230,n9231,n9329);
xor (n9231,n9232,n9281);
xor (n9232,n9233,n9257);
xor (n9233,n9234,n9254);
or (n9234,n9235,n9253);
and (n9235,n9236,n9245);
xor (n9236,n9237,n9243);
nand (n9237,n9238,n9239);
or (n9238,n9201,n7255);
nand (n9239,n9240,n7264);
nand (n9240,n9241,n9242);
or (n9241,n7173,n7252);
nand (n9242,n7252,n7173);
nand (n9243,n9244,n9173);
or (n9244,n7136,n7117);
nand (n9245,n9246,n9251);
or (n9246,n7467,n9247);
not (n9247,n9248);
nor (n9248,n9249,n9250);
and (n9249,n7244,n7147);
and (n9250,n7242,n7149);
or (n9251,n7150,n9252);
not (n9252,n9180);
and (n9253,n9237,n9243);
or (n9254,n9255,n9256);
and (n9255,n8958,n8979);
and (n9256,n8959,n8969);
xor (n9257,n9258,n9275);
xor (n9258,n9259,n9266);
nand (n9259,n9260,n9265);
or (n9260,n9000,n9261);
not (n9261,n9262);
nor (n9262,n9263,n9264);
and (n9263,n7250,n7852);
and (n9264,n7251,n7853);
nand (n9265,n7979,n9002);
nand (n9266,n9267,n9271);
or (n9267,n9268,n7998);
nor (n9268,n9269,n9270);
and (n9269,n8002,n7083);
and (n9270,n7084,n7859);
nand (n9271,n9272,n7749);
nor (n9272,n9273,n9274);
and (n9273,n8002,n7497);
and (n9274,n7859,n7496);
nand (n9275,n9276,n9277);
or (n9276,n9247,n7150);
nand (n9277,n7157,n9278);
nor (n9278,n9279,n9280);
and (n9279,n7919,n7147);
and (n9280,n7917,n7149);
or (n9281,n9282,n9328);
and (n9282,n9283,n9327);
xor (n9283,n9284,n9307);
or (n9284,n9285,n9306);
and (n9285,n9286,n9302);
xor (n9286,n9287,n9294);
nand (n9287,n9288,n9290);
or (n9288,n9289,n7207);
not (n9289,n9077);
nand (n9290,n7225,n9291);
nand (n9291,n9292,n9293);
or (n9292,n7557,n7205);
nand (n9293,n7205,n7557);
nand (n9294,n9295,n9298);
nand (n9295,n9296,n9297);
not (n9296,n9090);
not (n9297,n7998);
nand (n9298,n9299,n7749);
nor (n9299,n9300,n9301);
and (n9300,n8002,n7064);
and (n9301,n7859,n7063);
nand (n9302,n9303,n9305);
or (n9303,n9304,n7978);
not (n9304,n9084);
nand (n9305,n8996,n7756);
and (n9306,n9287,n9294);
xor (n9307,n9308,n9323);
xor (n9308,n9309,n9316);
nand (n9309,n9310,n9315);
or (n9310,n7095,n9311);
not (n9311,n9312);
nor (n9312,n9313,n9314);
and (n9313,n7463,n7092);
and (n9314,n7465,n7093);
or (n9315,n7088,n9038);
nand (n9316,n9317,n9319);
or (n9317,n9318,n7207);
not (n9318,n9291);
nand (n9319,n7225,n9320);
nand (n9320,n9321,n9322);
or (n9321,n7391,n7211);
nand (n9322,n7211,n7391);
nand (n9323,n9324,n9326);
or (n9324,n7998,n9325);
not (n9325,n9299);
or (n9326,n9268,n7750);
xor (n9327,n9236,n9245);
and (n9328,n9284,n9307);
xor (n9329,n9330,n9377);
xor (n9330,n9331,n9354);
xor (n9331,n9332,n9347);
xor (n9332,n9333,n9340);
nand (n9333,n9334,n9336);
or (n9334,n9335,n7184);
not (n9335,n9012);
nand (n9336,n9337,n7177);
nand (n9337,n9338,n9339);
or (n9338,n7867,n7188);
nand (n9339,n7188,n7867);
nand (n9340,n9341,n9343);
or (n9341,n9342,n7207);
not (n9342,n9320);
nand (n9343,n7225,n9344);
nor (n9344,n9345,n9346);
and (n9345,n7382,n7211);
and (n9346,n7383,n7205);
nand (n9347,n9348,n9350);
or (n9348,n9349,n7325);
not (n9349,n8966);
nand (n9350,n9351,n7327);
nor (n9351,n9352,n9353);
and (n9352,n8125,n7048);
and (n9353,n7194,n7049);
xor (n9354,n9355,n9370);
xor (n9355,n9356,n9364);
nand (n9356,n9357,n9359);
or (n9357,n9358,n7068);
not (n9358,n8954);
nand (n9359,n9360,n7075);
nand (n9360,n9361,n9363);
not (n9361,n9362);
and (n9362,n7146,n7065);
nand (n9363,n7067,n7145);
nand (n9364,n9365,n9366);
or (n9365,n9311,n7088);
nand (n9366,n9367,n7788);
nor (n9367,n9368,n9369);
and (n9368,n7470,n7093);
and (n9369,n7471,n7092);
nand (n9370,n9371,n9373);
or (n9371,n9372,n7255);
not (n9372,n9240);
nand (n9373,n9374,n7264);
nor (n9374,n9375,n9376);
and (n9375,n7557,n7252);
and (n9376,n7558,n7253);
xor (n9377,n9378,n9393);
xor (n9378,n9379,n9386);
nand (n9379,n9380,n9382);
or (n9380,n9381,n7475);
not (n9381,n8975);
nand (n9382,n7477,n9383);
nor (n9383,n9384,n9385);
and (n9384,n7234,n7483);
and (n9385,n7232,n7486);
nand (n9386,n9387,n9388);
or (n9387,n8981,n7523);
or (n9388,n9389,n7524);
nor (n9389,n9390,n9392);
and (n9390,n7077,n9391);
not (n9391,n7129);
and (n9392,n7129,n7078);
nand (n9393,n9394,n9396);
or (n9394,n9395,n7038);
not (n9395,n8944);
or (n9396,n7046,n9397);
not (n9397,n9398);
nor (n9398,n9399,n9400);
and (n9399,n7203,n7035);
and (n9400,n7204,n7036);
or (n9401,n9402,n9444);
and (n9402,n9403,n9412);
xor (n9403,n9404,n9411);
or (n9404,n9405,n9410);
and (n9405,n9406,n9409);
xor (n9406,n9407,n9408);
xor (n9407,n9286,n9302);
xnor (n9408,n9195,n9198);
xor (n9409,n9017,n9032);
and (n9410,n9407,n9408);
xor (n9411,n9283,n9327);
or (n9412,n9413,n9443);
and (n9413,n9414,n9430);
xor (n9414,n9415,n9416);
xor (n9415,n9211,n9219);
or (n9416,n9417,n9429);
and (n9417,n9418,n9425);
xor (n9418,n9419,n9422);
nand (n9419,n9420,n9421);
or (n9420,n7068,n7840);
nand (n9421,n7075,n9028);
nand (n9422,n9423,n9424);
or (n9423,n7990,n7088);
or (n9424,n9034,n7095);
nand (n9425,n9426,n9428);
or (n9426,n9427,n9061);
not (n9427,n9068);
nand (n9428,n9427,n9061);
and (n9429,n9419,n9422);
or (n9430,n9431,n9442);
and (n9431,n9432,n9439);
xor (n9432,n9433,n9436);
or (n9433,n9434,n9435);
and (n9434,n7903,n7920);
and (n9435,n7904,n7911);
or (n9436,n9437,n9438);
and (n9437,n8011,n8025);
and (n9438,n8012,n8018);
or (n9439,n9440,n9441);
and (n9440,n7878,n7893);
and (n9441,n7879,n7886);
and (n9442,n9433,n9436);
and (n9443,n9415,n9416);
and (n9444,n9404,n9411);
xor (n9445,n9446,n9453);
xor (n9446,n9447,n9450);
or (n9447,n9448,n9449);
and (n9448,n8928,n8991);
and (n9449,n8929,n8957);
or (n9450,n9451,n9452);
and (n9451,n9188,n9224);
and (n9452,n9189,n9192);
xor (n9453,n9454,n9461);
xor (n9454,n9455,n9458);
or (n9455,n9456,n9457);
and (n9456,n8992,n9015);
and (n9457,n8993,n9005);
or (n9458,n9459,n9460);
and (n9459,n9193,n9209);
and (n9460,n9194,n9206);
xor (n9461,n9462,n9466);
xor (n9462,n9006,n9463);
or (n9463,n9464,n9465);
and (n9464,n8930,n8947);
and (n9465,n8931,n8937);
or (n9466,n9467,n9468);
and (n9467,n9308,n9323);
and (n9468,n9309,n9316);
or (n9469,n9470,n9487);
and (n9470,n9471,n9486);
xor (n9471,n9472,n9473);
xor (n9472,n9403,n9412);
or (n9473,n9474,n9485);
and (n9474,n9475,n9484);
xor (n9475,n9476,n9483);
or (n9476,n9477,n9482);
and (n9477,n9478,n9481);
xor (n9478,n9479,n9480);
xor (n9479,n9147,n9163);
xor (n9480,n9096,n9108);
xor (n9481,n9121,n9136);
and (n9482,n9479,n9480);
xor (n9483,n9406,n9409);
xor (n9484,n9414,n9430);
and (n9485,n9476,n9483);
xor (n9486,n8926,n9187);
and (n9487,n9472,n9473);
or (n9488,n9489,n9540);
and (n9489,n9490,n9525);
xor (n9490,n9491,n9524);
or (n9491,n9492,n9523);
and (n9492,n9493,n9514);
xor (n9493,n9494,n9503);
or (n9494,n9495,n9502);
and (n9495,n9496,n9499);
xor (n9496,n9497,n9498);
xor (n9497,n9072,n9087);
xor (n9498,n9418,n9425);
or (n9499,n9500,n9501);
and (n9500,n7953,n7960);
and (n9501,n7954,n7957);
and (n9502,n9497,n9498);
or (n9503,n9504,n9513);
and (n9504,n9505,n9512);
xor (n9505,n9506,n9509);
or (n9506,n9507,n9508);
and (n9507,n7835,n7869);
and (n9508,n7836,n7843);
or (n9509,n9510,n9511);
and (n9510,n7876,n7927);
and (n9511,n7877,n7902);
xor (n9512,n9432,n9439);
and (n9513,n9506,n9509);
or (n9514,n9515,n9522);
and (n9515,n9516,n9521);
xor (n9516,n9517,n9518);
xor (n9517,n9047,n9054);
or (n9518,n9519,n9520);
and (n9519,n7966,n8010);
and (n9520,n7967,n7970);
xor (n9521,n9478,n9481);
and (n9522,n9517,n9518);
and (n9523,n9494,n9503);
xor (n9524,n9471,n9486);
or (n9525,n9526,n9539);
and (n9526,n9527,n9530);
xor (n9527,n9528,n9529);
xor (n9528,n9044,n9117);
xor (n9529,n9475,n9484);
or (n9530,n9531,n9538);
and (n9531,n9532,n9537);
xor (n9532,n9533,n9534);
xor (n9533,n9496,n9499);
or (n9534,n9535,n9536);
and (n9535,n7945,n7952);
and (n9536,n7946,n7949);
xor (n9537,n9516,n9521);
and (n9538,n9533,n9534);
and (n9539,n9528,n9529);
and (n9540,n9491,n9524);
nor (n9541,n9542,n9543);
xor (n9542,n9490,n9525);
or (n9543,n9544,n9559);
and (n9544,n9545,n9558);
xor (n9545,n9546,n9547);
xor (n9546,n9493,n9514);
or (n9547,n9548,n9557);
and (n9548,n9549,n9554);
xor (n9549,n9550,n9553);
or (n9550,n9551,n9552);
and (n9551,n7833,n7875);
and (n9552,n7834,n7872);
xor (n9553,n9505,n9512);
or (n9554,n9555,n9556);
and (n9555,n7964,n8035);
and (n9556,n7965,n8032);
and (n9557,n9550,n9553);
xor (n9558,n9527,n9530);
and (n9559,n9546,n9547);
nand (n9560,n9561,n9573);
not (n9561,n9562);
nor (n9562,n9563,n9564);
xor (n9563,n9545,n9558);
or (n9564,n9565,n9572);
and (n9565,n9566,n9569);
xor (n9566,n9567,n9568);
xor (n9567,n9532,n9537);
xor (n9568,n9549,n9554);
or (n9569,n9570,n9571);
and (n9570,n7831,n7963);
and (n9571,n7832,n7944);
and (n9572,n9567,n9568);
nand (n9573,n9574,n9576);
not (n9574,n9575);
xor (n9575,n9566,n9569);
not (n9576,n9577);
or (n9577,n9578,n9579);
and (n9578,n7020,n7830);
and (n9579,n7021,n7671);
nor (n9580,n9581,n9841);
nand (n9581,n9582,n9716);
nand (n9582,n9583,n9712);
not (n9583,n9584);
xor (n9584,n9585,n9709);
xor (n9585,n9586,n9682);
xor (n9586,n9587,n9679);
xor (n9587,n9588,n9634);
xor (n9588,n9589,n9612);
xor (n9589,n9590,n9593);
or (n9590,n9591,n9592);
and (n9591,n9378,n9393);
and (n9592,n9379,n9386);
xor (n9593,n9594,n9604);
xor (n9594,n9595,n9597);
nand (n9595,n9596,n9337);
or (n9596,n7177,n7185);
nand (n9597,n9598,n9600);
or (n9598,n9599,n7255);
not (n9599,n9374);
nand (n9600,n7264,n9601);
nor (n9601,n9602,n9603);
and (n9602,n7391,n7253);
and (n9603,n7390,n7252);
nand (n9604,n9605,n9607);
or (n9605,n7998,n9606);
not (n9606,n9272);
or (n9607,n9608,n7750);
not (n9608,n9609);
nor (n9609,n9610,n9611);
and (n9610,n7465,n7859);
and (n9611,n7463,n8002);
xor (n9612,n9613,n9628);
xor (n9613,n9614,n9621);
nand (n9614,n9615,n9617);
or (n9615,n9616,n7325);
not (n9616,n9351);
nand (n9617,n9618,n7327);
nor (n9618,n9619,n9620);
and (n9619,n7172,n7048);
and (n9620,n7173,n7049);
nand (n9621,n9622,n9624);
or (n9622,n7475,n9623);
not (n9623,n9383);
or (n9624,n7476,n9625);
nor (n9625,n9626,n9627);
and (n9626,n7244,n7486);
and (n9627,n7242,n7483);
nand (n9628,n9629,n9630);
or (n9629,n7523,n9389);
or (n9630,n7524,n9631);
nor (n9631,n9632,n9633);
and (n9632,n7077,n8977);
and (n9633,n7134,n7078);
xor (n9634,n9635,n9676);
xor (n9635,n9636,n9658);
xor (n9636,n9637,n9651);
xor (n9637,n9638,n9644);
nand (n9638,n9639,n9640);
or (n9639,n9397,n7038);
nand (n9640,n9641,n7057);
nor (n9641,n9642,n9643);
and (n9642,n7222,n7035);
and (n9643,n7223,n7036);
nand (n9644,n9645,n9647);
or (n9645,n9646,n7068);
not (n9646,n9360);
nand (n9647,n9648,n7075);
nor (n9648,n9649,n9650);
and (n9649,n7164,n7065);
and (n9650,n7165,n7067);
nand (n9651,n9652,n9654);
or (n9652,n7088,n9653);
not (n9653,n9367);
or (n9654,n9655,n7095);
nor (n9655,n9656,n9657);
and (n9656,n7092,n7310);
and (n9657,n7308,n7093);
xor (n9658,n9659,n9668);
xor (n9659,n9660,n9666);
nand (n9660,n9661,n9662);
or (n9661,n9261,n7978);
or (n9662,n9663,n9000);
nor (n9663,n9664,n9665);
and (n9664,n7270,n7852);
and (n9665,n7853,n7269);
nand (n9666,n9667,n9278);
or (n9667,n7157,n7151);
not (n9668,n9669);
nand (n9669,n9670,n9672);
or (n9670,n9671,n7207);
not (n9671,n9344);
nand (n9672,n7225,n9673);
nor (n9673,n9674,n9675);
and (n9674,n7744,n7211);
and (n9675,n7745,n7205);
or (n9676,n9677,n9678);
and (n9677,n9462,n9466);
and (n9678,n9006,n9463);
or (n9679,n9680,n9681);
and (n9680,n9454,n9461);
and (n9681,n9455,n9458);
xor (n9682,n9683,n9706);
xor (n9683,n9684,n9703);
xor (n9684,n9685,n9692);
xor (n9685,n9686,n9689);
or (n9686,n9687,n9688);
and (n9687,n9330,n9377);
and (n9688,n9331,n9354);
or (n9689,n9690,n9691);
and (n9690,n9233,n9257);
and (n9691,n9234,n9254);
xor (n9692,n9693,n9700);
xor (n9693,n9694,n9697);
or (n9694,n9695,n9696);
and (n9695,n9355,n9370);
and (n9696,n9356,n9364);
or (n9697,n9698,n9699);
and (n9698,n9258,n9275);
and (n9699,n9259,n9266);
or (n9700,n9701,n9702);
and (n9701,n9332,n9347);
and (n9702,n9333,n9340);
or (n9703,n9704,n9705);
and (n9704,n9231,n9329);
and (n9705,n9232,n9281);
or (n9706,n9707,n9708);
and (n9707,n9446,n9453);
and (n9708,n9447,n9450);
or (n9709,n9710,n9711);
and (n9710,n9229,n9445);
and (n9711,n9230,n9401);
not (n9712,n9713);
or (n9713,n9714,n9715);
and (n9714,n8923,n9469);
and (n9715,n8924,n9228);
nand (n9716,n9717,n9721);
not (n9717,n9718);
or (n9718,n9719,n9720);
and (n9719,n9585,n9709);
and (n9720,n9586,n9682);
not (n9721,n9722);
xor (n9722,n9723,n9838);
xor (n9723,n9724,n9727);
or (n9724,n9725,n9726);
and (n9725,n9587,n9679);
and (n9726,n9588,n9634);
xor (n9727,n9728,n9751);
xor (n9728,n9729,n9748);
xor (n9729,n9730,n9745);
xor (n9730,n9731,n9734);
or (n9731,n9732,n9733);
and (n9732,n9693,n9700);
and (n9733,n9694,n9697);
xor (n9734,n9735,n9742);
xor (n9735,n9736,n9669);
nand (n9736,n9737,n9738);
or (n9737,n7523,n9631);
or (n9738,n7524,n9739);
nor (n9739,n9740,n9741);
and (n9740,n7077,n7234);
and (n9741,n7232,n7078);
or (n9742,n9743,n9744);
and (n9743,n9613,n9628);
and (n9744,n9614,n9621);
or (n9745,n9746,n9747);
and (n9746,n9589,n9612);
and (n9747,n9590,n9593);
or (n9748,n9749,n9750);
and (n9749,n9685,n9692);
and (n9750,n9686,n9689);
xor (n9751,n9752,n9835);
xor (n9752,n9753,n9785);
xor (n9753,n9754,n9761);
xor (n9754,n9755,n9758);
or (n9755,n9756,n9757);
and (n9756,n9637,n9651);
and (n9757,n9638,n9644);
or (n9758,n9759,n9760);
and (n9759,n9594,n9604);
and (n9760,n9595,n9597);
xor (n9761,n9762,n9779);
xor (n9762,n9763,n9771);
nand (n9763,n9764,n9766);
or (n9764,n9765,n7068);
not (n9765,n9648);
nand (n9766,n9767,n7075);
nand (n9767,n9768,n9770);
not (n9768,n9769);
and (n9769,n7129,n7065);
nand (n9770,n7067,n9391);
nand (n9771,n9772,n9776);
or (n9772,n7095,n9773);
nor (n9773,n9774,n9775);
and (n9774,n7145,n7092);
and (n9775,n7146,n7093);
nand (n9776,n9777,n9778);
not (n9777,n9655);
not (n9778,n7088);
nand (n9779,n9780,n9781);
or (n9780,n7978,n9663);
or (n9781,n9782,n9000);
nor (n9782,n9783,n9784);
and (n9783,n7852,n7204);
and (n9784,n7853,n7203);
xor (n9785,n9786,n9832);
xor (n9786,n9787,n9808);
xor (n9787,n9788,n9802);
xor (n9788,n9789,n9795);
nand (n9789,n9790,n9791);
or (n9790,n9608,n7998);
nand (n9791,n9792,n7749);
nor (n9792,n9793,n9794);
and (n9793,n8002,n7471);
and (n9794,n7859,n7470);
nand (n9795,n9796,n9798);
or (n9796,n9797,n7325);
not (n9797,n9618);
nand (n9798,n9799,n7327);
nor (n9799,n9800,n9801);
and (n9800,n7557,n7048);
and (n9801,n7558,n7049);
nand (n9802,n9803,n9804);
or (n9803,n9625,n7475);
nand (n9804,n7477,n9805);
nor (n9805,n9806,n9807);
and (n9806,n7919,n7483);
and (n9807,n7917,n7486);
xor (n9808,n9809,n9824);
xor (n9809,n9810,n9817);
nand (n9810,n9811,n9813);
or (n9811,n9812,n7207);
not (n9812,n9673);
nand (n9813,n7225,n9814);
nand (n9814,n9815,n9816);
or (n9815,n7866,n7205);
nand (n9816,n7205,n7866);
nand (n9817,n9818,n9820);
or (n9818,n9819,n7255);
not (n9819,n9601);
nand (n9820,n7264,n9821);
nand (n9821,n9822,n9823);
or (n9822,n7383,n7252);
nand (n9823,n7252,n7383);
nand (n9824,n9825,n9827);
or (n9825,n7038,n9826);
not (n9826,n9641);
or (n9827,n7046,n9828);
not (n9828,n9829);
nand (n9829,n9830,n9831);
or (n9830,n7036,n8125);
nand (n9831,n7036,n8125);
or (n9832,n9833,n9834);
and (n9833,n9659,n9668);
and (n9834,n9660,n9666);
or (n9835,n9836,n9837);
and (n9836,n9635,n9676);
and (n9837,n9636,n9658);
or (n9838,n9839,n9840);
and (n9839,n9683,n9706);
and (n9840,n9684,n9703);
nand (n9841,n9842,n10048);
nor (n9842,n9843,n9952);
nor (n9843,n9844,n9847);
or (n9844,n9845,n9846);
and (n9845,n9723,n9838);
and (n9846,n9724,n9727);
xor (n9847,n9848,n9949);
xor (n9848,n9849,n9915);
xor (n9849,n9850,n9865);
xor (n9850,n9851,n9862);
xor (n9851,n9852,n9859);
xor (n9852,n9853,n9856);
nor (n9853,n9854,n9855);
and (n9854,n7207,n7226);
not (n9855,n9814);
or (n9856,n9857,n9858);
and (n9857,n9809,n9824);
and (n9858,n9810,n9817);
or (n9859,n9860,n9861);
and (n9860,n9762,n9779);
and (n9861,n9763,n9771);
or (n9862,n9863,n9864);
and (n9863,n9786,n9832);
and (n9864,n9787,n9808);
xor (n9865,n9866,n9893);
xor (n9866,n9867,n9870);
or (n9867,n9868,n9869);
and (n9868,n9788,n9802);
and (n9869,n9789,n9795);
xor (n9870,n9871,n9885);
xor (n9871,n9872,n9878);
nand (n9872,n9873,n9874);
or (n9873,n9828,n7038);
nand (n9874,n9875,n7057);
nor (n9875,n9876,n9877);
and (n9876,n7172,n7035);
and (n9877,n7173,n7036);
nand (n9878,n9879,n9881);
or (n9879,n7068,n9880);
not (n9880,n9767);
or (n9881,n7349,n9882);
nor (n9882,n9883,n9884);
and (n9883,n7067,n8977);
and (n9884,n7134,n7065);
nand (n9885,n9886,n9892);
or (n9886,n7095,n9887);
not (n9887,n9888);
nand (n9888,n9889,n9890);
or (n9889,n7093,n7165);
not (n9890,n9891);
and (n9891,n7165,n7093);
or (n9892,n7088,n9773);
xor (n9893,n9894,n9909);
xor (n9894,n9895,n9902);
nand (n9895,n9896,n9898);
or (n9896,n9897,n7255);
not (n9897,n9821);
nand (n9898,n7264,n9899);
nor (n9899,n9900,n9901);
and (n9900,n7744,n7252);
and (n9901,n7745,n7253);
nand (n9902,n9903,n9905);
or (n9903,n7998,n9904);
not (n9904,n9792);
or (n9905,n9906,n7750);
nor (n9906,n9907,n9908);
and (n9907,n7308,n7859);
and (n9908,n7310,n8002);
nand (n9909,n9910,n9911);
or (n9910,n7978,n9782);
or (n9911,n9000,n9912);
nor (n9912,n9913,n9914);
and (n9913,n7852,n7223);
and (n9914,n7853,n7222);
xor (n9915,n9916,n9946);
xor (n9916,n9917,n9943);
xor (n9917,n9918,n9940);
xor (n9918,n9919,n9937);
xor (n9919,n9920,n9931);
xor (n9920,n9921,n9928);
nand (n9921,n9922,n9924);
or (n9922,n9923,n7325);
not (n9923,n9799);
nand (n9924,n7327,n9925);
nor (n9925,n9926,n9927);
and (n9926,n7390,n7048);
and (n9927,n7391,n7049);
nand (n9928,n9929,n9805);
or (n9929,n7477,n9930);
not (n9930,n7475);
nand (n9931,n9932,n9933);
or (n9932,n7523,n9739);
or (n9933,n7524,n9934);
nor (n9934,n9935,n9936);
and (n9935,n7077,n7244);
and (n9936,n7242,n7078);
or (n9937,n9938,n9939);
and (n9938,n9735,n9742);
and (n9939,n9736,n9669);
or (n9940,n9941,n9942);
and (n9941,n9754,n9761);
and (n9942,n9755,n9758);
or (n9943,n9944,n9945);
and (n9944,n9730,n9745);
and (n9945,n9731,n9734);
or (n9946,n9947,n9948);
and (n9947,n9752,n9835);
and (n9948,n9753,n9785);
or (n9949,n9950,n9951);
and (n9950,n9728,n9751);
and (n9951,n9729,n9748);
nor (n9952,n9953,n9956);
or (n9953,n9954,n9955);
and (n9954,n9848,n9949);
and (n9955,n9849,n9915);
xor (n9956,n9957,n10045);
xor (n9957,n9958,n9977);
xor (n9958,n9959,n9966);
xor (n9959,n9960,n9963);
or (n9960,n9961,n9962);
and (n9961,n9852,n9859);
and (n9962,n9853,n9856);
or (n9963,n9964,n9965);
and (n9964,n9866,n9893);
and (n9965,n9867,n9870);
xor (n9966,n9967,n9974);
xor (n9967,n9968,n9971);
or (n9968,n9969,n9970);
and (n9969,n9871,n9885);
and (n9970,n9872,n9878);
or (n9971,n9972,n9973);
and (n9972,n9894,n9909);
and (n9973,n9895,n9902);
or (n9974,n9975,n9976);
and (n9975,n9920,n9931);
and (n9976,n9921,n9928);
xor (n9977,n9978,n10042);
xor (n9978,n9979,n10039);
xor (n9979,n9980,n10024);
xor (n9980,n9981,n10003);
xor (n9981,n9982,n9997);
xor (n9982,n9983,n9990);
nand (n9983,n9984,n9986);
or (n9984,n9985,n7255);
not (n9985,n9899);
nand (n9986,n7264,n9987);
nor (n9987,n9988,n9989);
and (n9988,n7866,n7252);
and (n9989,n7867,n7253);
nand (n9990,n9991,n9993);
or (n9991,n9992,n7325);
not (n9992,n9925);
nand (n9993,n9994,n7327);
nor (n9994,n9995,n9996);
and (n9995,n7382,n7048);
and (n9996,n7383,n7049);
nand (n9997,n9998,n9999);
or (n9998,n7978,n9912);
or (n9999,n10000,n9000);
nor (n10000,n10001,n10002);
and (n10001,n7852,n7194);
and (n10002,n7853,n8125);
xor (n10003,n10004,n10017);
xor (n10004,n10005,n10011);
nand (n10005,n10006,n10007);
or (n10006,n9906,n7998);
or (n10007,n10008,n7750);
nor (n10008,n10009,n10010);
and (n10009,n7145,n8002);
and (n10010,n7146,n7859);
nand (n10011,n10012,n10013);
or (n10012,n9934,n7523);
nand (n10013,n7525,n10014);
nor (n10014,n10015,n10016);
and (n10015,n7919,n7078);
and (n10016,n7917,n7077);
nand (n10017,n10018,n10020);
or (n10018,n7038,n10019);
not (n10019,n9875);
or (n10020,n7046,n10021);
nor (n10021,n10022,n10023);
and (n10022,n7035,n7558);
and (n10023,n7036,n7557);
xor (n10024,n10025,n10038);
xor (n10025,n10026,n10032);
nand (n10026,n10027,n10028);
or (n10027,n7068,n9882);
or (n10028,n7349,n10029);
nor (n10029,n10030,n10031);
and (n10030,n7067,n7234);
and (n10031,n7232,n7065);
nand (n10032,n10033,n10034);
or (n10033,n9887,n7088);
or (n10034,n10035,n7095);
nor (n10035,n10036,n10037);
and (n10036,n7092,n9391);
and (n10037,n7129,n7093);
not (n10038,n9853);
or (n10039,n10040,n10041);
and (n10040,n9918,n9940);
and (n10041,n9919,n9937);
or (n10042,n10043,n10044);
and (n10043,n9850,n9865);
and (n10044,n9851,n9862);
or (n10045,n10046,n10047);
and (n10046,n9916,n9946);
and (n10047,n9917,n9943);
not (n10048,n10049);
nand (n10049,n10050,n10133,n10313,n10320);
nand (n10050,n10051,n10055);
not (n10051,n10052);
or (n10052,n10053,n10054);
and (n10053,n9957,n10045);
and (n10054,n9958,n9977);
not (n10055,n10056);
xor (n10056,n10057,n10130);
xor (n10057,n10058,n10061);
or (n10058,n10059,n10060);
and (n10059,n9959,n9966);
and (n10060,n9960,n9963);
xor (n10061,n10062,n10109);
xor (n10062,n10063,n10106);
xor (n10063,n10064,n10090);
xor (n10064,n10065,n10068);
or (n10065,n10066,n10067);
and (n10066,n10004,n10017);
and (n10067,n10005,n10011);
xor (n10068,n10069,n10084);
xor (n10069,n10070,n10078);
nand (n10070,n10071,n10073);
or (n10071,n10072,n7325);
not (n10072,n9994);
nand (n10073,n10074,n7327);
not (n10074,n10075);
nor (n10075,n10076,n10077);
and (n10076,n7048,n7745);
and (n10077,n7049,n7744);
nand (n10078,n10079,n10080);
or (n10079,n7998,n10008);
or (n10080,n10081,n7750);
nor (n10081,n10082,n10083);
and (n10082,n8002,n7164);
and (n10083,n7165,n7859);
nand (n10084,n10085,n10086);
or (n10085,n7978,n10000);
or (n10086,n9000,n10087);
nor (n10087,n10088,n10089);
and (n10088,n7852,n7173);
and (n10089,n7853,n7172);
xor (n10090,n10091,n10100);
xor (n10091,n10092,n10094);
nand (n10092,n10093,n10014);
or (n10093,n7525,n7901);
nand (n10094,n10095,n10096);
or (n10095,n7038,n10021);
or (n10096,n7046,n10097);
nor (n10097,n10098,n10099);
and (n10098,n7035,n7391);
and (n10099,n7036,n7390);
nand (n10100,n10101,n10102);
or (n10101,n7068,n10029);
or (n10102,n7349,n10103);
nor (n10103,n10104,n10105);
and (n10104,n7067,n7244);
and (n10105,n7242,n7065);
or (n10106,n10107,n10108);
and (n10107,n9980,n10024);
and (n10108,n9981,n10003);
xor (n10109,n10110,n10127);
xor (n10110,n10111,n10114);
or (n10111,n10112,n10113);
and (n10112,n10025,n10038);
and (n10113,n10026,n10032);
xor (n10114,n10115,n10124);
xor (n10115,n10116,n10122);
nand (n10116,n10117,n10118);
or (n10117,n7088,n10035);
or (n10118,n10119,n7095);
nor (n10119,n10120,n10121);
and (n10120,n7092,n8977);
and (n10121,n7134,n7093);
and (n10122,n10123,n9987);
nand (n10123,n7255,n9205);
or (n10124,n10125,n10126);
and (n10125,n9982,n9997);
and (n10126,n9983,n9990);
or (n10127,n10128,n10129);
and (n10128,n9967,n9974);
and (n10129,n9968,n9971);
or (n10130,n10131,n10132);
and (n10131,n9978,n10042);
and (n10132,n9979,n10039);
nor (n10133,n10134,n10263);
nor (n10134,n10135,n10206);
or (n10135,n10136,n10205);
and (n10136,n10137,n10202);
xor (n10137,n10138,n10185);
xor (n10138,n10139,n10182);
xor (n10139,n10140,n10162);
xor (n10140,n10141,n10156);
xor (n10141,n10142,n10150);
nand (n10142,n10143,n10148);
or (n10143,n7095,n10144);
not (n10144,n10145);
nor (n10145,n10146,n10147);
and (n10146,n7234,n7093);
and (n10147,n7232,n7092);
nand (n10148,n10149,n9778);
not (n10149,n10119);
nand (n10150,n10151,n10152);
or (n10151,n7978,n10087);
or (n10152,n9000,n10153);
nor (n10153,n10154,n10155);
and (n10154,n7852,n7558);
and (n10155,n7853,n7557);
nand (n10156,n10157,n10158);
or (n10157,n7998,n10081);
or (n10158,n10159,n7750);
nor (n10159,n10160,n10161);
and (n10160,n8002,n9391);
and (n10161,n7129,n7859);
xor (n10162,n10163,n10176);
xor (n10163,n10164,n10170);
nand (n10164,n10165,n10166);
or (n10165,n7325,n10075);
or (n10166,n7326,n10167);
nor (n10167,n10168,n10169);
and (n10168,n7048,n7867);
and (n10169,n7049,n7866);
nand (n10170,n10171,n10172);
or (n10171,n7038,n10097);
or (n10172,n7046,n10173);
nor (n10173,n10174,n10175);
and (n10174,n7035,n7383);
and (n10175,n7036,n7382);
nand (n10176,n10177,n10178);
or (n10177,n7068,n10103);
or (n10178,n7349,n10179);
nor (n10179,n10180,n10181);
and (n10180,n7067,n7919);
and (n10181,n7917,n7065);
or (n10182,n10183,n10184);
and (n10183,n10115,n10124);
and (n10184,n10116,n10122);
xor (n10185,n10186,n10199);
xor (n10186,n10187,n10196);
xor (n10187,n10188,n10193);
xor (n10188,n10189,n10190);
not (n10189,n10122);
or (n10190,n10191,n10192);
and (n10191,n10069,n10084);
and (n10192,n10070,n10078);
or (n10193,n10194,n10195);
and (n10194,n10091,n10100);
and (n10195,n10092,n10094);
or (n10196,n10197,n10198);
and (n10197,n10064,n10090);
and (n10198,n10065,n10068);
or (n10199,n10200,n10201);
and (n10200,n10110,n10127);
and (n10201,n10111,n10114);
or (n10202,n10203,n10204);
and (n10203,n10062,n10109);
and (n10204,n10063,n10106);
and (n10205,n10138,n10185);
xor (n10206,n10207,n10260);
xor (n10207,n10208,n10211);
or (n10208,n10209,n10210);
and (n10209,n10139,n10182);
and (n10210,n10140,n10162);
xor (n10211,n10212,n10237);
xor (n10212,n10213,n10234);
xor (n10213,n10214,n10227);
xor (n10214,n10215,n10221);
nand (n10215,n10216,n10217);
or (n10216,n7998,n10159);
or (n10217,n10218,n7750);
nor (n10218,n10219,n10220);
and (n10219,n8002,n8977);
and (n10220,n7134,n7859);
nand (n10221,n10222,n10223);
or (n10222,n7978,n10153);
or (n10223,n9000,n10224);
nor (n10224,n10225,n10226);
and (n10225,n7852,n7391);
and (n10226,n7853,n7390);
not (n10227,n10228);
nand (n10228,n10229,n10230);
or (n10229,n7038,n10173);
or (n10230,n7046,n10231);
nor (n10231,n10232,n10233);
and (n10232,n7035,n7745);
and (n10233,n7036,n7744);
or (n10234,n10235,n10236);
and (n10235,n10188,n10193);
and (n10236,n10189,n10190);
xor (n10237,n10238,n10245);
xor (n10238,n10239,n10242);
or (n10239,n10240,n10241);
and (n10240,n10141,n10156);
and (n10241,n10142,n10150);
or (n10242,n10243,n10244);
and (n10243,n10163,n10176);
and (n10244,n10164,n10170);
xor (n10245,n10246,n10256);
xor (n10246,n10247,n10250);
nand (n10247,n10248,n10249);
or (n10248,n7075,n7069);
not (n10249,n10179);
nand (n10250,n10251,n10252);
or (n10251,n7088,n10144);
or (n10252,n10253,n7095);
nor (n10253,n10254,n10255);
and (n10254,n7092,n7244);
and (n10255,n7242,n7093);
nand (n10256,n10257,n10259);
or (n10257,n7327,n10258);
not (n10258,n7325);
not (n10259,n10167);
or (n10260,n10261,n10262);
and (n10261,n10186,n10199);
and (n10262,n10187,n10196);
nor (n10263,n10264,n10267);
or (n10264,n10265,n10266);
and (n10265,n10207,n10260);
and (n10266,n10208,n10211);
xor (n10267,n10268,n10310);
xor (n10268,n10269,n10272);
or (n10269,n10270,n10271);
and (n10270,n10238,n10245);
and (n10271,n10239,n10242);
xor (n10272,n10273,n10299);
xor (n10273,n10274,n10296);
xor (n10274,n10275,n10290);
xor (n10275,n10276,n10282);
nand (n10276,n10277,n10278);
or (n10277,n7038,n10231);
or (n10278,n7046,n10279);
nor (n10279,n10280,n10281);
and (n10280,n7035,n7867);
and (n10281,n7036,n7866);
nand (n10282,n10283,n10288);
or (n10283,n10284,n9000);
not (n10284,n10285);
nor (n10285,n10286,n10287);
and (n10286,n7382,n7852);
and (n10287,n7383,n7853);
nand (n10288,n10289,n7979);
not (n10289,n10224);
nand (n10290,n10291,n10292);
or (n10291,n7998,n10218);
or (n10292,n10293,n7750);
nor (n10293,n10294,n10295);
and (n10294,n8002,n7234);
and (n10295,n7232,n7859);
or (n10296,n10297,n10298);
and (n10297,n10214,n10227);
and (n10298,n10215,n10221);
xor (n10299,n10300,n10307);
xor (n10300,n10301,n10228);
nand (n10301,n10302,n10303);
or (n10302,n7088,n10253);
or (n10303,n10304,n7095);
nor (n10304,n10305,n10306);
and (n10305,n7092,n7919);
and (n10306,n7917,n7093);
or (n10307,n10308,n10309);
and (n10308,n10246,n10256);
and (n10309,n10247,n10250);
or (n10310,n10311,n10312);
and (n10311,n10212,n10237);
and (n10312,n10213,n10234);
nand (n10313,n10314,n10318);
not (n10314,n10315);
or (n10315,n10316,n10317);
and (n10316,n10057,n10130);
and (n10317,n10058,n10061);
not (n10318,n10319);
xor (n10319,n10137,n10202);
nor (n10320,n10321,n10360);
nor (n10321,n10322,n10325);
or (n10322,n10323,n10324);
and (n10323,n10268,n10310);
and (n10324,n10269,n10272);
xor (n10325,n10326,n10357);
xor (n10326,n10327,n10330);
or (n10327,n10328,n10329);
and (n10328,n10300,n10307);
and (n10329,n10301,n10228);
xor (n10330,n10331,n10340);
xor (n10331,n10332,n10337);
not (n10332,n10333);
nand (n10333,n10334,n10336);
or (n10334,n7057,n10335);
not (n10335,n7038);
not (n10336,n10279);
or (n10337,n10338,n10339);
and (n10338,n10275,n10290);
and (n10339,n10276,n10282);
xor (n10340,n10341,n10354);
xor (n10341,n10342,n10348);
nand (n10342,n10343,n10344);
or (n10343,n7998,n10293);
or (n10344,n10345,n7750);
nor (n10345,n10346,n10347);
and (n10346,n8002,n7244);
and (n10347,n7242,n7859);
nand (n10348,n10349,n10350);
or (n10349,n10284,n7978);
or (n10350,n9000,n10351);
nor (n10351,n10352,n10353);
and (n10352,n7852,n7745);
and (n10353,n7853,n7744);
nand (n10354,n10355,n10356);
or (n10355,n7788,n9778);
not (n10356,n10304);
or (n10357,n10358,n10359);
and (n10358,n10273,n10299);
and (n10359,n10274,n10296);
nand (n10360,n10361,n10387);
or (n10361,n10362,n10384);
xor (n10362,n10363,n10381);
xor (n10363,n10364,n10367);
or (n10364,n10365,n10366);
and (n10365,n10341,n10354);
and (n10366,n10342,n10348);
xor (n10367,n10368,n10333);
xor (n10368,n10369,n10375);
nand (n10369,n10370,n10371);
or (n10370,n7978,n10351);
or (n10371,n9000,n10372);
nor (n10372,n10373,n10374);
and (n10373,n7852,n7867);
and (n10374,n7853,n7866);
nand (n10375,n10376,n10377);
or (n10376,n7998,n10345);
or (n10377,n10378,n7750);
nor (n10378,n10379,n10380);
and (n10379,n8002,n7919);
and (n10380,n7917,n7859);
or (n10381,n10382,n10383);
and (n10382,n10331,n10340);
and (n10383,n10332,n10337);
or (n10384,n10385,n10386);
and (n10385,n10326,n10357);
and (n10386,n10327,n10330);
nand (n10387,n10388,n10392);
not (n10388,n10389);
or (n10389,n10390,n10391);
and (n10390,n10363,n10381);
and (n10391,n10364,n10367);
not (n10392,n10393);
xor (n10393,n10394,n10400);
xor (n10394,n10395,n10398);
nand (n10395,n10396,n10397);
or (n10396,n7979,n7756);
not (n10397,n10372);
nor (n10398,n10399,n10378);
and (n10399,n7998,n7750);
or (n10400,n10401,n10402);
and (n10401,n10368,n10333);
and (n10402,n10369,n10375);
nand (n10403,n10404,n9580);
nand (n10404,n10405,n10413);
or (n10405,n8919,n10406);
not (n10406,n10407);
nand (n10407,n10408,n10411);
or (n10408,n10409,n10410);
not (n10409,n9563);
not (n10410,n9564);
or (n10411,n9562,n10412);
nand (n10412,n9575,n9577);
nand (n10413,n10414,n10415);
not (n10414,n8921);
nand (n10415,n10416,n10419);
or (n10416,n10417,n10418);
not (n10417,n9488);
not (n10418,n8922);
nand (n10419,n9542,n9543);
nand (n10420,n10421,n10048);
or (n10421,n10422,n10428);
nor (n10422,n10423,n10427);
and (n10423,n10424,n10426);
nand (n10424,n9716,n10425);
nor (n10425,n9583,n9712);
nand (n10426,n9718,n9722);
not (n10427,n9842);
nor (n10428,n10429,n9952);
and (n10429,n10430,n10431);
nand (n10430,n9844,n9847);
nand (n10431,n9953,n9956);
nor (n10432,n10433,n10447);
and (n10433,n10434,n10320);
nand (n10434,n10435,n10443);
or (n10435,n10436,n10437);
not (n10436,n10133);
not (n10437,n10438);
nand (n10438,n10439,n10440);
or (n10439,n10318,n10314);
or (n10440,n10441,n10442);
not (n10441,n10313);
nand (n10442,n10052,n10056);
nor (n10443,n10444,n10446);
and (n10444,n10135,n10445,n10206);
not (n10445,n10263);
and (n10446,n10264,n10267);
nand (n10447,n10448,n10453);
or (n10448,n10449,n10452);
nor (n10449,n10450,n10451);
and (n10450,n10322,n10361,n10325);
and (n10451,n10384,n10362);
not (n10452,n10387);
or (n10453,n10388,n10392);
nor (n10454,n10455,n10460);
and (n10455,n10456,n10459);
or (n10456,n10457,n10458);
and (n10457,n10394,n10400);
and (n10458,n10395,n10398);
not (n10459,n10398);
and (n10460,n10461,n10398);
not (n10461,n10456);
nor (n10463,n10464,n10587);
and (n10464,n10465,n10568);
nand (n10465,n10466,n10490,n10496);
or (n10466,n10467,n10483);
nand (n10467,n10468,n10473,n10478);
not (n10468,n10469);
and (n10469,n10470,n10472);
not (n10470,n10471);
not (n10473,n10474);
and (n10474,n10475,n10477);
not (n10475,n10476);
not (n10478,n10479);
and (n10479,n10480,n10482);
not (n10480,n10481);
nor (n10483,n10484,n10488);
and (n10484,n10485,n10486);
not (n10486,n10487);
and (n10488,n10481,n10489);
not (n10489,n10482);
or (n10490,n10469,n10491);
nor (n10491,n10492,n10494);
and (n10492,n10476,n10493);
not (n10493,n10477);
and (n10494,n10471,n10495);
not (n10495,n10472);
nand (n10496,n10497,n10564,n10567);
or (n10497,n10498,n10558);
nor (n10498,n10499,n10544);
and (n10499,n10500,n10537);
nand (n10500,n10501,n10525,n10532);
or (n10501,n10502,n10523);
nor (n10502,n10503,n10505,n10522);
not (n10503,n10504);
nor (n10505,n10506,n10520);
and (n10506,n10507,n10519);
not (n10507,n10508);
or (n10508,n10509,n10513);
and (n10509,n10510,n10512);
not (n10510,n10511);
and (n10513,n10514,n10518);
and (n10514,n10515,n10517);
not (n10515,n10516);
xnor (n10518,n10512,n10511);
not (n10520,n10521);
nor (n10522,n10507,n10519);
not (n10523,n10524);
or (n10525,n10504,n10526);
not (n10526,n10527);
or (n10527,n10528,n10530);
and (n10528,n10529,n10521);
not (n10529,n10519);
and (n10530,n10508,n10531);
xnor (n10531,n10521,n10519);
not (n10532,n10533);
and (n10533,n10534,n10536);
not (n10534,n10535);
nor (n10537,n10538,n10540);
and (n10538,n10535,n10539);
not (n10539,n10536);
and (n10540,n10541,n10542);
not (n10542,n10543);
nand (n10544,n10545,n10550,n10555);
not (n10545,n10546);
and (n10546,n10547,n10549);
not (n10547,n10548);
not (n10550,n10551);
and (n10551,n10552,n10554);
not (n10552,n10553);
not (n10555,n10556);
and (n10556,n10557,n10543);
not (n10557,n10541);
nor (n10558,n10559,n10562);
and (n10559,n10560,n10554);
nand (n10560,n10548,n10553,n10561);
not (n10561,n10549);
nor (n10562,n10563,n10553);
and (n10563,n10548,n10561);
not (n10564,n10565);
and (n10565,n10566,n10487);
not (n10566,n10485);
not (n10567,n10467);
nor (n10568,n10569,n10573,n10583);
and (n10569,n10570,n10572);
not (n10570,n10571);
nand (n10573,n10574,n10579);
not (n10574,n10575);
and (n10575,n10576,n10578);
not (n10576,n10577);
nand (n10579,n10580,n10582);
not (n10580,n10581);
and (n10583,n10584,n10586);
not (n10584,n10585);
nand (n10587,n10588,n10595);
or (n10588,n10573,n10589);
nor (n10589,n10590,n10593);
and (n10590,n10591,n10571,n10592);
not (n10591,n10583);
not (n10592,n10572);
and (n10593,n10585,n10594);
not (n10594,n10586);
nor (n10595,n10596,n10598);
and (n10596,n10579,n10577,n10597);
not (n10597,n10578);
and (n10598,n10581,n10599);
not (n10599,n10582);
not (n10600,n10601);
nor (n10601,n10602,n10706,n10710);
and (n10602,n10603,n10687);
nand (n10603,n10604,n10677);
nand (n10604,n10605,n10658,n10671);
nand (n10605,n10606,n10610,n10614);
or (n10606,n10607,n10608);
not (n10608,n10609);
or (n10610,n10611,n10613);
not (n10611,n10612);
nand (n10614,n10615,n10651);
or (n10615,n10616,n10650);
and (n10616,n10617,n10647,n10648);
nand (n10617,n10618,n10645);
or (n10618,n10619,n10644);
or (n10619,n10620,n10624);
and (n10620,n10621,n10623);
not (n10621,n10622);
and (n10624,n10625,n10643);
or (n10625,n10626,n10630);
and (n10626,n10627,n10629);
not (n10627,n10628);
and (n10630,n10631,n10642);
not (n10631,n10632);
nand (n10632,n10633,n10639,n10640);
or (n10633,n10634,n10638);
and (n10634,n10635,n10636,n2);
not (n10636,n10637);
or (n10639,n2,n10635);
not (n10640,n10641);
and (n10641,n3,n10637);
xnor (n10642,n10628,n10629);
xnor (n10643,n10622,n10623);
not (n10645,n10646);
nand (n10647,n10619,n10644);
not (n10648,n10649);
nor (n10651,n10652,n10657);
and (n10652,n10653,n10649);
or (n10653,n10654,n10655);
and (n10654,n10645,n10644);
and (n10655,n10619,n10656);
xnor (n10656,n10646,n10644);
and (n10657,n10608,n10607);
nor (n10658,n10659,n10663,n10667);
and (n10659,n10660,n10662);
not (n10660,n10661);
and (n10663,n10664,n10666);
not (n10664,n10665);
and (n10667,n10668,n10670);
not (n10668,n10669);
nor (n10671,n10672,n10676);
and (n10672,n10673,n10675);
not (n10673,n10674);
and (n10676,n10611,n10613);
nor (n10677,n10678,n10682);
and (n10678,n10658,n10679);
nand (n10679,n10680,n10681);
or (n10680,n10675,n10673);
or (n10681,n10666,n10664);
and (n10682,n10683,n10685);
nand (n10683,n10684,n10668);
or (n10684,n10662,n10670,n10660);
nand (n10685,n10686,n10670);
or (n10686,n10662,n10660);
nor (n10687,n10688,n10692,n10702);
and (n10688,n10689,n10691);
not (n10689,n10690);
not (n10692,n10693);
nor (n10693,n10694,n10698);
and (n10694,n10695,n10697);
not (n10695,n10696);
and (n10698,n10699,n10701);
not (n10699,n10700);
and (n10702,n10703,n10705);
not (n10703,n10704);
and (n10706,n10693,n10707);
nand (n10707,n10708,n10709);
or (n10708,n10702,n10691,n10689);
or (n10709,n10705,n10703);
nand (n10710,n10711,n10712);
or (n10711,n10698,n10697,n10695);
or (n10712,n10701,n10699);
and (n10713,n10714,n10715);
nand (n10716,n4,n10717);
or (n10718,n10719,n22700);
and (n10719,n10720,n10713);
wire s0n10720,s1n10720,notn10720;
or (n10720,s0n10720,s1n10720);
not(notn10720,n10721);
and (s0n10720,notn10720,n3);
and (s1n10720,n10721,n10717);
and (n10721,n10600,n10722);
or (n10722,n10463,n10723);
and (n10723,n10724,n10462);
not (n10724,n10725);
and (n10725,n10726,n18719);
and (n10726,n10727,n14722);
not (n10727,n10728);
xor (n10728,n10729,n14510);
xor (n10729,n10730,n12641);
xor (n10730,n10731,n12088);
xor (n10731,n10732,n12639);
xor (n10732,n10733,n12083);
xor (n10733,n10734,n12632);
xor (n10734,n10735,n12077);
xor (n10735,n10736,n12620);
xor (n10736,n10737,n3953);
xor (n10737,n10738,n12603);
xor (n10738,n10739,n12066);
xor (n10739,n10740,n12581);
xor (n10740,n10741,n12060);
xor (n10741,n10742,n12554);
xor (n10742,n10743,n3792);
xor (n10743,n10744,n12522);
xor (n10744,n10745,n4259);
xor (n10745,n10746,n12485);
xor (n10746,n10747,n12044);
xor (n10747,n10748,n12443);
xor (n10748,n10749,n12038);
xor (n10749,n10750,n12396);
xor (n10750,n10751,n12032);
xor (n10751,n10752,n12344);
xor (n10752,n10753,n12026);
xor (n10753,n10754,n12287);
xor (n10754,n10755,n12020);
xor (n10755,n10756,n12225);
xor (n10756,n10757,n12014);
xor (n10757,n10758,n12158);
xor (n10758,n10759,n12008);
xor (n10759,n10760,n10822);
xor (n10760,n10761,n10820);
xor (n10761,n10762,n10821);
xor (n10762,n10763,n10820);
xor (n10763,n10764,n10819);
xor (n10764,n10765,n10818);
xor (n10765,n10766,n10817);
xor (n10766,n10767,n10816);
xor (n10767,n10768,n10815);
xor (n10768,n10769,n10814);
xor (n10769,n10770,n10813);
xor (n10770,n10771,n10812);
xor (n10771,n10772,n10811);
xor (n10772,n10773,n10810);
xor (n10773,n10774,n10809);
xor (n10774,n10775,n10808);
xor (n10775,n10776,n10807);
xor (n10776,n10777,n10806);
xor (n10777,n10778,n10805);
xor (n10778,n10779,n10804);
xor (n10779,n10780,n10803);
xor (n10780,n10781,n10802);
xor (n10781,n10782,n10801);
xor (n10782,n10783,n10800);
xor (n10783,n10784,n10799);
xor (n10784,n10785,n10798);
xor (n10785,n10786,n10797);
xor (n10786,n10787,n10796);
xor (n10787,n10788,n10795);
xor (n10788,n10789,n10794);
xor (n10789,n10790,n10793);
xor (n10790,n10791,n10792);
and (n10791,n3615,n4384);
and (n10792,n3615,n3867);
and (n10793,n10791,n10792);
and (n10794,n3615,n3866);
and (n10795,n10789,n10794);
and (n10796,n3615,n3603);
and (n10797,n10787,n10796);
and (n10798,n3615,n3602);
and (n10799,n10785,n10798);
and (n10800,n3615,n3611);
and (n10801,n10783,n10800);
and (n10802,n3615,n3828);
and (n10803,n10781,n10802);
and (n10804,n3615,n3632);
and (n10805,n10779,n10804);
and (n10806,n3615,n3633);
and (n10807,n10777,n10806);
and (n10808,n3615,n3624);
and (n10809,n10775,n10808);
and (n10810,n3615,n3687);
and (n10811,n10773,n10810);
and (n10812,n3615,n3573);
and (n10813,n10771,n10812);
and (n10814,n3615,n3575);
and (n10815,n10769,n10814);
and (n10816,n3615,n3581);
and (n10817,n10767,n10816);
and (n10818,n3615,n3783);
and (n10819,n10765,n10818);
and (n10820,n3615,n3790);
and (n10821,n10763,n10820);
or (n10822,n10823,n12089);
and (n10823,n10824,n12008);
xor (n10824,n10762,n10825);
or (n10825,n10826,n12009);
and (n10826,n10827,n12008);
xor (n10827,n10764,n10828);
or (n10828,n10829,n11926);
and (n10829,n10830,n11925);
xor (n10830,n10766,n10831);
or (n10831,n10832,n11845);
and (n10832,n10833,n11844);
xor (n10833,n10768,n10834);
or (n10834,n10835,n11762);
and (n10835,n10836,n11761);
xor (n10836,n10770,n10837);
or (n10837,n10838,n11686);
and (n10838,n10839,n11685);
xor (n10839,n10772,n10840);
or (n10840,n10841,n11603);
and (n10841,n10842,n11602);
xor (n10842,n10774,n10843);
or (n10843,n10844,n11522);
and (n10844,n10845,n11521);
xor (n10845,n10776,n10846);
or (n10846,n10847,n11439);
and (n10847,n10848,n11438);
xor (n10848,n10778,n10849);
or (n10849,n10850,n11357);
and (n10850,n10851,n11356);
xor (n10851,n10780,n10852);
or (n10852,n10853,n11274);
and (n10853,n10854,n11273);
xor (n10854,n10782,n10855);
or (n10855,n10856,n11194);
and (n10856,n10857,n11193);
xor (n10857,n10784,n10858);
or (n10858,n10859,n11111);
and (n10859,n10860,n11110);
xor (n10860,n10786,n10861);
or (n10861,n10862,n11030);
and (n10862,n10863,n11029);
xor (n10863,n10788,n10864);
or (n10864,n10865,n10947);
and (n10865,n10866,n10946);
xor (n10866,n10790,n10867);
or (n10867,n10868,n10870);
and (n10868,n10791,n10869);
and (n10869,n3843,n3867);
and (n10870,n10871,n10872);
xor (n10871,n10791,n10869);
or (n10872,n10873,n10876);
and (n10873,n10874,n10875);
and (n10874,n3843,n4384);
and (n10875,n3837,n3867);
and (n10876,n10877,n10878);
xor (n10877,n10874,n10875);
or (n10878,n10879,n10882);
and (n10879,n10880,n10881);
and (n10880,n3837,n4384);
and (n10881,n3641,n3867);
and (n10882,n10883,n10884);
xor (n10883,n10880,n10881);
or (n10884,n10885,n10888);
and (n10885,n10886,n10887);
and (n10886,n3641,n4384);
and (n10887,n3622,n3867);
and (n10888,n10889,n10890);
xor (n10889,n10886,n10887);
or (n10890,n10891,n10894);
and (n10891,n10892,n10893);
and (n10892,n3622,n4384);
and (n10893,n3695,n3867);
and (n10894,n10895,n10896);
xor (n10895,n10892,n10893);
or (n10896,n10897,n10899);
and (n10897,n10898,n6116);
and (n10898,n3695,n4384);
and (n10899,n10900,n10901);
xor (n10900,n10898,n6116);
or (n10901,n10902,n10904);
and (n10902,n10903,n6171);
and (n10903,n3680,n4384);
and (n10904,n10905,n10906);
xor (n10905,n10903,n6171);
or (n10906,n10907,n10910);
and (n10907,n10908,n10909);
and (n10908,n3723,n4384);
and (n10909,n3592,n3867);
and (n10910,n10911,n10912);
xor (n10911,n10908,n10909);
or (n10912,n10913,n10916);
and (n10913,n10914,n10915);
and (n10914,n3592,n4384);
and (n10915,n3586,n3867);
and (n10916,n10917,n10918);
xor (n10917,n10914,n10915);
or (n10918,n10919,n10921);
and (n10919,n10920,n6507);
and (n10920,n3586,n4384);
and (n10921,n10922,n10923);
xor (n10922,n10920,n6507);
or (n10923,n10924,n10926);
and (n10924,n10925,n6625);
and (n10925,n3800,n4384);
and (n10926,n10927,n10928);
xor (n10927,n10925,n6625);
or (n10928,n10929,n10931);
and (n10929,n10930,n6720);
and (n10930,n3959,n4384);
and (n10931,n10932,n10933);
xor (n10932,n10930,n6720);
or (n10933,n10934,n10936);
and (n10934,n10935,n6785);
and (n10935,n3952,n4384);
and (n10936,n10937,n10938);
xor (n10937,n10935,n6785);
or (n10938,n10939,n10941);
and (n10939,n10940,n6800);
and (n10940,n4350,n4384);
and (n10941,n10942,n10943);
xor (n10942,n10940,n6800);
and (n10943,n10944,n10945);
and (n10944,n4406,n4384);
and (n10945,n5233,n3867);
and (n10946,n3843,n3866);
and (n10947,n10948,n10949);
xor (n10948,n10866,n10946);
or (n10949,n10950,n10953);
and (n10950,n10951,n10952);
xor (n10951,n10871,n10872);
and (n10952,n3837,n3866);
and (n10953,n10954,n10955);
xor (n10954,n10951,n10952);
or (n10955,n10956,n10959);
and (n10956,n10957,n10958);
xor (n10957,n10877,n10878);
and (n10958,n3641,n3866);
and (n10959,n10960,n10961);
xor (n10960,n10957,n10958);
or (n10961,n10962,n10965);
and (n10962,n10963,n10964);
xor (n10963,n10883,n10884);
and (n10964,n3622,n3866);
and (n10965,n10966,n10967);
xor (n10966,n10963,n10964);
or (n10967,n10968,n10971);
and (n10968,n10969,n10970);
xor (n10969,n10889,n10890);
and (n10970,n3695,n3866);
and (n10971,n10972,n10973);
xor (n10972,n10969,n10970);
or (n10973,n10974,n10977);
and (n10974,n10975,n10976);
xor (n10975,n10895,n10896);
and (n10976,n3680,n3866);
and (n10977,n10978,n10979);
xor (n10978,n10975,n10976);
or (n10979,n10980,n10983);
and (n10980,n10981,n10982);
xor (n10981,n10900,n10901);
and (n10982,n3723,n3866);
and (n10983,n10984,n10985);
xor (n10984,n10981,n10982);
or (n10985,n10986,n10989);
and (n10986,n10987,n10988);
xor (n10987,n10905,n10906);
and (n10988,n3592,n3866);
and (n10989,n10990,n10991);
xor (n10990,n10987,n10988);
or (n10991,n10992,n10995);
and (n10992,n10993,n10994);
xor (n10993,n10911,n10912);
and (n10994,n3586,n3866);
and (n10995,n10996,n10997);
xor (n10996,n10993,n10994);
or (n10997,n10998,n11001);
and (n10998,n10999,n11000);
xor (n10999,n10917,n10918);
and (n11000,n3800,n3866);
and (n11001,n11002,n11003);
xor (n11002,n10999,n11000);
or (n11003,n11004,n11007);
and (n11004,n11005,n11006);
xor (n11005,n10922,n10923);
and (n11006,n3959,n3866);
and (n11007,n11008,n11009);
xor (n11008,n11005,n11006);
or (n11009,n11010,n11013);
and (n11010,n11011,n11012);
xor (n11011,n10927,n10928);
and (n11012,n3952,n3866);
and (n11013,n11014,n11015);
xor (n11014,n11011,n11012);
or (n11015,n11016,n11019);
and (n11016,n11017,n11018);
xor (n11017,n10932,n10933);
and (n11018,n4350,n3866);
and (n11019,n11020,n11021);
xor (n11020,n11017,n11018);
or (n11021,n11022,n11025);
and (n11022,n11023,n11024);
xor (n11023,n10937,n10938);
and (n11024,n4406,n3866);
and (n11025,n11026,n11027);
xor (n11026,n11023,n11024);
and (n11027,n11028,n6728);
xor (n11028,n10942,n10943);
and (n11029,n3843,n3603);
and (n11030,n11031,n11032);
xor (n11031,n10863,n11029);
or (n11032,n11033,n11036);
and (n11033,n11034,n11035);
xor (n11034,n10948,n10949);
and (n11035,n3837,n3603);
and (n11036,n11037,n11038);
xor (n11037,n11034,n11035);
or (n11038,n11039,n11042);
and (n11039,n11040,n11041);
xor (n11040,n10954,n10955);
and (n11041,n3641,n3603);
and (n11042,n11043,n11044);
xor (n11043,n11040,n11041);
or (n11044,n11045,n11048);
and (n11045,n11046,n11047);
xor (n11046,n10960,n10961);
and (n11047,n3622,n3603);
and (n11048,n11049,n11050);
xor (n11049,n11046,n11047);
or (n11050,n11051,n11054);
and (n11051,n11052,n11053);
xor (n11052,n10966,n10967);
and (n11053,n3695,n3603);
and (n11054,n11055,n11056);
xor (n11055,n11052,n11053);
or (n11056,n11057,n11060);
and (n11057,n11058,n11059);
xor (n11058,n10972,n10973);
and (n11059,n3680,n3603);
and (n11060,n11061,n11062);
xor (n11061,n11058,n11059);
or (n11062,n11063,n11066);
and (n11063,n11064,n11065);
xor (n11064,n10978,n10979);
and (n11065,n3723,n3603);
and (n11066,n11067,n11068);
xor (n11067,n11064,n11065);
or (n11068,n11069,n11071);
and (n11069,n11070,n6049);
xor (n11070,n10984,n10985);
and (n11071,n11072,n11073);
xor (n11072,n11070,n6049);
or (n11073,n11074,n11077);
and (n11074,n11075,n11076);
xor (n11075,n10990,n10991);
and (n11076,n3586,n3603);
and (n11077,n11078,n11079);
xor (n11078,n11075,n11076);
or (n11079,n11080,n11082);
and (n11080,n11081,n6318);
xor (n11081,n10996,n10997);
and (n11082,n11083,n11084);
xor (n11083,n11081,n6318);
or (n11084,n11085,n11088);
and (n11085,n11086,n11087);
xor (n11086,n11002,n11003);
and (n11087,n3959,n3603);
and (n11088,n11089,n11090);
xor (n11089,n11086,n11087);
or (n11090,n11091,n11093);
and (n11091,n11092,n6519);
xor (n11092,n11008,n11009);
and (n11093,n11094,n11095);
xor (n11094,n11092,n6519);
or (n11095,n11096,n11099);
and (n11096,n11097,n11098);
xor (n11097,n11014,n11015);
and (n11098,n4350,n3603);
and (n11099,n11100,n11101);
xor (n11100,n11097,n11098);
or (n11101,n11102,n11105);
and (n11102,n11103,n11104);
xor (n11103,n11020,n11021);
and (n11104,n4406,n3603);
and (n11105,n11106,n11107);
xor (n11106,n11103,n11104);
and (n11107,n11108,n11109);
xor (n11108,n11026,n11027);
and (n11109,n5233,n3603);
and (n11110,n3843,n3602);
and (n11111,n11112,n11113);
xor (n11112,n10860,n11110);
or (n11113,n11114,n11117);
and (n11114,n11115,n11116);
xor (n11115,n11031,n11032);
and (n11116,n3837,n3602);
and (n11117,n11118,n11119);
xor (n11118,n11115,n11116);
or (n11119,n11120,n11123);
and (n11120,n11121,n11122);
xor (n11121,n11037,n11038);
and (n11122,n3641,n3602);
and (n11123,n11124,n11125);
xor (n11124,n11121,n11122);
or (n11125,n11126,n11129);
and (n11126,n11127,n11128);
xor (n11127,n11043,n11044);
and (n11128,n3622,n3602);
and (n11129,n11130,n11131);
xor (n11130,n11127,n11128);
or (n11131,n11132,n11135);
and (n11132,n11133,n11134);
xor (n11133,n11049,n11050);
and (n11134,n3695,n3602);
and (n11135,n11136,n11137);
xor (n11136,n11133,n11134);
or (n11137,n11138,n11141);
and (n11138,n11139,n11140);
xor (n11139,n11055,n11056);
and (n11140,n3680,n3602);
and (n11141,n11142,n11143);
xor (n11142,n11139,n11140);
or (n11143,n11144,n11147);
and (n11144,n11145,n11146);
xor (n11145,n11061,n11062);
and (n11146,n3723,n3602);
and (n11147,n11148,n11149);
xor (n11148,n11145,n11146);
or (n11149,n11150,n11153);
and (n11150,n11151,n11152);
xor (n11151,n11067,n11068);
and (n11152,n3592,n3602);
and (n11153,n11154,n11155);
xor (n11154,n11151,n11152);
or (n11155,n11156,n11159);
and (n11156,n11157,n11158);
xor (n11157,n11072,n11073);
and (n11158,n3586,n3602);
and (n11159,n11160,n11161);
xor (n11160,n11157,n11158);
or (n11161,n11162,n11165);
and (n11162,n11163,n11164);
xor (n11163,n11078,n11079);
and (n11164,n3800,n3602);
and (n11165,n11166,n11167);
xor (n11166,n11163,n11164);
or (n11167,n11168,n11171);
and (n11168,n11169,n11170);
xor (n11169,n11083,n11084);
and (n11170,n3959,n3602);
and (n11171,n11172,n11173);
xor (n11172,n11169,n11170);
or (n11173,n11174,n11177);
and (n11174,n11175,n11176);
xor (n11175,n11089,n11090);
and (n11176,n3952,n3602);
and (n11177,n11178,n11179);
xor (n11178,n11175,n11176);
or (n11179,n11180,n11183);
and (n11180,n11181,n11182);
xor (n11181,n11094,n11095);
and (n11182,n4350,n3602);
and (n11183,n11184,n11185);
xor (n11184,n11181,n11182);
or (n11185,n11186,n11189);
and (n11186,n11187,n11188);
xor (n11187,n11100,n11101);
and (n11188,n4406,n3602);
and (n11189,n11190,n11191);
xor (n11190,n11187,n11188);
and (n11191,n11192,n6614);
xor (n11192,n11106,n11107);
and (n11193,n3843,n3611);
and (n11194,n11195,n11196);
xor (n11195,n10857,n11193);
or (n11196,n11197,n11199);
and (n11197,n11198,n3852);
xor (n11198,n11112,n11113);
and (n11199,n11200,n11201);
xor (n11200,n11198,n3852);
or (n11201,n11202,n11204);
and (n11202,n11203,n4010);
xor (n11203,n11118,n11119);
and (n11204,n11205,n11206);
xor (n11205,n11203,n4010);
or (n11206,n11207,n11210);
and (n11207,n11208,n11209);
xor (n11208,n11124,n11125);
and (n11209,n3622,n3611);
and (n11210,n11211,n11212);
xor (n11211,n11208,n11209);
or (n11212,n11213,n11216);
and (n11213,n11214,n11215);
xor (n11214,n11130,n11131);
and (n11215,n3695,n3611);
and (n11216,n11217,n11218);
xor (n11217,n11214,n11215);
or (n11218,n11219,n11222);
and (n11219,n11220,n11221);
xor (n11220,n11136,n11137);
and (n11221,n3680,n3611);
and (n11222,n11223,n11224);
xor (n11223,n11220,n11221);
or (n11224,n11225,n11228);
and (n11225,n11226,n11227);
xor (n11226,n11142,n11143);
and (n11227,n3723,n3611);
and (n11228,n11229,n11230);
xor (n11229,n11226,n11227);
or (n11230,n11231,n11234);
and (n11231,n11232,n11233);
xor (n11232,n11148,n11149);
and (n11233,n3592,n3611);
and (n11234,n11235,n11236);
xor (n11235,n11232,n11233);
or (n11236,n11237,n11240);
and (n11237,n11238,n11239);
xor (n11238,n11154,n11155);
and (n11239,n3586,n3611);
and (n11240,n11241,n11242);
xor (n11241,n11238,n11239);
or (n11242,n11243,n11246);
and (n11243,n11244,n11245);
xor (n11244,n11160,n11161);
and (n11245,n3800,n3611);
and (n11246,n11247,n11248);
xor (n11247,n11244,n11245);
or (n11248,n11249,n11252);
and (n11249,n11250,n11251);
xor (n11250,n11166,n11167);
and (n11251,n3959,n3611);
and (n11252,n11253,n11254);
xor (n11253,n11250,n11251);
or (n11254,n11255,n11258);
and (n11255,n11256,n11257);
xor (n11256,n11172,n11173);
and (n11257,n3952,n3611);
and (n11258,n11259,n11260);
xor (n11259,n11256,n11257);
or (n11260,n11261,n11264);
and (n11261,n11262,n11263);
xor (n11262,n11178,n11179);
and (n11263,n4350,n3611);
and (n11264,n11265,n11266);
xor (n11265,n11262,n11263);
or (n11266,n11267,n11269);
and (n11267,n11268,n6541);
xor (n11268,n11184,n11185);
and (n11269,n11270,n11271);
xor (n11270,n11268,n6541);
and (n11271,n11272,n6682);
xor (n11272,n11190,n11191);
and (n11273,n3843,n3828);
and (n11274,n11275,n11276);
xor (n11275,n10854,n11273);
or (n11276,n11277,n11280);
and (n11277,n11278,n11279);
xor (n11278,n11195,n11196);
and (n11279,n3837,n3828);
and (n11280,n11281,n11282);
xor (n11281,n11278,n11279);
or (n11282,n11283,n11286);
and (n11283,n11284,n11285);
xor (n11284,n11200,n11201);
and (n11285,n3641,n3828);
and (n11286,n11287,n11288);
xor (n11287,n11284,n11285);
or (n11288,n11289,n11292);
and (n11289,n11290,n11291);
xor (n11290,n11205,n11206);
and (n11291,n3622,n3828);
and (n11292,n11293,n11294);
xor (n11293,n11290,n11291);
or (n11294,n11295,n11298);
and (n11295,n11296,n11297);
xor (n11296,n11211,n11212);
and (n11297,n3695,n3828);
and (n11298,n11299,n11300);
xor (n11299,n11296,n11297);
or (n11300,n11301,n11304);
and (n11301,n11302,n11303);
xor (n11302,n11217,n11218);
and (n11303,n3680,n3828);
and (n11304,n11305,n11306);
xor (n11305,n11302,n11303);
or (n11306,n11307,n11310);
and (n11307,n11308,n11309);
xor (n11308,n11223,n11224);
and (n11309,n3723,n3828);
and (n11310,n11311,n11312);
xor (n11311,n11308,n11309);
or (n11312,n11313,n11316);
and (n11313,n11314,n11315);
xor (n11314,n11229,n11230);
and (n11315,n3592,n3828);
and (n11316,n11317,n11318);
xor (n11317,n11314,n11315);
or (n11318,n11319,n11322);
and (n11319,n11320,n11321);
xor (n11320,n11235,n11236);
and (n11321,n3586,n3828);
and (n11322,n11323,n11324);
xor (n11323,n11320,n11321);
or (n11324,n11325,n11328);
and (n11325,n11326,n11327);
xor (n11326,n11241,n11242);
and (n11327,n3800,n3828);
and (n11328,n11329,n11330);
xor (n11329,n11326,n11327);
or (n11330,n11331,n11334);
and (n11331,n11332,n11333);
xor (n11332,n11247,n11248);
and (n11333,n3959,n3828);
and (n11334,n11335,n11336);
xor (n11335,n11332,n11333);
or (n11336,n11337,n11340);
and (n11337,n11338,n11339);
xor (n11338,n11253,n11254);
and (n11339,n3952,n3828);
and (n11340,n11341,n11342);
xor (n11341,n11338,n11339);
or (n11342,n11343,n11346);
and (n11343,n11344,n11345);
xor (n11344,n11259,n11260);
and (n11345,n4350,n3828);
and (n11346,n11347,n11348);
xor (n11347,n11344,n11345);
or (n11348,n11349,n11352);
and (n11349,n11350,n11351);
xor (n11350,n11265,n11266);
and (n11351,n4406,n3828);
and (n11352,n11353,n11354);
xor (n11353,n11350,n11351);
and (n11354,n11355,n6432);
xor (n11355,n11270,n11271);
and (n11356,n3843,n3632);
and (n11357,n11358,n11359);
xor (n11358,n10851,n11356);
or (n11359,n11360,n11363);
and (n11360,n11361,n11362);
xor (n11361,n11275,n11276);
and (n11362,n3837,n3632);
and (n11363,n11364,n11365);
xor (n11364,n11361,n11362);
or (n11365,n11366,n11369);
and (n11366,n11367,n11368);
xor (n11367,n11281,n11282);
and (n11368,n3641,n3632);
and (n11369,n11370,n11371);
xor (n11370,n11367,n11368);
or (n11371,n11372,n11375);
and (n11372,n11373,n11374);
xor (n11373,n11287,n11288);
and (n11374,n3622,n3632);
and (n11375,n11376,n11377);
xor (n11376,n11373,n11374);
or (n11377,n11378,n11381);
and (n11378,n11379,n11380);
xor (n11379,n11293,n11294);
and (n11380,n3695,n3632);
and (n11381,n11382,n11383);
xor (n11382,n11379,n11380);
or (n11383,n11384,n11386);
and (n11384,n11385,n4399);
xor (n11385,n11299,n11300);
and (n11386,n11387,n11388);
xor (n11387,n11385,n4399);
or (n11388,n11389,n11392);
and (n11389,n11390,n11391);
xor (n11390,n11305,n11306);
and (n11391,n3723,n3632);
and (n11392,n11393,n11394);
xor (n11393,n11390,n11391);
or (n11394,n11395,n11398);
and (n11395,n11396,n11397);
xor (n11396,n11311,n11312);
and (n11397,n3592,n3632);
and (n11398,n11399,n11400);
xor (n11399,n11396,n11397);
or (n11400,n11401,n11404);
and (n11401,n11402,n11403);
xor (n11402,n11317,n11318);
and (n11403,n3586,n3632);
and (n11404,n11405,n11406);
xor (n11405,n11402,n11403);
or (n11406,n11407,n11410);
and (n11407,n11408,n11409);
xor (n11408,n11323,n11324);
and (n11409,n3800,n3632);
and (n11410,n11411,n11412);
xor (n11411,n11408,n11409);
or (n11412,n11413,n11416);
and (n11413,n11414,n11415);
xor (n11414,n11329,n11330);
and (n11415,n3959,n3632);
and (n11416,n11417,n11418);
xor (n11417,n11414,n11415);
or (n11418,n11419,n11422);
and (n11419,n11420,n11421);
xor (n11420,n11335,n11336);
and (n11421,n3952,n3632);
and (n11422,n11423,n11424);
xor (n11423,n11420,n11421);
or (n11424,n11425,n11428);
and (n11425,n11426,n11427);
xor (n11426,n11341,n11342);
and (n11427,n4350,n3632);
and (n11428,n11429,n11430);
xor (n11429,n11426,n11427);
or (n11430,n11431,n11434);
and (n11431,n11432,n11433);
xor (n11432,n11347,n11348);
and (n11433,n4406,n3632);
and (n11434,n11435,n11436);
xor (n11435,n11432,n11433);
and (n11436,n11437,n6446);
xor (n11437,n11353,n11354);
and (n11438,n3843,n3633);
and (n11439,n11440,n11441);
xor (n11440,n10848,n11438);
or (n11441,n11442,n11445);
and (n11442,n11443,n11444);
xor (n11443,n11358,n11359);
and (n11444,n3837,n3633);
and (n11445,n11446,n11447);
xor (n11446,n11443,n11444);
or (n11447,n11448,n11451);
and (n11448,n11449,n11450);
xor (n11449,n11364,n11365);
and (n11450,n3641,n3633);
and (n11451,n11452,n11453);
xor (n11452,n11449,n11450);
or (n11453,n11454,n11457);
and (n11454,n11455,n11456);
xor (n11455,n11370,n11371);
and (n11456,n3622,n3633);
and (n11457,n11458,n11459);
xor (n11458,n11455,n11456);
or (n11459,n11460,n11463);
and (n11460,n11461,n11462);
xor (n11461,n11376,n11377);
and (n11462,n3695,n3633);
and (n11463,n11464,n11465);
xor (n11464,n11461,n11462);
or (n11465,n11466,n11469);
and (n11466,n11467,n11468);
xor (n11467,n11382,n11383);
and (n11468,n3680,n3633);
and (n11469,n11470,n11471);
xor (n11470,n11467,n11468);
or (n11471,n11472,n11475);
and (n11472,n11473,n11474);
xor (n11473,n11387,n11388);
and (n11474,n3723,n3633);
and (n11475,n11476,n11477);
xor (n11476,n11473,n11474);
or (n11477,n11478,n11481);
and (n11478,n11479,n11480);
xor (n11479,n11393,n11394);
and (n11480,n3592,n3633);
and (n11481,n11482,n11483);
xor (n11482,n11479,n11480);
or (n11483,n11484,n11487);
and (n11484,n11485,n11486);
xor (n11485,n11399,n11400);
and (n11486,n3586,n3633);
and (n11487,n11488,n11489);
xor (n11488,n11485,n11486);
or (n11489,n11490,n11493);
and (n11490,n11491,n11492);
xor (n11491,n11405,n11406);
and (n11492,n3800,n3633);
and (n11493,n11494,n11495);
xor (n11494,n11491,n11492);
or (n11495,n11496,n11499);
and (n11496,n11497,n11498);
xor (n11497,n11411,n11412);
and (n11498,n3959,n3633);
and (n11499,n11500,n11501);
xor (n11500,n11497,n11498);
or (n11501,n11502,n11505);
and (n11502,n11503,n11504);
xor (n11503,n11417,n11418);
and (n11504,n3952,n3633);
and (n11505,n11506,n11507);
xor (n11506,n11503,n11504);
or (n11507,n11508,n11511);
and (n11508,n11509,n11510);
xor (n11509,n11423,n11424);
and (n11510,n4350,n3633);
and (n11511,n11512,n11513);
xor (n11512,n11509,n11510);
or (n11513,n11514,n11517);
and (n11514,n11515,n11516);
xor (n11515,n11429,n11430);
and (n11516,n4406,n3633);
and (n11517,n11518,n11519);
xor (n11518,n11515,n11516);
and (n11519,n11520,n6224);
xor (n11520,n11435,n11436);
and (n11521,n3843,n3624);
and (n11522,n11523,n11524);
xor (n11523,n10845,n11521);
or (n11524,n11525,n11528);
and (n11525,n11526,n11527);
xor (n11526,n11440,n11441);
and (n11527,n3837,n3624);
and (n11528,n11529,n11530);
xor (n11529,n11526,n11527);
or (n11530,n11531,n11533);
and (n11531,n11532,n3640);
xor (n11532,n11446,n11447);
and (n11533,n11534,n11535);
xor (n11534,n11532,n3640);
or (n11535,n11536,n11539);
and (n11536,n11537,n11538);
xor (n11537,n11452,n11453);
and (n11538,n3622,n3624);
and (n11539,n11540,n11541);
xor (n11540,n11537,n11538);
or (n11541,n11542,n11545);
and (n11542,n11543,n11544);
xor (n11543,n11458,n11459);
and (n11544,n3695,n3624);
and (n11545,n11546,n11547);
xor (n11546,n11543,n11544);
or (n11547,n11548,n11551);
and (n11548,n11549,n11550);
xor (n11549,n11464,n11465);
and (n11550,n3680,n3624);
and (n11551,n11552,n11553);
xor (n11552,n11549,n11550);
or (n11553,n11554,n11556);
and (n11554,n11555,n4000);
xor (n11555,n11470,n11471);
and (n11556,n11557,n11558);
xor (n11557,n11555,n4000);
or (n11558,n11559,n11562);
and (n11559,n11560,n11561);
xor (n11560,n11476,n11477);
and (n11561,n3592,n3624);
and (n11562,n11563,n11564);
xor (n11563,n11560,n11561);
or (n11564,n11565,n11568);
and (n11565,n11566,n11567);
xor (n11566,n11482,n11483);
and (n11567,n3586,n3624);
and (n11568,n11569,n11570);
xor (n11569,n11566,n11567);
or (n11570,n11571,n11573);
and (n11571,n11572,n5364);
xor (n11572,n11488,n11489);
and (n11573,n11574,n11575);
xor (n11574,n11572,n5364);
or (n11575,n11576,n11579);
and (n11576,n11577,n11578);
xor (n11577,n11494,n11495);
and (n11578,n3959,n3624);
and (n11579,n11580,n11581);
xor (n11580,n11577,n11578);
or (n11581,n11582,n11585);
and (n11582,n11583,n11584);
xor (n11583,n11500,n11501);
and (n11584,n3952,n3624);
and (n11585,n11586,n11587);
xor (n11586,n11583,n11584);
or (n11587,n11588,n11591);
and (n11588,n11589,n11590);
xor (n11589,n11506,n11507);
and (n11590,n4350,n3624);
and (n11591,n11592,n11593);
xor (n11592,n11589,n11590);
or (n11593,n11594,n11597);
and (n11594,n11595,n11596);
xor (n11595,n11512,n11513);
and (n11596,n4406,n3624);
and (n11597,n11598,n11599);
xor (n11598,n11595,n11596);
and (n11599,n11600,n11601);
xor (n11600,n11518,n11519);
and (n11601,n5233,n3624);
and (n11602,n3843,n3687);
and (n11603,n11604,n11605);
xor (n11604,n10842,n11602);
or (n11605,n11606,n11609);
and (n11606,n11607,n11608);
xor (n11607,n11523,n11524);
and (n11608,n3837,n3687);
and (n11609,n11610,n11611);
xor (n11610,n11607,n11608);
or (n11611,n11612,n11615);
and (n11612,n11613,n11614);
xor (n11613,n11529,n11530);
and (n11614,n3641,n3687);
and (n11615,n11616,n11617);
xor (n11616,n11613,n11614);
or (n11617,n11618,n11621);
and (n11618,n11619,n11620);
xor (n11619,n11534,n11535);
and (n11620,n3622,n3687);
and (n11621,n11622,n11623);
xor (n11622,n11619,n11620);
or (n11623,n11624,n11627);
and (n11624,n11625,n11626);
xor (n11625,n11540,n11541);
and (n11626,n3695,n3687);
and (n11627,n11628,n11629);
xor (n11628,n11625,n11626);
or (n11629,n11630,n11633);
and (n11630,n11631,n11632);
xor (n11631,n11546,n11547);
and (n11632,n3680,n3687);
and (n11633,n11634,n11635);
xor (n11634,n11631,n11632);
or (n11635,n11636,n11639);
and (n11636,n11637,n11638);
xor (n11637,n11552,n11553);
and (n11638,n3723,n3687);
and (n11639,n11640,n11641);
xor (n11640,n11637,n11638);
or (n11641,n11642,n11645);
and (n11642,n11643,n11644);
xor (n11643,n11557,n11558);
and (n11644,n3592,n3687);
and (n11645,n11646,n11647);
xor (n11646,n11643,n11644);
or (n11647,n11648,n11651);
and (n11648,n11649,n11650);
xor (n11649,n11563,n11564);
and (n11650,n3586,n3687);
and (n11651,n11652,n11653);
xor (n11652,n11649,n11650);
or (n11653,n11654,n11657);
and (n11654,n11655,n11656);
xor (n11655,n11569,n11570);
and (n11656,n3800,n3687);
and (n11657,n11658,n11659);
xor (n11658,n11655,n11656);
or (n11659,n11660,n11663);
and (n11660,n11661,n11662);
xor (n11661,n11574,n11575);
and (n11662,n3959,n3687);
and (n11663,n11664,n11665);
xor (n11664,n11661,n11662);
or (n11665,n11666,n11669);
and (n11666,n11667,n11668);
xor (n11667,n11580,n11581);
and (n11668,n3952,n3687);
and (n11669,n11670,n11671);
xor (n11670,n11667,n11668);
or (n11671,n11672,n11675);
and (n11672,n11673,n11674);
xor (n11673,n11586,n11587);
and (n11674,n4350,n3687);
and (n11675,n11676,n11677);
xor (n11676,n11673,n11674);
or (n11677,n11678,n11681);
and (n11678,n11679,n11680);
xor (n11679,n11592,n11593);
and (n11680,n4406,n3687);
and (n11681,n11682,n11683);
xor (n11682,n11679,n11680);
and (n11683,n11684,n5979);
xor (n11684,n11598,n11599);
and (n11685,n3843,n3573);
and (n11686,n11687,n11688);
xor (n11687,n10839,n11685);
or (n11688,n11689,n11691);
and (n11689,n11690,n4661);
xor (n11690,n11604,n11605);
and (n11691,n11692,n11693);
xor (n11692,n11690,n4661);
or (n11693,n11694,n11696);
and (n11694,n11695,n4593);
xor (n11695,n11610,n11611);
and (n11696,n11697,n11698);
xor (n11697,n11695,n4593);
or (n11698,n11699,n11701);
and (n11699,n11700,n4278);
xor (n11700,n11616,n11617);
and (n11701,n11702,n11703);
xor (n11702,n11700,n4278);
or (n11703,n11704,n11707);
and (n11704,n11705,n11706);
xor (n11705,n11622,n11623);
and (n11706,n3695,n3573);
and (n11707,n11708,n11709);
xor (n11708,n11705,n11706);
or (n11709,n11710,n11713);
and (n11710,n11711,n11712);
xor (n11711,n11628,n11629);
and (n11712,n3680,n3573);
and (n11713,n11714,n11715);
xor (n11714,n11711,n11712);
or (n11715,n11716,n11719);
and (n11716,n11717,n11718);
xor (n11717,n11634,n11635);
and (n11718,n3723,n3573);
and (n11719,n11720,n11721);
xor (n11720,n11717,n11718);
or (n11721,n11722,n11724);
and (n11722,n11723,n4059);
xor (n11723,n11640,n11641);
and (n11724,n11725,n11726);
xor (n11725,n11723,n4059);
or (n11726,n11727,n11730);
and (n11727,n11728,n11729);
xor (n11728,n11646,n11647);
and (n11729,n3586,n3573);
and (n11730,n11731,n11732);
xor (n11731,n11728,n11729);
or (n11732,n11733,n11736);
and (n11733,n11734,n11735);
xor (n11734,n11652,n11653);
and (n11735,n3800,n3573);
and (n11736,n11737,n11738);
xor (n11737,n11734,n11735);
or (n11738,n11739,n11741);
and (n11739,n11740,n5169);
xor (n11740,n11658,n11659);
and (n11741,n11742,n11743);
xor (n11742,n11740,n5169);
or (n11743,n11744,n11746);
and (n11744,n11745,n5401);
xor (n11745,n11664,n11665);
and (n11746,n11747,n11748);
xor (n11747,n11745,n5401);
or (n11748,n11749,n11751);
and (n11749,n11750,n5614);
xor (n11750,n11670,n11671);
and (n11751,n11752,n11753);
xor (n11752,n11750,n5614);
or (n11753,n11754,n11757);
and (n11754,n11755,n11756);
xor (n11755,n11676,n11677);
and (n11756,n4406,n3573);
and (n11757,n11758,n11759);
xor (n11758,n11755,n11756);
and (n11759,n11760,n5935);
xor (n11760,n11682,n11683);
and (n11761,n3843,n3575);
and (n11762,n11763,n11764);
xor (n11763,n10836,n11761);
or (n11764,n11765,n11768);
and (n11765,n11766,n11767);
xor (n11766,n11687,n11688);
and (n11767,n3837,n3575);
and (n11768,n11769,n11770);
xor (n11769,n11766,n11767);
or (n11770,n11771,n11774);
and (n11771,n11772,n11773);
xor (n11772,n11692,n11693);
and (n11773,n3641,n3575);
and (n11774,n11775,n11776);
xor (n11775,n11772,n11773);
or (n11776,n11777,n11780);
and (n11777,n11778,n11779);
xor (n11778,n11697,n11698);
and (n11779,n3622,n3575);
and (n11780,n11781,n11782);
xor (n11781,n11778,n11779);
or (n11782,n11783,n11786);
and (n11783,n11784,n11785);
xor (n11784,n11702,n11703);
and (n11785,n3695,n3575);
and (n11786,n11787,n11788);
xor (n11787,n11784,n11785);
or (n11788,n11789,n11792);
and (n11789,n11790,n11791);
xor (n11790,n11708,n11709);
and (n11791,n3680,n3575);
and (n11792,n11793,n11794);
xor (n11793,n11790,n11791);
or (n11794,n11795,n11798);
and (n11795,n11796,n11797);
xor (n11796,n11714,n11715);
and (n11797,n3723,n3575);
and (n11798,n11799,n11800);
xor (n11799,n11796,n11797);
or (n11800,n11801,n11804);
and (n11801,n11802,n11803);
xor (n11802,n11720,n11721);
and (n11803,n3592,n3575);
and (n11804,n11805,n11806);
xor (n11805,n11802,n11803);
or (n11806,n11807,n11810);
and (n11807,n11808,n11809);
xor (n11808,n11725,n11726);
and (n11809,n3586,n3575);
and (n11810,n11811,n11812);
xor (n11811,n11808,n11809);
or (n11812,n11813,n11816);
and (n11813,n11814,n11815);
xor (n11814,n11731,n11732);
and (n11815,n3800,n3575);
and (n11816,n11817,n11818);
xor (n11817,n11814,n11815);
or (n11818,n11819,n11822);
and (n11819,n11820,n11821);
xor (n11820,n11737,n11738);
and (n11821,n3959,n3575);
and (n11822,n11823,n11824);
xor (n11823,n11820,n11821);
or (n11824,n11825,n11828);
and (n11825,n11826,n11827);
xor (n11826,n11742,n11743);
and (n11827,n3952,n3575);
and (n11828,n11829,n11830);
xor (n11829,n11826,n11827);
or (n11830,n11831,n11834);
and (n11831,n11832,n11833);
xor (n11832,n11747,n11748);
and (n11833,n4350,n3575);
and (n11834,n11835,n11836);
xor (n11835,n11832,n11833);
or (n11836,n11837,n11840);
and (n11837,n11838,n11839);
xor (n11838,n11752,n11753);
and (n11839,n4406,n3575);
and (n11840,n11841,n11842);
xor (n11841,n11838,n11839);
and (n11842,n11843,n5528);
xor (n11843,n11758,n11759);
and (n11844,n3843,n3581);
and (n11845,n11846,n11847);
xor (n11846,n10833,n11844);
or (n11847,n11848,n11851);
and (n11848,n11849,n11850);
xor (n11849,n11763,n11764);
and (n11850,n3837,n3581);
and (n11851,n11852,n11853);
xor (n11852,n11849,n11850);
or (n11853,n11854,n11857);
and (n11854,n11855,n11856);
xor (n11855,n11769,n11770);
and (n11856,n3641,n3581);
and (n11857,n11858,n11859);
xor (n11858,n11855,n11856);
or (n11859,n11860,n11863);
and (n11860,n11861,n11862);
xor (n11861,n11775,n11776);
and (n11862,n3622,n3581);
and (n11863,n11864,n11865);
xor (n11864,n11861,n11862);
or (n11865,n11866,n11868);
and (n11866,n11867,n4542);
xor (n11867,n11781,n11782);
and (n11868,n11869,n11870);
xor (n11869,n11867,n4542);
or (n11870,n11871,n11874);
and (n11871,n11872,n11873);
xor (n11872,n11787,n11788);
and (n11873,n3680,n3581);
and (n11874,n11875,n11876);
xor (n11875,n11872,n11873);
or (n11876,n11877,n11880);
and (n11877,n11878,n11879);
xor (n11878,n11793,n11794);
and (n11879,n3723,n3581);
and (n11880,n11881,n11882);
xor (n11881,n11878,n11879);
or (n11882,n11883,n11886);
and (n11883,n11884,n11885);
xor (n11884,n11799,n11800);
and (n11885,n3592,n3581);
and (n11886,n11887,n11888);
xor (n11887,n11884,n11885);
or (n11888,n11889,n11892);
and (n11889,n11890,n11891);
xor (n11890,n11805,n11806);
and (n11891,n3586,n3581);
and (n11892,n11893,n11894);
xor (n11893,n11890,n11891);
or (n11894,n11895,n11898);
and (n11895,n11896,n11897);
xor (n11896,n11811,n11812);
and (n11897,n3800,n3581);
and (n11898,n11899,n11900);
xor (n11899,n11896,n11897);
or (n11900,n11901,n11904);
and (n11901,n11902,n11903);
xor (n11902,n11817,n11818);
and (n11903,n3959,n3581);
and (n11904,n11905,n11906);
xor (n11905,n11902,n11903);
or (n11906,n11907,n11909);
and (n11907,n11908,n4501);
xor (n11908,n11823,n11824);
and (n11909,n11910,n11911);
xor (n11910,n11908,n4501);
or (n11911,n11912,n11915);
and (n11912,n11913,n11914);
xor (n11913,n11829,n11830);
and (n11914,n4350,n3581);
and (n11915,n11916,n11917);
xor (n11916,n11913,n11914);
or (n11917,n11918,n11920);
and (n11918,n11919,n5483);
xor (n11919,n11835,n11836);
and (n11920,n11921,n11922);
xor (n11921,n11919,n5483);
and (n11922,n11923,n11924);
xor (n11923,n11841,n11842);
and (n11924,n5233,n3581);
and (n11925,n3843,n3783);
and (n11926,n11927,n11928);
xor (n11927,n10830,n11925);
or (n11928,n11929,n11932);
and (n11929,n11930,n11931);
xor (n11930,n11846,n11847);
and (n11931,n3837,n3783);
and (n11932,n11933,n11934);
xor (n11933,n11930,n11931);
or (n11934,n11935,n11938);
and (n11935,n11936,n11937);
xor (n11936,n11852,n11853);
and (n11937,n3641,n3783);
and (n11938,n11939,n11940);
xor (n11939,n11936,n11937);
or (n11940,n11941,n11944);
and (n11941,n11942,n11943);
xor (n11942,n11858,n11859);
and (n11943,n3622,n3783);
and (n11944,n11945,n11946);
xor (n11945,n11942,n11943);
or (n11946,n11947,n11950);
and (n11947,n11948,n11949);
xor (n11948,n11864,n11865);
and (n11949,n3695,n3783);
and (n11950,n11951,n11952);
xor (n11951,n11948,n11949);
or (n11952,n11953,n11956);
and (n11953,n11954,n11955);
xor (n11954,n11869,n11870);
and (n11955,n3680,n3783);
and (n11956,n11957,n11958);
xor (n11957,n11954,n11955);
or (n11958,n11959,n11962);
and (n11959,n11960,n11961);
xor (n11960,n11875,n11876);
and (n11961,n3723,n3783);
and (n11962,n11963,n11964);
xor (n11963,n11960,n11961);
or (n11964,n11965,n11968);
and (n11965,n11966,n11967);
xor (n11966,n11881,n11882);
and (n11967,n3592,n3783);
and (n11968,n11969,n11970);
xor (n11969,n11966,n11967);
or (n11970,n11971,n11974);
and (n11971,n11972,n11973);
xor (n11972,n11887,n11888);
and (n11973,n3586,n3783);
and (n11974,n11975,n11976);
xor (n11975,n11972,n11973);
or (n11976,n11977,n11980);
and (n11977,n11978,n11979);
xor (n11978,n11893,n11894);
and (n11979,n3800,n3783);
and (n11980,n11981,n11982);
xor (n11981,n11978,n11979);
or (n11982,n11983,n11986);
and (n11983,n11984,n11985);
xor (n11984,n11899,n11900);
and (n11985,n3959,n3783);
and (n11986,n11987,n11988);
xor (n11987,n11984,n11985);
or (n11988,n11989,n11992);
and (n11989,n11990,n11991);
xor (n11990,n11905,n11906);
and (n11991,n3952,n3783);
and (n11992,n11993,n11994);
xor (n11993,n11990,n11991);
or (n11994,n11995,n11998);
and (n11995,n11996,n11997);
xor (n11996,n11910,n11911);
and (n11997,n4350,n3783);
and (n11998,n11999,n12000);
xor (n11999,n11996,n11997);
or (n12000,n12001,n12004);
and (n12001,n12002,n12003);
xor (n12002,n11916,n11917);
and (n12003,n4406,n3783);
and (n12004,n12005,n12006);
xor (n12005,n12002,n12003);
and (n12006,n12007,n5232);
xor (n12007,n11921,n11922);
and (n12008,n3843,n3790);
and (n12009,n12010,n12011);
xor (n12010,n10827,n12008);
or (n12011,n12012,n12015);
and (n12012,n12013,n12014);
xor (n12013,n11927,n11928);
and (n12014,n3837,n3790);
and (n12015,n12016,n12017);
xor (n12016,n12013,n12014);
or (n12017,n12018,n12021);
and (n12018,n12019,n12020);
xor (n12019,n11933,n11934);
and (n12020,n3641,n3790);
and (n12021,n12022,n12023);
xor (n12022,n12019,n12020);
or (n12023,n12024,n12027);
and (n12024,n12025,n12026);
xor (n12025,n11939,n11940);
and (n12026,n3622,n3790);
and (n12027,n12028,n12029);
xor (n12028,n12025,n12026);
or (n12029,n12030,n12033);
and (n12030,n12031,n12032);
xor (n12031,n11945,n11946);
and (n12032,n3695,n3790);
and (n12033,n12034,n12035);
xor (n12034,n12031,n12032);
or (n12035,n12036,n12039);
and (n12036,n12037,n12038);
xor (n12037,n11951,n11952);
and (n12038,n3680,n3790);
and (n12039,n12040,n12041);
xor (n12040,n12037,n12038);
or (n12041,n12042,n12045);
and (n12042,n12043,n12044);
xor (n12043,n11957,n11958);
and (n12044,n3723,n3790);
and (n12045,n12046,n12047);
xor (n12046,n12043,n12044);
or (n12047,n12048,n12050);
and (n12048,n12049,n4259);
xor (n12049,n11963,n11964);
and (n12050,n12051,n12052);
xor (n12051,n12049,n4259);
or (n12052,n12053,n12055);
and (n12053,n12054,n3792);
xor (n12054,n11969,n11970);
and (n12055,n12056,n12057);
xor (n12056,n12054,n3792);
or (n12057,n12058,n12061);
and (n12058,n12059,n12060);
xor (n12059,n11975,n11976);
and (n12060,n3800,n3790);
and (n12061,n12062,n12063);
xor (n12062,n12059,n12060);
or (n12063,n12064,n12067);
and (n12064,n12065,n12066);
xor (n12065,n11981,n11982);
and (n12066,n3959,n3790);
and (n12067,n12068,n12069);
xor (n12068,n12065,n12066);
or (n12069,n12070,n12072);
and (n12070,n12071,n3953);
xor (n12071,n11987,n11988);
and (n12072,n12073,n12074);
xor (n12073,n12071,n3953);
or (n12074,n12075,n12078);
and (n12075,n12076,n12077);
xor (n12076,n11993,n11994);
and (n12077,n4350,n3790);
and (n12078,n12079,n12080);
xor (n12079,n12076,n12077);
or (n12080,n12081,n12084);
and (n12081,n12082,n12083);
xor (n12082,n11999,n12000);
and (n12083,n4406,n3790);
and (n12084,n12085,n12086);
xor (n12085,n12082,n12083);
and (n12086,n12087,n12088);
xor (n12087,n12005,n12006);
and (n12088,n5233,n3790);
and (n12089,n12090,n12091);
xor (n12090,n10824,n12008);
or (n12091,n12092,n12094);
and (n12092,n12093,n12014);
xor (n12093,n12010,n12011);
and (n12094,n12095,n12096);
xor (n12095,n12093,n12014);
or (n12096,n12097,n12099);
and (n12097,n12098,n12020);
xor (n12098,n12016,n12017);
and (n12099,n12100,n12101);
xor (n12100,n12098,n12020);
or (n12101,n12102,n12104);
and (n12102,n12103,n12026);
xor (n12103,n12022,n12023);
and (n12104,n12105,n12106);
xor (n12105,n12103,n12026);
or (n12106,n12107,n12109);
and (n12107,n12108,n12032);
xor (n12108,n12028,n12029);
and (n12109,n12110,n12111);
xor (n12110,n12108,n12032);
or (n12111,n12112,n12114);
and (n12112,n12113,n12038);
xor (n12113,n12034,n12035);
and (n12114,n12115,n12116);
xor (n12115,n12113,n12038);
or (n12116,n12117,n12119);
and (n12117,n12118,n12044);
xor (n12118,n12040,n12041);
and (n12119,n12120,n12121);
xor (n12120,n12118,n12044);
or (n12121,n12122,n12124);
and (n12122,n12123,n4259);
xor (n12123,n12046,n12047);
and (n12124,n12125,n12126);
xor (n12125,n12123,n4259);
or (n12126,n12127,n12129);
and (n12127,n12128,n3792);
xor (n12128,n12051,n12052);
and (n12129,n12130,n12131);
xor (n12130,n12128,n3792);
or (n12131,n12132,n12134);
and (n12132,n12133,n12060);
xor (n12133,n12056,n12057);
and (n12134,n12135,n12136);
xor (n12135,n12133,n12060);
or (n12136,n12137,n12139);
and (n12137,n12138,n12066);
xor (n12138,n12062,n12063);
and (n12139,n12140,n12141);
xor (n12140,n12138,n12066);
or (n12141,n12142,n12144);
and (n12142,n12143,n3953);
xor (n12143,n12068,n12069);
and (n12144,n12145,n12146);
xor (n12145,n12143,n3953);
or (n12146,n12147,n12149);
and (n12147,n12148,n12077);
xor (n12148,n12073,n12074);
and (n12149,n12150,n12151);
xor (n12150,n12148,n12077);
or (n12151,n12152,n12154);
and (n12152,n12153,n12083);
xor (n12153,n12079,n12080);
and (n12154,n12155,n12156);
xor (n12155,n12153,n12083);
and (n12156,n12157,n12088);
xor (n12157,n12085,n12086);
or (n12158,n12159,n12161);
and (n12159,n12160,n12014);
xor (n12160,n12090,n12091);
and (n12161,n12162,n12163);
xor (n12162,n12160,n12014);
or (n12163,n12164,n12166);
and (n12164,n12165,n12020);
xor (n12165,n12095,n12096);
and (n12166,n12167,n12168);
xor (n12167,n12165,n12020);
or (n12168,n12169,n12171);
and (n12169,n12170,n12026);
xor (n12170,n12100,n12101);
and (n12171,n12172,n12173);
xor (n12172,n12170,n12026);
or (n12173,n12174,n12176);
and (n12174,n12175,n12032);
xor (n12175,n12105,n12106);
and (n12176,n12177,n12178);
xor (n12177,n12175,n12032);
or (n12178,n12179,n12181);
and (n12179,n12180,n12038);
xor (n12180,n12110,n12111);
and (n12181,n12182,n12183);
xor (n12182,n12180,n12038);
or (n12183,n12184,n12186);
and (n12184,n12185,n12044);
xor (n12185,n12115,n12116);
and (n12186,n12187,n12188);
xor (n12187,n12185,n12044);
or (n12188,n12189,n12191);
and (n12189,n12190,n4259);
xor (n12190,n12120,n12121);
and (n12191,n12192,n12193);
xor (n12192,n12190,n4259);
or (n12193,n12194,n12196);
and (n12194,n12195,n3792);
xor (n12195,n12125,n12126);
and (n12196,n12197,n12198);
xor (n12197,n12195,n3792);
or (n12198,n12199,n12201);
and (n12199,n12200,n12060);
xor (n12200,n12130,n12131);
and (n12201,n12202,n12203);
xor (n12202,n12200,n12060);
or (n12203,n12204,n12206);
and (n12204,n12205,n12066);
xor (n12205,n12135,n12136);
and (n12206,n12207,n12208);
xor (n12207,n12205,n12066);
or (n12208,n12209,n12211);
and (n12209,n12210,n3953);
xor (n12210,n12140,n12141);
and (n12211,n12212,n12213);
xor (n12212,n12210,n3953);
or (n12213,n12214,n12216);
and (n12214,n12215,n12077);
xor (n12215,n12145,n12146);
and (n12216,n12217,n12218);
xor (n12217,n12215,n12077);
or (n12218,n12219,n12221);
and (n12219,n12220,n12083);
xor (n12220,n12150,n12151);
and (n12221,n12222,n12223);
xor (n12222,n12220,n12083);
and (n12223,n12224,n12088);
xor (n12224,n12155,n12156);
or (n12225,n12226,n12228);
and (n12226,n12227,n12020);
xor (n12227,n12162,n12163);
and (n12228,n12229,n12230);
xor (n12229,n12227,n12020);
or (n12230,n12231,n12233);
and (n12231,n12232,n12026);
xor (n12232,n12167,n12168);
and (n12233,n12234,n12235);
xor (n12234,n12232,n12026);
or (n12235,n12236,n12238);
and (n12236,n12237,n12032);
xor (n12237,n12172,n12173);
and (n12238,n12239,n12240);
xor (n12239,n12237,n12032);
or (n12240,n12241,n12243);
and (n12241,n12242,n12038);
xor (n12242,n12177,n12178);
and (n12243,n12244,n12245);
xor (n12244,n12242,n12038);
or (n12245,n12246,n12248);
and (n12246,n12247,n12044);
xor (n12247,n12182,n12183);
and (n12248,n12249,n12250);
xor (n12249,n12247,n12044);
or (n12250,n12251,n12253);
and (n12251,n12252,n4259);
xor (n12252,n12187,n12188);
and (n12253,n12254,n12255);
xor (n12254,n12252,n4259);
or (n12255,n12256,n12258);
and (n12256,n12257,n3792);
xor (n12257,n12192,n12193);
and (n12258,n12259,n12260);
xor (n12259,n12257,n3792);
or (n12260,n12261,n12263);
and (n12261,n12262,n12060);
xor (n12262,n12197,n12198);
and (n12263,n12264,n12265);
xor (n12264,n12262,n12060);
or (n12265,n12266,n12268);
and (n12266,n12267,n12066);
xor (n12267,n12202,n12203);
and (n12268,n12269,n12270);
xor (n12269,n12267,n12066);
or (n12270,n12271,n12273);
and (n12271,n12272,n3953);
xor (n12272,n12207,n12208);
and (n12273,n12274,n12275);
xor (n12274,n12272,n3953);
or (n12275,n12276,n12278);
and (n12276,n12277,n12077);
xor (n12277,n12212,n12213);
and (n12278,n12279,n12280);
xor (n12279,n12277,n12077);
or (n12280,n12281,n12283);
and (n12281,n12282,n12083);
xor (n12282,n12217,n12218);
and (n12283,n12284,n12285);
xor (n12284,n12282,n12083);
and (n12285,n12286,n12088);
xor (n12286,n12222,n12223);
or (n12287,n12288,n12290);
and (n12288,n12289,n12026);
xor (n12289,n12229,n12230);
and (n12290,n12291,n12292);
xor (n12291,n12289,n12026);
or (n12292,n12293,n12295);
and (n12293,n12294,n12032);
xor (n12294,n12234,n12235);
and (n12295,n12296,n12297);
xor (n12296,n12294,n12032);
or (n12297,n12298,n12300);
and (n12298,n12299,n12038);
xor (n12299,n12239,n12240);
and (n12300,n12301,n12302);
xor (n12301,n12299,n12038);
or (n12302,n12303,n12305);
and (n12303,n12304,n12044);
xor (n12304,n12244,n12245);
and (n12305,n12306,n12307);
xor (n12306,n12304,n12044);
or (n12307,n12308,n12310);
and (n12308,n12309,n4259);
xor (n12309,n12249,n12250);
and (n12310,n12311,n12312);
xor (n12311,n12309,n4259);
or (n12312,n12313,n12315);
and (n12313,n12314,n3792);
xor (n12314,n12254,n12255);
and (n12315,n12316,n12317);
xor (n12316,n12314,n3792);
or (n12317,n12318,n12320);
and (n12318,n12319,n12060);
xor (n12319,n12259,n12260);
and (n12320,n12321,n12322);
xor (n12321,n12319,n12060);
or (n12322,n12323,n12325);
and (n12323,n12324,n12066);
xor (n12324,n12264,n12265);
and (n12325,n12326,n12327);
xor (n12326,n12324,n12066);
or (n12327,n12328,n12330);
and (n12328,n12329,n3953);
xor (n12329,n12269,n12270);
and (n12330,n12331,n12332);
xor (n12331,n12329,n3953);
or (n12332,n12333,n12335);
and (n12333,n12334,n12077);
xor (n12334,n12274,n12275);
and (n12335,n12336,n12337);
xor (n12336,n12334,n12077);
or (n12337,n12338,n12340);
and (n12338,n12339,n12083);
xor (n12339,n12279,n12280);
and (n12340,n12341,n12342);
xor (n12341,n12339,n12083);
and (n12342,n12343,n12088);
xor (n12343,n12284,n12285);
or (n12344,n12345,n12347);
and (n12345,n12346,n12032);
xor (n12346,n12291,n12292);
and (n12347,n12348,n12349);
xor (n12348,n12346,n12032);
or (n12349,n12350,n12352);
and (n12350,n12351,n12038);
xor (n12351,n12296,n12297);
and (n12352,n12353,n12354);
xor (n12353,n12351,n12038);
or (n12354,n12355,n12357);
and (n12355,n12356,n12044);
xor (n12356,n12301,n12302);
and (n12357,n12358,n12359);
xor (n12358,n12356,n12044);
or (n12359,n12360,n12362);
and (n12360,n12361,n4259);
xor (n12361,n12306,n12307);
and (n12362,n12363,n12364);
xor (n12363,n12361,n4259);
or (n12364,n12365,n12367);
and (n12365,n12366,n3792);
xor (n12366,n12311,n12312);
and (n12367,n12368,n12369);
xor (n12368,n12366,n3792);
or (n12369,n12370,n12372);
and (n12370,n12371,n12060);
xor (n12371,n12316,n12317);
and (n12372,n12373,n12374);
xor (n12373,n12371,n12060);
or (n12374,n12375,n12377);
and (n12375,n12376,n12066);
xor (n12376,n12321,n12322);
and (n12377,n12378,n12379);
xor (n12378,n12376,n12066);
or (n12379,n12380,n12382);
and (n12380,n12381,n3953);
xor (n12381,n12326,n12327);
and (n12382,n12383,n12384);
xor (n12383,n12381,n3953);
or (n12384,n12385,n12387);
and (n12385,n12386,n12077);
xor (n12386,n12331,n12332);
and (n12387,n12388,n12389);
xor (n12388,n12386,n12077);
or (n12389,n12390,n12392);
and (n12390,n12391,n12083);
xor (n12391,n12336,n12337);
and (n12392,n12393,n12394);
xor (n12393,n12391,n12083);
and (n12394,n12395,n12088);
xor (n12395,n12341,n12342);
or (n12396,n12397,n12399);
and (n12397,n12398,n12038);
xor (n12398,n12348,n12349);
and (n12399,n12400,n12401);
xor (n12400,n12398,n12038);
or (n12401,n12402,n12404);
and (n12402,n12403,n12044);
xor (n12403,n12353,n12354);
and (n12404,n12405,n12406);
xor (n12405,n12403,n12044);
or (n12406,n12407,n12409);
and (n12407,n12408,n4259);
xor (n12408,n12358,n12359);
and (n12409,n12410,n12411);
xor (n12410,n12408,n4259);
or (n12411,n12412,n12414);
and (n12412,n12413,n3792);
xor (n12413,n12363,n12364);
and (n12414,n12415,n12416);
xor (n12415,n12413,n3792);
or (n12416,n12417,n12419);
and (n12417,n12418,n12060);
xor (n12418,n12368,n12369);
and (n12419,n12420,n12421);
xor (n12420,n12418,n12060);
or (n12421,n12422,n12424);
and (n12422,n12423,n12066);
xor (n12423,n12373,n12374);
and (n12424,n12425,n12426);
xor (n12425,n12423,n12066);
or (n12426,n12427,n12429);
and (n12427,n12428,n3953);
xor (n12428,n12378,n12379);
and (n12429,n12430,n12431);
xor (n12430,n12428,n3953);
or (n12431,n12432,n12434);
and (n12432,n12433,n12077);
xor (n12433,n12383,n12384);
and (n12434,n12435,n12436);
xor (n12435,n12433,n12077);
or (n12436,n12437,n12439);
and (n12437,n12438,n12083);
xor (n12438,n12388,n12389);
and (n12439,n12440,n12441);
xor (n12440,n12438,n12083);
and (n12441,n12442,n12088);
xor (n12442,n12393,n12394);
or (n12443,n12444,n12446);
and (n12444,n12445,n12044);
xor (n12445,n12400,n12401);
and (n12446,n12447,n12448);
xor (n12447,n12445,n12044);
or (n12448,n12449,n12451);
and (n12449,n12450,n4259);
xor (n12450,n12405,n12406);
and (n12451,n12452,n12453);
xor (n12452,n12450,n4259);
or (n12453,n12454,n12456);
and (n12454,n12455,n3792);
xor (n12455,n12410,n12411);
and (n12456,n12457,n12458);
xor (n12457,n12455,n3792);
or (n12458,n12459,n12461);
and (n12459,n12460,n12060);
xor (n12460,n12415,n12416);
and (n12461,n12462,n12463);
xor (n12462,n12460,n12060);
or (n12463,n12464,n12466);
and (n12464,n12465,n12066);
xor (n12465,n12420,n12421);
and (n12466,n12467,n12468);
xor (n12467,n12465,n12066);
or (n12468,n12469,n12471);
and (n12469,n12470,n3953);
xor (n12470,n12425,n12426);
and (n12471,n12472,n12473);
xor (n12472,n12470,n3953);
or (n12473,n12474,n12476);
and (n12474,n12475,n12077);
xor (n12475,n12430,n12431);
and (n12476,n12477,n12478);
xor (n12477,n12475,n12077);
or (n12478,n12479,n12481);
and (n12479,n12480,n12083);
xor (n12480,n12435,n12436);
and (n12481,n12482,n12483);
xor (n12482,n12480,n12083);
and (n12483,n12484,n12088);
xor (n12484,n12440,n12441);
or (n12485,n12486,n12488);
and (n12486,n12487,n4259);
xor (n12487,n12447,n12448);
and (n12488,n12489,n12490);
xor (n12489,n12487,n4259);
or (n12490,n12491,n12493);
and (n12491,n12492,n3792);
xor (n12492,n12452,n12453);
and (n12493,n12494,n12495);
xor (n12494,n12492,n3792);
or (n12495,n12496,n12498);
and (n12496,n12497,n12060);
xor (n12497,n12457,n12458);
and (n12498,n12499,n12500);
xor (n12499,n12497,n12060);
or (n12500,n12501,n12503);
and (n12501,n12502,n12066);
xor (n12502,n12462,n12463);
and (n12503,n12504,n12505);
xor (n12504,n12502,n12066);
or (n12505,n12506,n12508);
and (n12506,n12507,n3953);
xor (n12507,n12467,n12468);
and (n12508,n12509,n12510);
xor (n12509,n12507,n3953);
or (n12510,n12511,n12513);
and (n12511,n12512,n12077);
xor (n12512,n12472,n12473);
and (n12513,n12514,n12515);
xor (n12514,n12512,n12077);
or (n12515,n12516,n12518);
and (n12516,n12517,n12083);
xor (n12517,n12477,n12478);
and (n12518,n12519,n12520);
xor (n12519,n12517,n12083);
and (n12520,n12521,n12088);
xor (n12521,n12482,n12483);
or (n12522,n12523,n12525);
and (n12523,n12524,n3792);
xor (n12524,n12489,n12490);
and (n12525,n12526,n12527);
xor (n12526,n12524,n3792);
or (n12527,n12528,n12530);
and (n12528,n12529,n12060);
xor (n12529,n12494,n12495);
and (n12530,n12531,n12532);
xor (n12531,n12529,n12060);
or (n12532,n12533,n12535);
and (n12533,n12534,n12066);
xor (n12534,n12499,n12500);
and (n12535,n12536,n12537);
xor (n12536,n12534,n12066);
or (n12537,n12538,n12540);
and (n12538,n12539,n3953);
xor (n12539,n12504,n12505);
and (n12540,n12541,n12542);
xor (n12541,n12539,n3953);
or (n12542,n12543,n12545);
and (n12543,n12544,n12077);
xor (n12544,n12509,n12510);
and (n12545,n12546,n12547);
xor (n12546,n12544,n12077);
or (n12547,n12548,n12550);
and (n12548,n12549,n12083);
xor (n12549,n12514,n12515);
and (n12550,n12551,n12552);
xor (n12551,n12549,n12083);
and (n12552,n12553,n12088);
xor (n12553,n12519,n12520);
or (n12554,n12555,n12557);
and (n12555,n12556,n12060);
xor (n12556,n12526,n12527);
and (n12557,n12558,n12559);
xor (n12558,n12556,n12060);
or (n12559,n12560,n12562);
and (n12560,n12561,n12066);
xor (n12561,n12531,n12532);
and (n12562,n12563,n12564);
xor (n12563,n12561,n12066);
or (n12564,n12565,n12567);
and (n12565,n12566,n3953);
xor (n12566,n12536,n12537);
and (n12567,n12568,n12569);
xor (n12568,n12566,n3953);
or (n12569,n12570,n12572);
and (n12570,n12571,n12077);
xor (n12571,n12541,n12542);
and (n12572,n12573,n12574);
xor (n12573,n12571,n12077);
or (n12574,n12575,n12577);
and (n12575,n12576,n12083);
xor (n12576,n12546,n12547);
and (n12577,n12578,n12579);
xor (n12578,n12576,n12083);
and (n12579,n12580,n12088);
xor (n12580,n12551,n12552);
or (n12581,n12582,n12584);
and (n12582,n12583,n12066);
xor (n12583,n12558,n12559);
and (n12584,n12585,n12586);
xor (n12585,n12583,n12066);
or (n12586,n12587,n12589);
and (n12587,n12588,n3953);
xor (n12588,n12563,n12564);
and (n12589,n12590,n12591);
xor (n12590,n12588,n3953);
or (n12591,n12592,n12594);
and (n12592,n12593,n12077);
xor (n12593,n12568,n12569);
and (n12594,n12595,n12596);
xor (n12595,n12593,n12077);
or (n12596,n12597,n12599);
and (n12597,n12598,n12083);
xor (n12598,n12573,n12574);
and (n12599,n12600,n12601);
xor (n12600,n12598,n12083);
and (n12601,n12602,n12088);
xor (n12602,n12578,n12579);
or (n12603,n12604,n12606);
and (n12604,n12605,n3953);
xor (n12605,n12585,n12586);
and (n12606,n12607,n12608);
xor (n12607,n12605,n3953);
or (n12608,n12609,n12611);
and (n12609,n12610,n12077);
xor (n12610,n12590,n12591);
and (n12611,n12612,n12613);
xor (n12612,n12610,n12077);
or (n12613,n12614,n12616);
and (n12614,n12615,n12083);
xor (n12615,n12595,n12596);
and (n12616,n12617,n12618);
xor (n12617,n12615,n12083);
and (n12618,n12619,n12088);
xor (n12619,n12600,n12601);
or (n12620,n12621,n12623);
and (n12621,n12622,n12077);
xor (n12622,n12607,n12608);
and (n12623,n12624,n12625);
xor (n12624,n12622,n12077);
or (n12625,n12626,n12628);
and (n12626,n12627,n12083);
xor (n12627,n12612,n12613);
and (n12628,n12629,n12630);
xor (n12629,n12627,n12083);
and (n12630,n12631,n12088);
xor (n12631,n12617,n12618);
or (n12632,n12633,n12635);
and (n12633,n12634,n12083);
xor (n12634,n12624,n12625);
and (n12635,n12636,n12637);
xor (n12636,n12634,n12083);
and (n12637,n12638,n12088);
xor (n12638,n12629,n12630);
and (n12639,n12640,n12088);
xor (n12640,n12636,n12637);
not (n12641,n12642);
xor (n12642,n12643,n5270);
xor (n12643,n12644,n14508);
xor (n12644,n12645,n4412);
xor (n12645,n12646,n14501);
xor (n12646,n12647,n4343);
xor (n12647,n12648,n14489);
xor (n12648,n12649,n3934);
xor (n12649,n12650,n14472);
xor (n12650,n12651,n13938);
xor (n12651,n12652,n14450);
xor (n12652,n12653,n3669);
xor (n12653,n12654,n14423);
xor (n12654,n12655,n13927);
xor (n12655,n12656,n14391);
xor (n12656,n12657,n4269);
xor (n12657,n12658,n14354);
xor (n12658,n12659,n4572);
xor (n12659,n12660,n14312);
xor (n12660,n12661,n13911);
xor (n12661,n12662,n14265);
xor (n12662,n12663,n4756);
xor (n12663,n12664,n14213);
xor (n12664,n12665,n4834);
xor (n12665,n12666,n14156);
xor (n12666,n12667,n4894);
xor (n12667,n12668,n14094);
xor (n12668,n12669,n4966);
xor (n12669,n12670,n14027);
xor (n12670,n12671,n5016);
xor (n12671,n12672,n12729);
xor (n12672,n12673,n5050);
xor (n12673,n12674,n12728);
xor (n12674,n12675,n5050);
xor (n12675,n12676,n12727);
xor (n12676,n12677,n12726);
xor (n12677,n12678,n12725);
xor (n12678,n12679,n4977);
xor (n12679,n12680,n12724);
xor (n12680,n12681,n12723);
xor (n12681,n12682,n12722);
xor (n12682,n12683,n4855);
xor (n12683,n12684,n12721);
xor (n12684,n12685,n12720);
xor (n12685,n12686,n12719);
xor (n12686,n12687,n12718);
xor (n12687,n12688,n12717);
xor (n12688,n12689,n12716);
xor (n12689,n12690,n12715);
xor (n12690,n12691,n12714);
xor (n12691,n12692,n12713);
xor (n12692,n12693,n12712);
xor (n12693,n12694,n12711);
xor (n12694,n12695,n3819);
xor (n12695,n12696,n12710);
xor (n12696,n12697,n12709);
xor (n12697,n12698,n12708);
xor (n12698,n12699,n12707);
xor (n12699,n12700,n12706);
xor (n12700,n12701,n12705);
xor (n12701,n12702,n12704);
xor (n12702,n12703,n4430);
and (n12703,n3820,n4423);
and (n12704,n12703,n4430);
and (n12705,n3820,n4025);
and (n12706,n12701,n12705);
not (n12707,n4038);
and (n12708,n12699,n12707);
and (n12709,n3820,n3806);
and (n12710,n12697,n12709);
and (n12711,n12695,n3819);
and (n12712,n3820,n3529);
and (n12713,n12693,n12712);
not (n12714,n4285);
and (n12715,n12691,n12714);
and (n12716,n3820,n3554);
and (n12717,n12689,n12716);
and (n12718,n3820,n3546);
and (n12719,n12687,n12718);
and (n12720,n3820,n3741);
and (n12721,n12685,n12720);
and (n12722,n12683,n4855);
and (n12723,n3820,n3756);
and (n12724,n12681,n12723);
and (n12725,n12679,n4977);
and (n12726,n3820,n3657);
and (n12727,n12677,n12726);
and (n12728,n12675,n5050);
or (n12729,n12730,n13958);
and (n12730,n12731,n5016);
xor (n12731,n12674,n12732);
or (n12732,n12733,n13886);
and (n12733,n12734,n5016);
xor (n12734,n12676,n12735);
or (n12735,n12736,n13803);
and (n12736,n12737,n13802);
xor (n12737,n12678,n12738);
or (n12738,n12739,n13729);
and (n12739,n12740,n4930);
xor (n12740,n12680,n12741);
or (n12741,n12742,n13646);
and (n12742,n12743,n13645);
xor (n12743,n12682,n12744);
or (n12744,n12745,n13571);
and (n12745,n12746,n4780);
xor (n12746,n12684,n12747);
or (n12747,n12748,n13488);
and (n12748,n12749,n13487);
xor (n12749,n12686,n12750);
or (n12750,n12751,n13414);
and (n12751,n12752,n4603);
xor (n12752,n12688,n12753);
or (n12753,n12754,n13331);
and (n12754,n12755,n13330);
xor (n12755,n12690,n12756);
or (n12756,n12757,n13255);
and (n12757,n12758,n13254);
xor (n12758,n12692,n12759);
or (n12759,n12760,n13171);
and (n12760,n12761,n13170);
xor (n12761,n12694,n12762);
or (n12762,n12763,n13093);
and (n12763,n12764,n4141);
xor (n12764,n12696,n12765);
or (n12765,n12766,n13010);
and (n12766,n12767,n13009);
xor (n12767,n12698,n12768);
or (n12768,n12769,n12934);
and (n12769,n12770,n12933);
xor (n12770,n12700,n12771);
or (n12771,n12772,n12850);
and (n12772,n12773,n12849);
xor (n12773,n12702,n12774);
or (n12774,n12775,n12776);
and (n12775,n12703,n5143);
and (n12776,n12777,n12778);
xor (n12777,n12703,n5143);
or (n12778,n12779,n12781);
and (n12779,n12780,n5357);
and (n12780,n3704,n4423);
and (n12781,n12782,n12783);
xor (n12782,n12780,n5357);
or (n12783,n12784,n12786);
and (n12784,n12785,n5570);
and (n12785,n3537,n4423);
and (n12786,n12787,n12788);
xor (n12787,n12785,n5570);
or (n12788,n12789,n12791);
and (n12789,n12790,n5709);
and (n12790,n3518,n4423);
and (n12791,n12792,n12793);
xor (n12792,n12790,n5709);
or (n12793,n12794,n12796);
and (n12794,n12795,n5884);
and (n12795,n3566,n4423);
and (n12796,n12797,n12798);
xor (n12797,n12795,n5884);
or (n12798,n12799,n12801);
and (n12799,n12800,n6163);
and (n12800,n3545,n4423);
and (n12801,n12802,n12803);
xor (n12802,n12800,n6163);
or (n12803,n12804,n12807);
and (n12804,n12805,n12806);
and (n12805,n3732,n4423);
and (n12806,n3763,n4032);
and (n12807,n12808,n12809);
xor (n12808,n12805,n12806);
or (n12809,n12810,n12812);
and (n12810,n12811,n6336);
and (n12811,n3763,n4423);
and (n12812,n12813,n12814);
xor (n12813,n12811,n6336);
or (n12814,n12815,n12817);
and (n12815,n12816,n6490);
and (n12816,n3774,n4423);
and (n12817,n12818,n12819);
xor (n12818,n12816,n6490);
or (n12819,n12820,n12823);
and (n12820,n12821,n12822);
and (n12821,n3651,n4423);
and (n12822,n3670,n4032);
and (n12823,n12824,n12825);
xor (n12824,n12821,n12822);
or (n12825,n12826,n12828);
and (n12826,n12827,n6602);
and (n12827,n3670,n4423);
and (n12828,n12829,n12830);
xor (n12829,n12827,n6602);
or (n12830,n12831,n12833);
and (n12831,n12832,n6662);
and (n12832,n3929,n4423);
and (n12833,n12834,n12835);
xor (n12834,n12832,n6662);
or (n12835,n12836,n12838);
and (n12836,n12837,n6764);
and (n12837,n3935,n4423);
and (n12838,n12839,n12840);
xor (n12839,n12837,n6764);
or (n12840,n12841,n12844);
and (n12841,n12842,n12843);
and (n12842,n4342,n4423);
and (n12843,n4413,n4032);
and (n12844,n12845,n12846);
xor (n12845,n12842,n12843);
and (n12846,n12847,n12848);
and (n12847,n4413,n4423);
and (n12848,n5241,n4032);
and (n12849,n3704,n4025);
and (n12850,n12851,n12852);
xor (n12851,n12773,n12849);
or (n12852,n12853,n12856);
and (n12853,n12854,n12855);
xor (n12854,n12777,n12778);
and (n12855,n3537,n4025);
and (n12856,n12857,n12858);
xor (n12857,n12854,n12855);
or (n12858,n12859,n12862);
and (n12859,n12860,n12861);
xor (n12860,n12782,n12783);
and (n12861,n3518,n4025);
and (n12862,n12863,n12864);
xor (n12863,n12860,n12861);
or (n12864,n12865,n12868);
and (n12865,n12866,n12867);
xor (n12866,n12787,n12788);
and (n12867,n3566,n4025);
and (n12868,n12869,n12870);
xor (n12869,n12866,n12867);
or (n12870,n12871,n12874);
and (n12871,n12872,n12873);
xor (n12872,n12792,n12793);
and (n12873,n3545,n4025);
and (n12874,n12875,n12876);
xor (n12875,n12872,n12873);
or (n12876,n12877,n12880);
and (n12877,n12878,n12879);
xor (n12878,n12797,n12798);
and (n12879,n3732,n4025);
and (n12880,n12881,n12882);
xor (n12881,n12878,n12879);
or (n12882,n12883,n12886);
and (n12883,n12884,n12885);
xor (n12884,n12802,n12803);
and (n12885,n3763,n4025);
and (n12886,n12887,n12888);
xor (n12887,n12884,n12885);
or (n12888,n12889,n12892);
and (n12889,n12890,n12891);
xor (n12890,n12808,n12809);
and (n12891,n3774,n4025);
and (n12892,n12893,n12894);
xor (n12893,n12890,n12891);
or (n12894,n12895,n12898);
and (n12895,n12896,n12897);
xor (n12896,n12813,n12814);
and (n12897,n3651,n4025);
and (n12898,n12899,n12900);
xor (n12899,n12896,n12897);
or (n12900,n12901,n12904);
and (n12901,n12902,n12903);
xor (n12902,n12818,n12819);
and (n12903,n3670,n4025);
and (n12904,n12905,n12906);
xor (n12905,n12902,n12903);
or (n12906,n12907,n12910);
and (n12907,n12908,n12909);
xor (n12908,n12824,n12825);
and (n12909,n3929,n4025);
and (n12910,n12911,n12912);
xor (n12911,n12908,n12909);
or (n12912,n12913,n12916);
and (n12913,n12914,n12915);
xor (n12914,n12829,n12830);
and (n12915,n3935,n4025);
and (n12916,n12917,n12918);
xor (n12917,n12914,n12915);
or (n12918,n12919,n12922);
and (n12919,n12920,n12921);
xor (n12920,n12834,n12835);
and (n12921,n4342,n4025);
and (n12922,n12923,n12924);
xor (n12923,n12920,n12921);
or (n12924,n12925,n12928);
and (n12925,n12926,n12927);
xor (n12926,n12839,n12840);
and (n12927,n4413,n4025);
and (n12928,n12929,n12930);
xor (n12929,n12926,n12927);
and (n12930,n12931,n12932);
xor (n12931,n12845,n12846);
and (n12932,n5241,n4025);
and (n12933,n3704,n3808);
and (n12934,n12935,n12936);
xor (n12935,n12770,n12933);
or (n12936,n12937,n12940);
and (n12937,n12938,n12939);
xor (n12938,n12851,n12852);
and (n12939,n3537,n3808);
and (n12940,n12941,n12942);
xor (n12941,n12938,n12939);
or (n12942,n12943,n12945);
and (n12943,n12944,n5152);
xor (n12944,n12857,n12858);
and (n12945,n12946,n12947);
xor (n12946,n12944,n5152);
or (n12947,n12948,n12951);
and (n12948,n12949,n12950);
xor (n12949,n12863,n12864);
and (n12950,n3566,n3808);
and (n12951,n12952,n12953);
xor (n12952,n12949,n12950);
or (n12953,n12954,n12956);
and (n12954,n12955,n5586);
xor (n12955,n12869,n12870);
and (n12956,n12957,n12958);
xor (n12957,n12955,n5586);
or (n12958,n12959,n12961);
and (n12959,n12960,n5720);
xor (n12960,n12875,n12876);
and (n12961,n12962,n12963);
xor (n12962,n12960,n5720);
or (n12963,n12964,n12966);
and (n12964,n12965,n5893);
xor (n12965,n12881,n12882);
and (n12966,n12967,n12968);
xor (n12967,n12965,n5893);
or (n12968,n12969,n12971);
and (n12969,n12970,n6071);
xor (n12970,n12887,n12888);
and (n12971,n12972,n12973);
xor (n12972,n12970,n6071);
or (n12973,n12974,n12977);
and (n12974,n12975,n12976);
xor (n12975,n12893,n12894);
and (n12976,n3651,n3808);
and (n12977,n12978,n12979);
xor (n12978,n12975,n12976);
or (n12979,n12980,n12983);
and (n12980,n12981,n12982);
xor (n12981,n12899,n12900);
and (n12982,n3670,n3808);
and (n12983,n12984,n12985);
xor (n12984,n12981,n12982);
or (n12985,n12986,n12989);
and (n12986,n12987,n12988);
xor (n12987,n12905,n12906);
and (n12988,n3929,n3808);
and (n12989,n12990,n12991);
xor (n12990,n12987,n12988);
or (n12991,n12992,n12994);
and (n12992,n12993,n6549);
xor (n12993,n12911,n12912);
and (n12994,n12995,n12996);
xor (n12995,n12993,n6549);
or (n12996,n12997,n13000);
and (n12997,n12998,n12999);
xor (n12998,n12917,n12918);
and (n12999,n4342,n3808);
and (n13000,n13001,n13002);
xor (n13001,n12998,n12999);
or (n13002,n13003,n13005);
and (n13003,n13004,n6714);
xor (n13004,n12923,n12924);
and (n13005,n13006,n13007);
xor (n13006,n13004,n6714);
and (n13007,n13008,n6771);
xor (n13008,n12929,n12930);
and (n13009,n3704,n3806);
and (n13010,n13011,n13012);
xor (n13011,n12767,n13009);
or (n13012,n13013,n13016);
and (n13013,n13014,n13015);
xor (n13014,n12935,n12936);
and (n13015,n3537,n3806);
and (n13016,n13017,n13018);
xor (n13017,n13014,n13015);
or (n13018,n13019,n13022);
and (n13019,n13020,n13021);
xor (n13020,n12941,n12942);
and (n13021,n3518,n3806);
and (n13022,n13023,n13024);
xor (n13023,n13020,n13021);
or (n13024,n13025,n13028);
and (n13025,n13026,n13027);
xor (n13026,n12946,n12947);
and (n13027,n3566,n3806);
and (n13028,n13029,n13030);
xor (n13029,n13026,n13027);
or (n13030,n13031,n13034);
and (n13031,n13032,n13033);
xor (n13032,n12952,n12953);
and (n13033,n3545,n3806);
and (n13034,n13035,n13036);
xor (n13035,n13032,n13033);
or (n13036,n13037,n13040);
and (n13037,n13038,n13039);
xor (n13038,n12957,n12958);
and (n13039,n3732,n3806);
and (n13040,n13041,n13042);
xor (n13041,n13038,n13039);
or (n13042,n13043,n13046);
and (n13043,n13044,n13045);
xor (n13044,n12962,n12963);
and (n13045,n3763,n3806);
and (n13046,n13047,n13048);
xor (n13047,n13044,n13045);
or (n13048,n13049,n13052);
and (n13049,n13050,n13051);
xor (n13050,n12967,n12968);
and (n13051,n3774,n3806);
and (n13052,n13053,n13054);
xor (n13053,n13050,n13051);
or (n13054,n13055,n13058);
and (n13055,n13056,n13057);
xor (n13056,n12972,n12973);
and (n13057,n3651,n3806);
and (n13058,n13059,n13060);
xor (n13059,n13056,n13057);
or (n13060,n13061,n13064);
and (n13061,n13062,n13063);
xor (n13062,n12978,n12979);
and (n13063,n3670,n3806);
and (n13064,n13065,n13066);
xor (n13065,n13062,n13063);
or (n13066,n13067,n13070);
and (n13067,n13068,n13069);
xor (n13068,n12984,n12985);
and (n13069,n3929,n3806);
and (n13070,n13071,n13072);
xor (n13071,n13068,n13069);
or (n13072,n13073,n13076);
and (n13073,n13074,n13075);
xor (n13074,n12990,n12991);
and (n13075,n3935,n3806);
and (n13076,n13077,n13078);
xor (n13077,n13074,n13075);
or (n13078,n13079,n13082);
and (n13079,n13080,n13081);
xor (n13080,n12995,n12996);
and (n13081,n4342,n3806);
and (n13082,n13083,n13084);
xor (n13083,n13080,n13081);
or (n13084,n13085,n13088);
and (n13085,n13086,n13087);
xor (n13086,n13001,n13002);
and (n13087,n4413,n3806);
and (n13088,n13089,n13090);
xor (n13089,n13086,n13087);
and (n13090,n13091,n13092);
xor (n13091,n13006,n13007);
and (n13092,n5241,n3806);
and (n13093,n13094,n13095);
xor (n13094,n12764,n4141);
or (n13095,n13096,n13099);
and (n13096,n13097,n13098);
xor (n13097,n13011,n13012);
not (n13098,n4048);
and (n13099,n13100,n13101);
xor (n13100,n13097,n13098);
or (n13101,n13102,n13105);
and (n13102,n13103,n13104);
xor (n13103,n13017,n13018);
not (n13104,n4044);
and (n13105,n13106,n13107);
xor (n13106,n13103,n13104);
or (n13107,n13108,n13110);
and (n13108,n13109,n4459);
xor (n13109,n13023,n13024);
and (n13110,n13111,n13112);
xor (n13111,n13109,n4459);
or (n13112,n13113,n13115);
and (n13113,n13114,n5176);
xor (n13114,n13029,n13030);
and (n13115,n13116,n13117);
xor (n13116,n13114,n5176);
or (n13117,n13118,n13121);
and (n13118,n13119,n13120);
xor (n13119,n13035,n13036);
and (n13120,n3732,n3528);
and (n13121,n13122,n13123);
xor (n13122,n13119,n13120);
or (n13123,n13124,n13126);
and (n13124,n13125,n5599);
xor (n13125,n13041,n13042);
and (n13126,n13127,n13128);
xor (n13127,n13125,n5599);
or (n13128,n13129,n13131);
and (n13129,n13130,n5735);
xor (n13130,n13047,n13048);
and (n13131,n13132,n13133);
xor (n13132,n13130,n5735);
or (n13133,n13134,n13136);
and (n13134,n13135,n5911);
xor (n13135,n13053,n13054);
and (n13136,n13137,n13138);
xor (n13137,n13135,n5911);
or (n13138,n13139,n13142);
and (n13139,n13140,n13141);
xor (n13140,n13059,n13060);
and (n13141,n3670,n3528);
and (n13142,n13143,n13144);
xor (n13143,n13140,n13141);
or (n13144,n13145,n13148);
and (n13145,n13146,n13147);
xor (n13146,n13065,n13066);
and (n13147,n3929,n3528);
and (n13148,n13149,n13150);
xor (n13149,n13146,n13147);
or (n13150,n13151,n13154);
and (n13151,n13152,n13153);
xor (n13152,n13071,n13072);
and (n13153,n3935,n3528);
and (n13154,n13155,n13156);
xor (n13155,n13152,n13153);
or (n13156,n13157,n13160);
and (n13157,n13158,n13159);
xor (n13158,n13077,n13078);
and (n13159,n4342,n3528);
and (n13160,n13161,n13162);
xor (n13161,n13158,n13159);
or (n13162,n13163,n13166);
and (n13163,n13164,n13165);
xor (n13164,n13083,n13084);
and (n13165,n4413,n3528);
and (n13166,n13167,n13168);
xor (n13167,n13164,n13165);
and (n13168,n13169,n6697);
xor (n13169,n13089,n13090);
and (n13170,n3704,n3529);
and (n13171,n13172,n13173);
xor (n13172,n12761,n13170);
or (n13173,n13174,n13177);
and (n13174,n13175,n13176);
xor (n13175,n13094,n13095);
and (n13176,n3537,n3529);
and (n13177,n13178,n13179);
xor (n13178,n13175,n13176);
or (n13179,n13180,n13183);
and (n13180,n13181,n13182);
xor (n13181,n13100,n13101);
and (n13182,n3518,n3529);
and (n13183,n13184,n13185);
xor (n13184,n13181,n13182);
or (n13185,n13186,n13189);
and (n13186,n13187,n13188);
xor (n13187,n13106,n13107);
and (n13188,n3566,n3529);
and (n13189,n13190,n13191);
xor (n13190,n13187,n13188);
or (n13191,n13192,n13195);
and (n13192,n13193,n13194);
xor (n13193,n13111,n13112);
and (n13194,n3545,n3529);
and (n13195,n13196,n13197);
xor (n13196,n13193,n13194);
or (n13197,n13198,n13201);
and (n13198,n13199,n13200);
xor (n13199,n13116,n13117);
and (n13200,n3732,n3529);
and (n13201,n13202,n13203);
xor (n13202,n13199,n13200);
or (n13203,n13204,n13207);
and (n13204,n13205,n13206);
xor (n13205,n13122,n13123);
and (n13206,n3763,n3529);
and (n13207,n13208,n13209);
xor (n13208,n13205,n13206);
or (n13209,n13210,n13213);
and (n13210,n13211,n13212);
xor (n13211,n13127,n13128);
and (n13212,n3774,n3529);
and (n13213,n13214,n13215);
xor (n13214,n13211,n13212);
or (n13215,n13216,n13219);
and (n13216,n13217,n13218);
xor (n13217,n13132,n13133);
and (n13218,n3651,n3529);
and (n13219,n13220,n13221);
xor (n13220,n13217,n13218);
or (n13221,n13222,n13225);
and (n13222,n13223,n13224);
xor (n13223,n13137,n13138);
and (n13224,n3670,n3529);
and (n13225,n13226,n13227);
xor (n13226,n13223,n13224);
or (n13227,n13228,n13231);
and (n13228,n13229,n13230);
xor (n13229,n13143,n13144);
and (n13230,n3929,n3529);
and (n13231,n13232,n13233);
xor (n13232,n13229,n13230);
or (n13233,n13234,n13237);
and (n13234,n13235,n13236);
xor (n13235,n13149,n13150);
and (n13236,n3935,n3529);
and (n13237,n13238,n13239);
xor (n13238,n13235,n13236);
or (n13239,n13240,n13243);
and (n13240,n13241,n13242);
xor (n13241,n13155,n13156);
and (n13242,n4342,n3529);
and (n13243,n13244,n13245);
xor (n13244,n13241,n13242);
or (n13245,n13246,n13249);
and (n13246,n13247,n13248);
xor (n13247,n13161,n13162);
and (n13248,n4413,n3529);
and (n13249,n13250,n13251);
xor (n13250,n13247,n13248);
and (n13251,n13252,n13253);
xor (n13252,n13167,n13168);
and (n13253,n5241,n3529);
and (n13254,n3704,n3519);
and (n13255,n13256,n13257);
xor (n13256,n12758,n13254);
or (n13257,n13258,n13261);
and (n13258,n13259,n13260);
xor (n13259,n13172,n13173);
not (n13260,n3538);
and (n13261,n13262,n13263);
xor (n13262,n13259,n13260);
or (n13263,n13264,n13266);
and (n13264,n13265,n3517);
xor (n13265,n13178,n13179);
and (n13266,n13267,n13268);
xor (n13267,n13265,n3517);
or (n13268,n13269,n13271);
and (n13269,n13270,n4073);
xor (n13270,n13184,n13185);
and (n13271,n13272,n13273);
xor (n13272,n13270,n4073);
or (n13273,n13274,n13277);
and (n13274,n13275,n13276);
xor (n13275,n13190,n13191);
not (n13276,n4069);
and (n13277,n13278,n13279);
xor (n13278,n13275,n13276);
or (n13279,n13280,n13283);
and (n13280,n13281,n13282);
xor (n13281,n13196,n13197);
and (n13282,n3732,n3519);
and (n13283,n13284,n13285);
xor (n13284,n13281,n13282);
or (n13285,n13286,n13289);
and (n13286,n13287,n13288);
xor (n13287,n13202,n13203);
and (n13288,n3763,n3519);
and (n13289,n13290,n13291);
xor (n13290,n13287,n13288);
or (n13291,n13292,n13294);
and (n13292,n13293,n5408);
xor (n13293,n13208,n13209);
and (n13294,n13295,n13296);
xor (n13295,n13293,n5408);
or (n13296,n13297,n13299);
and (n13297,n13298,n5625);
xor (n13298,n13214,n13215);
and (n13299,n13300,n13301);
xor (n13300,n13298,n5625);
or (n13301,n13302,n13305);
and (n13302,n13303,n13304);
xor (n13303,n13220,n13221);
and (n13304,n3670,n3519);
and (n13305,n13306,n13307);
xor (n13306,n13303,n13304);
or (n13307,n13308,n13310);
and (n13308,n13309,n5919);
xor (n13309,n13226,n13227);
and (n13310,n13311,n13312);
xor (n13311,n13309,n5919);
or (n13312,n13313,n13315);
and (n13313,n13314,n6100);
xor (n13314,n13232,n13233);
and (n13315,n13316,n13317);
xor (n13316,n13314,n6100);
or (n13317,n13318,n13320);
and (n13318,n13319,n6208);
xor (n13319,n13238,n13239);
and (n13320,n13321,n13322);
xor (n13321,n13319,n6208);
or (n13322,n13323,n13326);
and (n13323,n13324,n13325);
xor (n13324,n13244,n13245);
and (n13325,n4413,n3519);
and (n13326,n13327,n13328);
xor (n13327,n13324,n13325);
and (n13328,n13329,n6465);
xor (n13329,n13250,n13251);
and (n13330,n3704,n3554);
and (n13331,n13332,n13333);
xor (n13332,n12755,n13330);
or (n13333,n13334,n13337);
and (n13334,n13335,n13336);
xor (n13335,n13256,n13257);
and (n13336,n3537,n3554);
and (n13337,n13338,n13339);
xor (n13338,n13335,n13336);
or (n13339,n13340,n13343);
and (n13340,n13341,n13342);
xor (n13341,n13262,n13263);
and (n13342,n3518,n3554);
and (n13343,n13344,n13345);
xor (n13344,n13341,n13342);
or (n13345,n13346,n13349);
and (n13346,n13347,n13348);
xor (n13347,n13267,n13268);
and (n13348,n3566,n3554);
and (n13349,n13350,n13351);
xor (n13350,n13347,n13348);
or (n13351,n13352,n13355);
and (n13352,n13353,n13354);
xor (n13353,n13272,n13273);
and (n13354,n3545,n3554);
and (n13355,n13356,n13357);
xor (n13356,n13353,n13354);
or (n13357,n13358,n13361);
and (n13358,n13359,n13360);
xor (n13359,n13278,n13279);
and (n13360,n3732,n3554);
and (n13361,n13362,n13363);
xor (n13362,n13359,n13360);
or (n13363,n13364,n13367);
and (n13364,n13365,n13366);
xor (n13365,n13284,n13285);
and (n13366,n3763,n3554);
and (n13367,n13368,n13369);
xor (n13368,n13365,n13366);
or (n13369,n13370,n13373);
and (n13370,n13371,n13372);
xor (n13371,n13290,n13291);
and (n13372,n3774,n3554);
and (n13373,n13374,n13375);
xor (n13374,n13371,n13372);
or (n13375,n13376,n13379);
and (n13376,n13377,n13378);
xor (n13377,n13295,n13296);
and (n13378,n3651,n3554);
and (n13379,n13380,n13381);
xor (n13380,n13377,n13378);
or (n13381,n13382,n13385);
and (n13382,n13383,n13384);
xor (n13383,n13300,n13301);
and (n13384,n3670,n3554);
and (n13385,n13386,n13387);
xor (n13386,n13383,n13384);
or (n13387,n13388,n13391);
and (n13388,n13389,n13390);
xor (n13389,n13306,n13307);
and (n13390,n3929,n3554);
and (n13391,n13392,n13393);
xor (n13392,n13389,n13390);
or (n13393,n13394,n13397);
and (n13394,n13395,n13396);
xor (n13395,n13311,n13312);
and (n13396,n3935,n3554);
and (n13397,n13398,n13399);
xor (n13398,n13395,n13396);
or (n13399,n13400,n13403);
and (n13400,n13401,n13402);
xor (n13401,n13316,n13317);
and (n13402,n4342,n3554);
and (n13403,n13404,n13405);
xor (n13404,n13401,n13402);
or (n13405,n13406,n13409);
and (n13406,n13407,n13408);
xor (n13407,n13321,n13322);
and (n13408,n4413,n3554);
and (n13409,n13410,n13411);
xor (n13410,n13407,n13408);
and (n13411,n13412,n13413);
xor (n13412,n13327,n13328);
and (n13413,n5241,n3554);
and (n13414,n13415,n13416);
xor (n13415,n12752,n4603);
or (n13416,n13417,n13419);
and (n13417,n13418,n4172);
xor (n13418,n13332,n13333);
and (n13419,n13420,n13421);
xor (n13420,n13418,n4172);
or (n13421,n13422,n13424);
and (n13422,n13423,n3712);
xor (n13423,n13338,n13339);
and (n13424,n13425,n13426);
xor (n13425,n13423,n3712);
or (n13426,n13427,n13429);
and (n13427,n13428,n3567);
xor (n13428,n13344,n13345);
and (n13429,n13430,n13431);
xor (n13430,n13428,n3567);
or (n13431,n13432,n13435);
and (n13432,n13433,n13434);
xor (n13433,n13350,n13351);
and (n13434,n3545,n3546);
and (n13435,n13436,n13437);
xor (n13436,n13433,n13434);
or (n13437,n13438,n13441);
and (n13438,n13439,n13440);
xor (n13439,n13356,n13357);
and (n13440,n3732,n3546);
and (n13441,n13442,n13443);
xor (n13442,n13439,n13440);
or (n13443,n13444,n13447);
and (n13444,n13445,n13446);
xor (n13445,n13362,n13363);
and (n13446,n3763,n3546);
and (n13447,n13448,n13449);
xor (n13448,n13445,n13446);
or (n13449,n13450,n13453);
and (n13450,n13451,n13452);
xor (n13451,n13368,n13369);
and (n13452,n3774,n3546);
and (n13453,n13454,n13455);
xor (n13454,n13451,n13452);
or (n13455,n13456,n13458);
and (n13456,n13457,n5200);
xor (n13457,n13374,n13375);
and (n13458,n13459,n13460);
xor (n13459,n13457,n5200);
or (n13460,n13461,n13463);
and (n13461,n13462,n5415);
xor (n13462,n13380,n13381);
and (n13463,n13464,n13465);
xor (n13464,n13462,n5415);
or (n13465,n13466,n13468);
and (n13466,n13467,n5634);
xor (n13467,n13386,n13387);
and (n13468,n13469,n13470);
xor (n13469,n13467,n5634);
or (n13470,n13471,n13473);
and (n13471,n13472,n5760);
xor (n13472,n13392,n13393);
and (n13473,n13474,n13475);
xor (n13474,n13472,n5760);
or (n13475,n13476,n13478);
and (n13476,n13477,n5942);
xor (n13477,n13398,n13399);
and (n13478,n13479,n13480);
xor (n13479,n13477,n5942);
or (n13480,n13481,n13483);
and (n13481,n13482,n6109);
xor (n13482,n13404,n13405);
and (n13483,n13484,n13485);
xor (n13484,n13482,n6109);
and (n13485,n13486,n6215);
xor (n13486,n13410,n13411);
and (n13487,n3704,n3741);
and (n13488,n13489,n13490);
xor (n13489,n12749,n13487);
or (n13490,n13491,n13494);
and (n13491,n13492,n13493);
xor (n13492,n13415,n13416);
and (n13493,n3537,n3741);
and (n13494,n13495,n13496);
xor (n13495,n13492,n13493);
or (n13496,n13497,n13500);
and (n13497,n13498,n13499);
xor (n13498,n13420,n13421);
and (n13499,n3518,n3741);
and (n13500,n13501,n13502);
xor (n13501,n13498,n13499);
or (n13502,n13503,n13506);
and (n13503,n13504,n13505);
xor (n13504,n13425,n13426);
and (n13505,n3566,n3741);
and (n13506,n13507,n13508);
xor (n13507,n13504,n13505);
or (n13508,n13509,n13512);
and (n13509,n13510,n13511);
xor (n13510,n13430,n13431);
and (n13511,n3545,n3741);
and (n13512,n13513,n13514);
xor (n13513,n13510,n13511);
or (n13514,n13515,n13518);
and (n13515,n13516,n13517);
xor (n13516,n13436,n13437);
and (n13517,n3732,n3741);
and (n13518,n13519,n13520);
xor (n13519,n13516,n13517);
or (n13520,n13521,n13524);
and (n13521,n13522,n13523);
xor (n13522,n13442,n13443);
and (n13523,n3763,n3741);
and (n13524,n13525,n13526);
xor (n13525,n13522,n13523);
or (n13526,n13527,n13530);
and (n13527,n13528,n13529);
xor (n13528,n13448,n13449);
and (n13529,n3774,n3741);
and (n13530,n13531,n13532);
xor (n13531,n13528,n13529);
or (n13532,n13533,n13536);
and (n13533,n13534,n13535);
xor (n13534,n13454,n13455);
and (n13535,n3651,n3741);
and (n13536,n13537,n13538);
xor (n13537,n13534,n13535);
or (n13538,n13539,n13542);
and (n13539,n13540,n13541);
xor (n13540,n13459,n13460);
and (n13541,n3670,n3741);
and (n13542,n13543,n13544);
xor (n13543,n13540,n13541);
or (n13544,n13545,n13548);
and (n13545,n13546,n13547);
xor (n13546,n13464,n13465);
and (n13547,n3929,n3741);
and (n13548,n13549,n13550);
xor (n13549,n13546,n13547);
or (n13550,n13551,n13554);
and (n13551,n13552,n13553);
xor (n13552,n13469,n13470);
and (n13553,n3935,n3741);
and (n13554,n13555,n13556);
xor (n13555,n13552,n13553);
or (n13556,n13557,n13560);
and (n13557,n13558,n13559);
xor (n13558,n13474,n13475);
and (n13559,n4342,n3741);
and (n13560,n13561,n13562);
xor (n13561,n13558,n13559);
or (n13562,n13563,n13566);
and (n13563,n13564,n13565);
xor (n13564,n13479,n13480);
and (n13565,n4413,n3741);
and (n13566,n13567,n13568);
xor (n13567,n13564,n13565);
and (n13568,n13569,n13570);
xor (n13569,n13484,n13485);
and (n13570,n5241,n3741);
and (n13571,n13572,n13573);
xor (n13572,n12746,n4780);
or (n13573,n13574,n13576);
and (n13574,n13575,n4701);
xor (n13575,n13489,n13490);
and (n13576,n13577,n13578);
xor (n13577,n13575,n4701);
or (n13578,n13579,n13581);
and (n13579,n13580,n4549);
xor (n13580,n13495,n13496);
and (n13581,n13582,n13583);
xor (n13582,n13580,n4549);
or (n13583,n13584,n13586);
and (n13584,n13585,n4245);
xor (n13585,n13501,n13502);
and (n13586,n13587,n13588);
xor (n13587,n13585,n4245);
or (n13588,n13589,n13591);
and (n13589,n13590,n3750);
xor (n13590,n13507,n13508);
and (n13591,n13592,n13593);
xor (n13592,n13590,n3750);
or (n13593,n13594,n13596);
and (n13594,n13595,n3731);
xor (n13595,n13513,n13514);
and (n13596,n13597,n13598);
xor (n13597,n13595,n3731);
or (n13598,n13599,n13601);
and (n13599,n13600,n3890);
xor (n13600,n13519,n13520);
and (n13601,n13602,n13603);
xor (n13602,n13600,n3890);
or (n13603,n13604,n13607);
and (n13604,n13605,n13606);
xor (n13605,n13525,n13526);
not (n13606,n3897);
and (n13607,n13608,n13609);
xor (n13608,n13605,n13606);
or (n13609,n13610,n13613);
and (n13610,n13611,n13612);
xor (n13611,n13531,n13532);
and (n13612,n3651,n3733);
and (n13613,n13614,n13615);
xor (n13614,n13611,n13612);
or (n13615,n13616,n13618);
and (n13616,n13617,n5109);
xor (n13617,n13537,n13538);
and (n13618,n13619,n13620);
xor (n13619,n13617,n5109);
or (n13620,n13621,n13624);
and (n13621,n13622,n13623);
xor (n13622,n13543,n13544);
and (n13623,n3929,n3733);
and (n13624,n13625,n13626);
xor (n13625,n13622,n13623);
or (n13626,n13627,n13630);
and (n13627,n13628,n13629);
xor (n13628,n13549,n13550);
and (n13629,n3935,n3733);
and (n13630,n13631,n13632);
xor (n13631,n13628,n13629);
or (n13632,n13633,n13635);
and (n13633,n13634,n5771);
xor (n13634,n13555,n13556);
and (n13635,n13636,n13637);
xor (n13636,n13634,n5771);
or (n13637,n13638,n13640);
and (n13638,n13639,n5803);
xor (n13639,n13561,n13562);
and (n13640,n13641,n13642);
xor (n13641,n13639,n5803);
and (n13642,n13643,n13644);
xor (n13643,n13567,n13568);
and (n13644,n5241,n3733);
and (n13645,n3704,n3756);
and (n13646,n13647,n13648);
xor (n13647,n12743,n13645);
or (n13648,n13649,n13652);
and (n13649,n13650,n13651);
xor (n13650,n13572,n13573);
and (n13651,n3537,n3756);
and (n13652,n13653,n13654);
xor (n13653,n13650,n13651);
or (n13654,n13655,n13658);
and (n13655,n13656,n13657);
xor (n13656,n13577,n13578);
and (n13657,n3518,n3756);
and (n13658,n13659,n13660);
xor (n13659,n13656,n13657);
or (n13660,n13661,n13664);
and (n13661,n13662,n13663);
xor (n13662,n13582,n13583);
and (n13663,n3566,n3756);
and (n13664,n13665,n13666);
xor (n13665,n13662,n13663);
or (n13666,n13667,n13670);
and (n13667,n13668,n13669);
xor (n13668,n13587,n13588);
and (n13669,n3545,n3756);
and (n13670,n13671,n13672);
xor (n13671,n13668,n13669);
or (n13672,n13673,n13676);
and (n13673,n13674,n13675);
xor (n13674,n13592,n13593);
and (n13675,n3732,n3756);
and (n13676,n13677,n13678);
xor (n13677,n13674,n13675);
or (n13678,n13679,n13682);
and (n13679,n13680,n13681);
xor (n13680,n13597,n13598);
and (n13681,n3763,n3756);
and (n13682,n13683,n13684);
xor (n13683,n13680,n13681);
or (n13684,n13685,n13688);
and (n13685,n13686,n13687);
xor (n13686,n13602,n13603);
and (n13687,n3774,n3756);
and (n13688,n13689,n13690);
xor (n13689,n13686,n13687);
or (n13690,n13691,n13694);
and (n13691,n13692,n13693);
xor (n13692,n13608,n13609);
and (n13693,n3651,n3756);
and (n13694,n13695,n13696);
xor (n13695,n13692,n13693);
or (n13696,n13697,n13700);
and (n13697,n13698,n13699);
xor (n13698,n13614,n13615);
and (n13699,n3670,n3756);
and (n13700,n13701,n13702);
xor (n13701,n13698,n13699);
or (n13702,n13703,n13706);
and (n13703,n13704,n13705);
xor (n13704,n13619,n13620);
and (n13705,n3929,n3756);
and (n13706,n13707,n13708);
xor (n13707,n13704,n13705);
or (n13708,n13709,n13712);
and (n13709,n13710,n13711);
xor (n13710,n13625,n13626);
and (n13711,n3935,n3756);
and (n13712,n13713,n13714);
xor (n13713,n13710,n13711);
or (n13714,n13715,n13718);
and (n13715,n13716,n13717);
xor (n13716,n13631,n13632);
and (n13717,n4342,n3756);
and (n13718,n13719,n13720);
xor (n13719,n13716,n13717);
or (n13720,n13721,n13724);
and (n13721,n13722,n13723);
xor (n13722,n13636,n13637);
and (n13723,n4413,n3756);
and (n13724,n13725,n13726);
xor (n13725,n13722,n13723);
and (n13726,n13727,n13728);
xor (n13727,n13641,n13642);
and (n13728,n5241,n3756);
and (n13729,n13730,n13731);
xor (n13730,n12740,n4930);
or (n13731,n13732,n13735);
and (n13732,n13733,n13734);
xor (n13733,n13647,n13648);
and (n13734,n3537,n3659);
and (n13735,n13736,n13737);
xor (n13736,n13733,n13734);
or (n13737,n13738,n13740);
and (n13738,n13739,n4796);
xor (n13739,n13653,n13654);
and (n13740,n13741,n13742);
xor (n13741,n13739,n4796);
or (n13742,n13743,n13745);
and (n13743,n13744,n4707);
xor (n13744,n13659,n13660);
and (n13745,n13746,n13747);
xor (n13746,n13744,n4707);
or (n13747,n13748,n13750);
and (n13748,n13749,n4555);
xor (n13749,n13665,n13666);
and (n13750,n13751,n13752);
xor (n13751,n13749,n4555);
or (n13752,n13753,n13755);
and (n13753,n13754,n4252);
xor (n13754,n13671,n13672);
and (n13755,n13756,n13757);
xor (n13756,n13754,n4252);
or (n13757,n13758,n13761);
and (n13758,n13759,n13760);
xor (n13759,n13677,n13678);
and (n13760,n3763,n3659);
and (n13761,n13762,n13763);
xor (n13762,n13759,n13760);
or (n13763,n13764,n13767);
and (n13764,n13765,n13766);
xor (n13765,n13683,n13684);
not (n13766,n3775);
and (n13767,n13768,n13769);
xor (n13768,n13765,n13766);
or (n13769,n13770,n13773);
and (n13770,n13771,n13772);
xor (n13771,n13689,n13690);
not (n13772,n3907);
and (n13773,n13774,n13775);
xor (n13774,n13771,n13772);
or (n13775,n13776,n13778);
and (n13776,n13777,n3911);
xor (n13777,n13695,n13696);
and (n13778,n13779,n13780);
xor (n13779,n13777,n3911);
or (n13780,n13781,n13783);
and (n13781,n13782,n3985);
xor (n13782,n13701,n13702);
and (n13783,n13784,n13785);
xor (n13784,n13782,n3985);
or (n13785,n13786,n13788);
and (n13786,n13787,n5117);
xor (n13787,n13707,n13708);
and (n13788,n13789,n13790);
xor (n13789,n13787,n5117);
or (n13790,n13791,n13793);
and (n13791,n13792,n5264);
xor (n13792,n13713,n13714);
and (n13793,n13794,n13795);
xor (n13794,n13792,n5264);
or (n13795,n13796,n13798);
and (n13796,n13797,n5497);
xor (n13797,n13719,n13720);
and (n13798,n13799,n13800);
xor (n13799,n13797,n5497);
and (n13800,n13801,n5777);
xor (n13801,n13725,n13726);
and (n13802,n3704,n3657);
and (n13803,n13804,n13805);
xor (n13804,n12737,n13802);
or (n13805,n13806,n13809);
and (n13806,n13807,n13808);
xor (n13807,n13730,n13731);
and (n13808,n3537,n3657);
and (n13809,n13810,n13811);
xor (n13810,n13807,n13808);
or (n13811,n13812,n13815);
and (n13812,n13813,n13814);
xor (n13813,n13736,n13737);
and (n13814,n3518,n3657);
and (n13815,n13816,n13817);
xor (n13816,n13813,n13814);
or (n13817,n13818,n13821);
and (n13818,n13819,n13820);
xor (n13819,n13741,n13742);
and (n13820,n3566,n3657);
and (n13821,n13822,n13823);
xor (n13822,n13819,n13820);
or (n13823,n13824,n13827);
and (n13824,n13825,n13826);
xor (n13825,n13746,n13747);
and (n13826,n3545,n3657);
and (n13827,n13828,n13829);
xor (n13828,n13825,n13826);
or (n13829,n13830,n13833);
and (n13830,n13831,n13832);
xor (n13831,n13751,n13752);
and (n13832,n3732,n3657);
and (n13833,n13834,n13835);
xor (n13834,n13831,n13832);
or (n13835,n13836,n13839);
and (n13836,n13837,n13838);
xor (n13837,n13756,n13757);
and (n13838,n3763,n3657);
and (n13839,n13840,n13841);
xor (n13840,n13837,n13838);
or (n13841,n13842,n13845);
and (n13842,n13843,n13844);
xor (n13843,n13762,n13763);
and (n13844,n3774,n3657);
and (n13845,n13846,n13847);
xor (n13846,n13843,n13844);
or (n13847,n13848,n13851);
and (n13848,n13849,n13850);
xor (n13849,n13768,n13769);
and (n13850,n3651,n3657);
and (n13851,n13852,n13853);
xor (n13852,n13849,n13850);
or (n13853,n13854,n13857);
and (n13854,n13855,n13856);
xor (n13855,n13774,n13775);
and (n13856,n3670,n3657);
and (n13857,n13858,n13859);
xor (n13858,n13855,n13856);
or (n13859,n13860,n13863);
and (n13860,n13861,n13862);
xor (n13861,n13779,n13780);
and (n13862,n3929,n3657);
and (n13863,n13864,n13865);
xor (n13864,n13861,n13862);
or (n13865,n13866,n13869);
and (n13866,n13867,n13868);
xor (n13867,n13784,n13785);
and (n13868,n3935,n3657);
and (n13869,n13870,n13871);
xor (n13870,n13867,n13868);
or (n13871,n13872,n13875);
and (n13872,n13873,n13874);
xor (n13873,n13789,n13790);
and (n13874,n4342,n3657);
and (n13875,n13876,n13877);
xor (n13876,n13873,n13874);
or (n13877,n13878,n13881);
and (n13878,n13879,n13880);
xor (n13879,n13794,n13795);
and (n13880,n4413,n3657);
and (n13881,n13882,n13883);
xor (n13882,n13879,n13880);
and (n13883,n13884,n13885);
xor (n13884,n13799,n13800);
and (n13885,n5241,n3657);
and (n13886,n13887,n13888);
xor (n13887,n12734,n5016);
or (n13888,n13889,n13891);
and (n13889,n13890,n4966);
xor (n13890,n13804,n13805);
and (n13891,n13892,n13893);
xor (n13892,n13890,n4966);
or (n13893,n13894,n13896);
and (n13894,n13895,n4894);
xor (n13895,n13810,n13811);
and (n13896,n13897,n13898);
xor (n13897,n13895,n4894);
or (n13898,n13899,n13901);
and (n13899,n13900,n4834);
xor (n13900,n13816,n13817);
and (n13901,n13902,n13903);
xor (n13902,n13900,n4834);
or (n13903,n13904,n13906);
and (n13904,n13905,n4756);
xor (n13905,n13822,n13823);
and (n13906,n13907,n13908);
xor (n13907,n13905,n4756);
or (n13908,n13909,n13912);
and (n13909,n13910,n13911);
xor (n13910,n13828,n13829);
not (n13911,n4676);
and (n13912,n13913,n13914);
xor (n13913,n13910,n13911);
or (n13914,n13915,n13917);
and (n13915,n13916,n4572);
xor (n13916,n13834,n13835);
and (n13917,n13918,n13919);
xor (n13918,n13916,n4572);
or (n13919,n13920,n13922);
and (n13920,n13921,n4269);
xor (n13921,n13840,n13841);
and (n13922,n13923,n13924);
xor (n13923,n13921,n4269);
or (n13924,n13925,n13928);
and (n13925,n13926,n13927);
xor (n13926,n13846,n13847);
and (n13927,n3651,n3650);
and (n13928,n13929,n13930);
xor (n13929,n13926,n13927);
or (n13930,n13931,n13933);
and (n13931,n13932,n3669);
xor (n13932,n13852,n13853);
and (n13933,n13934,n13935);
xor (n13934,n13932,n3669);
or (n13935,n13936,n13939);
and (n13936,n13937,n13938);
xor (n13937,n13858,n13859);
not (n13938,n3930);
and (n13939,n13940,n13941);
xor (n13940,n13937,n13938);
or (n13941,n13942,n13944);
and (n13942,n13943,n3934);
xor (n13943,n13864,n13865);
and (n13944,n13945,n13946);
xor (n13945,n13943,n3934);
or (n13946,n13947,n13949);
and (n13947,n13948,n4343);
xor (n13948,n13870,n13871);
and (n13949,n13950,n13951);
xor (n13950,n13948,n4343);
or (n13951,n13952,n13954);
and (n13952,n13953,n4412);
xor (n13953,n13876,n13877);
and (n13954,n13955,n13956);
xor (n13955,n13953,n4412);
and (n13956,n13957,n5270);
xor (n13957,n13882,n13883);
and (n13958,n13959,n13960);
xor (n13959,n12731,n5016);
or (n13960,n13961,n13963);
and (n13961,n13962,n4966);
xor (n13962,n13887,n13888);
and (n13963,n13964,n13965);
xor (n13964,n13962,n4966);
or (n13965,n13966,n13968);
and (n13966,n13967,n4894);
xor (n13967,n13892,n13893);
and (n13968,n13969,n13970);
xor (n13969,n13967,n4894);
or (n13970,n13971,n13973);
and (n13971,n13972,n4834);
xor (n13972,n13897,n13898);
and (n13973,n13974,n13975);
xor (n13974,n13972,n4834);
or (n13975,n13976,n13978);
and (n13976,n13977,n4756);
xor (n13977,n13902,n13903);
and (n13978,n13979,n13980);
xor (n13979,n13977,n4756);
or (n13980,n13981,n13983);
and (n13981,n13982,n13911);
xor (n13982,n13907,n13908);
and (n13983,n13984,n13985);
xor (n13984,n13982,n13911);
or (n13985,n13986,n13988);
and (n13986,n13987,n4572);
xor (n13987,n13913,n13914);
and (n13988,n13989,n13990);
xor (n13989,n13987,n4572);
or (n13990,n13991,n13993);
and (n13991,n13992,n4269);
xor (n13992,n13918,n13919);
and (n13993,n13994,n13995);
xor (n13994,n13992,n4269);
or (n13995,n13996,n13998);
and (n13996,n13997,n13927);
xor (n13997,n13923,n13924);
and (n13998,n13999,n14000);
xor (n13999,n13997,n13927);
or (n14000,n14001,n14003);
and (n14001,n14002,n3669);
xor (n14002,n13929,n13930);
and (n14003,n14004,n14005);
xor (n14004,n14002,n3669);
or (n14005,n14006,n14008);
and (n14006,n14007,n13938);
xor (n14007,n13934,n13935);
and (n14008,n14009,n14010);
xor (n14009,n14007,n13938);
or (n14010,n14011,n14013);
and (n14011,n14012,n3934);
xor (n14012,n13940,n13941);
and (n14013,n14014,n14015);
xor (n14014,n14012,n3934);
or (n14015,n14016,n14018);
and (n14016,n14017,n4343);
xor (n14017,n13945,n13946);
and (n14018,n14019,n14020);
xor (n14019,n14017,n4343);
or (n14020,n14021,n14023);
and (n14021,n14022,n4412);
xor (n14022,n13950,n13951);
and (n14023,n14024,n14025);
xor (n14024,n14022,n4412);
and (n14025,n14026,n5270);
xor (n14026,n13955,n13956);
or (n14027,n14028,n14030);
and (n14028,n14029,n4966);
xor (n14029,n13959,n13960);
and (n14030,n14031,n14032);
xor (n14031,n14029,n4966);
or (n14032,n14033,n14035);
and (n14033,n14034,n4894);
xor (n14034,n13964,n13965);
and (n14035,n14036,n14037);
xor (n14036,n14034,n4894);
or (n14037,n14038,n14040);
and (n14038,n14039,n4834);
xor (n14039,n13969,n13970);
and (n14040,n14041,n14042);
xor (n14041,n14039,n4834);
or (n14042,n14043,n14045);
and (n14043,n14044,n4756);
xor (n14044,n13974,n13975);
and (n14045,n14046,n14047);
xor (n14046,n14044,n4756);
or (n14047,n14048,n14050);
and (n14048,n14049,n13911);
xor (n14049,n13979,n13980);
and (n14050,n14051,n14052);
xor (n14051,n14049,n13911);
or (n14052,n14053,n14055);
and (n14053,n14054,n4572);
xor (n14054,n13984,n13985);
and (n14055,n14056,n14057);
xor (n14056,n14054,n4572);
or (n14057,n14058,n14060);
and (n14058,n14059,n4269);
xor (n14059,n13989,n13990);
and (n14060,n14061,n14062);
xor (n14061,n14059,n4269);
or (n14062,n14063,n14065);
and (n14063,n14064,n13927);
xor (n14064,n13994,n13995);
and (n14065,n14066,n14067);
xor (n14066,n14064,n13927);
or (n14067,n14068,n14070);
and (n14068,n14069,n3669);
xor (n14069,n13999,n14000);
and (n14070,n14071,n14072);
xor (n14071,n14069,n3669);
or (n14072,n14073,n14075);
and (n14073,n14074,n13938);
xor (n14074,n14004,n14005);
and (n14075,n14076,n14077);
xor (n14076,n14074,n13938);
or (n14077,n14078,n14080);
and (n14078,n14079,n3934);
xor (n14079,n14009,n14010);
and (n14080,n14081,n14082);
xor (n14081,n14079,n3934);
or (n14082,n14083,n14085);
and (n14083,n14084,n4343);
xor (n14084,n14014,n14015);
and (n14085,n14086,n14087);
xor (n14086,n14084,n4343);
or (n14087,n14088,n14090);
and (n14088,n14089,n4412);
xor (n14089,n14019,n14020);
and (n14090,n14091,n14092);
xor (n14091,n14089,n4412);
and (n14092,n14093,n5270);
xor (n14093,n14024,n14025);
or (n14094,n14095,n14097);
and (n14095,n14096,n4894);
xor (n14096,n14031,n14032);
and (n14097,n14098,n14099);
xor (n14098,n14096,n4894);
or (n14099,n14100,n14102);
and (n14100,n14101,n4834);
xor (n14101,n14036,n14037);
and (n14102,n14103,n14104);
xor (n14103,n14101,n4834);
or (n14104,n14105,n14107);
and (n14105,n14106,n4756);
xor (n14106,n14041,n14042);
and (n14107,n14108,n14109);
xor (n14108,n14106,n4756);
or (n14109,n14110,n14112);
and (n14110,n14111,n13911);
xor (n14111,n14046,n14047);
and (n14112,n14113,n14114);
xor (n14113,n14111,n13911);
or (n14114,n14115,n14117);
and (n14115,n14116,n4572);
xor (n14116,n14051,n14052);
and (n14117,n14118,n14119);
xor (n14118,n14116,n4572);
or (n14119,n14120,n14122);
and (n14120,n14121,n4269);
xor (n14121,n14056,n14057);
and (n14122,n14123,n14124);
xor (n14123,n14121,n4269);
or (n14124,n14125,n14127);
and (n14125,n14126,n13927);
xor (n14126,n14061,n14062);
and (n14127,n14128,n14129);
xor (n14128,n14126,n13927);
or (n14129,n14130,n14132);
and (n14130,n14131,n3669);
xor (n14131,n14066,n14067);
and (n14132,n14133,n14134);
xor (n14133,n14131,n3669);
or (n14134,n14135,n14137);
and (n14135,n14136,n13938);
xor (n14136,n14071,n14072);
and (n14137,n14138,n14139);
xor (n14138,n14136,n13938);
or (n14139,n14140,n14142);
and (n14140,n14141,n3934);
xor (n14141,n14076,n14077);
and (n14142,n14143,n14144);
xor (n14143,n14141,n3934);
or (n14144,n14145,n14147);
and (n14145,n14146,n4343);
xor (n14146,n14081,n14082);
and (n14147,n14148,n14149);
xor (n14148,n14146,n4343);
or (n14149,n14150,n14152);
and (n14150,n14151,n4412);
xor (n14151,n14086,n14087);
and (n14152,n14153,n14154);
xor (n14153,n14151,n4412);
and (n14154,n14155,n5270);
xor (n14155,n14091,n14092);
or (n14156,n14157,n14159);
and (n14157,n14158,n4834);
xor (n14158,n14098,n14099);
and (n14159,n14160,n14161);
xor (n14160,n14158,n4834);
or (n14161,n14162,n14164);
and (n14162,n14163,n4756);
xor (n14163,n14103,n14104);
and (n14164,n14165,n14166);
xor (n14165,n14163,n4756);
or (n14166,n14167,n14169);
and (n14167,n14168,n13911);
xor (n14168,n14108,n14109);
and (n14169,n14170,n14171);
xor (n14170,n14168,n13911);
or (n14171,n14172,n14174);
and (n14172,n14173,n4572);
xor (n14173,n14113,n14114);
and (n14174,n14175,n14176);
xor (n14175,n14173,n4572);
or (n14176,n14177,n14179);
and (n14177,n14178,n4269);
xor (n14178,n14118,n14119);
and (n14179,n14180,n14181);
xor (n14180,n14178,n4269);
or (n14181,n14182,n14184);
and (n14182,n14183,n13927);
xor (n14183,n14123,n14124);
and (n14184,n14185,n14186);
xor (n14185,n14183,n13927);
or (n14186,n14187,n14189);
and (n14187,n14188,n3669);
xor (n14188,n14128,n14129);
and (n14189,n14190,n14191);
xor (n14190,n14188,n3669);
or (n14191,n14192,n14194);
and (n14192,n14193,n13938);
xor (n14193,n14133,n14134);
and (n14194,n14195,n14196);
xor (n14195,n14193,n13938);
or (n14196,n14197,n14199);
and (n14197,n14198,n3934);
xor (n14198,n14138,n14139);
and (n14199,n14200,n14201);
xor (n14200,n14198,n3934);
or (n14201,n14202,n14204);
and (n14202,n14203,n4343);
xor (n14203,n14143,n14144);
and (n14204,n14205,n14206);
xor (n14205,n14203,n4343);
or (n14206,n14207,n14209);
and (n14207,n14208,n4412);
xor (n14208,n14148,n14149);
and (n14209,n14210,n14211);
xor (n14210,n14208,n4412);
and (n14211,n14212,n5270);
xor (n14212,n14153,n14154);
or (n14213,n14214,n14216);
and (n14214,n14215,n4756);
xor (n14215,n14160,n14161);
and (n14216,n14217,n14218);
xor (n14217,n14215,n4756);
or (n14218,n14219,n14221);
and (n14219,n14220,n13911);
xor (n14220,n14165,n14166);
and (n14221,n14222,n14223);
xor (n14222,n14220,n13911);
or (n14223,n14224,n14226);
and (n14224,n14225,n4572);
xor (n14225,n14170,n14171);
and (n14226,n14227,n14228);
xor (n14227,n14225,n4572);
or (n14228,n14229,n14231);
and (n14229,n14230,n4269);
xor (n14230,n14175,n14176);
and (n14231,n14232,n14233);
xor (n14232,n14230,n4269);
or (n14233,n14234,n14236);
and (n14234,n14235,n13927);
xor (n14235,n14180,n14181);
and (n14236,n14237,n14238);
xor (n14237,n14235,n13927);
or (n14238,n14239,n14241);
and (n14239,n14240,n3669);
xor (n14240,n14185,n14186);
and (n14241,n14242,n14243);
xor (n14242,n14240,n3669);
or (n14243,n14244,n14246);
and (n14244,n14245,n13938);
xor (n14245,n14190,n14191);
and (n14246,n14247,n14248);
xor (n14247,n14245,n13938);
or (n14248,n14249,n14251);
and (n14249,n14250,n3934);
xor (n14250,n14195,n14196);
and (n14251,n14252,n14253);
xor (n14252,n14250,n3934);
or (n14253,n14254,n14256);
and (n14254,n14255,n4343);
xor (n14255,n14200,n14201);
and (n14256,n14257,n14258);
xor (n14257,n14255,n4343);
or (n14258,n14259,n14261);
and (n14259,n14260,n4412);
xor (n14260,n14205,n14206);
and (n14261,n14262,n14263);
xor (n14262,n14260,n4412);
and (n14263,n14264,n5270);
xor (n14264,n14210,n14211);
or (n14265,n14266,n14268);
and (n14266,n14267,n13911);
xor (n14267,n14217,n14218);
and (n14268,n14269,n14270);
xor (n14269,n14267,n13911);
or (n14270,n14271,n14273);
and (n14271,n14272,n4572);
xor (n14272,n14222,n14223);
and (n14273,n14274,n14275);
xor (n14274,n14272,n4572);
or (n14275,n14276,n14278);
and (n14276,n14277,n4269);
xor (n14277,n14227,n14228);
and (n14278,n14279,n14280);
xor (n14279,n14277,n4269);
or (n14280,n14281,n14283);
and (n14281,n14282,n13927);
xor (n14282,n14232,n14233);
and (n14283,n14284,n14285);
xor (n14284,n14282,n13927);
or (n14285,n14286,n14288);
and (n14286,n14287,n3669);
xor (n14287,n14237,n14238);
and (n14288,n14289,n14290);
xor (n14289,n14287,n3669);
or (n14290,n14291,n14293);
and (n14291,n14292,n13938);
xor (n14292,n14242,n14243);
and (n14293,n14294,n14295);
xor (n14294,n14292,n13938);
or (n14295,n14296,n14298);
and (n14296,n14297,n3934);
xor (n14297,n14247,n14248);
and (n14298,n14299,n14300);
xor (n14299,n14297,n3934);
or (n14300,n14301,n14303);
and (n14301,n14302,n4343);
xor (n14302,n14252,n14253);
and (n14303,n14304,n14305);
xor (n14304,n14302,n4343);
or (n14305,n14306,n14308);
and (n14306,n14307,n4412);
xor (n14307,n14257,n14258);
and (n14308,n14309,n14310);
xor (n14309,n14307,n4412);
and (n14310,n14311,n5270);
xor (n14311,n14262,n14263);
or (n14312,n14313,n14315);
and (n14313,n14314,n4572);
xor (n14314,n14269,n14270);
and (n14315,n14316,n14317);
xor (n14316,n14314,n4572);
or (n14317,n14318,n14320);
and (n14318,n14319,n4269);
xor (n14319,n14274,n14275);
and (n14320,n14321,n14322);
xor (n14321,n14319,n4269);
or (n14322,n14323,n14325);
and (n14323,n14324,n13927);
xor (n14324,n14279,n14280);
and (n14325,n14326,n14327);
xor (n14326,n14324,n13927);
or (n14327,n14328,n14330);
and (n14328,n14329,n3669);
xor (n14329,n14284,n14285);
and (n14330,n14331,n14332);
xor (n14331,n14329,n3669);
or (n14332,n14333,n14335);
and (n14333,n14334,n13938);
xor (n14334,n14289,n14290);
and (n14335,n14336,n14337);
xor (n14336,n14334,n13938);
or (n14337,n14338,n14340);
and (n14338,n14339,n3934);
xor (n14339,n14294,n14295);
and (n14340,n14341,n14342);
xor (n14341,n14339,n3934);
or (n14342,n14343,n14345);
and (n14343,n14344,n4343);
xor (n14344,n14299,n14300);
and (n14345,n14346,n14347);
xor (n14346,n14344,n4343);
or (n14347,n14348,n14350);
and (n14348,n14349,n4412);
xor (n14349,n14304,n14305);
and (n14350,n14351,n14352);
xor (n14351,n14349,n4412);
and (n14352,n14353,n5270);
xor (n14353,n14309,n14310);
or (n14354,n14355,n14357);
and (n14355,n14356,n4269);
xor (n14356,n14316,n14317);
and (n14357,n14358,n14359);
xor (n14358,n14356,n4269);
or (n14359,n14360,n14362);
and (n14360,n14361,n13927);
xor (n14361,n14321,n14322);
and (n14362,n14363,n14364);
xor (n14363,n14361,n13927);
or (n14364,n14365,n14367);
and (n14365,n14366,n3669);
xor (n14366,n14326,n14327);
and (n14367,n14368,n14369);
xor (n14368,n14366,n3669);
or (n14369,n14370,n14372);
and (n14370,n14371,n13938);
xor (n14371,n14331,n14332);
and (n14372,n14373,n14374);
xor (n14373,n14371,n13938);
or (n14374,n14375,n14377);
and (n14375,n14376,n3934);
xor (n14376,n14336,n14337);
and (n14377,n14378,n14379);
xor (n14378,n14376,n3934);
or (n14379,n14380,n14382);
and (n14380,n14381,n4343);
xor (n14381,n14341,n14342);
and (n14382,n14383,n14384);
xor (n14383,n14381,n4343);
or (n14384,n14385,n14387);
and (n14385,n14386,n4412);
xor (n14386,n14346,n14347);
and (n14387,n14388,n14389);
xor (n14388,n14386,n4412);
and (n14389,n14390,n5270);
xor (n14390,n14351,n14352);
or (n14391,n14392,n14394);
and (n14392,n14393,n13927);
xor (n14393,n14358,n14359);
and (n14394,n14395,n14396);
xor (n14395,n14393,n13927);
or (n14396,n14397,n14399);
and (n14397,n14398,n3669);
xor (n14398,n14363,n14364);
and (n14399,n14400,n14401);
xor (n14400,n14398,n3669);
or (n14401,n14402,n14404);
and (n14402,n14403,n13938);
xor (n14403,n14368,n14369);
and (n14404,n14405,n14406);
xor (n14405,n14403,n13938);
or (n14406,n14407,n14409);
and (n14407,n14408,n3934);
xor (n14408,n14373,n14374);
and (n14409,n14410,n14411);
xor (n14410,n14408,n3934);
or (n14411,n14412,n14414);
and (n14412,n14413,n4343);
xor (n14413,n14378,n14379);
and (n14414,n14415,n14416);
xor (n14415,n14413,n4343);
or (n14416,n14417,n14419);
and (n14417,n14418,n4412);
xor (n14418,n14383,n14384);
and (n14419,n14420,n14421);
xor (n14420,n14418,n4412);
and (n14421,n14422,n5270);
xor (n14422,n14388,n14389);
or (n14423,n14424,n14426);
and (n14424,n14425,n3669);
xor (n14425,n14395,n14396);
and (n14426,n14427,n14428);
xor (n14427,n14425,n3669);
or (n14428,n14429,n14431);
and (n14429,n14430,n13938);
xor (n14430,n14400,n14401);
and (n14431,n14432,n14433);
xor (n14432,n14430,n13938);
or (n14433,n14434,n14436);
and (n14434,n14435,n3934);
xor (n14435,n14405,n14406);
and (n14436,n14437,n14438);
xor (n14437,n14435,n3934);
or (n14438,n14439,n14441);
and (n14439,n14440,n4343);
xor (n14440,n14410,n14411);
and (n14441,n14442,n14443);
xor (n14442,n14440,n4343);
or (n14443,n14444,n14446);
and (n14444,n14445,n4412);
xor (n14445,n14415,n14416);
and (n14446,n14447,n14448);
xor (n14447,n14445,n4412);
and (n14448,n14449,n5270);
xor (n14449,n14420,n14421);
or (n14450,n14451,n14453);
and (n14451,n14452,n13938);
xor (n14452,n14427,n14428);
and (n14453,n14454,n14455);
xor (n14454,n14452,n13938);
or (n14455,n14456,n14458);
and (n14456,n14457,n3934);
xor (n14457,n14432,n14433);
and (n14458,n14459,n14460);
xor (n14459,n14457,n3934);
or (n14460,n14461,n14463);
and (n14461,n14462,n4343);
xor (n14462,n14437,n14438);
and (n14463,n14464,n14465);
xor (n14464,n14462,n4343);
or (n14465,n14466,n14468);
and (n14466,n14467,n4412);
xor (n14467,n14442,n14443);
and (n14468,n14469,n14470);
xor (n14469,n14467,n4412);
and (n14470,n14471,n5270);
xor (n14471,n14447,n14448);
or (n14472,n14473,n14475);
and (n14473,n14474,n3934);
xor (n14474,n14454,n14455);
and (n14475,n14476,n14477);
xor (n14476,n14474,n3934);
or (n14477,n14478,n14480);
and (n14478,n14479,n4343);
xor (n14479,n14459,n14460);
and (n14480,n14481,n14482);
xor (n14481,n14479,n4343);
or (n14482,n14483,n14485);
and (n14483,n14484,n4412);
xor (n14484,n14464,n14465);
and (n14485,n14486,n14487);
xor (n14486,n14484,n4412);
and (n14487,n14488,n5270);
xor (n14488,n14469,n14470);
or (n14489,n14490,n14492);
and (n14490,n14491,n4343);
xor (n14491,n14476,n14477);
and (n14492,n14493,n14494);
xor (n14493,n14491,n4343);
or (n14494,n14495,n14497);
and (n14495,n14496,n4412);
xor (n14496,n14481,n14482);
and (n14497,n14498,n14499);
xor (n14498,n14496,n4412);
and (n14499,n14500,n5270);
xor (n14500,n14486,n14487);
or (n14501,n14502,n14504);
and (n14502,n14503,n4412);
xor (n14503,n14493,n14494);
and (n14504,n14505,n14506);
xor (n14505,n14503,n4412);
and (n14506,n14507,n5270);
xor (n14507,n14498,n14499);
and (n14508,n14509,n5270);
xor (n14509,n14505,n14506);
or (n14510,n14511,n14515,n14721);
and (n14511,n14512,n14513);
xor (n14512,n12640,n12088);
not (n14513,n14514);
xor (n14514,n14509,n5270);
and (n14515,n14513,n14516);
or (n14516,n14517,n14521,n14720);
and (n14517,n14518,n14519);
xor (n14518,n12638,n12088);
not (n14519,n14520);
xor (n14520,n14507,n5270);
and (n14521,n14519,n14522);
or (n14522,n14523,n14527,n14719);
and (n14523,n14524,n14525);
xor (n14524,n12631,n12088);
not (n14525,n14526);
xor (n14526,n14500,n5270);
and (n14527,n14525,n14528);
or (n14528,n14529,n14533,n14718);
and (n14529,n14530,n14531);
xor (n14530,n12619,n12088);
not (n14531,n14532);
xor (n14532,n14488,n5270);
and (n14533,n14531,n14534);
or (n14534,n14535,n14539,n14717);
and (n14535,n14536,n14537);
xor (n14536,n12602,n12088);
not (n14537,n14538);
xor (n14538,n14471,n5270);
and (n14539,n14537,n14540);
or (n14540,n14541,n14545,n14716);
and (n14541,n14542,n14543);
xor (n14542,n12580,n12088);
not (n14543,n14544);
xor (n14544,n14449,n5270);
and (n14545,n14543,n14546);
or (n14546,n14547,n14551,n14715);
and (n14547,n14548,n14549);
xor (n14548,n12553,n12088);
not (n14549,n14550);
xor (n14550,n14422,n5270);
and (n14551,n14549,n14552);
or (n14552,n14553,n14557,n14714);
and (n14553,n14554,n14555);
xor (n14554,n12521,n12088);
not (n14555,n14556);
xor (n14556,n14390,n5270);
and (n14557,n14555,n14558);
or (n14558,n14559,n14563,n14713);
and (n14559,n14560,n14561);
xor (n14560,n12484,n12088);
not (n14561,n14562);
xor (n14562,n14353,n5270);
and (n14563,n14561,n14564);
or (n14564,n14565,n14569,n14712);
and (n14565,n14566,n14567);
xor (n14566,n12442,n12088);
not (n14567,n14568);
xor (n14568,n14311,n5270);
and (n14569,n14567,n14570);
or (n14570,n14571,n14575,n14711);
and (n14571,n14572,n14573);
xor (n14572,n12395,n12088);
not (n14573,n14574);
xor (n14574,n14264,n5270);
and (n14575,n14573,n14576);
or (n14576,n14577,n14581,n14710);
and (n14577,n14578,n14579);
xor (n14578,n12343,n12088);
not (n14579,n14580);
xor (n14580,n14212,n5270);
and (n14581,n14579,n14582);
or (n14582,n14583,n14587,n14709);
and (n14583,n14584,n14585);
xor (n14584,n12286,n12088);
not (n14585,n14586);
xor (n14586,n14155,n5270);
and (n14587,n14585,n14588);
or (n14588,n14589,n14593,n14708);
and (n14589,n14590,n14591);
xor (n14590,n12224,n12088);
not (n14591,n14592);
xor (n14592,n14093,n5270);
and (n14593,n14591,n14594);
or (n14594,n14595,n14599,n14707);
and (n14595,n14596,n14597);
xor (n14596,n12157,n12088);
not (n14597,n14598);
xor (n14598,n14026,n5270);
and (n14599,n14597,n14600);
or (n14600,n14601,n14605,n14706);
and (n14601,n14602,n14603);
xor (n14602,n12087,n12088);
not (n14603,n14604);
xor (n14604,n13957,n5270);
and (n14605,n14603,n14606);
or (n14606,n14607,n14611,n14705);
and (n14607,n14608,n14609);
xor (n14608,n12007,n5232);
not (n14609,n14610);
xor (n14610,n13884,n13885);
and (n14611,n14609,n14612);
or (n14612,n14613,n14617,n14704);
and (n14613,n14614,n14615);
xor (n14614,n11923,n11924);
not (n14615,n14616);
xor (n14616,n13801,n5777);
and (n14617,n14615,n14618);
or (n14618,n14619,n14623,n14703);
and (n14619,n14620,n14621);
xor (n14620,n11843,n5528);
not (n14621,n14622);
xor (n14622,n13727,n13728);
and (n14623,n14621,n14624);
or (n14624,n14625,n14629,n14702);
and (n14625,n14626,n14627);
xor (n14626,n11760,n5935);
not (n14627,n14628);
xor (n14628,n13643,n13644);
and (n14629,n14627,n14630);
or (n14630,n14631,n14635,n14701);
and (n14631,n14632,n14633);
xor (n14632,n11684,n5979);
not (n14633,n14634);
xor (n14634,n13569,n13570);
and (n14635,n14633,n14636);
or (n14636,n14637,n14641,n14700);
and (n14637,n14638,n14639);
xor (n14638,n11600,n11601);
not (n14639,n14640);
xor (n14640,n13486,n6215);
and (n14641,n14639,n14642);
or (n14642,n14643,n14647,n14699);
and (n14643,n14644,n14645);
xor (n14644,n11520,n6224);
not (n14645,n14646);
xor (n14646,n13412,n13413);
and (n14647,n14645,n14648);
or (n14648,n14649,n14653,n14698);
and (n14649,n14650,n14651);
xor (n14650,n11437,n6446);
not (n14651,n14652);
xor (n14652,n13329,n6465);
and (n14653,n14651,n14654);
or (n14654,n14655,n14659,n14697);
and (n14655,n14656,n14657);
xor (n14656,n11355,n6432);
not (n14657,n14658);
xor (n14658,n13252,n13253);
and (n14659,n14657,n14660);
or (n14660,n14661,n14665,n14696);
and (n14661,n14662,n14663);
xor (n14662,n11272,n6682);
not (n14663,n14664);
xor (n14664,n13169,n6697);
and (n14665,n14663,n14666);
or (n14666,n14667,n14671,n14695);
and (n14667,n14668,n14669);
xor (n14668,n11192,n6614);
not (n14669,n14670);
xor (n14670,n13091,n13092);
and (n14671,n14669,n14672);
or (n14672,n14673,n14677,n14694);
and (n14673,n14674,n14675);
xor (n14674,n11108,n11109);
not (n14675,n14676);
xor (n14676,n13008,n6771);
and (n14677,n14675,n14678);
or (n14678,n14679,n14683,n14693);
and (n14679,n14680,n14681);
xor (n14680,n11028,n6728);
not (n14681,n14682);
xor (n14682,n12931,n12932);
and (n14683,n14681,n14684);
or (n14684,n14685,n14689,n14692);
and (n14685,n14686,n14687);
xor (n14686,n10944,n10945);
not (n14687,n14688);
xor (n14688,n12847,n12848);
and (n14689,n14687,n14690);
or (n14690,n6831,n14691);
not (n14691,n6844);
and (n14692,n14686,n14690);
and (n14693,n14680,n14684);
and (n14694,n14674,n14678);
and (n14695,n14668,n14672);
and (n14696,n14662,n14666);
and (n14697,n14656,n14660);
and (n14698,n14650,n14654);
and (n14699,n14644,n14648);
and (n14700,n14638,n14642);
and (n14701,n14632,n14636);
and (n14702,n14626,n14630);
and (n14703,n14620,n14624);
and (n14704,n14614,n14618);
and (n14705,n14608,n14612);
and (n14706,n14602,n14606);
and (n14707,n14596,n14600);
and (n14708,n14590,n14594);
and (n14709,n14584,n14588);
and (n14710,n14578,n14582);
and (n14711,n14572,n14576);
and (n14712,n14566,n14570);
and (n14713,n14560,n14564);
and (n14714,n14554,n14558);
and (n14715,n14548,n14552);
and (n14716,n14542,n14546);
and (n14717,n14536,n14540);
and (n14718,n14530,n14534);
and (n14719,n14524,n14528);
and (n14720,n14518,n14522);
and (n14721,n14512,n14516);
not (n14722,n14723);
xor (n14723,n14724,n18507);
xor (n14724,n14725,n16632);
xor (n14725,n14726,n16079);
xor (n14726,n14727,n16630);
xor (n14727,n14728,n16074);
xor (n14728,n14729,n16623);
xor (n14729,n14730,n16068);
xor (n14730,n14731,n16611);
xor (n14731,n14732,n1107);
xor (n14732,n14733,n16594);
xor (n14733,n14734,n1457);
xor (n14734,n14735,n16572);
xor (n14735,n14736,n16052);
xor (n14736,n14737,n16545);
xor (n14737,n14738,n1797);
xor (n14738,n14739,n16513);
xor (n14739,n14740,n16041);
xor (n14740,n14741,n16476);
xor (n14741,n14742,n16035);
xor (n14742,n14743,n16434);
xor (n14743,n14744,n16029);
xor (n14744,n14745,n16387);
xor (n14745,n14746,n16023);
xor (n14746,n14747,n16335);
xor (n14747,n14748,n16017);
xor (n14748,n14749,n16278);
xor (n14749,n14750,n16011);
xor (n14750,n14751,n16216);
xor (n14751,n14752,n16005);
xor (n14752,n14753,n16149);
xor (n14753,n14754,n15999);
xor (n14754,n14755,n14815);
xor (n14755,n14756,n14813);
xor (n14756,n14757,n14814);
xor (n14757,n14758,n14813);
xor (n14758,n14759,n14812);
xor (n14759,n14760,n14811);
xor (n14760,n14761,n14810);
xor (n14761,n14762,n14809);
xor (n14762,n14763,n14808);
xor (n14763,n14764,n14807);
xor (n14764,n14765,n14806);
xor (n14765,n14766,n14805);
xor (n14766,n14767,n14804);
xor (n14767,n14768,n14803);
xor (n14768,n14769,n14802);
xor (n14769,n14770,n2119);
xor (n14770,n14771,n14801);
xor (n14771,n14772,n14800);
xor (n14772,n14773,n14799);
xor (n14773,n14774,n1947);
xor (n14774,n14775,n14798);
xor (n14775,n14776,n14797);
xor (n14776,n14777,n14796);
xor (n14777,n14778,n14795);
xor (n14778,n14779,n14794);
xor (n14779,n14780,n14793);
xor (n14780,n14781,n14792);
xor (n14781,n14782,n14791);
xor (n14782,n14783,n14790);
xor (n14783,n14784,n14789);
xor (n14784,n14785,n14788);
xor (n14785,n14786,n14787);
and (n14786,n203,n196);
and (n14787,n203,n179);
and (n14788,n14786,n14787);
and (n14789,n203,n180);
and (n14790,n14784,n14789);
and (n14791,n203,n174);
and (n14792,n14782,n14791);
and (n14793,n203,n335);
and (n14794,n14780,n14793);
and (n14795,n203,n37);
and (n14796,n14778,n14795);
and (n14797,n203,n38);
and (n14798,n14776,n14797);
and (n14799,n14774,n1947);
and (n14800,n203,n257);
and (n14801,n14772,n14800);
and (n14802,n14770,n2119);
and (n14803,n203,n368);
and (n14804,n14768,n14803);
and (n14805,n203,n360);
and (n14806,n14766,n14805);
and (n14807,n203,n517);
and (n14808,n14764,n14807);
and (n14809,n203,n76);
and (n14810,n14762,n14809);
and (n14811,n203,n69);
and (n14812,n14760,n14811);
and (n14813,n203,n62);
and (n14814,n14758,n14813);
or (n14815,n14816,n16080);
and (n14816,n14817,n15999);
xor (n14817,n14757,n14818);
or (n14818,n14819,n16000);
and (n14819,n14820,n15999);
xor (n14820,n14759,n14821);
or (n14821,n14822,n15917);
and (n14822,n14823,n15916);
xor (n14823,n14761,n14824);
or (n14824,n14825,n15836);
and (n14825,n14826,n15835);
xor (n14826,n14763,n14827);
or (n14827,n14828,n15753);
and (n14828,n14829,n15752);
xor (n14829,n14765,n14830);
or (n14830,n14831,n15675);
and (n14831,n14832,n15674);
xor (n14832,n14767,n14833);
or (n14833,n14834,n15591);
and (n14834,n14835,n15590);
xor (n14835,n14769,n14836);
or (n14836,n14837,n15513);
and (n14837,n14838,n2032);
xor (n14838,n14771,n14839);
or (n14839,n14840,n15431);
and (n14840,n14841,n15430);
xor (n14841,n14773,n14842);
or (n14842,n14843,n15350);
and (n14843,n14844,n1811);
xor (n14844,n14775,n14845);
or (n14845,n14846,n15268);
and (n14846,n14847,n15267);
xor (n14847,n14777,n14848);
or (n14848,n14849,n15188);
and (n14849,n14850,n15187);
xor (n14850,n14779,n14851);
or (n14851,n14852,n15105);
and (n14852,n14853,n15104);
xor (n14853,n14781,n14854);
or (n14854,n14855,n15025);
and (n14855,n14856,n15024);
xor (n14856,n14783,n14857);
or (n14857,n14858,n14942);
and (n14858,n14859,n14941);
xor (n14859,n14785,n14860);
or (n14860,n14861,n14863);
and (n14861,n14786,n14862);
and (n14862,n192,n179);
and (n14863,n14864,n14865);
xor (n14864,n14786,n14862);
or (n14865,n14866,n14869);
and (n14866,n14867,n14868);
and (n14867,n192,n196);
and (n14868,n173,n179);
and (n14869,n14870,n14871);
xor (n14870,n14867,n14868);
or (n14871,n14872,n14875);
and (n14872,n14873,n14874);
and (n14873,n173,n196);
and (n14874,n496,n179);
and (n14875,n14876,n14877);
xor (n14876,n14873,n14874);
or (n14877,n14878,n14881);
and (n14878,n14879,n14880);
and (n14879,n496,n196);
and (n14880,n490,n179);
and (n14881,n14882,n14883);
xor (n14882,n14879,n14880);
or (n14883,n14884,n14887);
and (n14884,n14885,n14886);
and (n14885,n490,n196);
and (n14886,n43,n179);
and (n14887,n14888,n14889);
xor (n14888,n14885,n14886);
or (n14889,n14890,n14893);
and (n14890,n14891,n14892);
and (n14891,n43,n196);
and (n14892,n53,n179);
and (n14893,n14894,n14895);
xor (n14894,n14891,n14892);
or (n14895,n14896,n14899);
and (n14896,n14897,n14898);
and (n14897,n53,n196);
and (n14898,n223,n179);
and (n14899,n14900,n14901);
xor (n14900,n14897,n14898);
or (n14901,n14902,n14904);
and (n14902,n14903,n2825);
and (n14903,n223,n196);
and (n14904,n14905,n14906);
xor (n14905,n14903,n2825);
or (n14906,n14907,n14910);
and (n14907,n14908,n14909);
and (n14908,n217,n196);
and (n14909,n267,n179);
and (n14910,n14911,n14912);
xor (n14911,n14908,n14909);
or (n14912,n14913,n14915);
and (n14913,n14914,n3021);
and (n14914,n267,n196);
and (n14915,n14916,n14917);
xor (n14916,n14914,n3021);
or (n14917,n14918,n14921);
and (n14918,n14919,n14920);
and (n14919,n249,n196);
and (n14920,n376,n179);
and (n14921,n14922,n14923);
xor (n14922,n14919,n14920);
or (n14923,n14924,n14926);
and (n14924,n14925,n3189);
and (n14925,n376,n196);
and (n14926,n14927,n14928);
xor (n14927,n14925,n3189);
or (n14928,n14929,n14931);
and (n14929,n14930,n3278);
and (n14930,n358,n196);
and (n14931,n14932,n14933);
xor (n14932,n14930,n3278);
or (n14933,n14934,n14936);
and (n14934,n14935,n3293);
and (n14935,n81,n196);
and (n14936,n14937,n14938);
xor (n14937,n14935,n3293);
and (n14938,n14939,n14940);
and (n14939,n63,n196);
and (n14940,n452,n179);
and (n14941,n192,n180);
and (n14942,n14943,n14944);
xor (n14943,n14859,n14941);
or (n14944,n14945,n14948);
and (n14945,n14946,n14947);
xor (n14946,n14864,n14865);
and (n14947,n173,n180);
and (n14948,n14949,n14950);
xor (n14949,n14946,n14947);
or (n14950,n14951,n14954);
and (n14951,n14952,n14953);
xor (n14952,n14870,n14871);
and (n14953,n496,n180);
and (n14954,n14955,n14956);
xor (n14955,n14952,n14953);
or (n14956,n14957,n14960);
and (n14957,n14958,n14959);
xor (n14958,n14876,n14877);
and (n14959,n490,n180);
and (n14960,n14961,n14962);
xor (n14961,n14958,n14959);
or (n14962,n14963,n14966);
and (n14963,n14964,n14965);
xor (n14964,n14882,n14883);
and (n14965,n43,n180);
and (n14966,n14967,n14968);
xor (n14967,n14964,n14965);
or (n14968,n14969,n14972);
and (n14969,n14970,n14971);
xor (n14970,n14888,n14889);
and (n14971,n53,n180);
and (n14972,n14973,n14974);
xor (n14973,n14970,n14971);
or (n14974,n14975,n14978);
and (n14975,n14976,n14977);
xor (n14976,n14894,n14895);
and (n14977,n223,n180);
and (n14978,n14979,n14980);
xor (n14979,n14976,n14977);
or (n14980,n14981,n14984);
and (n14981,n14982,n14983);
xor (n14982,n14900,n14901);
and (n14983,n217,n180);
and (n14984,n14985,n14986);
xor (n14985,n14982,n14983);
or (n14986,n14987,n14990);
and (n14987,n14988,n14989);
xor (n14988,n14905,n14906);
and (n14989,n267,n180);
and (n14990,n14991,n14992);
xor (n14991,n14988,n14989);
or (n14992,n14993,n14996);
and (n14993,n14994,n14995);
xor (n14994,n14911,n14912);
and (n14995,n249,n180);
and (n14996,n14997,n14998);
xor (n14997,n14994,n14995);
or (n14998,n14999,n15002);
and (n14999,n15000,n15001);
xor (n15000,n14916,n14917);
and (n15001,n376,n180);
and (n15002,n15003,n15004);
xor (n15003,n15000,n15001);
or (n15004,n15005,n15008);
and (n15005,n15006,n15007);
xor (n15006,n14922,n14923);
and (n15007,n358,n180);
and (n15008,n15009,n15010);
xor (n15009,n15006,n15007);
or (n15010,n15011,n15014);
and (n15011,n15012,n15013);
xor (n15012,n14927,n14928);
and (n15013,n81,n180);
and (n15014,n15015,n15016);
xor (n15015,n15012,n15013);
or (n15016,n15017,n15020);
and (n15017,n15018,n15019);
xor (n15018,n14932,n14933);
and (n15019,n63,n180);
and (n15020,n15021,n15022);
xor (n15021,n15018,n15019);
and (n15022,n15023,n3198);
xor (n15023,n14937,n14938);
and (n15024,n192,n174);
and (n15025,n15026,n15027);
xor (n15026,n14856,n15024);
or (n15027,n15028,n15031);
and (n15028,n15029,n15030);
xor (n15029,n14943,n14944);
and (n15030,n173,n174);
and (n15031,n15032,n15033);
xor (n15032,n15029,n15030);
or (n15033,n15034,n15037);
and (n15034,n15035,n15036);
xor (n15035,n14949,n14950);
and (n15036,n496,n174);
and (n15037,n15038,n15039);
xor (n15038,n15035,n15036);
or (n15039,n15040,n15043);
and (n15040,n15041,n15042);
xor (n15041,n14955,n14956);
and (n15042,n490,n174);
and (n15043,n15044,n15045);
xor (n15044,n15041,n15042);
or (n15045,n15046,n15049);
and (n15046,n15047,n15048);
xor (n15047,n14961,n14962);
and (n15048,n43,n174);
and (n15049,n15050,n15051);
xor (n15050,n15047,n15048);
or (n15051,n15052,n15055);
and (n15052,n15053,n15054);
xor (n15053,n14967,n14968);
and (n15054,n53,n174);
and (n15055,n15056,n15057);
xor (n15056,n15053,n15054);
or (n15057,n15058,n15060);
and (n15058,n15059,n1366);
xor (n15059,n14973,n14974);
and (n15060,n15061,n15062);
xor (n15061,n15059,n1366);
or (n15062,n15063,n15065);
and (n15063,n15064,n2569);
xor (n15064,n14979,n14980);
and (n15065,n15066,n15067);
xor (n15066,n15064,n2569);
or (n15067,n15068,n15071);
and (n15068,n15069,n15070);
xor (n15069,n14985,n14986);
and (n15070,n267,n174);
and (n15071,n15072,n15073);
xor (n15072,n15069,n15070);
or (n15073,n15074,n15076);
and (n15074,n15075,n2833);
xor (n15075,n14991,n14992);
and (n15076,n15077,n15078);
xor (n15077,n15075,n2833);
or (n15078,n15079,n15082);
and (n15079,n15080,n15081);
xor (n15080,n14997,n14998);
and (n15081,n376,n174);
and (n15082,n15083,n15084);
xor (n15083,n15080,n15081);
or (n15084,n15085,n15088);
and (n15085,n15086,n15087);
xor (n15086,n15003,n15004);
and (n15087,n358,n174);
and (n15088,n15089,n15090);
xor (n15089,n15086,n15087);
or (n15090,n15091,n15094);
and (n15091,n15092,n15093);
xor (n15092,n15009,n15010);
and (n15093,n81,n174);
and (n15094,n15095,n15096);
xor (n15095,n15092,n15093);
or (n15096,n15097,n15100);
and (n15097,n15098,n15099);
xor (n15098,n15015,n15016);
and (n15099,n63,n174);
and (n15100,n15101,n15102);
xor (n15101,n15098,n15099);
and (n15102,n15103,n3244);
xor (n15103,n15021,n15022);
and (n15104,n192,n335);
and (n15105,n15106,n15107);
xor (n15106,n14853,n15104);
or (n15107,n15108,n15111);
and (n15108,n15109,n15110);
xor (n15109,n15026,n15027);
and (n15110,n173,n335);
and (n15111,n15112,n15113);
xor (n15112,n15109,n15110);
or (n15113,n15114,n15117);
and (n15114,n15115,n15116);
xor (n15115,n15032,n15033);
and (n15116,n496,n335);
and (n15117,n15118,n15119);
xor (n15118,n15115,n15116);
or (n15119,n15120,n15123);
and (n15120,n15121,n15122);
xor (n15121,n15038,n15039);
and (n15122,n490,n335);
and (n15123,n15124,n15125);
xor (n15124,n15121,n15122);
or (n15125,n15126,n15129);
and (n15126,n15127,n15128);
xor (n15127,n15044,n15045);
and (n15128,n43,n335);
and (n15129,n15130,n15131);
xor (n15130,n15127,n15128);
or (n15131,n15132,n15135);
and (n15132,n15133,n15134);
xor (n15133,n15050,n15051);
and (n15134,n53,n335);
and (n15135,n15136,n15137);
xor (n15136,n15133,n15134);
or (n15137,n15138,n15141);
and (n15138,n15139,n15140);
xor (n15139,n15056,n15057);
and (n15140,n223,n335);
and (n15141,n15142,n15143);
xor (n15142,n15139,n15140);
or (n15143,n15144,n15147);
and (n15144,n15145,n15146);
xor (n15145,n15061,n15062);
and (n15146,n217,n335);
and (n15147,n15148,n15149);
xor (n15148,n15145,n15146);
or (n15149,n15150,n15153);
and (n15150,n15151,n15152);
xor (n15151,n15066,n15067);
and (n15152,n267,n335);
and (n15153,n15154,n15155);
xor (n15154,n15151,n15152);
or (n15155,n15156,n15159);
and (n15156,n15157,n15158);
xor (n15157,n15072,n15073);
and (n15158,n249,n335);
and (n15159,n15160,n15161);
xor (n15160,n15157,n15158);
or (n15161,n15162,n15165);
and (n15162,n15163,n15164);
xor (n15163,n15077,n15078);
and (n15164,n376,n335);
and (n15165,n15166,n15167);
xor (n15166,n15163,n15164);
or (n15167,n15168,n15171);
and (n15168,n15169,n15170);
xor (n15169,n15083,n15084);
and (n15170,n358,n335);
and (n15171,n15172,n15173);
xor (n15172,n15169,n15170);
or (n15173,n15174,n15177);
and (n15174,n15175,n15176);
xor (n15175,n15089,n15090);
and (n15176,n81,n335);
and (n15177,n15178,n15179);
xor (n15178,n15175,n15176);
or (n15179,n15180,n15183);
and (n15180,n15181,n15182);
xor (n15181,n15095,n15096);
and (n15182,n63,n335);
and (n15183,n15184,n15185);
xor (n15184,n15181,n15182);
and (n15185,n15186,n3124);
xor (n15186,n15101,n15102);
and (n15187,n192,n37);
and (n15188,n15189,n15190);
xor (n15189,n14850,n15187);
or (n15190,n15191,n15194);
and (n15191,n15192,n15193);
xor (n15192,n15106,n15107);
and (n15193,n173,n37);
and (n15194,n15195,n15196);
xor (n15195,n15192,n15193);
or (n15196,n15197,n15200);
and (n15197,n15198,n15199);
xor (n15198,n15112,n15113);
and (n15199,n496,n37);
and (n15200,n15201,n15202);
xor (n15201,n15198,n15199);
or (n15202,n15203,n15206);
and (n15203,n15204,n15205);
xor (n15204,n15118,n15119);
and (n15205,n490,n37);
and (n15206,n15207,n15208);
xor (n15207,n15204,n15205);
or (n15208,n15209,n15212);
and (n15209,n15210,n15211);
xor (n15210,n15124,n15125);
and (n15211,n43,n37);
and (n15212,n15213,n15214);
xor (n15213,n15210,n15211);
or (n15214,n15215,n15218);
and (n15215,n15216,n15217);
xor (n15216,n15130,n15131);
and (n15217,n53,n37);
and (n15218,n15219,n15220);
xor (n15219,n15216,n15217);
or (n15220,n15221,n15224);
and (n15221,n15222,n15223);
xor (n15222,n15136,n15137);
and (n15223,n223,n37);
and (n15224,n15225,n15226);
xor (n15225,n15222,n15223);
or (n15226,n15227,n15229);
and (n15227,n15228,n1242);
xor (n15228,n15142,n15143);
and (n15229,n15230,n15231);
xor (n15230,n15228,n1242);
or (n15231,n15232,n15235);
and (n15232,n15233,n15234);
xor (n15233,n15148,n15149);
and (n15234,n267,n37);
and (n15235,n15236,n15237);
xor (n15236,n15233,n15234);
or (n15237,n15238,n15240);
and (n15238,n15239,n2670);
xor (n15239,n15154,n15155);
and (n15240,n15241,n15242);
xor (n15241,n15239,n2670);
or (n15242,n15243,n15245);
and (n15243,n15244,n2694);
xor (n15244,n15160,n15161);
and (n15245,n15246,n15247);
xor (n15246,n15244,n2694);
or (n15247,n15248,n15251);
and (n15248,n15249,n15250);
xor (n15249,n15166,n15167);
and (n15250,n358,n37);
and (n15251,n15252,n15253);
xor (n15252,n15249,n15250);
or (n15253,n15254,n15257);
and (n15254,n15255,n15256);
xor (n15255,n15172,n15173);
and (n15256,n81,n37);
and (n15257,n15258,n15259);
xor (n15258,n15255,n15256);
or (n15259,n15260,n15262);
and (n15260,n15261,n3055);
xor (n15261,n15178,n15179);
and (n15262,n15263,n15264);
xor (n15263,n15261,n3055);
and (n15264,n15265,n15266);
xor (n15265,n15184,n15185);
and (n15266,n452,n37);
and (n15267,n192,n38);
and (n15268,n15269,n15270);
xor (n15269,n14847,n15267);
or (n15270,n15271,n15274);
and (n15271,n15272,n15273);
xor (n15272,n15189,n15190);
and (n15273,n173,n38);
and (n15274,n15275,n15276);
xor (n15275,n15272,n15273);
or (n15276,n15277,n15280);
and (n15277,n15278,n15279);
xor (n15278,n15195,n15196);
and (n15279,n496,n38);
and (n15280,n15281,n15282);
xor (n15281,n15278,n15279);
or (n15282,n15283,n15286);
and (n15283,n15284,n15285);
xor (n15284,n15201,n15202);
and (n15285,n490,n38);
and (n15286,n15287,n15288);
xor (n15287,n15284,n15285);
or (n15288,n15289,n15292);
and (n15289,n15290,n15291);
xor (n15290,n15207,n15208);
and (n15291,n43,n38);
and (n15292,n15293,n15294);
xor (n15293,n15290,n15291);
or (n15294,n15295,n15298);
and (n15295,n15296,n15297);
xor (n15296,n15213,n15214);
and (n15297,n53,n38);
and (n15298,n15299,n15300);
xor (n15299,n15296,n15297);
or (n15300,n15301,n15304);
and (n15301,n15302,n15303);
xor (n15302,n15219,n15220);
and (n15303,n223,n38);
and (n15304,n15305,n15306);
xor (n15305,n15302,n15303);
or (n15306,n15307,n15310);
and (n15307,n15308,n15309);
xor (n15308,n15225,n15226);
and (n15309,n217,n38);
and (n15310,n15311,n15312);
xor (n15311,n15308,n15309);
or (n15312,n15313,n15316);
and (n15313,n15314,n15315);
xor (n15314,n15230,n15231);
and (n15315,n267,n38);
and (n15316,n15317,n15318);
xor (n15317,n15314,n15315);
or (n15318,n15319,n15322);
and (n15319,n15320,n15321);
xor (n15320,n15236,n15237);
and (n15321,n249,n38);
and (n15322,n15323,n15324);
xor (n15323,n15320,n15321);
or (n15324,n15325,n15328);
and (n15325,n15326,n15327);
xor (n15326,n15241,n15242);
and (n15327,n376,n38);
and (n15328,n15329,n15330);
xor (n15329,n15326,n15327);
or (n15330,n15331,n15334);
and (n15331,n15332,n15333);
xor (n15332,n15246,n15247);
and (n15333,n358,n38);
and (n15334,n15335,n15336);
xor (n15335,n15332,n15333);
or (n15336,n15337,n15340);
and (n15337,n15338,n15339);
xor (n15338,n15252,n15253);
and (n15339,n81,n38);
and (n15340,n15341,n15342);
xor (n15341,n15338,n15339);
or (n15342,n15343,n15346);
and (n15343,n15344,n15345);
xor (n15344,n15258,n15259);
and (n15345,n63,n38);
and (n15346,n15347,n15348);
xor (n15347,n15344,n15345);
and (n15348,n15349,n2947);
xor (n15349,n15263,n15264);
and (n15350,n15351,n15352);
xor (n15351,n14844,n1811);
or (n15352,n15353,n15356);
and (n15353,n15354,n15355);
xor (n15354,n15269,n15270);
and (n15355,n173,n45);
and (n15356,n15357,n15358);
xor (n15357,n15354,n15355);
or (n15358,n15359,n15362);
and (n15359,n15360,n15361);
xor (n15360,n15275,n15276);
and (n15361,n496,n45);
and (n15362,n15363,n15364);
xor (n15363,n15360,n15361);
or (n15364,n15365,n15368);
and (n15365,n15366,n15367);
xor (n15366,n15281,n15282);
and (n15367,n490,n45);
and (n15368,n15369,n15370);
xor (n15369,n15366,n15367);
or (n15370,n15371,n15374);
and (n15371,n15372,n15373);
xor (n15372,n15287,n15288);
and (n15373,n43,n45);
and (n15374,n15375,n15376);
xor (n15375,n15372,n15373);
or (n15376,n15377,n15379);
and (n15377,n15378,n52);
xor (n15378,n15293,n15294);
and (n15379,n15380,n15381);
xor (n15380,n15378,n52);
or (n15381,n15382,n15385);
and (n15382,n15383,n15384);
xor (n15383,n15299,n15300);
and (n15384,n223,n45);
and (n15385,n15386,n15387);
xor (n15386,n15383,n15384);
or (n15387,n15388,n15391);
and (n15388,n15389,n15390);
xor (n15389,n15305,n15306);
and (n15390,n217,n45);
and (n15391,n15392,n15393);
xor (n15392,n15389,n15390);
or (n15393,n15394,n15397);
and (n15394,n15395,n15396);
xor (n15395,n15311,n15312);
and (n15396,n267,n45);
and (n15397,n15398,n15399);
xor (n15398,n15395,n15396);
or (n15399,n15400,n15403);
and (n15400,n15401,n15402);
xor (n15401,n15317,n15318);
and (n15402,n249,n45);
and (n15403,n15404,n15405);
xor (n15404,n15401,n15402);
or (n15405,n15406,n15409);
and (n15406,n15407,n15408);
xor (n15407,n15323,n15324);
and (n15408,n376,n45);
and (n15409,n15410,n15411);
xor (n15410,n15407,n15408);
or (n15411,n15412,n15414);
and (n15412,n15413,n2577);
xor (n15413,n15329,n15330);
and (n15414,n15415,n15416);
xor (n15415,n15413,n2577);
or (n15416,n15417,n15420);
and (n15417,n15418,n15419);
xor (n15418,n15335,n15336);
and (n15419,n81,n45);
and (n15420,n15421,n15422);
xor (n15421,n15418,n15419);
or (n15422,n15423,n15426);
and (n15423,n15424,n15425);
xor (n15424,n15341,n15342);
and (n15425,n63,n45);
and (n15426,n15427,n15428);
xor (n15427,n15424,n15425);
and (n15428,n15429,n2960);
xor (n15429,n15347,n15348);
and (n15430,n192,n257);
and (n15431,n15432,n15433);
xor (n15432,n14841,n15430);
or (n15433,n15434,n15437);
and (n15434,n15435,n15436);
xor (n15435,n15351,n15352);
and (n15436,n173,n257);
and (n15437,n15438,n15439);
xor (n15438,n15435,n15436);
or (n15439,n15440,n15443);
and (n15440,n15441,n15442);
xor (n15441,n15357,n15358);
and (n15442,n496,n257);
and (n15443,n15444,n15445);
xor (n15444,n15441,n15442);
or (n15445,n15446,n15449);
and (n15446,n15447,n15448);
xor (n15447,n15363,n15364);
and (n15448,n490,n257);
and (n15449,n15450,n15451);
xor (n15450,n15447,n15448);
or (n15451,n15452,n15455);
and (n15452,n15453,n15454);
xor (n15453,n15369,n15370);
and (n15454,n43,n257);
and (n15455,n15456,n15457);
xor (n15456,n15453,n15454);
or (n15457,n15458,n15461);
and (n15458,n15459,n15460);
xor (n15459,n15375,n15376);
and (n15460,n53,n257);
and (n15461,n15462,n15463);
xor (n15462,n15459,n15460);
or (n15463,n15464,n15467);
and (n15464,n15465,n15466);
xor (n15465,n15380,n15381);
and (n15466,n223,n257);
and (n15467,n15468,n15469);
xor (n15468,n15465,n15466);
or (n15469,n15470,n15473);
and (n15470,n15471,n15472);
xor (n15471,n15386,n15387);
and (n15472,n217,n257);
and (n15473,n15474,n15475);
xor (n15474,n15471,n15472);
or (n15475,n15476,n15479);
and (n15476,n15477,n15478);
xor (n15477,n15392,n15393);
and (n15478,n267,n257);
and (n15479,n15480,n15481);
xor (n15480,n15477,n15478);
or (n15481,n15482,n15485);
and (n15482,n15483,n15484);
xor (n15483,n15398,n15399);
and (n15484,n249,n257);
and (n15485,n15486,n15487);
xor (n15486,n15483,n15484);
or (n15487,n15488,n15491);
and (n15488,n15489,n15490);
xor (n15489,n15404,n15405);
and (n15490,n376,n257);
and (n15491,n15492,n15493);
xor (n15492,n15489,n15490);
or (n15493,n15494,n15497);
and (n15494,n15495,n15496);
xor (n15495,n15410,n15411);
and (n15496,n358,n257);
and (n15497,n15498,n15499);
xor (n15498,n15495,n15496);
or (n15499,n15500,n15503);
and (n15500,n15501,n15502);
xor (n15501,n15415,n15416);
and (n15502,n81,n257);
and (n15503,n15504,n15505);
xor (n15504,n15501,n15502);
or (n15505,n15506,n15509);
and (n15506,n15507,n15508);
xor (n15507,n15421,n15422);
and (n15508,n63,n257);
and (n15509,n15510,n15511);
xor (n15510,n15507,n15508);
and (n15511,n15512,n2739);
xor (n15512,n15427,n15428);
and (n15513,n15514,n15515);
xor (n15514,n14838,n2032);
or (n15515,n15516,n15518);
and (n15516,n15517,n1953);
xor (n15517,n15432,n15433);
and (n15518,n15519,n15520);
xor (n15519,n15517,n1953);
or (n15520,n15521,n15523);
and (n15521,n15522,n1735);
xor (n15522,n15438,n15439);
and (n15523,n15524,n15525);
xor (n15524,n15522,n1735);
or (n15525,n15526,n15528);
and (n15526,n15527,n1621);
xor (n15527,n15444,n15445);
and (n15528,n15529,n15530);
xor (n15529,n15527,n1621);
or (n15530,n15531,n15534);
and (n15531,n15532,n15533);
xor (n15532,n15450,n15451);
and (n15533,n43,n251);
and (n15534,n15535,n15536);
xor (n15535,n15532,n15533);
or (n15536,n15537,n15540);
and (n15537,n15538,n15539);
xor (n15538,n15456,n15457);
and (n15539,n53,n251);
and (n15540,n15541,n15542);
xor (n15541,n15538,n15539);
or (n15542,n15543,n15546);
and (n15543,n15544,n15545);
xor (n15544,n15462,n15463);
and (n15545,n223,n251);
and (n15546,n15547,n15548);
xor (n15547,n15544,n15545);
or (n15548,n15549,n15552);
and (n15549,n15550,n15551);
xor (n15550,n15468,n15469);
and (n15551,n217,n251);
and (n15552,n15553,n15554);
xor (n15553,n15550,n15551);
or (n15554,n15555,n15558);
and (n15555,n15556,n15557);
xor (n15556,n15474,n15475);
and (n15557,n267,n251);
and (n15558,n15559,n15560);
xor (n15559,n15556,n15557);
or (n15560,n15561,n15563);
and (n15561,n15562,n252);
xor (n15562,n15480,n15481);
and (n15563,n15564,n15565);
xor (n15564,n15562,n252);
or (n15565,n15566,n15569);
and (n15566,n15567,n15568);
xor (n15567,n15486,n15487);
and (n15568,n376,n251);
and (n15569,n15570,n15571);
xor (n15570,n15567,n15568);
or (n15571,n15572,n15574);
and (n15572,n15573,n840);
xor (n15573,n15492,n15493);
and (n15574,n15575,n15576);
xor (n15575,n15573,n840);
or (n15576,n15577,n15579);
and (n15577,n15578,n1280);
xor (n15578,n15498,n15499);
and (n15579,n15580,n15581);
xor (n15580,n15578,n1280);
or (n15581,n15582,n15585);
and (n15582,n15583,n15584);
xor (n15583,n15504,n15505);
and (n15584,n63,n251);
and (n15585,n15586,n15587);
xor (n15586,n15583,n15584);
and (n15587,n15588,n15589);
xor (n15588,n15510,n15511);
and (n15589,n452,n251);
and (n15590,n192,n368);
and (n15591,n15592,n15593);
xor (n15592,n14835,n15590);
or (n15593,n15594,n15597);
and (n15594,n15595,n15596);
xor (n15595,n15514,n15515);
and (n15596,n173,n368);
and (n15597,n15598,n15599);
xor (n15598,n15595,n15596);
or (n15599,n15600,n15603);
and (n15600,n15601,n15602);
xor (n15601,n15519,n15520);
and (n15602,n496,n368);
and (n15603,n15604,n15605);
xor (n15604,n15601,n15602);
or (n15605,n15606,n15609);
and (n15606,n15607,n15608);
xor (n15607,n15524,n15525);
and (n15608,n490,n368);
and (n15609,n15610,n15611);
xor (n15610,n15607,n15608);
or (n15611,n15612,n15615);
and (n15612,n15613,n15614);
xor (n15613,n15529,n15530);
and (n15614,n43,n368);
and (n15615,n15616,n15617);
xor (n15616,n15613,n15614);
or (n15617,n15618,n15621);
and (n15618,n15619,n15620);
xor (n15619,n15535,n15536);
and (n15620,n53,n368);
and (n15621,n15622,n15623);
xor (n15622,n15619,n15620);
or (n15623,n15624,n15627);
and (n15624,n15625,n15626);
xor (n15625,n15541,n15542);
and (n15626,n223,n368);
and (n15627,n15628,n15629);
xor (n15628,n15625,n15626);
or (n15629,n15630,n15633);
and (n15630,n15631,n15632);
xor (n15631,n15547,n15548);
and (n15632,n217,n368);
and (n15633,n15634,n15635);
xor (n15634,n15631,n15632);
or (n15635,n15636,n15639);
and (n15636,n15637,n15638);
xor (n15637,n15553,n15554);
and (n15638,n267,n368);
and (n15639,n15640,n15641);
xor (n15640,n15637,n15638);
or (n15641,n15642,n15645);
and (n15642,n15643,n15644);
xor (n15643,n15559,n15560);
and (n15644,n249,n368);
and (n15645,n15646,n15647);
xor (n15646,n15643,n15644);
or (n15647,n15648,n15651);
and (n15648,n15649,n15650);
xor (n15649,n15564,n15565);
and (n15650,n376,n368);
and (n15651,n15652,n15653);
xor (n15652,n15649,n15650);
or (n15653,n15654,n15657);
and (n15654,n15655,n15656);
xor (n15655,n15570,n15571);
and (n15656,n358,n368);
and (n15657,n15658,n15659);
xor (n15658,n15655,n15656);
or (n15659,n15660,n15663);
and (n15660,n15661,n15662);
xor (n15661,n15575,n15576);
and (n15662,n81,n368);
and (n15663,n15664,n15665);
xor (n15664,n15661,n15662);
or (n15665,n15666,n15669);
and (n15666,n15667,n15668);
xor (n15667,n15580,n15581);
and (n15668,n63,n368);
and (n15669,n15670,n15671);
xor (n15670,n15667,n15668);
and (n15671,n15672,n15673);
xor (n15672,n15586,n15587);
not (n15673,n1355);
and (n15674,n192,n360);
and (n15675,n15676,n15677);
xor (n15676,n14832,n15674);
or (n15677,n15678,n15680);
and (n15678,n15679,n2125);
xor (n15679,n15592,n15593);
and (n15680,n15681,n15682);
xor (n15681,n15679,n2125);
or (n15682,n15683,n15686);
and (n15683,n15684,n15685);
xor (n15684,n15598,n15599);
and (n15685,n496,n360);
and (n15686,n15687,n15688);
xor (n15687,n15684,n15685);
or (n15688,n15689,n15691);
and (n15689,n15690,n1932);
xor (n15690,n15604,n15605);
and (n15691,n15692,n15693);
xor (n15692,n15690,n1932);
or (n15693,n15694,n15697);
and (n15694,n15695,n15696);
xor (n15695,n15610,n15611);
and (n15696,n43,n360);
and (n15697,n15698,n15699);
xor (n15698,n15695,n15696);
or (n15699,n15700,n15703);
and (n15700,n15701,n15702);
xor (n15701,n15616,n15617);
and (n15702,n53,n360);
and (n15703,n15704,n15705);
xor (n15704,n15701,n15702);
or (n15705,n15706,n15708);
and (n15706,n15707,n1433);
xor (n15707,n15622,n15623);
and (n15708,n15709,n15710);
xor (n15709,n15707,n1433);
or (n15710,n15711,n15713);
and (n15711,n15712,n1079);
xor (n15712,n15628,n15629);
and (n15713,n15714,n15715);
xor (n15714,n15712,n1079);
or (n15715,n15716,n15719);
and (n15716,n15717,n15718);
xor (n15717,n15634,n15635);
and (n15718,n267,n360);
and (n15719,n15720,n15721);
xor (n15720,n15717,n15718);
or (n15721,n15722,n15725);
and (n15722,n15723,n15724);
xor (n15723,n15640,n15641);
and (n15724,n249,n360);
and (n15725,n15726,n15727);
xor (n15726,n15723,n15724);
or (n15727,n15728,n15731);
and (n15728,n15729,n15730);
xor (n15729,n15646,n15647);
and (n15730,n376,n360);
and (n15731,n15732,n15733);
xor (n15732,n15729,n15730);
or (n15733,n15734,n15737);
and (n15734,n15735,n15736);
xor (n15735,n15652,n15653);
and (n15736,n358,n360);
and (n15737,n15738,n15739);
xor (n15738,n15735,n15736);
or (n15739,n15740,n15742);
and (n15740,n15741,n879);
xor (n15741,n15658,n15659);
and (n15742,n15743,n15744);
xor (n15743,n15741,n879);
or (n15744,n15745,n15748);
and (n15745,n15746,n15747);
xor (n15746,n15664,n15665);
and (n15747,n63,n360);
and (n15748,n15749,n15750);
xor (n15749,n15746,n15747);
and (n15750,n15751,n1310);
xor (n15751,n15670,n15671);
and (n15752,n192,n517);
and (n15753,n15754,n15755);
xor (n15754,n14829,n15752);
or (n15755,n15756,n15759);
and (n15756,n15757,n15758);
xor (n15757,n15676,n15677);
and (n15758,n173,n517);
and (n15759,n15760,n15761);
xor (n15760,n15757,n15758);
or (n15761,n15762,n15765);
and (n15762,n15763,n15764);
xor (n15763,n15681,n15682);
and (n15764,n496,n517);
and (n15765,n15766,n15767);
xor (n15766,n15763,n15764);
or (n15767,n15768,n15771);
and (n15768,n15769,n15770);
xor (n15769,n15687,n15688);
and (n15770,n490,n517);
and (n15771,n15772,n15773);
xor (n15772,n15769,n15770);
or (n15773,n15774,n15777);
and (n15774,n15775,n15776);
xor (n15775,n15692,n15693);
and (n15776,n43,n517);
and (n15777,n15778,n15779);
xor (n15778,n15775,n15776);
or (n15779,n15780,n15783);
and (n15780,n15781,n15782);
xor (n15781,n15698,n15699);
and (n15782,n53,n517);
and (n15783,n15784,n15785);
xor (n15784,n15781,n15782);
or (n15785,n15786,n15789);
and (n15786,n15787,n15788);
xor (n15787,n15704,n15705);
and (n15788,n223,n517);
and (n15789,n15790,n15791);
xor (n15790,n15787,n15788);
or (n15791,n15792,n15795);
and (n15792,n15793,n15794);
xor (n15793,n15709,n15710);
and (n15794,n217,n517);
and (n15795,n15796,n15797);
xor (n15796,n15793,n15794);
or (n15797,n15798,n15801);
and (n15798,n15799,n15800);
xor (n15799,n15714,n15715);
and (n15800,n267,n517);
and (n15801,n15802,n15803);
xor (n15802,n15799,n15800);
or (n15803,n15804,n15807);
and (n15804,n15805,n15806);
xor (n15805,n15720,n15721);
and (n15806,n249,n517);
and (n15807,n15808,n15809);
xor (n15808,n15805,n15806);
or (n15809,n15810,n15813);
and (n15810,n15811,n15812);
xor (n15811,n15726,n15727);
and (n15812,n376,n517);
and (n15813,n15814,n15815);
xor (n15814,n15811,n15812);
or (n15815,n15816,n15819);
and (n15816,n15817,n15818);
xor (n15817,n15732,n15733);
and (n15818,n358,n517);
and (n15819,n15820,n15821);
xor (n15820,n15817,n15818);
or (n15821,n15822,n15825);
and (n15822,n15823,n15824);
xor (n15823,n15738,n15739);
and (n15824,n81,n517);
and (n15825,n15826,n15827);
xor (n15826,n15823,n15824);
or (n15827,n15828,n15831);
and (n15828,n15829,n15830);
xor (n15829,n15743,n15744);
and (n15830,n63,n517);
and (n15831,n15832,n15833);
xor (n15832,n15829,n15830);
and (n15833,n15834,n915);
xor (n15834,n15749,n15750);
and (n15835,n192,n76);
and (n15836,n15837,n15838);
xor (n15837,n14826,n15835);
or (n15838,n15839,n15842);
and (n15839,n15840,n15841);
xor (n15840,n15754,n15755);
and (n15841,n173,n76);
and (n15842,n15843,n15844);
xor (n15843,n15840,n15841);
or (n15844,n15845,n15848);
and (n15845,n15846,n15847);
xor (n15846,n15760,n15761);
and (n15847,n496,n76);
and (n15848,n15849,n15850);
xor (n15849,n15846,n15847);
or (n15850,n15851,n15854);
and (n15851,n15852,n15853);
xor (n15852,n15766,n15767);
and (n15853,n490,n76);
and (n15854,n15855,n15856);
xor (n15855,n15852,n15853);
or (n15856,n15857,n15859);
and (n15857,n15858,n2009);
xor (n15858,n15772,n15773);
and (n15859,n15860,n15861);
xor (n15860,n15858,n2009);
or (n15861,n15862,n15865);
and (n15862,n15863,n15864);
xor (n15863,n15778,n15779);
and (n15864,n53,n76);
and (n15865,n15866,n15867);
xor (n15866,n15863,n15864);
or (n15867,n15868,n15870);
and (n15868,n15869,n1774);
xor (n15869,n15784,n15785);
and (n15870,n15871,n15872);
xor (n15871,n15869,n1774);
or (n15872,n15873,n15876);
and (n15873,n15874,n15875);
xor (n15874,n15790,n15791);
and (n15875,n217,n76);
and (n15876,n15877,n15878);
xor (n15877,n15874,n15875);
or (n15878,n15879,n15882);
and (n15879,n15880,n15881);
xor (n15880,n15796,n15797);
and (n15881,n267,n76);
and (n15882,n15883,n15884);
xor (n15883,n15880,n15881);
or (n15884,n15885,n15888);
and (n15885,n15886,n15887);
xor (n15886,n15802,n15803);
and (n15887,n249,n76);
and (n15888,n15889,n15890);
xor (n15889,n15886,n15887);
or (n15890,n15891,n15894);
and (n15891,n15892,n15893);
xor (n15892,n15808,n15809);
and (n15893,n376,n76);
and (n15894,n15895,n15896);
xor (n15895,n15892,n15893);
or (n15896,n15897,n15900);
and (n15897,n15898,n15899);
xor (n15898,n15814,n15815);
and (n15899,n358,n76);
and (n15900,n15901,n15902);
xor (n15901,n15898,n15899);
or (n15902,n15903,n15906);
and (n15903,n15904,n15905);
xor (n15904,n15820,n15821);
and (n15905,n81,n76);
and (n15906,n15907,n15908);
xor (n15907,n15904,n15905);
or (n15908,n15909,n15911);
and (n15909,n15910,n663);
xor (n15910,n15826,n15827);
and (n15911,n15912,n15913);
xor (n15912,n15910,n663);
and (n15913,n15914,n15915);
xor (n15914,n15832,n15833);
and (n15915,n452,n76);
and (n15916,n192,n69);
and (n15917,n15918,n15919);
xor (n15918,n14823,n15916);
or (n15919,n15920,n15923);
and (n15920,n15921,n15922);
xor (n15921,n15837,n15838);
and (n15922,n173,n69);
and (n15923,n15924,n15925);
xor (n15924,n15921,n15922);
or (n15925,n15926,n15929);
and (n15926,n15927,n15928);
xor (n15927,n15843,n15844);
and (n15928,n496,n69);
and (n15929,n15930,n15931);
xor (n15930,n15927,n15928);
or (n15931,n15932,n15935);
and (n15932,n15933,n15934);
xor (n15933,n15849,n15850);
and (n15934,n490,n69);
and (n15935,n15936,n15937);
xor (n15936,n15933,n15934);
or (n15937,n15938,n15941);
and (n15938,n15939,n15940);
xor (n15939,n15855,n15856);
and (n15940,n43,n69);
and (n15941,n15942,n15943);
xor (n15942,n15939,n15940);
or (n15943,n15944,n15947);
and (n15944,n15945,n15946);
xor (n15945,n15860,n15861);
and (n15946,n53,n69);
and (n15947,n15948,n15949);
xor (n15948,n15945,n15946);
or (n15949,n15950,n15953);
and (n15950,n15951,n15952);
xor (n15951,n15866,n15867);
and (n15952,n223,n69);
and (n15953,n15954,n15955);
xor (n15954,n15951,n15952);
or (n15955,n15956,n15959);
and (n15956,n15957,n15958);
xor (n15957,n15871,n15872);
and (n15958,n217,n69);
and (n15959,n15960,n15961);
xor (n15960,n15957,n15958);
or (n15961,n15962,n15965);
and (n15962,n15963,n15964);
xor (n15963,n15877,n15878);
and (n15964,n267,n69);
and (n15965,n15966,n15967);
xor (n15966,n15963,n15964);
or (n15967,n15968,n15971);
and (n15968,n15969,n15970);
xor (n15969,n15883,n15884);
and (n15970,n249,n69);
and (n15971,n15972,n15973);
xor (n15972,n15969,n15970);
or (n15973,n15974,n15977);
and (n15974,n15975,n15976);
xor (n15975,n15889,n15890);
and (n15976,n376,n69);
and (n15977,n15978,n15979);
xor (n15978,n15975,n15976);
or (n15979,n15980,n15983);
and (n15980,n15981,n15982);
xor (n15981,n15895,n15896);
and (n15982,n358,n69);
and (n15983,n15984,n15985);
xor (n15984,n15981,n15982);
or (n15985,n15986,n15989);
and (n15986,n15987,n15988);
xor (n15987,n15901,n15902);
and (n15988,n81,n69);
and (n15989,n15990,n15991);
xor (n15990,n15987,n15988);
or (n15991,n15992,n15995);
and (n15992,n15993,n15994);
xor (n15993,n15907,n15908);
and (n15994,n63,n69);
and (n15995,n15996,n15997);
xor (n15996,n15993,n15994);
and (n15997,n15998,n451);
xor (n15998,n15912,n15913);
and (n15999,n192,n62);
and (n16000,n16001,n16002);
xor (n16001,n14820,n15999);
or (n16002,n16003,n16006);
and (n16003,n16004,n16005);
xor (n16004,n15918,n15919);
and (n16005,n173,n62);
and (n16006,n16007,n16008);
xor (n16007,n16004,n16005);
or (n16008,n16009,n16012);
and (n16009,n16010,n16011);
xor (n16010,n15924,n15925);
and (n16011,n496,n62);
and (n16012,n16013,n16014);
xor (n16013,n16010,n16011);
or (n16014,n16015,n16018);
and (n16015,n16016,n16017);
xor (n16016,n15930,n15931);
and (n16017,n490,n62);
and (n16018,n16019,n16020);
xor (n16019,n16016,n16017);
or (n16020,n16021,n16024);
and (n16021,n16022,n16023);
xor (n16022,n15936,n15937);
and (n16023,n43,n62);
and (n16024,n16025,n16026);
xor (n16025,n16022,n16023);
or (n16026,n16027,n16030);
and (n16027,n16028,n16029);
xor (n16028,n15942,n15943);
and (n16029,n53,n62);
and (n16030,n16031,n16032);
xor (n16031,n16028,n16029);
or (n16032,n16033,n16036);
and (n16033,n16034,n16035);
xor (n16034,n15948,n15949);
and (n16035,n223,n62);
and (n16036,n16037,n16038);
xor (n16037,n16034,n16035);
or (n16038,n16039,n16042);
and (n16039,n16040,n16041);
xor (n16040,n15954,n15955);
and (n16041,n217,n62);
and (n16042,n16043,n16044);
xor (n16043,n16040,n16041);
or (n16044,n16045,n16047);
and (n16045,n16046,n1797);
xor (n16046,n15960,n15961);
and (n16047,n16048,n16049);
xor (n16048,n16046,n1797);
or (n16049,n16050,n16053);
and (n16050,n16051,n16052);
xor (n16051,n15966,n15967);
and (n16052,n249,n62);
and (n16053,n16054,n16055);
xor (n16054,n16051,n16052);
or (n16055,n16056,n16058);
and (n16056,n16057,n1457);
xor (n16057,n15972,n15973);
and (n16058,n16059,n16060);
xor (n16059,n16057,n1457);
or (n16060,n16061,n16063);
and (n16061,n16062,n1107);
xor (n16062,n15978,n15979);
and (n16063,n16064,n16065);
xor (n16064,n16062,n1107);
or (n16065,n16066,n16069);
and (n16066,n16067,n16068);
xor (n16067,n15984,n15985);
and (n16068,n81,n62);
and (n16069,n16070,n16071);
xor (n16070,n16067,n16068);
or (n16071,n16072,n16075);
and (n16072,n16073,n16074);
xor (n16073,n15990,n15991);
and (n16074,n63,n62);
and (n16075,n16076,n16077);
xor (n16076,n16073,n16074);
and (n16077,n16078,n16079);
xor (n16078,n15996,n15997);
and (n16079,n452,n62);
and (n16080,n16081,n16082);
xor (n16081,n14817,n15999);
or (n16082,n16083,n16085);
and (n16083,n16084,n16005);
xor (n16084,n16001,n16002);
and (n16085,n16086,n16087);
xor (n16086,n16084,n16005);
or (n16087,n16088,n16090);
and (n16088,n16089,n16011);
xor (n16089,n16007,n16008);
and (n16090,n16091,n16092);
xor (n16091,n16089,n16011);
or (n16092,n16093,n16095);
and (n16093,n16094,n16017);
xor (n16094,n16013,n16014);
and (n16095,n16096,n16097);
xor (n16096,n16094,n16017);
or (n16097,n16098,n16100);
and (n16098,n16099,n16023);
xor (n16099,n16019,n16020);
and (n16100,n16101,n16102);
xor (n16101,n16099,n16023);
or (n16102,n16103,n16105);
and (n16103,n16104,n16029);
xor (n16104,n16025,n16026);
and (n16105,n16106,n16107);
xor (n16106,n16104,n16029);
or (n16107,n16108,n16110);
and (n16108,n16109,n16035);
xor (n16109,n16031,n16032);
and (n16110,n16111,n16112);
xor (n16111,n16109,n16035);
or (n16112,n16113,n16115);
and (n16113,n16114,n16041);
xor (n16114,n16037,n16038);
and (n16115,n16116,n16117);
xor (n16116,n16114,n16041);
or (n16117,n16118,n16120);
and (n16118,n16119,n1797);
xor (n16119,n16043,n16044);
and (n16120,n16121,n16122);
xor (n16121,n16119,n1797);
or (n16122,n16123,n16125);
and (n16123,n16124,n16052);
xor (n16124,n16048,n16049);
and (n16125,n16126,n16127);
xor (n16126,n16124,n16052);
or (n16127,n16128,n16130);
and (n16128,n16129,n1457);
xor (n16129,n16054,n16055);
and (n16130,n16131,n16132);
xor (n16131,n16129,n1457);
or (n16132,n16133,n16135);
and (n16133,n16134,n1107);
xor (n16134,n16059,n16060);
and (n16135,n16136,n16137);
xor (n16136,n16134,n1107);
or (n16137,n16138,n16140);
and (n16138,n16139,n16068);
xor (n16139,n16064,n16065);
and (n16140,n16141,n16142);
xor (n16141,n16139,n16068);
or (n16142,n16143,n16145);
and (n16143,n16144,n16074);
xor (n16144,n16070,n16071);
and (n16145,n16146,n16147);
xor (n16146,n16144,n16074);
and (n16147,n16148,n16079);
xor (n16148,n16076,n16077);
or (n16149,n16150,n16152);
and (n16150,n16151,n16005);
xor (n16151,n16081,n16082);
and (n16152,n16153,n16154);
xor (n16153,n16151,n16005);
or (n16154,n16155,n16157);
and (n16155,n16156,n16011);
xor (n16156,n16086,n16087);
and (n16157,n16158,n16159);
xor (n16158,n16156,n16011);
or (n16159,n16160,n16162);
and (n16160,n16161,n16017);
xor (n16161,n16091,n16092);
and (n16162,n16163,n16164);
xor (n16163,n16161,n16017);
or (n16164,n16165,n16167);
and (n16165,n16166,n16023);
xor (n16166,n16096,n16097);
and (n16167,n16168,n16169);
xor (n16168,n16166,n16023);
or (n16169,n16170,n16172);
and (n16170,n16171,n16029);
xor (n16171,n16101,n16102);
and (n16172,n16173,n16174);
xor (n16173,n16171,n16029);
or (n16174,n16175,n16177);
and (n16175,n16176,n16035);
xor (n16176,n16106,n16107);
and (n16177,n16178,n16179);
xor (n16178,n16176,n16035);
or (n16179,n16180,n16182);
and (n16180,n16181,n16041);
xor (n16181,n16111,n16112);
and (n16182,n16183,n16184);
xor (n16183,n16181,n16041);
or (n16184,n16185,n16187);
and (n16185,n16186,n1797);
xor (n16186,n16116,n16117);
and (n16187,n16188,n16189);
xor (n16188,n16186,n1797);
or (n16189,n16190,n16192);
and (n16190,n16191,n16052);
xor (n16191,n16121,n16122);
and (n16192,n16193,n16194);
xor (n16193,n16191,n16052);
or (n16194,n16195,n16197);
and (n16195,n16196,n1457);
xor (n16196,n16126,n16127);
and (n16197,n16198,n16199);
xor (n16198,n16196,n1457);
or (n16199,n16200,n16202);
and (n16200,n16201,n1107);
xor (n16201,n16131,n16132);
and (n16202,n16203,n16204);
xor (n16203,n16201,n1107);
or (n16204,n16205,n16207);
and (n16205,n16206,n16068);
xor (n16206,n16136,n16137);
and (n16207,n16208,n16209);
xor (n16208,n16206,n16068);
or (n16209,n16210,n16212);
and (n16210,n16211,n16074);
xor (n16211,n16141,n16142);
and (n16212,n16213,n16214);
xor (n16213,n16211,n16074);
and (n16214,n16215,n16079);
xor (n16215,n16146,n16147);
or (n16216,n16217,n16219);
and (n16217,n16218,n16011);
xor (n16218,n16153,n16154);
and (n16219,n16220,n16221);
xor (n16220,n16218,n16011);
or (n16221,n16222,n16224);
and (n16222,n16223,n16017);
xor (n16223,n16158,n16159);
and (n16224,n16225,n16226);
xor (n16225,n16223,n16017);
or (n16226,n16227,n16229);
and (n16227,n16228,n16023);
xor (n16228,n16163,n16164);
and (n16229,n16230,n16231);
xor (n16230,n16228,n16023);
or (n16231,n16232,n16234);
and (n16232,n16233,n16029);
xor (n16233,n16168,n16169);
and (n16234,n16235,n16236);
xor (n16235,n16233,n16029);
or (n16236,n16237,n16239);
and (n16237,n16238,n16035);
xor (n16238,n16173,n16174);
and (n16239,n16240,n16241);
xor (n16240,n16238,n16035);
or (n16241,n16242,n16244);
and (n16242,n16243,n16041);
xor (n16243,n16178,n16179);
and (n16244,n16245,n16246);
xor (n16245,n16243,n16041);
or (n16246,n16247,n16249);
and (n16247,n16248,n1797);
xor (n16248,n16183,n16184);
and (n16249,n16250,n16251);
xor (n16250,n16248,n1797);
or (n16251,n16252,n16254);
and (n16252,n16253,n16052);
xor (n16253,n16188,n16189);
and (n16254,n16255,n16256);
xor (n16255,n16253,n16052);
or (n16256,n16257,n16259);
and (n16257,n16258,n1457);
xor (n16258,n16193,n16194);
and (n16259,n16260,n16261);
xor (n16260,n16258,n1457);
or (n16261,n16262,n16264);
and (n16262,n16263,n1107);
xor (n16263,n16198,n16199);
and (n16264,n16265,n16266);
xor (n16265,n16263,n1107);
or (n16266,n16267,n16269);
and (n16267,n16268,n16068);
xor (n16268,n16203,n16204);
and (n16269,n16270,n16271);
xor (n16270,n16268,n16068);
or (n16271,n16272,n16274);
and (n16272,n16273,n16074);
xor (n16273,n16208,n16209);
and (n16274,n16275,n16276);
xor (n16275,n16273,n16074);
and (n16276,n16277,n16079);
xor (n16277,n16213,n16214);
or (n16278,n16279,n16281);
and (n16279,n16280,n16017);
xor (n16280,n16220,n16221);
and (n16281,n16282,n16283);
xor (n16282,n16280,n16017);
or (n16283,n16284,n16286);
and (n16284,n16285,n16023);
xor (n16285,n16225,n16226);
and (n16286,n16287,n16288);
xor (n16287,n16285,n16023);
or (n16288,n16289,n16291);
and (n16289,n16290,n16029);
xor (n16290,n16230,n16231);
and (n16291,n16292,n16293);
xor (n16292,n16290,n16029);
or (n16293,n16294,n16296);
and (n16294,n16295,n16035);
xor (n16295,n16235,n16236);
and (n16296,n16297,n16298);
xor (n16297,n16295,n16035);
or (n16298,n16299,n16301);
and (n16299,n16300,n16041);
xor (n16300,n16240,n16241);
and (n16301,n16302,n16303);
xor (n16302,n16300,n16041);
or (n16303,n16304,n16306);
and (n16304,n16305,n1797);
xor (n16305,n16245,n16246);
and (n16306,n16307,n16308);
xor (n16307,n16305,n1797);
or (n16308,n16309,n16311);
and (n16309,n16310,n16052);
xor (n16310,n16250,n16251);
and (n16311,n16312,n16313);
xor (n16312,n16310,n16052);
or (n16313,n16314,n16316);
and (n16314,n16315,n1457);
xor (n16315,n16255,n16256);
and (n16316,n16317,n16318);
xor (n16317,n16315,n1457);
or (n16318,n16319,n16321);
and (n16319,n16320,n1107);
xor (n16320,n16260,n16261);
and (n16321,n16322,n16323);
xor (n16322,n16320,n1107);
or (n16323,n16324,n16326);
and (n16324,n16325,n16068);
xor (n16325,n16265,n16266);
and (n16326,n16327,n16328);
xor (n16327,n16325,n16068);
or (n16328,n16329,n16331);
and (n16329,n16330,n16074);
xor (n16330,n16270,n16271);
and (n16331,n16332,n16333);
xor (n16332,n16330,n16074);
and (n16333,n16334,n16079);
xor (n16334,n16275,n16276);
or (n16335,n16336,n16338);
and (n16336,n16337,n16023);
xor (n16337,n16282,n16283);
and (n16338,n16339,n16340);
xor (n16339,n16337,n16023);
or (n16340,n16341,n16343);
and (n16341,n16342,n16029);
xor (n16342,n16287,n16288);
and (n16343,n16344,n16345);
xor (n16344,n16342,n16029);
or (n16345,n16346,n16348);
and (n16346,n16347,n16035);
xor (n16347,n16292,n16293);
and (n16348,n16349,n16350);
xor (n16349,n16347,n16035);
or (n16350,n16351,n16353);
and (n16351,n16352,n16041);
xor (n16352,n16297,n16298);
and (n16353,n16354,n16355);
xor (n16354,n16352,n16041);
or (n16355,n16356,n16358);
and (n16356,n16357,n1797);
xor (n16357,n16302,n16303);
and (n16358,n16359,n16360);
xor (n16359,n16357,n1797);
or (n16360,n16361,n16363);
and (n16361,n16362,n16052);
xor (n16362,n16307,n16308);
and (n16363,n16364,n16365);
xor (n16364,n16362,n16052);
or (n16365,n16366,n16368);
and (n16366,n16367,n1457);
xor (n16367,n16312,n16313);
and (n16368,n16369,n16370);
xor (n16369,n16367,n1457);
or (n16370,n16371,n16373);
and (n16371,n16372,n1107);
xor (n16372,n16317,n16318);
and (n16373,n16374,n16375);
xor (n16374,n16372,n1107);
or (n16375,n16376,n16378);
and (n16376,n16377,n16068);
xor (n16377,n16322,n16323);
and (n16378,n16379,n16380);
xor (n16379,n16377,n16068);
or (n16380,n16381,n16383);
and (n16381,n16382,n16074);
xor (n16382,n16327,n16328);
and (n16383,n16384,n16385);
xor (n16384,n16382,n16074);
and (n16385,n16386,n16079);
xor (n16386,n16332,n16333);
or (n16387,n16388,n16390);
and (n16388,n16389,n16029);
xor (n16389,n16339,n16340);
and (n16390,n16391,n16392);
xor (n16391,n16389,n16029);
or (n16392,n16393,n16395);
and (n16393,n16394,n16035);
xor (n16394,n16344,n16345);
and (n16395,n16396,n16397);
xor (n16396,n16394,n16035);
or (n16397,n16398,n16400);
and (n16398,n16399,n16041);
xor (n16399,n16349,n16350);
and (n16400,n16401,n16402);
xor (n16401,n16399,n16041);
or (n16402,n16403,n16405);
and (n16403,n16404,n1797);
xor (n16404,n16354,n16355);
and (n16405,n16406,n16407);
xor (n16406,n16404,n1797);
or (n16407,n16408,n16410);
and (n16408,n16409,n16052);
xor (n16409,n16359,n16360);
and (n16410,n16411,n16412);
xor (n16411,n16409,n16052);
or (n16412,n16413,n16415);
and (n16413,n16414,n1457);
xor (n16414,n16364,n16365);
and (n16415,n16416,n16417);
xor (n16416,n16414,n1457);
or (n16417,n16418,n16420);
and (n16418,n16419,n1107);
xor (n16419,n16369,n16370);
and (n16420,n16421,n16422);
xor (n16421,n16419,n1107);
or (n16422,n16423,n16425);
and (n16423,n16424,n16068);
xor (n16424,n16374,n16375);
and (n16425,n16426,n16427);
xor (n16426,n16424,n16068);
or (n16427,n16428,n16430);
and (n16428,n16429,n16074);
xor (n16429,n16379,n16380);
and (n16430,n16431,n16432);
xor (n16431,n16429,n16074);
and (n16432,n16433,n16079);
xor (n16433,n16384,n16385);
or (n16434,n16435,n16437);
and (n16435,n16436,n16035);
xor (n16436,n16391,n16392);
and (n16437,n16438,n16439);
xor (n16438,n16436,n16035);
or (n16439,n16440,n16442);
and (n16440,n16441,n16041);
xor (n16441,n16396,n16397);
and (n16442,n16443,n16444);
xor (n16443,n16441,n16041);
or (n16444,n16445,n16447);
and (n16445,n16446,n1797);
xor (n16446,n16401,n16402);
and (n16447,n16448,n16449);
xor (n16448,n16446,n1797);
or (n16449,n16450,n16452);
and (n16450,n16451,n16052);
xor (n16451,n16406,n16407);
and (n16452,n16453,n16454);
xor (n16453,n16451,n16052);
or (n16454,n16455,n16457);
and (n16455,n16456,n1457);
xor (n16456,n16411,n16412);
and (n16457,n16458,n16459);
xor (n16458,n16456,n1457);
or (n16459,n16460,n16462);
and (n16460,n16461,n1107);
xor (n16461,n16416,n16417);
and (n16462,n16463,n16464);
xor (n16463,n16461,n1107);
or (n16464,n16465,n16467);
and (n16465,n16466,n16068);
xor (n16466,n16421,n16422);
and (n16467,n16468,n16469);
xor (n16468,n16466,n16068);
or (n16469,n16470,n16472);
and (n16470,n16471,n16074);
xor (n16471,n16426,n16427);
and (n16472,n16473,n16474);
xor (n16473,n16471,n16074);
and (n16474,n16475,n16079);
xor (n16475,n16431,n16432);
or (n16476,n16477,n16479);
and (n16477,n16478,n16041);
xor (n16478,n16438,n16439);
and (n16479,n16480,n16481);
xor (n16480,n16478,n16041);
or (n16481,n16482,n16484);
and (n16482,n16483,n1797);
xor (n16483,n16443,n16444);
and (n16484,n16485,n16486);
xor (n16485,n16483,n1797);
or (n16486,n16487,n16489);
and (n16487,n16488,n16052);
xor (n16488,n16448,n16449);
and (n16489,n16490,n16491);
xor (n16490,n16488,n16052);
or (n16491,n16492,n16494);
and (n16492,n16493,n1457);
xor (n16493,n16453,n16454);
and (n16494,n16495,n16496);
xor (n16495,n16493,n1457);
or (n16496,n16497,n16499);
and (n16497,n16498,n1107);
xor (n16498,n16458,n16459);
and (n16499,n16500,n16501);
xor (n16500,n16498,n1107);
or (n16501,n16502,n16504);
and (n16502,n16503,n16068);
xor (n16503,n16463,n16464);
and (n16504,n16505,n16506);
xor (n16505,n16503,n16068);
or (n16506,n16507,n16509);
and (n16507,n16508,n16074);
xor (n16508,n16468,n16469);
and (n16509,n16510,n16511);
xor (n16510,n16508,n16074);
and (n16511,n16512,n16079);
xor (n16512,n16473,n16474);
or (n16513,n16514,n16516);
and (n16514,n16515,n1797);
xor (n16515,n16480,n16481);
and (n16516,n16517,n16518);
xor (n16517,n16515,n1797);
or (n16518,n16519,n16521);
and (n16519,n16520,n16052);
xor (n16520,n16485,n16486);
and (n16521,n16522,n16523);
xor (n16522,n16520,n16052);
or (n16523,n16524,n16526);
and (n16524,n16525,n1457);
xor (n16525,n16490,n16491);
and (n16526,n16527,n16528);
xor (n16527,n16525,n1457);
or (n16528,n16529,n16531);
and (n16529,n16530,n1107);
xor (n16530,n16495,n16496);
and (n16531,n16532,n16533);
xor (n16532,n16530,n1107);
or (n16533,n16534,n16536);
and (n16534,n16535,n16068);
xor (n16535,n16500,n16501);
and (n16536,n16537,n16538);
xor (n16537,n16535,n16068);
or (n16538,n16539,n16541);
and (n16539,n16540,n16074);
xor (n16540,n16505,n16506);
and (n16541,n16542,n16543);
xor (n16542,n16540,n16074);
and (n16543,n16544,n16079);
xor (n16544,n16510,n16511);
or (n16545,n16546,n16548);
and (n16546,n16547,n16052);
xor (n16547,n16517,n16518);
and (n16548,n16549,n16550);
xor (n16549,n16547,n16052);
or (n16550,n16551,n16553);
and (n16551,n16552,n1457);
xor (n16552,n16522,n16523);
and (n16553,n16554,n16555);
xor (n16554,n16552,n1457);
or (n16555,n16556,n16558);
and (n16556,n16557,n1107);
xor (n16557,n16527,n16528);
and (n16558,n16559,n16560);
xor (n16559,n16557,n1107);
or (n16560,n16561,n16563);
and (n16561,n16562,n16068);
xor (n16562,n16532,n16533);
and (n16563,n16564,n16565);
xor (n16564,n16562,n16068);
or (n16565,n16566,n16568);
and (n16566,n16567,n16074);
xor (n16567,n16537,n16538);
and (n16568,n16569,n16570);
xor (n16569,n16567,n16074);
and (n16570,n16571,n16079);
xor (n16571,n16542,n16543);
or (n16572,n16573,n16575);
and (n16573,n16574,n1457);
xor (n16574,n16549,n16550);
and (n16575,n16576,n16577);
xor (n16576,n16574,n1457);
or (n16577,n16578,n16580);
and (n16578,n16579,n1107);
xor (n16579,n16554,n16555);
and (n16580,n16581,n16582);
xor (n16581,n16579,n1107);
or (n16582,n16583,n16585);
and (n16583,n16584,n16068);
xor (n16584,n16559,n16560);
and (n16585,n16586,n16587);
xor (n16586,n16584,n16068);
or (n16587,n16588,n16590);
and (n16588,n16589,n16074);
xor (n16589,n16564,n16565);
and (n16590,n16591,n16592);
xor (n16591,n16589,n16074);
and (n16592,n16593,n16079);
xor (n16593,n16569,n16570);
or (n16594,n16595,n16597);
and (n16595,n16596,n1107);
xor (n16596,n16576,n16577);
and (n16597,n16598,n16599);
xor (n16598,n16596,n1107);
or (n16599,n16600,n16602);
and (n16600,n16601,n16068);
xor (n16601,n16581,n16582);
and (n16602,n16603,n16604);
xor (n16603,n16601,n16068);
or (n16604,n16605,n16607);
and (n16605,n16606,n16074);
xor (n16606,n16586,n16587);
and (n16607,n16608,n16609);
xor (n16608,n16606,n16074);
and (n16609,n16610,n16079);
xor (n16610,n16591,n16592);
or (n16611,n16612,n16614);
and (n16612,n16613,n16068);
xor (n16613,n16598,n16599);
and (n16614,n16615,n16616);
xor (n16615,n16613,n16068);
or (n16616,n16617,n16619);
and (n16617,n16618,n16074);
xor (n16618,n16603,n16604);
and (n16619,n16620,n16621);
xor (n16620,n16618,n16074);
and (n16621,n16622,n16079);
xor (n16622,n16608,n16609);
or (n16623,n16624,n16626);
and (n16624,n16625,n16074);
xor (n16625,n16615,n16616);
and (n16626,n16627,n16628);
xor (n16627,n16625,n16074);
and (n16628,n16629,n16079);
xor (n16629,n16620,n16621);
and (n16630,n16631,n16079);
xor (n16631,n16627,n16628);
not (n16632,n16633);
xor (n16633,n16634,n644);
xor (n16634,n16635,n18505);
xor (n16635,n16636,n103);
xor (n16636,n16637,n18498);
xor (n16637,n16638,n109);
xor (n16638,n16639,n18486);
xor (n16639,n16640,n1101);
xor (n16640,n16641,n18469);
xor (n16641,n16642,n1534);
xor (n16642,n16643,n18447);
xor (n16643,n16644,n1538);
xor (n16644,n16645,n18420);
xor (n16645,n16646,n17925);
xor (n16646,n16647,n18388);
xor (n16647,n16648,n17919);
xor (n16648,n16649,n18351);
xor (n16649,n16650,n2040);
xor (n16650,n16651,n18309);
xor (n16651,n16652,n17908);
xor (n16652,n16653,n18262);
xor (n16653,n16654,n2218);
xor (n16654,n16655,n18210);
xor (n16655,n16656,n2295);
xor (n16656,n16657,n18153);
xor (n16657,n16658,n2397);
xor (n16658,n16659,n18091);
xor (n16659,n16660,n2401);
xor (n16660,n16661,n18024);
xor (n16661,n16662,n2457);
xor (n16662,n16663,n16721);
xor (n16663,n16664,n2494);
xor (n16664,n16665,n16720);
xor (n16665,n16666,n2494);
xor (n16666,n16667,n16719);
xor (n16667,n16668,n16718);
xor (n16668,n16669,n16717);
xor (n16669,n16670,n2424);
xor (n16670,n16671,n16716);
xor (n16671,n16672,n16715);
xor (n16672,n16673,n16714);
xor (n16673,n16674,n2316);
xor (n16674,n16675,n16713);
xor (n16675,n16676,n16712);
xor (n16676,n16677,n16711);
xor (n16677,n16678,n16710);
xor (n16678,n16679,n16709);
xor (n16679,n16680,n16708);
xor (n16680,n16681,n16707);
xor (n16681,n16682,n16706);
xor (n16682,n16683,n16705);
xor (n16683,n16684,n16704);
xor (n16684,n16685,n16703);
xor (n16685,n16686,n16702);
xor (n16686,n16687,n16701);
xor (n16687,n16688,n16700);
xor (n16688,n16689,n16699);
xor (n16689,n16690,n16698);
xor (n16690,n16691,n16697);
xor (n16691,n16692,n16696);
xor (n16692,n16693,n16695);
xor (n16693,n16694,n558);
and (n16694,n556,n229);
and (n16695,n16694,n558);
and (n16696,n556,n288);
and (n16697,n16692,n16696);
not (n16698,n1066);
and (n16699,n16690,n16698);
and (n16700,n556,n314);
and (n16701,n16688,n16700);
and (n16702,n556,n307);
and (n16703,n16686,n16702);
and (n16704,n556,n392);
and (n16705,n16684,n16704);
and (n16706,n556,n385);
and (n16707,n16682,n16706);
and (n16708,n556,n416);
and (n16709,n16680,n16708);
and (n16710,n556,n126);
and (n16711,n16678,n16710);
and (n16712,n556,n120);
and (n16713,n16676,n16712);
and (n16714,n16674,n2316);
and (n16715,n556,n147);
and (n16716,n16672,n16715);
and (n16717,n16670,n2424);
and (n16718,n556,n92);
and (n16719,n16668,n16718);
and (n16720,n16666,n2494);
or (n16721,n16722,n17955);
and (n16722,n16723,n2457);
xor (n16723,n16665,n16724);
or (n16724,n16725,n17883);
and (n16725,n16726,n2457);
xor (n16726,n16667,n16727);
or (n16727,n16728,n17800);
and (n16728,n16729,n17799);
xor (n16729,n16669,n16730);
or (n16730,n16731,n17727);
and (n16731,n16732,n2367);
xor (n16732,n16671,n16733);
or (n16733,n16734,n17644);
and (n16734,n16735,n17643);
xor (n16735,n16673,n16736);
or (n16736,n16737,n17567);
and (n16737,n16738,n2241);
xor (n16738,n16675,n16739);
or (n16739,n16740,n17484);
and (n16740,n16741,n17483);
xor (n16741,n16677,n16742);
or (n16742,n16743,n17408);
and (n16743,n16744,n2068);
xor (n16744,n16679,n16745);
or (n16745,n16746,n17325);
and (n16746,n16747,n17324);
xor (n16747,n16681,n16748);
or (n16748,n16749,n17248);
and (n16749,n16750,n17247);
xor (n16750,n16683,n16751);
or (n16751,n16752,n17164);
and (n16752,n16753,n17163);
xor (n16753,n16685,n16754);
or (n16754,n16755,n17086);
and (n16755,n16756,n1514);
xor (n16756,n16687,n16757);
or (n16757,n16758,n17003);
and (n16758,n16759,n17002);
xor (n16759,n16689,n16760);
or (n16760,n16761,n16927);
and (n16761,n16762,n16926);
xor (n16762,n16691,n16763);
or (n16763,n16764,n16843);
and (n16764,n16765,n16842);
xor (n16765,n16693,n16766);
or (n16766,n16767,n16768);
and (n16767,n16694,n242);
and (n16768,n16769,n16770);
xor (n16769,n16694,n242);
or (n16770,n16771,n16773);
and (n16771,n16772,n236);
and (n16772,n240,n229);
and (n16773,n16774,n16775);
xor (n16774,n16772,n236);
or (n16775,n16776,n16778);
and (n16776,n16777,n813);
and (n16777,n234,n229);
and (n16778,n16779,n16780);
xor (n16779,n16777,n813);
or (n16780,n16781,n16783);
and (n16781,n16782,n819);
and (n16782,n297,n229);
and (n16783,n16784,n16785);
xor (n16784,n16782,n819);
or (n16785,n16786,n16789);
and (n16786,n16787,n16788);
and (n16787,n278,n229);
and (n16788,n323,n230);
and (n16789,n16790,n16791);
xor (n16790,n16787,n16788);
or (n16791,n16792,n16794);
and (n16792,n16793,n2678);
and (n16793,n323,n229);
and (n16794,n16795,n16796);
xor (n16795,n16793,n2678);
or (n16796,n16797,n16800);
and (n16797,n16798,n16799);
and (n16798,n306,n229);
and (n16799,n384,n230);
and (n16800,n16801,n16802);
xor (n16801,n16798,n16799);
or (n16802,n16803,n16805);
and (n16803,n16804,n2850);
and (n16804,n384,n229);
and (n16805,n16806,n16807);
xor (n16806,n16804,n2850);
or (n16807,n16808,n16810);
and (n16808,n16809,n3004);
and (n16809,n403,n229);
and (n16810,n16811,n16812);
xor (n16811,n16809,n3004);
or (n16812,n16813,n16815);
and (n16813,n16814,n3048);
and (n16814,n138,n229);
and (n16815,n16816,n16817);
xor (n16816,n16814,n3048);
or (n16817,n16818,n16821);
and (n16818,n16819,n16820);
and (n16819,n131,n229);
and (n16820,n163,n230);
and (n16821,n16822,n16823);
xor (n16822,n16819,n16820);
or (n16823,n16824,n16826);
and (n16824,n16825,n3223);
and (n16825,n163,n229);
and (n16826,n16827,n16828);
xor (n16827,n16825,n3223);
or (n16828,n16829,n16832);
and (n16829,n16830,n16831);
and (n16830,n156,n229);
and (n16831,n108,n230);
and (n16832,n16833,n16834);
xor (n16833,n16830,n16831);
or (n16834,n16835,n16838);
and (n16835,n16836,n16837);
and (n16836,n108,n229);
and (n16837,n102,n230);
and (n16838,n16839,n16840);
xor (n16839,n16836,n16837);
and (n16840,n16841,n3331);
and (n16841,n102,n229);
and (n16842,n240,n288);
and (n16843,n16844,n16845);
xor (n16844,n16765,n16842);
or (n16845,n16846,n16849);
and (n16846,n16847,n16848);
xor (n16847,n16769,n16770);
and (n16848,n234,n288);
and (n16849,n16850,n16851);
xor (n16850,n16847,n16848);
or (n16851,n16852,n16855);
and (n16852,n16853,n16854);
xor (n16853,n16774,n16775);
and (n16854,n297,n288);
and (n16855,n16856,n16857);
xor (n16856,n16853,n16854);
or (n16857,n16858,n16861);
and (n16858,n16859,n16860);
xor (n16859,n16779,n16780);
and (n16860,n278,n288);
and (n16861,n16862,n16863);
xor (n16862,n16859,n16860);
or (n16863,n16864,n16867);
and (n16864,n16865,n16866);
xor (n16865,n16784,n16785);
and (n16866,n323,n288);
and (n16867,n16868,n16869);
xor (n16868,n16865,n16866);
or (n16869,n16870,n16873);
and (n16870,n16871,n16872);
xor (n16871,n16790,n16791);
and (n16872,n306,n288);
and (n16873,n16874,n16875);
xor (n16874,n16871,n16872);
or (n16875,n16876,n16879);
and (n16876,n16877,n16878);
xor (n16877,n16795,n16796);
and (n16878,n384,n288);
and (n16879,n16880,n16881);
xor (n16880,n16877,n16878);
or (n16881,n16882,n16885);
and (n16882,n16883,n16884);
xor (n16883,n16801,n16802);
and (n16884,n403,n288);
and (n16885,n16886,n16887);
xor (n16886,n16883,n16884);
or (n16887,n16888,n16891);
and (n16888,n16889,n16890);
xor (n16889,n16806,n16807);
and (n16890,n138,n288);
and (n16891,n16892,n16893);
xor (n16892,n16889,n16890);
or (n16893,n16894,n16897);
and (n16894,n16895,n16896);
xor (n16895,n16811,n16812);
and (n16896,n131,n288);
and (n16897,n16898,n16899);
xor (n16898,n16895,n16896);
or (n16899,n16900,n16903);
and (n16900,n16901,n16902);
xor (n16901,n16816,n16817);
and (n16902,n163,n288);
and (n16903,n16904,n16905);
xor (n16904,n16901,n16902);
or (n16905,n16906,n16909);
and (n16906,n16907,n16908);
xor (n16907,n16822,n16823);
and (n16908,n156,n288);
and (n16909,n16910,n16911);
xor (n16910,n16907,n16908);
or (n16911,n16912,n16915);
and (n16912,n16913,n16914);
xor (n16913,n16827,n16828);
and (n16914,n108,n288);
and (n16915,n16916,n16917);
xor (n16916,n16913,n16914);
or (n16917,n16918,n16921);
and (n16918,n16919,n16920);
xor (n16919,n16833,n16834);
and (n16920,n102,n288);
and (n16921,n16922,n16923);
xor (n16922,n16919,n16920);
and (n16923,n16924,n16925);
xor (n16924,n16839,n16840);
and (n16925,n460,n288);
and (n16926,n240,n280);
and (n16927,n16928,n16929);
xor (n16928,n16762,n16926);
or (n16929,n16930,n16933);
and (n16930,n16931,n16932);
xor (n16931,n16844,n16845);
and (n16932,n234,n280);
and (n16933,n16934,n16935);
xor (n16934,n16931,n16932);
or (n16935,n16936,n16938);
and (n16936,n16937,n299);
xor (n16937,n16850,n16851);
and (n16938,n16939,n16940);
xor (n16939,n16937,n299);
or (n16940,n16941,n16944);
and (n16941,n16942,n16943);
xor (n16942,n16856,n16857);
and (n16943,n278,n280);
and (n16944,n16945,n16946);
xor (n16945,n16942,n16943);
or (n16946,n16947,n16949);
and (n16947,n16948,n830);
xor (n16948,n16862,n16863);
and (n16949,n16950,n16951);
xor (n16950,n16948,n830);
or (n16951,n16952,n16954);
and (n16952,n16953,n834);
xor (n16953,n16868,n16869);
and (n16954,n16955,n16956);
xor (n16955,n16953,n834);
or (n16956,n16957,n16959);
and (n16957,n16958,n1268);
xor (n16958,n16874,n16875);
and (n16959,n16960,n16961);
xor (n16960,n16958,n1268);
or (n16961,n16962,n16964);
and (n16962,n16963,n2589);
xor (n16963,n16880,n16881);
and (n16964,n16965,n16966);
xor (n16965,n16963,n2589);
or (n16966,n16967,n16970);
and (n16967,n16968,n16969);
xor (n16968,n16886,n16887);
and (n16969,n138,n280);
and (n16970,n16971,n16972);
xor (n16971,n16968,n16969);
or (n16972,n16973,n16976);
and (n16973,n16974,n16975);
xor (n16974,n16892,n16893);
and (n16975,n131,n280);
and (n16976,n16977,n16978);
xor (n16977,n16974,n16975);
or (n16978,n16979,n16982);
and (n16979,n16980,n16981);
xor (n16980,n16898,n16899);
and (n16981,n163,n280);
and (n16982,n16983,n16984);
xor (n16983,n16980,n16981);
or (n16984,n16985,n16987);
and (n16985,n16986,n3061);
xor (n16986,n16904,n16905);
and (n16987,n16988,n16989);
xor (n16988,n16986,n3061);
or (n16989,n16990,n16993);
and (n16990,n16991,n16992);
xor (n16991,n16910,n16911);
and (n16992,n108,n280);
and (n16993,n16994,n16995);
xor (n16994,n16991,n16992);
or (n16995,n16996,n16998);
and (n16996,n16997,n3182);
xor (n16997,n16916,n16917);
and (n16998,n16999,n17000);
xor (n16999,n16997,n3182);
and (n17000,n17001,n3257);
xor (n17001,n16922,n16923);
and (n17002,n240,n314);
and (n17003,n17004,n17005);
xor (n17004,n16759,n17002);
or (n17005,n17006,n17009);
and (n17006,n17007,n17008);
xor (n17007,n16928,n16929);
and (n17008,n234,n314);
and (n17009,n17010,n17011);
xor (n17010,n17007,n17008);
or (n17011,n17012,n17015);
and (n17012,n17013,n17014);
xor (n17013,n16934,n16935);
and (n17014,n297,n314);
and (n17015,n17016,n17017);
xor (n17016,n17013,n17014);
or (n17017,n17018,n17021);
and (n17018,n17019,n17020);
xor (n17019,n16939,n16940);
and (n17020,n278,n314);
and (n17021,n17022,n17023);
xor (n17022,n17019,n17020);
or (n17023,n17024,n17027);
and (n17024,n17025,n17026);
xor (n17025,n16945,n16946);
and (n17026,n323,n314);
and (n17027,n17028,n17029);
xor (n17028,n17025,n17026);
or (n17029,n17030,n17033);
and (n17030,n17031,n17032);
xor (n17031,n16950,n16951);
and (n17032,n306,n314);
and (n17033,n17034,n17035);
xor (n17034,n17031,n17032);
or (n17035,n17036,n17039);
and (n17036,n17037,n17038);
xor (n17037,n16955,n16956);
and (n17038,n384,n314);
and (n17039,n17040,n17041);
xor (n17040,n17037,n17038);
or (n17041,n17042,n17045);
and (n17042,n17043,n17044);
xor (n17043,n16960,n16961);
and (n17044,n403,n314);
and (n17045,n17046,n17047);
xor (n17046,n17043,n17044);
or (n17047,n17048,n17051);
and (n17048,n17049,n17050);
xor (n17049,n16965,n16966);
and (n17050,n138,n314);
and (n17051,n17052,n17053);
xor (n17052,n17049,n17050);
or (n17053,n17054,n17057);
and (n17054,n17055,n17056);
xor (n17055,n16971,n16972);
and (n17056,n131,n314);
and (n17057,n17058,n17059);
xor (n17058,n17055,n17056);
or (n17059,n17060,n17063);
and (n17060,n17061,n17062);
xor (n17061,n16977,n16978);
and (n17062,n163,n314);
and (n17063,n17064,n17065);
xor (n17064,n17061,n17062);
or (n17065,n17066,n17069);
and (n17066,n17067,n17068);
xor (n17067,n16983,n16984);
and (n17068,n156,n314);
and (n17069,n17070,n17071);
xor (n17070,n17067,n17068);
or (n17071,n17072,n17075);
and (n17072,n17073,n17074);
xor (n17073,n16988,n16989);
and (n17074,n108,n314);
and (n17075,n17076,n17077);
xor (n17076,n17073,n17074);
or (n17077,n17078,n17081);
and (n17078,n17079,n17080);
xor (n17079,n16994,n16995);
and (n17080,n102,n314);
and (n17081,n17082,n17083);
xor (n17082,n17079,n17080);
and (n17083,n17084,n17085);
xor (n17084,n16999,n17000);
and (n17085,n460,n314);
and (n17086,n17087,n17088);
xor (n17087,n16756,n1514);
or (n17088,n17089,n17092);
and (n17089,n17090,n17091);
xor (n17090,n17004,n17005);
not (n17091,n1073);
and (n17092,n17093,n17094);
xor (n17093,n17090,n17091);
or (n17094,n17095,n17098);
and (n17095,n17096,n17097);
xor (n17096,n17010,n17011);
not (n17097,n738);
and (n17098,n17099,n17100);
xor (n17099,n17096,n17097);
or (n17100,n17101,n17103);
and (n17101,n17102,n607);
xor (n17102,n17016,n17017);
and (n17103,n17104,n17105);
xor (n17104,n17102,n607);
or (n17105,n17106,n17108);
and (n17106,n17107,n325);
xor (n17107,n17022,n17023);
and (n17108,n17109,n17110);
xor (n17109,n17107,n325);
or (n17110,n17111,n17114);
and (n17111,n17112,n17113);
xor (n17112,n17028,n17029);
and (n17113,n306,n307);
and (n17114,n17115,n17116);
xor (n17115,n17112,n17113);
or (n17116,n17117,n17119);
and (n17117,n17118,n850);
xor (n17118,n17034,n17035);
and (n17119,n17120,n17121);
xor (n17120,n17118,n850);
or (n17121,n17122,n17124);
and (n17122,n17123,n855);
xor (n17123,n17040,n17041);
and (n17124,n17125,n17126);
xor (n17125,n17123,n855);
or (n17126,n17127,n17130);
and (n17127,n17128,n17129);
xor (n17128,n17046,n17047);
and (n17129,n138,n307);
and (n17130,n17131,n17132);
xor (n17131,n17128,n17129);
or (n17132,n17133,n17136);
and (n17133,n17134,n17135);
xor (n17134,n17052,n17053);
and (n17135,n131,n307);
and (n17136,n17137,n17138);
xor (n17137,n17134,n17135);
or (n17138,n17139,n17142);
and (n17139,n17140,n17141);
xor (n17140,n17058,n17059);
and (n17141,n163,n307);
and (n17142,n17143,n17144);
xor (n17143,n17140,n17141);
or (n17144,n17145,n17148);
and (n17145,n17146,n17147);
xor (n17146,n17064,n17065);
and (n17147,n156,n307);
and (n17148,n17149,n17150);
xor (n17149,n17146,n17147);
or (n17150,n17151,n17154);
and (n17151,n17152,n17153);
xor (n17152,n17070,n17071);
and (n17153,n108,n307);
and (n17154,n17155,n17156);
xor (n17155,n17152,n17153);
or (n17156,n17157,n17159);
and (n17157,n17158,n3094);
xor (n17158,n17076,n17077);
and (n17159,n17160,n17161);
xor (n17160,n17158,n3094);
and (n17161,n17162,n3175);
xor (n17162,n17082,n17083);
and (n17163,n240,n392);
and (n17164,n17165,n17166);
xor (n17165,n16753,n17163);
or (n17166,n17167,n17170);
and (n17167,n17168,n17169);
xor (n17168,n17087,n17088);
and (n17169,n234,n392);
and (n17170,n17171,n17172);
xor (n17171,n17168,n17169);
or (n17172,n17173,n17176);
and (n17173,n17174,n17175);
xor (n17174,n17093,n17094);
and (n17175,n297,n392);
and (n17176,n17177,n17178);
xor (n17177,n17174,n17175);
or (n17178,n17179,n17182);
and (n17179,n17180,n17181);
xor (n17180,n17099,n17100);
and (n17181,n278,n392);
and (n17182,n17183,n17184);
xor (n17183,n17180,n17181);
or (n17184,n17185,n17188);
and (n17185,n17186,n17187);
xor (n17186,n17104,n17105);
and (n17187,n323,n392);
and (n17188,n17189,n17190);
xor (n17189,n17186,n17187);
or (n17190,n17191,n17194);
and (n17191,n17192,n17193);
xor (n17192,n17109,n17110);
and (n17193,n306,n392);
and (n17194,n17195,n17196);
xor (n17195,n17192,n17193);
or (n17196,n17197,n17200);
and (n17197,n17198,n17199);
xor (n17198,n17115,n17116);
and (n17199,n384,n392);
and (n17200,n17201,n17202);
xor (n17201,n17198,n17199);
or (n17202,n17203,n17206);
and (n17203,n17204,n17205);
xor (n17204,n17120,n17121);
and (n17205,n403,n392);
and (n17206,n17207,n17208);
xor (n17207,n17204,n17205);
or (n17208,n17209,n17212);
and (n17209,n17210,n17211);
xor (n17210,n17125,n17126);
and (n17211,n138,n392);
and (n17212,n17213,n17214);
xor (n17213,n17210,n17211);
or (n17214,n17215,n17218);
and (n17215,n17216,n17217);
xor (n17216,n17131,n17132);
and (n17217,n131,n392);
and (n17218,n17219,n17220);
xor (n17219,n17216,n17217);
or (n17220,n17221,n17224);
and (n17221,n17222,n17223);
xor (n17222,n17137,n17138);
and (n17223,n163,n392);
and (n17224,n17225,n17226);
xor (n17225,n17222,n17223);
or (n17226,n17227,n17230);
and (n17227,n17228,n17229);
xor (n17228,n17143,n17144);
and (n17229,n156,n392);
and (n17230,n17231,n17232);
xor (n17231,n17228,n17229);
or (n17232,n17233,n17236);
and (n17233,n17234,n17235);
xor (n17234,n17149,n17150);
and (n17235,n108,n392);
and (n17236,n17237,n17238);
xor (n17237,n17234,n17235);
or (n17238,n17239,n17242);
and (n17239,n17240,n17241);
xor (n17240,n17155,n17156);
and (n17241,n102,n392);
and (n17242,n17243,n17244);
xor (n17243,n17240,n17241);
and (n17244,n17245,n17246);
xor (n17245,n17160,n17161);
and (n17246,n460,n392);
and (n17247,n240,n385);
and (n17248,n17249,n17250);
xor (n17249,n16750,n17247);
or (n17250,n17251,n17254);
and (n17251,n17252,n17253);
xor (n17252,n17165,n17166);
not (n17253,n1630);
and (n17254,n17255,n17256);
xor (n17255,n17252,n17253);
or (n17256,n17257,n17260);
and (n17257,n17258,n17259);
xor (n17258,n17171,n17172);
and (n17259,n297,n385);
and (n17260,n17261,n17262);
xor (n17261,n17258,n17259);
or (n17262,n17263,n17265);
and (n17263,n17264,n1160);
xor (n17264,n17177,n17178);
and (n17265,n17266,n17267);
xor (n17266,n17264,n1160);
or (n17267,n17268,n17271);
and (n17268,n17269,n17270);
xor (n17269,n17183,n17184);
not (n17270,n693);
and (n17271,n17272,n17273);
xor (n17272,n17269,n17270);
or (n17273,n17274,n17277);
and (n17274,n17275,n17276);
xor (n17275,n17189,n17190);
and (n17276,n306,n385);
and (n17277,n17278,n17279);
xor (n17278,n17275,n17276);
or (n17279,n17280,n17283);
and (n17280,n17281,n17282);
xor (n17281,n17195,n17196);
and (n17282,n384,n385);
and (n17283,n17284,n17285);
xor (n17284,n17281,n17282);
or (n17285,n17286,n17288);
and (n17286,n17287,n402);
xor (n17287,n17201,n17202);
and (n17288,n17289,n17290);
xor (n17289,n17287,n402);
or (n17290,n17291,n17294);
and (n17291,n17292,n17293);
xor (n17292,n17207,n17208);
and (n17293,n138,n385);
and (n17294,n17295,n17296);
xor (n17295,n17292,n17293);
or (n17296,n17297,n17300);
and (n17297,n17298,n17299);
xor (n17298,n17213,n17214);
and (n17299,n131,n385);
and (n17300,n17301,n17302);
xor (n17301,n17298,n17299);
or (n17302,n17303,n17305);
and (n17303,n17304,n1294);
xor (n17304,n17219,n17220);
and (n17305,n17306,n17307);
xor (n17306,n17304,n1294);
or (n17307,n17308,n17310);
and (n17308,n17309,n2618);
xor (n17309,n17225,n17226);
and (n17310,n17311,n17312);
xor (n17311,n17309,n2618);
or (n17312,n17313,n17315);
and (n17313,n17314,n2723);
xor (n17314,n17231,n17232);
and (n17315,n17316,n17317);
xor (n17316,n17314,n2723);
or (n17317,n17318,n17320);
and (n17318,n17319,n2886);
xor (n17319,n17237,n17238);
and (n17320,n17321,n17322);
xor (n17321,n17319,n2886);
and (n17322,n17323,n2979);
xor (n17323,n17243,n17244);
and (n17324,n240,n416);
and (n17325,n17326,n17327);
xor (n17326,n16747,n17324);
or (n17327,n17328,n17331);
and (n17328,n17329,n17330);
xor (n17329,n17249,n17250);
and (n17330,n234,n416);
and (n17331,n17332,n17333);
xor (n17332,n17329,n17330);
or (n17333,n17334,n17337);
and (n17334,n17335,n17336);
xor (n17335,n17255,n17256);
and (n17336,n297,n416);
and (n17337,n17338,n17339);
xor (n17338,n17335,n17336);
or (n17339,n17340,n17343);
and (n17340,n17341,n17342);
xor (n17341,n17261,n17262);
and (n17342,n278,n416);
and (n17343,n17344,n17345);
xor (n17344,n17341,n17342);
or (n17345,n17346,n17349);
and (n17346,n17347,n17348);
xor (n17347,n17266,n17267);
and (n17348,n323,n416);
and (n17349,n17350,n17351);
xor (n17350,n17347,n17348);
or (n17351,n17352,n17355);
and (n17352,n17353,n17354);
xor (n17353,n17272,n17273);
and (n17354,n306,n416);
and (n17355,n17356,n17357);
xor (n17356,n17353,n17354);
or (n17357,n17358,n17361);
and (n17358,n17359,n17360);
xor (n17359,n17278,n17279);
and (n17360,n384,n416);
and (n17361,n17362,n17363);
xor (n17362,n17359,n17360);
or (n17363,n17364,n17367);
and (n17364,n17365,n17366);
xor (n17365,n17284,n17285);
and (n17366,n403,n416);
and (n17367,n17368,n17369);
xor (n17368,n17365,n17366);
or (n17369,n17370,n17373);
and (n17370,n17371,n17372);
xor (n17371,n17289,n17290);
and (n17372,n138,n416);
and (n17373,n17374,n17375);
xor (n17374,n17371,n17372);
or (n17375,n17376,n17379);
and (n17376,n17377,n17378);
xor (n17377,n17295,n17296);
and (n17378,n131,n416);
and (n17379,n17380,n17381);
xor (n17380,n17377,n17378);
or (n17381,n17382,n17385);
and (n17382,n17383,n17384);
xor (n17383,n17301,n17302);
and (n17384,n163,n416);
and (n17385,n17386,n17387);
xor (n17386,n17383,n17384);
or (n17387,n17388,n17391);
and (n17388,n17389,n17390);
xor (n17389,n17306,n17307);
and (n17390,n156,n416);
and (n17391,n17392,n17393);
xor (n17392,n17389,n17390);
or (n17393,n17394,n17397);
and (n17394,n17395,n17396);
xor (n17395,n17311,n17312);
and (n17396,n108,n416);
and (n17397,n17398,n17399);
xor (n17398,n17395,n17396);
or (n17399,n17400,n17403);
and (n17400,n17401,n17402);
xor (n17401,n17316,n17317);
and (n17402,n102,n416);
and (n17403,n17404,n17405);
xor (n17404,n17401,n17402);
and (n17405,n17406,n17407);
xor (n17406,n17321,n17322);
and (n17407,n460,n416);
and (n17408,n17409,n17410);
xor (n17409,n16744,n2068);
or (n17410,n17411,n17413);
and (n17411,n17412,n1875);
xor (n17412,n17326,n17327);
and (n17413,n17414,n17415);
xor (n17414,n17412,n1875);
or (n17415,n17416,n17418);
and (n17416,n17417,n1764);
xor (n17417,n17332,n17333);
and (n17418,n17419,n17420);
xor (n17419,n17417,n1764);
or (n17420,n17421,n17424);
and (n17421,n17422,n17423);
xor (n17422,n17338,n17339);
and (n17423,n278,n126);
and (n17424,n17425,n17426);
xor (n17425,n17422,n17423);
or (n17426,n17427,n17430);
and (n17427,n17428,n17429);
xor (n17428,n17344,n17345);
and (n17429,n323,n126);
and (n17430,n17431,n17432);
xor (n17431,n17428,n17429);
or (n17432,n17433,n17436);
and (n17433,n17434,n17435);
xor (n17434,n17350,n17351);
and (n17435,n306,n126);
and (n17436,n17437,n17438);
xor (n17437,n17434,n17435);
or (n17438,n17439,n17442);
and (n17439,n17440,n17441);
xor (n17440,n17356,n17357);
and (n17441,n384,n126);
and (n17442,n17443,n17444);
xor (n17443,n17440,n17441);
or (n17444,n17445,n17448);
and (n17445,n17446,n17447);
xor (n17446,n17362,n17363);
and (n17447,n403,n126);
and (n17448,n17449,n17450);
xor (n17449,n17446,n17447);
or (n17450,n17451,n17453);
and (n17451,n17452,n428);
xor (n17452,n17368,n17369);
and (n17453,n17454,n17455);
xor (n17454,n17452,n428);
or (n17455,n17456,n17459);
and (n17456,n17457,n17458);
xor (n17457,n17374,n17375);
and (n17458,n131,n126);
and (n17459,n17460,n17461);
xor (n17460,n17457,n17458);
or (n17461,n17462,n17464);
and (n17462,n17463,n890);
xor (n17463,n17380,n17381);
and (n17464,n17465,n17466);
xor (n17465,n17463,n890);
or (n17466,n17467,n17469);
and (n17467,n17468,n886);
xor (n17468,n17386,n17387);
and (n17469,n17470,n17471);
xor (n17470,n17468,n886);
or (n17471,n17472,n17474);
and (n17472,n17473,n1318);
xor (n17473,n17392,n17393);
and (n17474,n17475,n17476);
xor (n17475,n17473,n1318);
or (n17476,n17477,n17479);
and (n17477,n17478,n2625);
xor (n17478,n17398,n17399);
and (n17479,n17480,n17481);
xor (n17480,n17478,n2625);
and (n17481,n17482,n2729);
xor (n17482,n17404,n17405);
and (n17483,n240,n120);
and (n17484,n17485,n17486);
xor (n17485,n16741,n17483);
or (n17486,n17487,n17490);
and (n17487,n17488,n17489);
xor (n17488,n17409,n17410);
and (n17489,n234,n120);
and (n17490,n17491,n17492);
xor (n17491,n17488,n17489);
or (n17492,n17493,n17496);
and (n17493,n17494,n17495);
xor (n17494,n17414,n17415);
and (n17495,n297,n120);
and (n17496,n17497,n17498);
xor (n17497,n17494,n17495);
or (n17498,n17499,n17502);
and (n17499,n17500,n17501);
xor (n17500,n17419,n17420);
and (n17501,n278,n120);
and (n17502,n17503,n17504);
xor (n17503,n17500,n17501);
or (n17504,n17505,n17508);
and (n17505,n17506,n17507);
xor (n17506,n17425,n17426);
and (n17507,n323,n120);
and (n17508,n17509,n17510);
xor (n17509,n17506,n17507);
or (n17510,n17511,n17514);
and (n17511,n17512,n17513);
xor (n17512,n17431,n17432);
and (n17513,n306,n120);
and (n17514,n17515,n17516);
xor (n17515,n17512,n17513);
or (n17516,n17517,n17520);
and (n17517,n17518,n17519);
xor (n17518,n17437,n17438);
and (n17519,n384,n120);
and (n17520,n17521,n17522);
xor (n17521,n17518,n17519);
or (n17522,n17523,n17526);
and (n17523,n17524,n17525);
xor (n17524,n17443,n17444);
and (n17525,n403,n120);
and (n17526,n17527,n17528);
xor (n17527,n17524,n17525);
or (n17528,n17529,n17532);
and (n17529,n17530,n17531);
xor (n17530,n17449,n17450);
and (n17531,n138,n120);
and (n17532,n17533,n17534);
xor (n17533,n17530,n17531);
or (n17534,n17535,n17538);
and (n17535,n17536,n17537);
xor (n17536,n17454,n17455);
and (n17537,n131,n120);
and (n17538,n17539,n17540);
xor (n17539,n17536,n17537);
or (n17540,n17541,n17544);
and (n17541,n17542,n17543);
xor (n17542,n17460,n17461);
and (n17543,n163,n120);
and (n17544,n17545,n17546);
xor (n17545,n17542,n17543);
or (n17546,n17547,n17550);
and (n17547,n17548,n17549);
xor (n17548,n17465,n17466);
and (n17549,n156,n120);
and (n17550,n17551,n17552);
xor (n17551,n17548,n17549);
or (n17552,n17553,n17556);
and (n17553,n17554,n17555);
xor (n17554,n17470,n17471);
and (n17555,n108,n120);
and (n17556,n17557,n17558);
xor (n17557,n17554,n17555);
or (n17558,n17559,n17562);
and (n17559,n17560,n17561);
xor (n17560,n17475,n17476);
and (n17561,n102,n120);
and (n17562,n17563,n17564);
xor (n17563,n17560,n17561);
and (n17564,n17565,n17566);
xor (n17565,n17480,n17481);
and (n17566,n460,n120);
and (n17567,n17568,n17569);
xor (n17568,n16738,n2241);
or (n17569,n17570,n17572);
and (n17570,n17571,n2163);
xor (n17571,n17485,n17486);
and (n17572,n17573,n17574);
xor (n17573,n17571,n2163);
or (n17574,n17575,n17578);
and (n17575,n17576,n17577);
xor (n17576,n17491,n17492);
and (n17577,n297,n119);
and (n17578,n17579,n17580);
xor (n17579,n17576,n17577);
or (n17580,n17581,n17584);
and (n17581,n17582,n17583);
xor (n17582,n17497,n17498);
not (n17583,n1903);
and (n17584,n17585,n17586);
xor (n17585,n17582,n17583);
or (n17586,n17587,n17590);
and (n17587,n17588,n17589);
xor (n17588,n17503,n17504);
not (n17589,n1781);
and (n17590,n17591,n17592);
xor (n17591,n17588,n17589);
or (n17592,n17593,n17595);
and (n17593,n17594,n1607);
xor (n17594,n17509,n17510);
and (n17595,n17596,n17597);
xor (n17596,n17594,n1607);
or (n17597,n17598,n17600);
and (n17598,n17599,n1423);
xor (n17599,n17515,n17516);
and (n17600,n17601,n17602);
xor (n17601,n17599,n1423);
or (n17602,n17603,n17606);
and (n17603,n17604,n17605);
xor (n17604,n17521,n17522);
not (n17605,n1141);
and (n17606,n17607,n17608);
xor (n17607,n17604,n17605);
or (n17608,n17609,n17612);
and (n17609,n17610,n17611);
xor (n17610,n17527,n17528);
and (n17611,n138,n119);
and (n17612,n17613,n17614);
xor (n17613,n17610,n17611);
or (n17614,n17615,n17617);
and (n17615,n17616,n132);
xor (n17616,n17533,n17534);
and (n17617,n17618,n17619);
xor (n17618,n17616,n132);
or (n17619,n17620,n17623);
and (n17620,n17621,n17622);
xor (n17621,n17539,n17540);
and (n17622,n163,n119);
and (n17623,n17624,n17625);
xor (n17624,n17621,n17622);
or (n17625,n17626,n17629);
and (n17626,n17627,n17628);
xor (n17627,n17545,n17546);
and (n17628,n156,n119);
and (n17629,n17630,n17631);
xor (n17630,n17627,n17628);
or (n17631,n17632,n17634);
and (n17632,n17633,n901);
xor (n17633,n17551,n17552);
and (n17634,n17635,n17636);
xor (n17635,n17633,n901);
or (n17636,n17637,n17639);
and (n17637,n17638,n1020);
xor (n17638,n17557,n17558);
and (n17639,n17640,n17641);
xor (n17640,n17638,n1020);
and (n17641,n17642,n1326);
xor (n17642,n17563,n17564);
and (n17643,n240,n147);
and (n17644,n17645,n17646);
xor (n17645,n16735,n17643);
or (n17646,n17647,n17650);
and (n17647,n17648,n17649);
xor (n17648,n17568,n17569);
and (n17649,n234,n147);
and (n17650,n17651,n17652);
xor (n17651,n17648,n17649);
or (n17652,n17653,n17656);
and (n17653,n17654,n17655);
xor (n17654,n17573,n17574);
and (n17655,n297,n147);
and (n17656,n17657,n17658);
xor (n17657,n17654,n17655);
or (n17658,n17659,n17662);
and (n17659,n17660,n17661);
xor (n17660,n17579,n17580);
and (n17661,n278,n147);
and (n17662,n17663,n17664);
xor (n17663,n17660,n17661);
or (n17664,n17665,n17668);
and (n17665,n17666,n17667);
xor (n17666,n17585,n17586);
and (n17667,n323,n147);
and (n17668,n17669,n17670);
xor (n17669,n17666,n17667);
or (n17670,n17671,n17674);
and (n17671,n17672,n17673);
xor (n17672,n17591,n17592);
and (n17673,n306,n147);
and (n17674,n17675,n17676);
xor (n17675,n17672,n17673);
or (n17676,n17677,n17680);
and (n17677,n17678,n17679);
xor (n17678,n17596,n17597);
and (n17679,n384,n147);
and (n17680,n17681,n17682);
xor (n17681,n17678,n17679);
or (n17682,n17683,n17686);
and (n17683,n17684,n17685);
xor (n17684,n17601,n17602);
and (n17685,n403,n147);
and (n17686,n17687,n17688);
xor (n17687,n17684,n17685);
or (n17688,n17689,n17692);
and (n17689,n17690,n17691);
xor (n17690,n17607,n17608);
and (n17691,n138,n147);
and (n17692,n17693,n17694);
xor (n17693,n17690,n17691);
or (n17694,n17695,n17698);
and (n17695,n17696,n17697);
xor (n17696,n17613,n17614);
and (n17697,n131,n147);
and (n17698,n17699,n17700);
xor (n17699,n17696,n17697);
or (n17700,n17701,n17704);
and (n17701,n17702,n17703);
xor (n17702,n17618,n17619);
and (n17703,n163,n147);
and (n17704,n17705,n17706);
xor (n17705,n17702,n17703);
or (n17706,n17707,n17710);
and (n17707,n17708,n17709);
xor (n17708,n17624,n17625);
and (n17709,n156,n147);
and (n17710,n17711,n17712);
xor (n17711,n17708,n17709);
or (n17712,n17713,n17716);
and (n17713,n17714,n17715);
xor (n17714,n17630,n17631);
and (n17715,n108,n147);
and (n17716,n17717,n17718);
xor (n17717,n17714,n17715);
or (n17718,n17719,n17722);
and (n17719,n17720,n17721);
xor (n17720,n17635,n17636);
and (n17721,n102,n147);
and (n17722,n17723,n17724);
xor (n17723,n17720,n17721);
and (n17724,n17725,n17726);
xor (n17725,n17640,n17641);
and (n17726,n460,n147);
and (n17727,n17728,n17729);
xor (n17728,n16732,n2367);
or (n17729,n17730,n17732);
and (n17730,n17731,n2283);
xor (n17731,n17645,n17646);
and (n17732,n17733,n17734);
xor (n17733,n17731,n2283);
or (n17734,n17735,n17737);
and (n17735,n17736,n2256);
xor (n17736,n17651,n17652);
and (n17737,n17738,n17739);
xor (n17738,n17736,n2256);
or (n17739,n17740,n17742);
and (n17740,n17741,n2169);
xor (n17741,n17657,n17658);
and (n17742,n17743,n17744);
xor (n17743,n17741,n2169);
or (n17744,n17745,n17747);
and (n17745,n17746,n2023);
xor (n17746,n17663,n17664);
and (n17747,n17748,n17749);
xor (n17748,n17746,n2023);
or (n17749,n17750,n17753);
and (n17750,n17751,n17752);
xor (n17751,n17669,n17670);
and (n17752,n306,n91);
and (n17753,n17754,n17755);
xor (n17754,n17751,n17752);
or (n17755,n17756,n17759);
and (n17756,n17757,n17758);
xor (n17757,n17675,n17676);
and (n17758,n384,n91);
and (n17759,n17760,n17761);
xor (n17760,n17757,n17758);
or (n17761,n17762,n17765);
and (n17762,n17763,n17764);
xor (n17763,n17681,n17682);
not (n17764,n1614);
and (n17765,n17766,n17767);
xor (n17766,n17763,n17764);
or (n17767,n17768,n17770);
and (n17768,n17769,n1560);
xor (n17769,n17687,n17688);
and (n17770,n17771,n17772);
xor (n17771,n17769,n1560);
or (n17772,n17773,n17775);
and (n17773,n17774,n1148);
xor (n17774,n17693,n17694);
and (n17775,n17776,n17777);
xor (n17776,n17774,n1148);
or (n17777,n17778,n17780);
and (n17778,n17779,n164);
xor (n17779,n17699,n17700);
and (n17780,n17781,n17782);
xor (n17781,n17779,n164);
or (n17782,n17783,n17785);
and (n17783,n17784,n158);
xor (n17784,n17705,n17706);
and (n17785,n17786,n17787);
xor (n17786,n17784,n158);
or (n17787,n17788,n17790);
and (n17788,n17789,n638);
xor (n17789,n17711,n17712);
and (n17790,n17791,n17792);
xor (n17791,n17789,n638);
or (n17792,n17793,n17795);
and (n17793,n17794,n677);
xor (n17794,n17717,n17718);
and (n17795,n17796,n17797);
xor (n17796,n17794,n677);
and (n17797,n17798,n907);
xor (n17798,n17723,n17724);
and (n17799,n240,n92);
and (n17800,n17801,n17802);
xor (n17801,n16729,n17799);
or (n17802,n17803,n17806);
and (n17803,n17804,n17805);
xor (n17804,n17728,n17729);
and (n17805,n234,n92);
and (n17806,n17807,n17808);
xor (n17807,n17804,n17805);
or (n17808,n17809,n17812);
and (n17809,n17810,n17811);
xor (n17810,n17733,n17734);
and (n17811,n297,n92);
and (n17812,n17813,n17814);
xor (n17813,n17810,n17811);
or (n17814,n17815,n17818);
and (n17815,n17816,n17817);
xor (n17816,n17738,n17739);
and (n17817,n278,n92);
and (n17818,n17819,n17820);
xor (n17819,n17816,n17817);
or (n17820,n17821,n17824);
and (n17821,n17822,n17823);
xor (n17822,n17743,n17744);
and (n17823,n323,n92);
and (n17824,n17825,n17826);
xor (n17825,n17822,n17823);
or (n17826,n17827,n17830);
and (n17827,n17828,n17829);
xor (n17828,n17748,n17749);
and (n17829,n306,n92);
and (n17830,n17831,n17832);
xor (n17831,n17828,n17829);
or (n17832,n17833,n17836);
and (n17833,n17834,n17835);
xor (n17834,n17754,n17755);
and (n17835,n384,n92);
and (n17836,n17837,n17838);
xor (n17837,n17834,n17835);
or (n17838,n17839,n17842);
and (n17839,n17840,n17841);
xor (n17840,n17760,n17761);
and (n17841,n403,n92);
and (n17842,n17843,n17844);
xor (n17843,n17840,n17841);
or (n17844,n17845,n17848);
and (n17845,n17846,n17847);
xor (n17846,n17766,n17767);
and (n17847,n138,n92);
and (n17848,n17849,n17850);
xor (n17849,n17846,n17847);
or (n17850,n17851,n17854);
and (n17851,n17852,n17853);
xor (n17852,n17771,n17772);
and (n17853,n131,n92);
and (n17854,n17855,n17856);
xor (n17855,n17852,n17853);
or (n17856,n17857,n17860);
and (n17857,n17858,n17859);
xor (n17858,n17776,n17777);
and (n17859,n163,n92);
and (n17860,n17861,n17862);
xor (n17861,n17858,n17859);
or (n17862,n17863,n17866);
and (n17863,n17864,n17865);
xor (n17864,n17781,n17782);
and (n17865,n156,n92);
and (n17866,n17867,n17868);
xor (n17867,n17864,n17865);
or (n17868,n17869,n17872);
and (n17869,n17870,n17871);
xor (n17870,n17786,n17787);
and (n17871,n108,n92);
and (n17872,n17873,n17874);
xor (n17873,n17870,n17871);
or (n17874,n17875,n17878);
and (n17875,n17876,n17877);
xor (n17876,n17791,n17792);
and (n17877,n102,n92);
and (n17878,n17879,n17880);
xor (n17879,n17876,n17877);
and (n17880,n17881,n17882);
xor (n17881,n17796,n17797);
and (n17882,n460,n92);
and (n17883,n17884,n17885);
xor (n17884,n16726,n2457);
or (n17885,n17886,n17888);
and (n17886,n17887,n2401);
xor (n17887,n17801,n17802);
and (n17888,n17889,n17890);
xor (n17889,n17887,n2401);
or (n17890,n17891,n17893);
and (n17891,n17892,n2397);
xor (n17892,n17807,n17808);
and (n17893,n17894,n17895);
xor (n17894,n17892,n2397);
or (n17895,n17896,n17898);
and (n17896,n17897,n2295);
xor (n17897,n17813,n17814);
and (n17898,n17899,n17900);
xor (n17899,n17897,n2295);
or (n17900,n17901,n17903);
and (n17901,n17902,n2218);
xor (n17902,n17819,n17820);
and (n17903,n17904,n17905);
xor (n17904,n17902,n2218);
or (n17905,n17906,n17909);
and (n17906,n17907,n17908);
xor (n17907,n17825,n17826);
and (n17908,n306,n97);
and (n17909,n17910,n17911);
xor (n17910,n17907,n17908);
or (n17911,n17912,n17914);
and (n17912,n17913,n2040);
xor (n17913,n17831,n17832);
and (n17914,n17915,n17916);
xor (n17915,n17913,n2040);
or (n17916,n17917,n17920);
and (n17917,n17918,n17919);
xor (n17918,n17837,n17838);
and (n17919,n403,n97);
and (n17920,n17921,n17922);
xor (n17921,n17918,n17919);
or (n17922,n17923,n17926);
and (n17923,n17924,n17925);
xor (n17924,n17843,n17844);
and (n17925,n138,n97);
and (n17926,n17927,n17928);
xor (n17927,n17924,n17925);
or (n17928,n17929,n17931);
and (n17929,n17930,n1538);
xor (n17930,n17849,n17850);
and (n17931,n17932,n17933);
xor (n17932,n17930,n1538);
or (n17933,n17934,n17936);
and (n17934,n17935,n1534);
xor (n17935,n17855,n17856);
and (n17936,n17937,n17938);
xor (n17937,n17935,n1534);
or (n17938,n17939,n17941);
and (n17939,n17940,n1101);
xor (n17940,n17861,n17862);
and (n17941,n17942,n17943);
xor (n17942,n17940,n1101);
or (n17943,n17944,n17946);
and (n17944,n17945,n109);
xor (n17945,n17867,n17868);
and (n17946,n17947,n17948);
xor (n17947,n17945,n109);
or (n17948,n17949,n17951);
and (n17949,n17950,n103);
xor (n17950,n17873,n17874);
and (n17951,n17952,n17953);
xor (n17952,n17950,n103);
and (n17953,n17954,n644);
xor (n17954,n17879,n17880);
and (n17955,n17956,n17957);
xor (n17956,n16723,n2457);
or (n17957,n17958,n17960);
and (n17958,n17959,n2401);
xor (n17959,n17884,n17885);
and (n17960,n17961,n17962);
xor (n17961,n17959,n2401);
or (n17962,n17963,n17965);
and (n17963,n17964,n2397);
xor (n17964,n17889,n17890);
and (n17965,n17966,n17967);
xor (n17966,n17964,n2397);
or (n17967,n17968,n17970);
and (n17968,n17969,n2295);
xor (n17969,n17894,n17895);
and (n17970,n17971,n17972);
xor (n17971,n17969,n2295);
or (n17972,n17973,n17975);
and (n17973,n17974,n2218);
xor (n17974,n17899,n17900);
and (n17975,n17976,n17977);
xor (n17976,n17974,n2218);
or (n17977,n17978,n17980);
and (n17978,n17979,n17908);
xor (n17979,n17904,n17905);
and (n17980,n17981,n17982);
xor (n17981,n17979,n17908);
or (n17982,n17983,n17985);
and (n17983,n17984,n2040);
xor (n17984,n17910,n17911);
and (n17985,n17986,n17987);
xor (n17986,n17984,n2040);
or (n17987,n17988,n17990);
and (n17988,n17989,n17919);
xor (n17989,n17915,n17916);
and (n17990,n17991,n17992);
xor (n17991,n17989,n17919);
or (n17992,n17993,n17995);
and (n17993,n17994,n17925);
xor (n17994,n17921,n17922);
and (n17995,n17996,n17997);
xor (n17996,n17994,n17925);
or (n17997,n17998,n18000);
and (n17998,n17999,n1538);
xor (n17999,n17927,n17928);
and (n18000,n18001,n18002);
xor (n18001,n17999,n1538);
or (n18002,n18003,n18005);
and (n18003,n18004,n1534);
xor (n18004,n17932,n17933);
and (n18005,n18006,n18007);
xor (n18006,n18004,n1534);
or (n18007,n18008,n18010);
and (n18008,n18009,n1101);
xor (n18009,n17937,n17938);
and (n18010,n18011,n18012);
xor (n18011,n18009,n1101);
or (n18012,n18013,n18015);
and (n18013,n18014,n109);
xor (n18014,n17942,n17943);
and (n18015,n18016,n18017);
xor (n18016,n18014,n109);
or (n18017,n18018,n18020);
and (n18018,n18019,n103);
xor (n18019,n17947,n17948);
and (n18020,n18021,n18022);
xor (n18021,n18019,n103);
and (n18022,n18023,n644);
xor (n18023,n17952,n17953);
or (n18024,n18025,n18027);
and (n18025,n18026,n2401);
xor (n18026,n17956,n17957);
and (n18027,n18028,n18029);
xor (n18028,n18026,n2401);
or (n18029,n18030,n18032);
and (n18030,n18031,n2397);
xor (n18031,n17961,n17962);
and (n18032,n18033,n18034);
xor (n18033,n18031,n2397);
or (n18034,n18035,n18037);
and (n18035,n18036,n2295);
xor (n18036,n17966,n17967);
and (n18037,n18038,n18039);
xor (n18038,n18036,n2295);
or (n18039,n18040,n18042);
and (n18040,n18041,n2218);
xor (n18041,n17971,n17972);
and (n18042,n18043,n18044);
xor (n18043,n18041,n2218);
or (n18044,n18045,n18047);
and (n18045,n18046,n17908);
xor (n18046,n17976,n17977);
and (n18047,n18048,n18049);
xor (n18048,n18046,n17908);
or (n18049,n18050,n18052);
and (n18050,n18051,n2040);
xor (n18051,n17981,n17982);
and (n18052,n18053,n18054);
xor (n18053,n18051,n2040);
or (n18054,n18055,n18057);
and (n18055,n18056,n17919);
xor (n18056,n17986,n17987);
and (n18057,n18058,n18059);
xor (n18058,n18056,n17919);
or (n18059,n18060,n18062);
and (n18060,n18061,n17925);
xor (n18061,n17991,n17992);
and (n18062,n18063,n18064);
xor (n18063,n18061,n17925);
or (n18064,n18065,n18067);
and (n18065,n18066,n1538);
xor (n18066,n17996,n17997);
and (n18067,n18068,n18069);
xor (n18068,n18066,n1538);
or (n18069,n18070,n18072);
and (n18070,n18071,n1534);
xor (n18071,n18001,n18002);
and (n18072,n18073,n18074);
xor (n18073,n18071,n1534);
or (n18074,n18075,n18077);
and (n18075,n18076,n1101);
xor (n18076,n18006,n18007);
and (n18077,n18078,n18079);
xor (n18078,n18076,n1101);
or (n18079,n18080,n18082);
and (n18080,n18081,n109);
xor (n18081,n18011,n18012);
and (n18082,n18083,n18084);
xor (n18083,n18081,n109);
or (n18084,n18085,n18087);
and (n18085,n18086,n103);
xor (n18086,n18016,n18017);
and (n18087,n18088,n18089);
xor (n18088,n18086,n103);
and (n18089,n18090,n644);
xor (n18090,n18021,n18022);
or (n18091,n18092,n18094);
and (n18092,n18093,n2397);
xor (n18093,n18028,n18029);
and (n18094,n18095,n18096);
xor (n18095,n18093,n2397);
or (n18096,n18097,n18099);
and (n18097,n18098,n2295);
xor (n18098,n18033,n18034);
and (n18099,n18100,n18101);
xor (n18100,n18098,n2295);
or (n18101,n18102,n18104);
and (n18102,n18103,n2218);
xor (n18103,n18038,n18039);
and (n18104,n18105,n18106);
xor (n18105,n18103,n2218);
or (n18106,n18107,n18109);
and (n18107,n18108,n17908);
xor (n18108,n18043,n18044);
and (n18109,n18110,n18111);
xor (n18110,n18108,n17908);
or (n18111,n18112,n18114);
and (n18112,n18113,n2040);
xor (n18113,n18048,n18049);
and (n18114,n18115,n18116);
xor (n18115,n18113,n2040);
or (n18116,n18117,n18119);
and (n18117,n18118,n17919);
xor (n18118,n18053,n18054);
and (n18119,n18120,n18121);
xor (n18120,n18118,n17919);
or (n18121,n18122,n18124);
and (n18122,n18123,n17925);
xor (n18123,n18058,n18059);
and (n18124,n18125,n18126);
xor (n18125,n18123,n17925);
or (n18126,n18127,n18129);
and (n18127,n18128,n1538);
xor (n18128,n18063,n18064);
and (n18129,n18130,n18131);
xor (n18130,n18128,n1538);
or (n18131,n18132,n18134);
and (n18132,n18133,n1534);
xor (n18133,n18068,n18069);
and (n18134,n18135,n18136);
xor (n18135,n18133,n1534);
or (n18136,n18137,n18139);
and (n18137,n18138,n1101);
xor (n18138,n18073,n18074);
and (n18139,n18140,n18141);
xor (n18140,n18138,n1101);
or (n18141,n18142,n18144);
and (n18142,n18143,n109);
xor (n18143,n18078,n18079);
and (n18144,n18145,n18146);
xor (n18145,n18143,n109);
or (n18146,n18147,n18149);
and (n18147,n18148,n103);
xor (n18148,n18083,n18084);
and (n18149,n18150,n18151);
xor (n18150,n18148,n103);
and (n18151,n18152,n644);
xor (n18152,n18088,n18089);
or (n18153,n18154,n18156);
and (n18154,n18155,n2295);
xor (n18155,n18095,n18096);
and (n18156,n18157,n18158);
xor (n18157,n18155,n2295);
or (n18158,n18159,n18161);
and (n18159,n18160,n2218);
xor (n18160,n18100,n18101);
and (n18161,n18162,n18163);
xor (n18162,n18160,n2218);
or (n18163,n18164,n18166);
and (n18164,n18165,n17908);
xor (n18165,n18105,n18106);
and (n18166,n18167,n18168);
xor (n18167,n18165,n17908);
or (n18168,n18169,n18171);
and (n18169,n18170,n2040);
xor (n18170,n18110,n18111);
and (n18171,n18172,n18173);
xor (n18172,n18170,n2040);
or (n18173,n18174,n18176);
and (n18174,n18175,n17919);
xor (n18175,n18115,n18116);
and (n18176,n18177,n18178);
xor (n18177,n18175,n17919);
or (n18178,n18179,n18181);
and (n18179,n18180,n17925);
xor (n18180,n18120,n18121);
and (n18181,n18182,n18183);
xor (n18182,n18180,n17925);
or (n18183,n18184,n18186);
and (n18184,n18185,n1538);
xor (n18185,n18125,n18126);
and (n18186,n18187,n18188);
xor (n18187,n18185,n1538);
or (n18188,n18189,n18191);
and (n18189,n18190,n1534);
xor (n18190,n18130,n18131);
and (n18191,n18192,n18193);
xor (n18192,n18190,n1534);
or (n18193,n18194,n18196);
and (n18194,n18195,n1101);
xor (n18195,n18135,n18136);
and (n18196,n18197,n18198);
xor (n18197,n18195,n1101);
or (n18198,n18199,n18201);
and (n18199,n18200,n109);
xor (n18200,n18140,n18141);
and (n18201,n18202,n18203);
xor (n18202,n18200,n109);
or (n18203,n18204,n18206);
and (n18204,n18205,n103);
xor (n18205,n18145,n18146);
and (n18206,n18207,n18208);
xor (n18207,n18205,n103);
and (n18208,n18209,n644);
xor (n18209,n18150,n18151);
or (n18210,n18211,n18213);
and (n18211,n18212,n2218);
xor (n18212,n18157,n18158);
and (n18213,n18214,n18215);
xor (n18214,n18212,n2218);
or (n18215,n18216,n18218);
and (n18216,n18217,n17908);
xor (n18217,n18162,n18163);
and (n18218,n18219,n18220);
xor (n18219,n18217,n17908);
or (n18220,n18221,n18223);
and (n18221,n18222,n2040);
xor (n18222,n18167,n18168);
and (n18223,n18224,n18225);
xor (n18224,n18222,n2040);
or (n18225,n18226,n18228);
and (n18226,n18227,n17919);
xor (n18227,n18172,n18173);
and (n18228,n18229,n18230);
xor (n18229,n18227,n17919);
or (n18230,n18231,n18233);
and (n18231,n18232,n17925);
xor (n18232,n18177,n18178);
and (n18233,n18234,n18235);
xor (n18234,n18232,n17925);
or (n18235,n18236,n18238);
and (n18236,n18237,n1538);
xor (n18237,n18182,n18183);
and (n18238,n18239,n18240);
xor (n18239,n18237,n1538);
or (n18240,n18241,n18243);
and (n18241,n18242,n1534);
xor (n18242,n18187,n18188);
and (n18243,n18244,n18245);
xor (n18244,n18242,n1534);
or (n18245,n18246,n18248);
and (n18246,n18247,n1101);
xor (n18247,n18192,n18193);
and (n18248,n18249,n18250);
xor (n18249,n18247,n1101);
or (n18250,n18251,n18253);
and (n18251,n18252,n109);
xor (n18252,n18197,n18198);
and (n18253,n18254,n18255);
xor (n18254,n18252,n109);
or (n18255,n18256,n18258);
and (n18256,n18257,n103);
xor (n18257,n18202,n18203);
and (n18258,n18259,n18260);
xor (n18259,n18257,n103);
and (n18260,n18261,n644);
xor (n18261,n18207,n18208);
or (n18262,n18263,n18265);
and (n18263,n18264,n17908);
xor (n18264,n18214,n18215);
and (n18265,n18266,n18267);
xor (n18266,n18264,n17908);
or (n18267,n18268,n18270);
and (n18268,n18269,n2040);
xor (n18269,n18219,n18220);
and (n18270,n18271,n18272);
xor (n18271,n18269,n2040);
or (n18272,n18273,n18275);
and (n18273,n18274,n17919);
xor (n18274,n18224,n18225);
and (n18275,n18276,n18277);
xor (n18276,n18274,n17919);
or (n18277,n18278,n18280);
and (n18278,n18279,n17925);
xor (n18279,n18229,n18230);
and (n18280,n18281,n18282);
xor (n18281,n18279,n17925);
or (n18282,n18283,n18285);
and (n18283,n18284,n1538);
xor (n18284,n18234,n18235);
and (n18285,n18286,n18287);
xor (n18286,n18284,n1538);
or (n18287,n18288,n18290);
and (n18288,n18289,n1534);
xor (n18289,n18239,n18240);
and (n18290,n18291,n18292);
xor (n18291,n18289,n1534);
or (n18292,n18293,n18295);
and (n18293,n18294,n1101);
xor (n18294,n18244,n18245);
and (n18295,n18296,n18297);
xor (n18296,n18294,n1101);
or (n18297,n18298,n18300);
and (n18298,n18299,n109);
xor (n18299,n18249,n18250);
and (n18300,n18301,n18302);
xor (n18301,n18299,n109);
or (n18302,n18303,n18305);
and (n18303,n18304,n103);
xor (n18304,n18254,n18255);
and (n18305,n18306,n18307);
xor (n18306,n18304,n103);
and (n18307,n18308,n644);
xor (n18308,n18259,n18260);
or (n18309,n18310,n18312);
and (n18310,n18311,n2040);
xor (n18311,n18266,n18267);
and (n18312,n18313,n18314);
xor (n18313,n18311,n2040);
or (n18314,n18315,n18317);
and (n18315,n18316,n17919);
xor (n18316,n18271,n18272);
and (n18317,n18318,n18319);
xor (n18318,n18316,n17919);
or (n18319,n18320,n18322);
and (n18320,n18321,n17925);
xor (n18321,n18276,n18277);
and (n18322,n18323,n18324);
xor (n18323,n18321,n17925);
or (n18324,n18325,n18327);
and (n18325,n18326,n1538);
xor (n18326,n18281,n18282);
and (n18327,n18328,n18329);
xor (n18328,n18326,n1538);
or (n18329,n18330,n18332);
and (n18330,n18331,n1534);
xor (n18331,n18286,n18287);
and (n18332,n18333,n18334);
xor (n18333,n18331,n1534);
or (n18334,n18335,n18337);
and (n18335,n18336,n1101);
xor (n18336,n18291,n18292);
and (n18337,n18338,n18339);
xor (n18338,n18336,n1101);
or (n18339,n18340,n18342);
and (n18340,n18341,n109);
xor (n18341,n18296,n18297);
and (n18342,n18343,n18344);
xor (n18343,n18341,n109);
or (n18344,n18345,n18347);
and (n18345,n18346,n103);
xor (n18346,n18301,n18302);
and (n18347,n18348,n18349);
xor (n18348,n18346,n103);
and (n18349,n18350,n644);
xor (n18350,n18306,n18307);
or (n18351,n18352,n18354);
and (n18352,n18353,n17919);
xor (n18353,n18313,n18314);
and (n18354,n18355,n18356);
xor (n18355,n18353,n17919);
or (n18356,n18357,n18359);
and (n18357,n18358,n17925);
xor (n18358,n18318,n18319);
and (n18359,n18360,n18361);
xor (n18360,n18358,n17925);
or (n18361,n18362,n18364);
and (n18362,n18363,n1538);
xor (n18363,n18323,n18324);
and (n18364,n18365,n18366);
xor (n18365,n18363,n1538);
or (n18366,n18367,n18369);
and (n18367,n18368,n1534);
xor (n18368,n18328,n18329);
and (n18369,n18370,n18371);
xor (n18370,n18368,n1534);
or (n18371,n18372,n18374);
and (n18372,n18373,n1101);
xor (n18373,n18333,n18334);
and (n18374,n18375,n18376);
xor (n18375,n18373,n1101);
or (n18376,n18377,n18379);
and (n18377,n18378,n109);
xor (n18378,n18338,n18339);
and (n18379,n18380,n18381);
xor (n18380,n18378,n109);
or (n18381,n18382,n18384);
and (n18382,n18383,n103);
xor (n18383,n18343,n18344);
and (n18384,n18385,n18386);
xor (n18385,n18383,n103);
and (n18386,n18387,n644);
xor (n18387,n18348,n18349);
or (n18388,n18389,n18391);
and (n18389,n18390,n17925);
xor (n18390,n18355,n18356);
and (n18391,n18392,n18393);
xor (n18392,n18390,n17925);
or (n18393,n18394,n18396);
and (n18394,n18395,n1538);
xor (n18395,n18360,n18361);
and (n18396,n18397,n18398);
xor (n18397,n18395,n1538);
or (n18398,n18399,n18401);
and (n18399,n18400,n1534);
xor (n18400,n18365,n18366);
and (n18401,n18402,n18403);
xor (n18402,n18400,n1534);
or (n18403,n18404,n18406);
and (n18404,n18405,n1101);
xor (n18405,n18370,n18371);
and (n18406,n18407,n18408);
xor (n18407,n18405,n1101);
or (n18408,n18409,n18411);
and (n18409,n18410,n109);
xor (n18410,n18375,n18376);
and (n18411,n18412,n18413);
xor (n18412,n18410,n109);
or (n18413,n18414,n18416);
and (n18414,n18415,n103);
xor (n18415,n18380,n18381);
and (n18416,n18417,n18418);
xor (n18417,n18415,n103);
and (n18418,n18419,n644);
xor (n18419,n18385,n18386);
or (n18420,n18421,n18423);
and (n18421,n18422,n1538);
xor (n18422,n18392,n18393);
and (n18423,n18424,n18425);
xor (n18424,n18422,n1538);
or (n18425,n18426,n18428);
and (n18426,n18427,n1534);
xor (n18427,n18397,n18398);
and (n18428,n18429,n18430);
xor (n18429,n18427,n1534);
or (n18430,n18431,n18433);
and (n18431,n18432,n1101);
xor (n18432,n18402,n18403);
and (n18433,n18434,n18435);
xor (n18434,n18432,n1101);
or (n18435,n18436,n18438);
and (n18436,n18437,n109);
xor (n18437,n18407,n18408);
and (n18438,n18439,n18440);
xor (n18439,n18437,n109);
or (n18440,n18441,n18443);
and (n18441,n18442,n103);
xor (n18442,n18412,n18413);
and (n18443,n18444,n18445);
xor (n18444,n18442,n103);
and (n18445,n18446,n644);
xor (n18446,n18417,n18418);
or (n18447,n18448,n18450);
and (n18448,n18449,n1534);
xor (n18449,n18424,n18425);
and (n18450,n18451,n18452);
xor (n18451,n18449,n1534);
or (n18452,n18453,n18455);
and (n18453,n18454,n1101);
xor (n18454,n18429,n18430);
and (n18455,n18456,n18457);
xor (n18456,n18454,n1101);
or (n18457,n18458,n18460);
and (n18458,n18459,n109);
xor (n18459,n18434,n18435);
and (n18460,n18461,n18462);
xor (n18461,n18459,n109);
or (n18462,n18463,n18465);
and (n18463,n18464,n103);
xor (n18464,n18439,n18440);
and (n18465,n18466,n18467);
xor (n18466,n18464,n103);
and (n18467,n18468,n644);
xor (n18468,n18444,n18445);
or (n18469,n18470,n18472);
and (n18470,n18471,n1101);
xor (n18471,n18451,n18452);
and (n18472,n18473,n18474);
xor (n18473,n18471,n1101);
or (n18474,n18475,n18477);
and (n18475,n18476,n109);
xor (n18476,n18456,n18457);
and (n18477,n18478,n18479);
xor (n18478,n18476,n109);
or (n18479,n18480,n18482);
and (n18480,n18481,n103);
xor (n18481,n18461,n18462);
and (n18482,n18483,n18484);
xor (n18483,n18481,n103);
and (n18484,n18485,n644);
xor (n18485,n18466,n18467);
or (n18486,n18487,n18489);
and (n18487,n18488,n109);
xor (n18488,n18473,n18474);
and (n18489,n18490,n18491);
xor (n18490,n18488,n109);
or (n18491,n18492,n18494);
and (n18492,n18493,n103);
xor (n18493,n18478,n18479);
and (n18494,n18495,n18496);
xor (n18495,n18493,n103);
and (n18496,n18497,n644);
xor (n18497,n18483,n18484);
or (n18498,n18499,n18501);
and (n18499,n18500,n103);
xor (n18500,n18490,n18491);
and (n18501,n18502,n18503);
xor (n18502,n18500,n103);
and (n18503,n18504,n644);
xor (n18504,n18495,n18496);
and (n18505,n18506,n644);
xor (n18506,n18502,n18503);
or (n18507,n18508,n18512,n18718);
and (n18508,n18509,n18510);
xor (n18509,n16631,n16079);
not (n18510,n18511);
xor (n18511,n18506,n644);
and (n18512,n18510,n18513);
or (n18513,n18514,n18518,n18717);
and (n18514,n18515,n18516);
xor (n18515,n16629,n16079);
not (n18516,n18517);
xor (n18517,n18504,n644);
and (n18518,n18516,n18519);
or (n18519,n18520,n18524,n18716);
and (n18520,n18521,n18522);
xor (n18521,n16622,n16079);
not (n18522,n18523);
xor (n18523,n18497,n644);
and (n18524,n18522,n18525);
or (n18525,n18526,n18530,n18715);
and (n18526,n18527,n18528);
xor (n18527,n16610,n16079);
not (n18528,n18529);
xor (n18529,n18485,n644);
and (n18530,n18528,n18531);
or (n18531,n18532,n18536,n18714);
and (n18532,n18533,n18534);
xor (n18533,n16593,n16079);
not (n18534,n18535);
xor (n18535,n18468,n644);
and (n18536,n18534,n18537);
or (n18537,n18538,n18542,n18713);
and (n18538,n18539,n18540);
xor (n18539,n16571,n16079);
not (n18540,n18541);
xor (n18541,n18446,n644);
and (n18542,n18540,n18543);
or (n18543,n18544,n18548,n18712);
and (n18544,n18545,n18546);
xor (n18545,n16544,n16079);
not (n18546,n18547);
xor (n18547,n18419,n644);
and (n18548,n18546,n18549);
or (n18549,n18550,n18554,n18711);
and (n18550,n18551,n18552);
xor (n18551,n16512,n16079);
not (n18552,n18553);
xor (n18553,n18387,n644);
and (n18554,n18552,n18555);
or (n18555,n18556,n18560,n18710);
and (n18556,n18557,n18558);
xor (n18557,n16475,n16079);
not (n18558,n18559);
xor (n18559,n18350,n644);
and (n18560,n18558,n18561);
or (n18561,n18562,n18566,n18709);
and (n18562,n18563,n18564);
xor (n18563,n16433,n16079);
not (n18564,n18565);
xor (n18565,n18308,n644);
and (n18566,n18564,n18567);
or (n18567,n18568,n18572,n18708);
and (n18568,n18569,n18570);
xor (n18569,n16386,n16079);
not (n18570,n18571);
xor (n18571,n18261,n644);
and (n18572,n18570,n18573);
or (n18573,n18574,n18578,n18707);
and (n18574,n18575,n18576);
xor (n18575,n16334,n16079);
not (n18576,n18577);
xor (n18577,n18209,n644);
and (n18578,n18576,n18579);
or (n18579,n18580,n18584,n18706);
and (n18580,n18581,n18582);
xor (n18581,n16277,n16079);
not (n18582,n18583);
xor (n18583,n18152,n644);
and (n18584,n18582,n18585);
or (n18585,n18586,n18590,n18705);
and (n18586,n18587,n18588);
xor (n18587,n16215,n16079);
not (n18588,n18589);
xor (n18589,n18090,n644);
and (n18590,n18588,n18591);
or (n18591,n18592,n18596,n18704);
and (n18592,n18593,n18594);
xor (n18593,n16148,n16079);
not (n18594,n18595);
xor (n18595,n18023,n644);
and (n18596,n18594,n18597);
or (n18597,n18598,n18602,n18703);
and (n18598,n18599,n18600);
xor (n18599,n16078,n16079);
not (n18600,n18601);
xor (n18601,n17954,n644);
and (n18602,n18600,n18603);
or (n18603,n18604,n18608,n18702);
and (n18604,n18605,n18606);
xor (n18605,n15998,n451);
not (n18606,n18607);
xor (n18607,n17881,n17882);
and (n18608,n18606,n18609);
or (n18609,n18610,n18614,n18701);
and (n18610,n18611,n18612);
xor (n18611,n15914,n15915);
not (n18612,n18613);
xor (n18613,n17798,n907);
and (n18614,n18612,n18615);
or (n18615,n18616,n18620,n18700);
and (n18616,n18617,n18618);
xor (n18617,n15834,n915);
not (n18618,n18619);
xor (n18619,n17725,n17726);
and (n18620,n18618,n18621);
or (n18621,n18622,n18626,n18699);
and (n18622,n18623,n18624);
xor (n18623,n15751,n1310);
not (n18624,n18625);
xor (n18625,n17642,n1326);
and (n18626,n18624,n18627);
or (n18627,n18628,n18632,n18698);
and (n18628,n18629,n18630);
xor (n18629,n15672,n15673);
not (n18630,n18631);
xor (n18631,n17565,n17566);
and (n18632,n18630,n18633);
or (n18633,n18634,n18638,n18697);
and (n18634,n18635,n18636);
xor (n18635,n15588,n15589);
not (n18636,n18637);
xor (n18637,n17482,n2729);
and (n18638,n18636,n18639);
or (n18639,n18640,n18644,n18696);
and (n18640,n18641,n18642);
xor (n18641,n15512,n2739);
not (n18642,n18643);
xor (n18643,n17406,n17407);
and (n18644,n18642,n18645);
or (n18645,n18646,n18650,n18695);
and (n18646,n18647,n18648);
xor (n18647,n15429,n2960);
not (n18648,n18649);
xor (n18649,n17323,n2979);
and (n18650,n18648,n18651);
or (n18651,n18652,n18656,n18694);
and (n18652,n18653,n18654);
xor (n18653,n15349,n2947);
not (n18654,n18655);
xor (n18655,n17245,n17246);
and (n18656,n18654,n18657);
or (n18657,n18658,n18662,n18693);
and (n18658,n18659,n18660);
xor (n18659,n15265,n15266);
not (n18660,n18661);
xor (n18661,n17162,n3175);
and (n18662,n18660,n18663);
or (n18663,n18664,n18668,n18692);
and (n18664,n18665,n18666);
xor (n18665,n15186,n3124);
not (n18666,n18667);
xor (n18667,n17084,n17085);
and (n18668,n18666,n18669);
or (n18669,n18670,n18674,n18691);
and (n18670,n18671,n18672);
xor (n18671,n15103,n3244);
not (n18672,n18673);
xor (n18673,n17001,n3257);
and (n18674,n18672,n18675);
or (n18675,n18676,n18680,n18690);
and (n18676,n18677,n18678);
xor (n18677,n15023,n3198);
not (n18678,n18679);
xor (n18679,n16924,n16925);
and (n18680,n18678,n18681);
or (n18681,n18682,n18686,n18689);
and (n18682,n18683,n18684);
xor (n18683,n14939,n14940);
not (n18684,n18685);
xor (n18685,n16841,n3331);
and (n18686,n18684,n18687);
or (n18687,n3324,n18688);
not (n18688,n3337);
and (n18689,n18683,n18687);
and (n18690,n18677,n18681);
and (n18691,n18671,n18675);
and (n18692,n18665,n18669);
and (n18693,n18659,n18663);
and (n18694,n18653,n18657);
and (n18695,n18647,n18651);
and (n18696,n18641,n18645);
and (n18697,n18635,n18639);
and (n18698,n18629,n18633);
and (n18699,n18623,n18627);
and (n18700,n18617,n18621);
and (n18701,n18611,n18615);
and (n18702,n18605,n18609);
and (n18703,n18599,n18603);
and (n18704,n18593,n18597);
and (n18705,n18587,n18591);
and (n18706,n18581,n18585);
and (n18707,n18575,n18579);
and (n18708,n18569,n18573);
and (n18709,n18563,n18567);
and (n18710,n18557,n18561);
and (n18711,n18551,n18555);
and (n18712,n18545,n18549);
and (n18713,n18539,n18543);
and (n18714,n18533,n18537);
and (n18715,n18527,n18531);
and (n18716,n18521,n18525);
and (n18717,n18515,n18519);
and (n18718,n18509,n18513);
not (n18719,n18720);
xor (n18720,n18721,n22487);
xor (n18721,n18722,n20616);
xor (n18722,n18723,n7977);
xor (n18723,n18724,n20614);
xor (n18724,n18725,n20059);
xor (n18725,n18726,n20607);
xor (n18726,n18727,n20053);
xor (n18727,n18728,n20595);
xor (n18728,n18729,n20047);
xor (n18729,n18730,n20578);
xor (n18730,n18731,n9004);
xor (n18731,n18732,n20556);
xor (n18732,n18733,n9264);
xor (n18733,n18734,n20529);
xor (n18734,n18735,n20031);
xor (n18735,n18736,n20497);
xor (n18736,n18737,n20025);
xor (n18737,n18738,n20460);
xor (n18738,n18739,n20019);
xor (n18739,n18740,n20418);
xor (n18740,n18741,n20013);
xor (n18741,n18742,n20371);
xor (n18742,n18743,n20007);
xor (n18743,n18744,n20319);
xor (n18744,n18745,n20001);
xor (n18745,n18746,n20262);
xor (n18746,n18747,n19995);
xor (n18747,n18748,n20200);
xor (n18748,n18749,n10287);
xor (n18749,n18750,n20133);
xor (n18750,n18751,n19984);
xor (n18751,n18752,n18812);
xor (n18752,n18753,n18810);
xor (n18753,n18754,n18811);
xor (n18754,n18755,n18810);
xor (n18755,n18756,n18809);
xor (n18756,n18757,n18808);
xor (n18757,n18758,n18807);
xor (n18758,n18759,n18806);
xor (n18759,n18760,n18805);
xor (n18760,n18761,n18804);
xor (n18761,n18762,n18803);
xor (n18762,n18763,n18802);
xor (n18763,n18764,n18801);
xor (n18764,n18765,n18800);
xor (n18765,n18766,n18799);
xor (n18766,n18767,n9989);
xor (n18767,n18768,n18798);
xor (n18768,n18769,n18797);
xor (n18769,n18770,n18796);
xor (n18770,n18771,n18795);
xor (n18771,n18772,n18794);
xor (n18772,n18773,n18793);
xor (n18773,n18774,n18792);
xor (n18774,n18775,n18791);
xor (n18775,n18776,n18790);
xor (n18776,n18777,n18789);
xor (n18777,n18778,n18788);
xor (n18778,n18779,n8936);
xor (n18779,n18780,n18787);
xor (n18780,n18781,n18786);
xor (n18781,n18782,n18785);
xor (n18782,n18783,n18784);
and (n18783,n7867,n7378);
and (n18784,n7867,n7385);
and (n18785,n18783,n18784);
and (n18786,n7867,n7595);
and (n18787,n18781,n18786);
and (n18788,n18779,n8936);
and (n18789,n7867,n7181);
and (n18790,n18777,n18789);
and (n18791,n7867,n7174);
and (n18792,n18775,n18791);
and (n18793,n7867,n7212);
and (n18794,n18773,n18793);
and (n18795,n7867,n7205);
and (n18796,n18771,n18795);
and (n18797,n7867,n7261);
and (n18798,n18769,n18797);
and (n18799,n18767,n9989);
and (n18800,n7867,n7330);
and (n18801,n18765,n18800);
and (n18802,n7867,n7049);
and (n18803,n18763,n18802);
and (n18804,n7867,n7042);
and (n18805,n18761,n18804);
and (n18806,n7867,n7036);
and (n18807,n18759,n18806);
and (n18808,n7867,n7758);
and (n18809,n18757,n18808);
and (n18810,n7867,n7853);
and (n18811,n18755,n18810);
or (n18812,n18813,n20064);
and (n18813,n18814,n19984);
xor (n18814,n18754,n18815);
or (n18815,n18816,n19985);
and (n18816,n18817,n19984);
xor (n18817,n18756,n18818);
or (n18818,n18819,n19902);
and (n18819,n18820,n19901);
xor (n18820,n18758,n18821);
or (n18821,n18822,n19825);
and (n18822,n18823,n19824);
xor (n18823,n18760,n18824);
or (n18824,n18825,n19742);
and (n18825,n18826,n19741);
xor (n18826,n18762,n18827);
or (n18827,n18828,n19665);
and (n18828,n18829,n19664);
xor (n18829,n18764,n18830);
or (n18830,n18831,n19582);
and (n18831,n18832,n19581);
xor (n18832,n18766,n18833);
or (n18833,n18834,n19505);
and (n18834,n18835,n9901);
xor (n18835,n18768,n18836);
or (n18836,n18837,n19423);
and (n18837,n18838,n19422);
xor (n18838,n18770,n18839);
or (n18839,n18840,n19343);
and (n18840,n18841,n9675);
xor (n18841,n18772,n18842);
or (n18842,n18843,n19261);
and (n18843,n18844,n19260);
xor (n18844,n18774,n18845);
or (n18845,n18846,n19180);
and (n18846,n18847,n9014);
xor (n18847,n18776,n18848);
or (n18848,n18849,n19098);
and (n18849,n18850,n19097);
xor (n18850,n18778,n18851);
or (n18851,n18852,n19020);
and (n18852,n18853,n9067);
xor (n18853,n18780,n18854);
or (n18854,n18855,n18938);
and (n18855,n18856,n18937);
xor (n18856,n18782,n18857);
or (n18857,n18858,n18860);
and (n18858,n18783,n18859);
and (n18859,n7745,n7385);
and (n18860,n18861,n18862);
xor (n18861,n18783,n18859);
or (n18862,n18863,n18865);
and (n18863,n18864,n7386);
and (n18864,n7745,n7378);
and (n18865,n18866,n18867);
xor (n18866,n18864,n7386);
or (n18867,n18868,n18870);
and (n18868,n18869,n7392);
and (n18869,n7383,n7378);
and (n18870,n18871,n18872);
xor (n18871,n18869,n7392);
or (n18872,n18873,n18875);
and (n18873,n18874,n7559);
and (n18874,n7391,n7378);
and (n18875,n18876,n18877);
xor (n18876,n18874,n7559);
or (n18877,n18878,n18881);
and (n18878,n18879,n18880);
and (n18879,n7558,n7378);
and (n18880,n7173,n7385);
and (n18881,n18882,n18883);
xor (n18882,n18879,n18880);
or (n18883,n18884,n18886);
and (n18884,n18885,n8126);
and (n18885,n7173,n7378);
and (n18886,n18887,n18888);
xor (n18887,n18885,n8126);
or (n18888,n18889,n18891);
and (n18889,n18890,n8181);
and (n18890,n7194,n7378);
and (n18891,n18892,n18893);
xor (n18892,n18890,n8181);
or (n18893,n18894,n18896);
and (n18894,n18895,n8323);
and (n18895,n7223,n7378);
and (n18896,n18897,n18898);
xor (n18897,n18895,n8323);
or (n18898,n18899,n18902);
and (n18899,n18900,n18901);
and (n18900,n7204,n7378);
and (n18901,n7270,n7385);
and (n18902,n18903,n18904);
xor (n18903,n18900,n18901);
or (n18904,n18905,n18908);
and (n18905,n18906,n18907);
and (n18906,n7270,n7378);
and (n18907,n7251,n7385);
and (n18908,n18909,n18910);
xor (n18909,n18906,n18907);
or (n18910,n18911,n18914);
and (n18911,n18912,n18913);
and (n18912,n7251,n7378);
and (n18913,n7289,n7385);
and (n18914,n18915,n18916);
xor (n18915,n18912,n18913);
or (n18916,n18917,n18920);
and (n18917,n18918,n18919);
and (n18918,n7289,n7378);
and (n18919,n7339,n7385);
and (n18920,n18921,n18922);
xor (n18921,n18918,n18919);
or (n18922,n18923,n18926);
and (n18923,n18924,n18925);
and (n18924,n7339,n7378);
and (n18925,n7055,n7385);
and (n18926,n18927,n18928);
xor (n18927,n18924,n18925);
or (n18928,n18929,n18932);
and (n18929,n18930,n18931);
and (n18930,n7055,n7378);
and (n18931,n7034,n7385);
and (n18932,n18933,n18934);
xor (n18933,n18930,n18931);
and (n18934,n18935,n18936);
and (n18935,n7034,n7378);
and (n18936,n7366,n7385);
and (n18937,n7745,n7595);
and (n18938,n18939,n18940);
xor (n18939,n18856,n18937);
or (n18940,n18941,n18944);
and (n18941,n18942,n18943);
xor (n18942,n18861,n18862);
and (n18943,n7383,n7595);
and (n18944,n18945,n18946);
xor (n18945,n18942,n18943);
or (n18946,n18947,n18950);
and (n18947,n18948,n18949);
xor (n18948,n18866,n18867);
and (n18949,n7391,n7595);
and (n18950,n18951,n18952);
xor (n18951,n18948,n18949);
or (n18952,n18953,n18956);
and (n18953,n18954,n18955);
xor (n18954,n18871,n18872);
and (n18955,n7558,n7595);
and (n18956,n18957,n18958);
xor (n18957,n18954,n18955);
or (n18958,n18959,n18962);
and (n18959,n18960,n18961);
xor (n18960,n18876,n18877);
and (n18961,n7173,n7595);
and (n18962,n18963,n18964);
xor (n18963,n18960,n18961);
or (n18964,n18965,n18968);
and (n18965,n18966,n18967);
xor (n18966,n18882,n18883);
and (n18967,n7194,n7595);
and (n18968,n18969,n18970);
xor (n18969,n18966,n18967);
or (n18970,n18971,n18974);
and (n18971,n18972,n18973);
xor (n18972,n18887,n18888);
and (n18973,n7223,n7595);
and (n18974,n18975,n18976);
xor (n18975,n18972,n18973);
or (n18976,n18977,n18980);
and (n18977,n18978,n18979);
xor (n18978,n18892,n18893);
and (n18979,n7204,n7595);
and (n18980,n18981,n18982);
xor (n18981,n18978,n18979);
or (n18982,n18983,n18986);
and (n18983,n18984,n18985);
xor (n18984,n18897,n18898);
and (n18985,n7270,n7595);
and (n18986,n18987,n18988);
xor (n18987,n18984,n18985);
or (n18988,n18989,n18992);
and (n18989,n18990,n18991);
xor (n18990,n18903,n18904);
and (n18991,n7251,n7595);
and (n18992,n18993,n18994);
xor (n18993,n18990,n18991);
or (n18994,n18995,n18998);
and (n18995,n18996,n18997);
xor (n18996,n18909,n18910);
and (n18997,n7289,n7595);
and (n18998,n18999,n19000);
xor (n18999,n18996,n18997);
or (n19000,n19001,n19004);
and (n19001,n19002,n19003);
xor (n19002,n18915,n18916);
and (n19003,n7339,n7595);
and (n19004,n19005,n19006);
xor (n19005,n19002,n19003);
or (n19006,n19007,n19010);
and (n19007,n19008,n19009);
xor (n19008,n18921,n18922);
and (n19009,n7055,n7595);
and (n19010,n19011,n19012);
xor (n19011,n19008,n19009);
or (n19012,n19013,n19016);
and (n19013,n19014,n19015);
xor (n19014,n18927,n18928);
and (n19015,n7034,n7595);
and (n19016,n19017,n19018);
xor (n19017,n19014,n19015);
and (n19018,n19019,n8745);
xor (n19019,n18933,n18934);
and (n19020,n19021,n19022);
xor (n19021,n18853,n9067);
or (n19022,n19023,n19026);
and (n19023,n19024,n19025);
xor (n19024,n18939,n18940);
and (n19025,n7383,n7180);
and (n19026,n19027,n19028);
xor (n19027,n19024,n19025);
or (n19028,n19029,n19031);
and (n19029,n19030,n7769);
xor (n19030,n18945,n18946);
and (n19031,n19032,n19033);
xor (n19032,n19030,n7769);
or (n19033,n19034,n19037);
and (n19034,n19035,n19036);
xor (n19035,n18951,n18952);
and (n19036,n7558,n7180);
and (n19037,n19038,n19039);
xor (n19038,n19035,n19036);
or (n19039,n19040,n19043);
and (n19040,n19041,n19042);
xor (n19041,n18957,n18958);
and (n19042,n7173,n7180);
and (n19043,n19044,n19045);
xor (n19044,n19041,n19042);
or (n19045,n19046,n19049);
and (n19046,n19047,n19048);
xor (n19047,n18963,n18964);
and (n19048,n7194,n7180);
and (n19049,n19050,n19051);
xor (n19050,n19047,n19048);
or (n19051,n19052,n19054);
and (n19052,n19053,n7590);
xor (n19053,n18969,n18970);
and (n19054,n19055,n19056);
xor (n19055,n19053,n7590);
or (n19056,n19057,n19059);
and (n19057,n19058,n8062);
xor (n19058,n18975,n18976);
and (n19059,n19060,n19061);
xor (n19060,n19058,n8062);
or (n19061,n19062,n19064);
and (n19062,n19063,n8244);
xor (n19063,n18981,n18982);
and (n19064,n19065,n19066);
xor (n19065,n19063,n8244);
or (n19066,n19067,n19070);
and (n19067,n19068,n19069);
xor (n19068,n18987,n18988);
and (n19069,n7251,n7180);
and (n19070,n19071,n19072);
xor (n19071,n19068,n19069);
or (n19072,n19073,n19075);
and (n19073,n19074,n8419);
xor (n19074,n18993,n18994);
and (n19075,n19076,n19077);
xor (n19076,n19074,n8419);
or (n19077,n19078,n19080);
and (n19078,n19079,n8555);
xor (n19079,n18999,n19000);
and (n19080,n19081,n19082);
xor (n19081,n19079,n8555);
or (n19082,n19083,n19086);
and (n19083,n19084,n19085);
xor (n19084,n19005,n19006);
and (n19085,n7055,n7180);
and (n19086,n19087,n19088);
xor (n19087,n19084,n19085);
or (n19088,n19089,n19092);
and (n19089,n19090,n19091);
xor (n19090,n19011,n19012);
and (n19091,n7034,n7180);
and (n19092,n19093,n19094);
xor (n19093,n19090,n19091);
and (n19094,n19095,n19096);
xor (n19095,n19017,n19018);
and (n19096,n7366,n7180);
and (n19097,n7745,n7181);
and (n19098,n19099,n19100);
xor (n19099,n18850,n19097);
or (n19100,n19101,n19104);
and (n19101,n19102,n19103);
xor (n19102,n19021,n19022);
and (n19103,n7383,n7181);
and (n19104,n19105,n19106);
xor (n19105,n19102,n19103);
or (n19106,n19107,n19110);
and (n19107,n19108,n19109);
xor (n19108,n19027,n19028);
and (n19109,n7391,n7181);
and (n19110,n19111,n19112);
xor (n19111,n19108,n19109);
or (n19112,n19113,n19116);
and (n19113,n19114,n19115);
xor (n19114,n19032,n19033);
and (n19115,n7558,n7181);
and (n19116,n19117,n19118);
xor (n19117,n19114,n19115);
or (n19118,n19119,n19122);
and (n19119,n19120,n19121);
xor (n19120,n19038,n19039);
and (n19121,n7173,n7181);
and (n19122,n19123,n19124);
xor (n19123,n19120,n19121);
or (n19124,n19125,n19128);
and (n19125,n19126,n19127);
xor (n19126,n19044,n19045);
and (n19127,n7194,n7181);
and (n19128,n19129,n19130);
xor (n19129,n19126,n19127);
or (n19130,n19131,n19134);
and (n19131,n19132,n19133);
xor (n19132,n19050,n19051);
and (n19133,n7223,n7181);
and (n19134,n19135,n19136);
xor (n19135,n19132,n19133);
or (n19136,n19137,n19140);
and (n19137,n19138,n19139);
xor (n19138,n19055,n19056);
and (n19139,n7204,n7181);
and (n19140,n19141,n19142);
xor (n19141,n19138,n19139);
or (n19142,n19143,n19146);
and (n19143,n19144,n19145);
xor (n19144,n19060,n19061);
and (n19145,n7270,n7181);
and (n19146,n19147,n19148);
xor (n19147,n19144,n19145);
or (n19148,n19149,n19152);
and (n19149,n19150,n19151);
xor (n19150,n19065,n19066);
and (n19151,n7251,n7181);
and (n19152,n19153,n19154);
xor (n19153,n19150,n19151);
or (n19154,n19155,n19158);
and (n19155,n19156,n19157);
xor (n19156,n19071,n19072);
and (n19157,n7289,n7181);
and (n19158,n19159,n19160);
xor (n19159,n19156,n19157);
or (n19160,n19161,n19164);
and (n19161,n19162,n19163);
xor (n19162,n19076,n19077);
and (n19163,n7339,n7181);
and (n19164,n19165,n19166);
xor (n19165,n19162,n19163);
or (n19166,n19167,n19170);
and (n19167,n19168,n19169);
xor (n19168,n19081,n19082);
and (n19169,n7055,n7181);
and (n19170,n19171,n19172);
xor (n19171,n19168,n19169);
or (n19172,n19173,n19176);
and (n19173,n19174,n19175);
xor (n19174,n19087,n19088);
and (n19175,n7034,n7181);
and (n19176,n19177,n19178);
xor (n19177,n19174,n19175);
and (n19178,n19179,n8670);
xor (n19179,n19093,n19094);
and (n19180,n19181,n19182);
xor (n19181,n18847,n9014);
or (n19182,n19183,n19186);
and (n19183,n19184,n19185);
xor (n19184,n19099,n19100);
and (n19185,n7383,n7174);
and (n19186,n19187,n19188);
xor (n19187,n19184,n19185);
or (n19188,n19189,n19192);
and (n19189,n19190,n19191);
xor (n19190,n19105,n19106);
and (n19191,n7391,n7174);
and (n19192,n19193,n19194);
xor (n19193,n19190,n19191);
or (n19194,n19195,n19198);
and (n19195,n19196,n19197);
xor (n19196,n19111,n19112);
and (n19197,n7558,n7174);
and (n19198,n19199,n19200);
xor (n19199,n19196,n19197);
or (n19200,n19201,n19204);
and (n19201,n19202,n19203);
xor (n19202,n19117,n19118);
and (n19203,n7173,n7174);
and (n19204,n19205,n19206);
xor (n19205,n19202,n19203);
or (n19206,n19207,n19210);
and (n19207,n19208,n19209);
xor (n19208,n19123,n19124);
and (n19209,n7194,n7174);
and (n19210,n19211,n19212);
xor (n19211,n19208,n19209);
or (n19212,n19213,n19216);
and (n19213,n19214,n19215);
xor (n19214,n19129,n19130);
and (n19215,n7223,n7174);
and (n19216,n19217,n19218);
xor (n19217,n19214,n19215);
or (n19218,n19219,n19222);
and (n19219,n19220,n19221);
xor (n19220,n19135,n19136);
and (n19221,n7204,n7174);
and (n19222,n19223,n19224);
xor (n19223,n19220,n19221);
or (n19224,n19225,n19228);
and (n19225,n19226,n19227);
xor (n19226,n19141,n19142);
and (n19227,n7270,n7174);
and (n19228,n19229,n19230);
xor (n19229,n19226,n19227);
or (n19230,n19231,n19233);
and (n19231,n19232,n8165);
xor (n19232,n19147,n19148);
and (n19233,n19234,n19235);
xor (n19234,n19232,n8165);
or (n19235,n19236,n19238);
and (n19236,n19237,n8187);
xor (n19237,n19153,n19154);
and (n19238,n19239,n19240);
xor (n19239,n19237,n8187);
or (n19240,n19241,n19243);
and (n19241,n19242,n8340);
xor (n19242,n19159,n19160);
and (n19243,n19244,n19245);
xor (n19244,n19242,n8340);
or (n19245,n19246,n19249);
and (n19246,n19247,n19248);
xor (n19247,n19165,n19166);
and (n19248,n7055,n7174);
and (n19249,n19250,n19251);
xor (n19250,n19247,n19248);
or (n19251,n19252,n19255);
and (n19252,n19253,n19254);
xor (n19253,n19171,n19172);
and (n19254,n7034,n7174);
and (n19255,n19256,n19257);
xor (n19256,n19253,n19254);
and (n19257,n19258,n19259);
xor (n19258,n19177,n19178);
and (n19259,n7366,n7174);
and (n19260,n7745,n7212);
and (n19261,n19262,n19263);
xor (n19262,n18844,n19260);
or (n19263,n19264,n19267);
and (n19264,n19265,n19266);
xor (n19265,n19181,n19182);
and (n19266,n7383,n7212);
and (n19267,n19268,n19269);
xor (n19268,n19265,n19266);
or (n19269,n19270,n19273);
and (n19270,n19271,n19272);
xor (n19271,n19187,n19188);
and (n19272,n7391,n7212);
and (n19273,n19274,n19275);
xor (n19274,n19271,n19272);
or (n19275,n19276,n19279);
and (n19276,n19277,n19278);
xor (n19277,n19193,n19194);
and (n19278,n7558,n7212);
and (n19279,n19280,n19281);
xor (n19280,n19277,n19278);
or (n19281,n19282,n19285);
and (n19282,n19283,n19284);
xor (n19283,n19199,n19200);
and (n19284,n7173,n7212);
and (n19285,n19286,n19287);
xor (n19286,n19283,n19284);
or (n19287,n19288,n19291);
and (n19288,n19289,n19290);
xor (n19289,n19205,n19206);
and (n19290,n7194,n7212);
and (n19291,n19292,n19293);
xor (n19292,n19289,n19290);
or (n19293,n19294,n19297);
and (n19294,n19295,n19296);
xor (n19295,n19211,n19212);
and (n19296,n7223,n7212);
and (n19297,n19298,n19299);
xor (n19298,n19295,n19296);
or (n19299,n19300,n19303);
and (n19300,n19301,n19302);
xor (n19301,n19217,n19218);
and (n19302,n7204,n7212);
and (n19303,n19304,n19305);
xor (n19304,n19301,n19302);
or (n19305,n19306,n19309);
and (n19306,n19307,n19308);
xor (n19307,n19223,n19224);
and (n19308,n7270,n7212);
and (n19309,n19310,n19311);
xor (n19310,n19307,n19308);
or (n19311,n19312,n19315);
and (n19312,n19313,n19314);
xor (n19313,n19229,n19230);
and (n19314,n7251,n7212);
and (n19315,n19316,n19317);
xor (n19316,n19313,n19314);
or (n19317,n19318,n19321);
and (n19318,n19319,n19320);
xor (n19319,n19234,n19235);
and (n19320,n7289,n7212);
and (n19321,n19322,n19323);
xor (n19322,n19319,n19320);
or (n19323,n19324,n19327);
and (n19324,n19325,n19326);
xor (n19325,n19239,n19240);
and (n19326,n7339,n7212);
and (n19327,n19328,n19329);
xor (n19328,n19325,n19326);
or (n19329,n19330,n19333);
and (n19330,n19331,n19332);
xor (n19331,n19244,n19245);
and (n19332,n7055,n7212);
and (n19333,n19334,n19335);
xor (n19334,n19331,n19332);
or (n19335,n19336,n19339);
and (n19336,n19337,n19338);
xor (n19337,n19250,n19251);
and (n19338,n7034,n7212);
and (n19339,n19340,n19341);
xor (n19340,n19337,n19338);
and (n19341,n19342,n8439);
xor (n19342,n19256,n19257);
and (n19343,n19344,n19345);
xor (n19344,n18841,n9675);
or (n19345,n19346,n19348);
and (n19346,n19347,n9346);
xor (n19347,n19262,n19263);
and (n19348,n19349,n19350);
xor (n19349,n19347,n9346);
or (n19350,n19351,n19354);
and (n19351,n19352,n19353);
xor (n19352,n19268,n19269);
and (n19353,n7391,n7205);
and (n19354,n19355,n19356);
xor (n19355,n19352,n19353);
or (n19356,n19357,n19360);
and (n19357,n19358,n19359);
xor (n19358,n19274,n19275);
and (n19359,n7558,n7205);
and (n19360,n19361,n19362);
xor (n19361,n19358,n19359);
or (n19362,n19363,n19366);
and (n19363,n19364,n19365);
xor (n19364,n19280,n19281);
and (n19365,n7173,n7205);
and (n19366,n19367,n19368);
xor (n19367,n19364,n19365);
or (n19368,n19369,n19372);
and (n19369,n19370,n19371);
xor (n19370,n19286,n19287);
and (n19371,n7194,n7205);
and (n19372,n19373,n19374);
xor (n19373,n19370,n19371);
or (n19374,n19375,n19377);
and (n19375,n19376,n7224);
xor (n19376,n19292,n19293);
and (n19377,n19378,n19379);
xor (n19378,n19376,n7224);
or (n19379,n19380,n19383);
and (n19380,n19381,n19382);
xor (n19381,n19298,n19299);
and (n19382,n7204,n7205);
and (n19383,n19384,n19385);
xor (n19384,n19381,n19382);
or (n19385,n19386,n19389);
and (n19386,n19387,n19388);
xor (n19387,n19304,n19305);
and (n19388,n7270,n7205);
and (n19389,n19390,n19391);
xor (n19390,n19387,n19388);
or (n19391,n19392,n19395);
and (n19392,n19393,n19394);
xor (n19393,n19310,n19311);
and (n19394,n7251,n7205);
and (n19395,n19396,n19397);
xor (n19396,n19393,n19394);
or (n19397,n19398,n19400);
and (n19398,n19399,n7417);
xor (n19399,n19316,n19317);
and (n19400,n19401,n19402);
xor (n19401,n19399,n7417);
or (n19402,n19403,n19406);
and (n19403,n19404,n19405);
xor (n19404,n19322,n19323);
and (n19405,n7339,n7205);
and (n19406,n19407,n19408);
xor (n19407,n19404,n19405);
or (n19408,n19409,n19412);
and (n19409,n19410,n19411);
xor (n19410,n19328,n19329);
and (n19411,n7055,n7205);
and (n19412,n19413,n19414);
xor (n19413,n19410,n19411);
or (n19414,n19415,n19417);
and (n19415,n19416,n8383);
xor (n19416,n19334,n19335);
and (n19417,n19418,n19419);
xor (n19418,n19416,n8383);
and (n19419,n19420,n19421);
xor (n19420,n19340,n19341);
and (n19421,n7366,n7205);
and (n19422,n7745,n7261);
and (n19423,n19424,n19425);
xor (n19424,n18838,n19422);
or (n19425,n19426,n19429);
and (n19426,n19427,n19428);
xor (n19427,n19344,n19345);
and (n19428,n7383,n7261);
and (n19429,n19430,n19431);
xor (n19430,n19427,n19428);
or (n19431,n19432,n19435);
and (n19432,n19433,n19434);
xor (n19433,n19349,n19350);
and (n19434,n7391,n7261);
and (n19435,n19436,n19437);
xor (n19436,n19433,n19434);
or (n19437,n19438,n19441);
and (n19438,n19439,n19440);
xor (n19439,n19355,n19356);
and (n19440,n7558,n7261);
and (n19441,n19442,n19443);
xor (n19442,n19439,n19440);
or (n19443,n19444,n19447);
and (n19444,n19445,n19446);
xor (n19445,n19361,n19362);
and (n19446,n7173,n7261);
and (n19447,n19448,n19449);
xor (n19448,n19445,n19446);
or (n19449,n19450,n19453);
and (n19450,n19451,n19452);
xor (n19451,n19367,n19368);
and (n19452,n7194,n7261);
and (n19453,n19454,n19455);
xor (n19454,n19451,n19452);
or (n19455,n19456,n19459);
and (n19456,n19457,n19458);
xor (n19457,n19373,n19374);
and (n19458,n7223,n7261);
and (n19459,n19460,n19461);
xor (n19460,n19457,n19458);
or (n19461,n19462,n19465);
and (n19462,n19463,n19464);
xor (n19463,n19378,n19379);
and (n19464,n7204,n7261);
and (n19465,n19466,n19467);
xor (n19466,n19463,n19464);
or (n19467,n19468,n19471);
and (n19468,n19469,n19470);
xor (n19469,n19384,n19385);
and (n19470,n7270,n7261);
and (n19471,n19472,n19473);
xor (n19472,n19469,n19470);
or (n19473,n19474,n19477);
and (n19474,n19475,n19476);
xor (n19475,n19390,n19391);
and (n19476,n7251,n7261);
and (n19477,n19478,n19479);
xor (n19478,n19475,n19476);
or (n19479,n19480,n19483);
and (n19480,n19481,n19482);
xor (n19481,n19396,n19397);
and (n19482,n7289,n7261);
and (n19483,n19484,n19485);
xor (n19484,n19481,n19482);
or (n19485,n19486,n19489);
and (n19486,n19487,n19488);
xor (n19487,n19401,n19402);
and (n19488,n7339,n7261);
and (n19489,n19490,n19491);
xor (n19490,n19487,n19488);
or (n19491,n19492,n19495);
and (n19492,n19493,n19494);
xor (n19493,n19407,n19408);
and (n19494,n7055,n7261);
and (n19495,n19496,n19497);
xor (n19496,n19493,n19494);
or (n19497,n19498,n19501);
and (n19498,n19499,n19500);
xor (n19499,n19413,n19414);
and (n19500,n7034,n7261);
and (n19501,n19502,n19503);
xor (n19502,n19499,n19500);
and (n19503,n19504,n8232);
xor (n19504,n19418,n19419);
and (n19505,n19506,n19507);
xor (n19506,n18835,n9901);
or (n19507,n19508,n19511);
and (n19508,n19509,n19510);
xor (n19509,n19424,n19425);
and (n19510,n7383,n7253);
and (n19511,n19512,n19513);
xor (n19512,n19509,n19510);
or (n19513,n19514,n19516);
and (n19514,n19515,n9602);
xor (n19515,n19430,n19431);
and (n19516,n19517,n19518);
xor (n19517,n19515,n9602);
or (n19518,n19519,n19521);
and (n19519,n19520,n9376);
xor (n19520,n19436,n19437);
and (n19521,n19522,n19523);
xor (n19522,n19520,n9376);
or (n19523,n19524,n19527);
and (n19524,n19525,n19526);
xor (n19525,n19442,n19443);
and (n19526,n7173,n7253);
and (n19527,n19528,n19529);
xor (n19528,n19525,n19526);
or (n19529,n19530,n19533);
and (n19530,n19531,n19532);
xor (n19531,n19448,n19449);
and (n19532,n7194,n7253);
and (n19533,n19534,n19535);
xor (n19534,n19531,n19532);
or (n19535,n19536,n19539);
and (n19536,n19537,n19538);
xor (n19537,n19454,n19455);
and (n19538,n7223,n7253);
and (n19539,n19540,n19541);
xor (n19540,n19537,n19538);
or (n19541,n19542,n19545);
and (n19542,n19543,n19544);
xor (n19543,n19460,n19461);
and (n19544,n7204,n7253);
and (n19545,n19546,n19547);
xor (n19546,n19543,n19544);
or (n19547,n19548,n19551);
and (n19548,n19549,n19550);
xor (n19549,n19466,n19467);
and (n19550,n7270,n7253);
and (n19551,n19552,n19553);
xor (n19552,n19549,n19550);
or (n19553,n19554,n19556);
and (n19554,n19555,n7254);
xor (n19555,n19472,n19473);
and (n19556,n19557,n19558);
xor (n19557,n19555,n7254);
or (n19558,n19559,n19561);
and (n19559,n19560,n7290);
xor (n19560,n19478,n19479);
and (n19561,n19562,n19563);
xor (n19562,n19560,n7290);
or (n19563,n19564,n19566);
and (n19564,n19565,n7456);
xor (n19565,n19484,n19485);
and (n19566,n19567,n19568);
xor (n19567,n19565,n7456);
or (n19568,n19569,n19571);
and (n19569,n19570,n7452);
xor (n19570,n19490,n19491);
and (n19571,n19572,n19573);
xor (n19572,n19570,n7452);
or (n19573,n19574,n19577);
and (n19574,n19575,n19576);
xor (n19575,n19496,n19497);
and (n19576,n7034,n7253);
and (n19577,n19578,n19579);
xor (n19578,n19575,n19576);
and (n19579,n19580,n8209);
xor (n19580,n19502,n19503);
and (n19581,n7745,n7330);
and (n19582,n19583,n19584);
xor (n19583,n18832,n19581);
or (n19584,n19585,n19588);
and (n19585,n19586,n19587);
xor (n19586,n19506,n19507);
and (n19587,n7383,n7330);
and (n19588,n19589,n19590);
xor (n19589,n19586,n19587);
or (n19590,n19591,n19594);
and (n19591,n19592,n19593);
xor (n19592,n19512,n19513);
and (n19593,n7391,n7330);
and (n19594,n19595,n19596);
xor (n19595,n19592,n19593);
or (n19596,n19597,n19600);
and (n19597,n19598,n19599);
xor (n19598,n19517,n19518);
and (n19599,n7558,n7330);
and (n19600,n19601,n19602);
xor (n19601,n19598,n19599);
or (n19602,n19603,n19606);
and (n19603,n19604,n19605);
xor (n19604,n19522,n19523);
and (n19605,n7173,n7330);
and (n19606,n19607,n19608);
xor (n19607,n19604,n19605);
or (n19608,n19609,n19612);
and (n19609,n19610,n19611);
xor (n19610,n19528,n19529);
and (n19611,n7194,n7330);
and (n19612,n19613,n19614);
xor (n19613,n19610,n19611);
or (n19614,n19615,n19618);
and (n19615,n19616,n19617);
xor (n19616,n19534,n19535);
and (n19617,n7223,n7330);
and (n19618,n19619,n19620);
xor (n19619,n19616,n19617);
or (n19620,n19621,n19624);
and (n19621,n19622,n19623);
xor (n19622,n19540,n19541);
and (n19623,n7204,n7330);
and (n19624,n19625,n19626);
xor (n19625,n19622,n19623);
or (n19626,n19627,n19630);
and (n19627,n19628,n19629);
xor (n19628,n19546,n19547);
and (n19629,n7270,n7330);
and (n19630,n19631,n19632);
xor (n19631,n19628,n19629);
or (n19632,n19633,n19636);
and (n19633,n19634,n19635);
xor (n19634,n19552,n19553);
and (n19635,n7251,n7330);
and (n19636,n19637,n19638);
xor (n19637,n19634,n19635);
or (n19638,n19639,n19642);
and (n19639,n19640,n19641);
xor (n19640,n19557,n19558);
and (n19641,n7289,n7330);
and (n19642,n19643,n19644);
xor (n19643,n19640,n19641);
or (n19644,n19645,n19648);
and (n19645,n19646,n19647);
xor (n19646,n19562,n19563);
and (n19647,n7339,n7330);
and (n19648,n19649,n19650);
xor (n19649,n19646,n19647);
or (n19650,n19651,n19654);
and (n19651,n19652,n19653);
xor (n19652,n19567,n19568);
and (n19653,n7055,n7330);
and (n19654,n19655,n19656);
xor (n19655,n19652,n19653);
or (n19656,n19657,n19660);
and (n19657,n19658,n19659);
xor (n19658,n19572,n19573);
and (n19659,n7034,n7330);
and (n19660,n19661,n19662);
xor (n19661,n19658,n19659);
and (n19662,n19663,n7577);
xor (n19663,n19578,n19579);
and (n19664,n7745,n7049);
and (n19665,n19666,n19667);
xor (n19666,n18829,n19664);
or (n19667,n19668,n19670);
and (n19668,n19669,n9996);
xor (n19669,n19583,n19584);
and (n19670,n19671,n19672);
xor (n19671,n19669,n9996);
or (n19672,n19673,n19675);
and (n19673,n19674,n9927);
xor (n19674,n19589,n19590);
and (n19675,n19676,n19677);
xor (n19676,n19674,n9927);
or (n19677,n19678,n19680);
and (n19678,n19679,n9801);
xor (n19679,n19595,n19596);
and (n19680,n19681,n19682);
xor (n19681,n19679,n9801);
or (n19682,n19683,n19685);
and (n19683,n19684,n9620);
xor (n19684,n19601,n19602);
and (n19685,n19686,n19687);
xor (n19686,n19684,n9620);
or (n19687,n19688,n19690);
and (n19688,n19689,n9353);
xor (n19689,n19607,n19608);
and (n19690,n19691,n19692);
xor (n19691,n19689,n9353);
or (n19692,n19693,n19696);
and (n19693,n19694,n19695);
xor (n19694,n19613,n19614);
and (n19695,n7223,n7049);
and (n19696,n19697,n19698);
xor (n19697,n19694,n19695);
or (n19698,n19699,n19702);
and (n19699,n19700,n19701);
xor (n19700,n19619,n19620);
and (n19701,n7204,n7049);
and (n19702,n19703,n19704);
xor (n19703,n19700,n19701);
or (n19704,n19705,n19707);
and (n19705,n19706,n9141);
xor (n19706,n19625,n19626);
and (n19707,n19708,n19709);
xor (n19708,n19706,n9141);
or (n19709,n19710,n19713);
and (n19710,n19711,n19712);
xor (n19711,n19631,n19632);
and (n19712,n7251,n7049);
and (n19713,n19714,n19715);
xor (n19714,n19711,n19712);
or (n19715,n19716,n19719);
and (n19716,n19717,n19718);
xor (n19717,n19637,n19638);
and (n19718,n7289,n7049);
and (n19719,n19720,n19721);
xor (n19720,n19717,n19718);
or (n19721,n19722,n19725);
and (n19722,n19723,n19724);
xor (n19723,n19643,n19644);
and (n19724,n7339,n7049);
and (n19725,n19726,n19727);
xor (n19726,n19723,n19724);
or (n19727,n19728,n19730);
and (n19728,n19729,n7324);
xor (n19729,n19649,n19650);
and (n19730,n19731,n19732);
xor (n19731,n19729,n7324);
or (n19732,n19733,n19736);
and (n19733,n19734,n19735);
xor (n19734,n19655,n19656);
and (n19735,n7034,n7049);
and (n19736,n19737,n19738);
xor (n19737,n19734,n19735);
and (n19738,n19739,n19740);
xor (n19739,n19661,n19662);
and (n19740,n7366,n7049);
and (n19741,n7745,n7042);
and (n19742,n19743,n19744);
xor (n19743,n18826,n19741);
or (n19744,n19745,n19748);
and (n19745,n19746,n19747);
xor (n19746,n19666,n19667);
and (n19747,n7383,n7042);
and (n19748,n19749,n19750);
xor (n19749,n19746,n19747);
or (n19750,n19751,n19754);
and (n19751,n19752,n19753);
xor (n19752,n19671,n19672);
and (n19753,n7391,n7042);
and (n19754,n19755,n19756);
xor (n19755,n19752,n19753);
or (n19756,n19757,n19760);
and (n19757,n19758,n19759);
xor (n19758,n19676,n19677);
and (n19759,n7558,n7042);
and (n19760,n19761,n19762);
xor (n19761,n19758,n19759);
or (n19762,n19763,n19766);
and (n19763,n19764,n19765);
xor (n19764,n19681,n19682);
and (n19765,n7173,n7042);
and (n19766,n19767,n19768);
xor (n19767,n19764,n19765);
or (n19768,n19769,n19772);
and (n19769,n19770,n19771);
xor (n19770,n19686,n19687);
and (n19771,n7194,n7042);
and (n19772,n19773,n19774);
xor (n19773,n19770,n19771);
or (n19774,n19775,n19778);
and (n19775,n19776,n19777);
xor (n19776,n19691,n19692);
and (n19777,n7223,n7042);
and (n19778,n19779,n19780);
xor (n19779,n19776,n19777);
or (n19780,n19781,n19784);
and (n19781,n19782,n19783);
xor (n19782,n19697,n19698);
and (n19783,n7204,n7042);
and (n19784,n19785,n19786);
xor (n19785,n19782,n19783);
or (n19786,n19787,n19790);
and (n19787,n19788,n19789);
xor (n19788,n19703,n19704);
and (n19789,n7270,n7042);
and (n19790,n19791,n19792);
xor (n19791,n19788,n19789);
or (n19792,n19793,n19796);
and (n19793,n19794,n19795);
xor (n19794,n19708,n19709);
and (n19795,n7251,n7042);
and (n19796,n19797,n19798);
xor (n19797,n19794,n19795);
or (n19798,n19799,n19802);
and (n19799,n19800,n19801);
xor (n19800,n19714,n19715);
and (n19801,n7289,n7042);
and (n19802,n19803,n19804);
xor (n19803,n19800,n19801);
or (n19804,n19805,n19808);
and (n19805,n19806,n19807);
xor (n19806,n19720,n19721);
and (n19807,n7339,n7042);
and (n19808,n19809,n19810);
xor (n19809,n19806,n19807);
or (n19810,n19811,n19814);
and (n19811,n19812,n19813);
xor (n19812,n19726,n19727);
and (n19813,n7055,n7042);
and (n19814,n19815,n19816);
xor (n19815,n19812,n19813);
or (n19816,n19817,n19820);
and (n19817,n19818,n19819);
xor (n19818,n19731,n19732);
and (n19819,n7034,n7042);
and (n19820,n19821,n19822);
xor (n19821,n19818,n19819);
and (n19822,n19823,n7365);
xor (n19823,n19737,n19738);
and (n19824,n7745,n7036);
and (n19825,n19826,n19827);
xor (n19826,n18823,n19824);
or (n19827,n19828,n19831);
and (n19828,n19829,n19830);
xor (n19829,n19743,n19744);
and (n19830,n7383,n7036);
and (n19831,n19832,n19833);
xor (n19832,n19829,n19830);
or (n19833,n19834,n19837);
and (n19834,n19835,n19836);
xor (n19835,n19749,n19750);
and (n19836,n7391,n7036);
and (n19837,n19838,n19839);
xor (n19838,n19835,n19836);
or (n19839,n19840,n19843);
and (n19840,n19841,n19842);
xor (n19841,n19755,n19756);
and (n19842,n7558,n7036);
and (n19843,n19844,n19845);
xor (n19844,n19841,n19842);
or (n19845,n19846,n19848);
and (n19846,n19847,n9877);
xor (n19847,n19761,n19762);
and (n19848,n19849,n19850);
xor (n19849,n19847,n9877);
or (n19850,n19851,n19854);
and (n19851,n19852,n19853);
xor (n19852,n19767,n19768);
and (n19853,n7194,n7036);
and (n19854,n19855,n19856);
xor (n19855,n19852,n19853);
or (n19856,n19857,n19859);
and (n19857,n19858,n9643);
xor (n19858,n19773,n19774);
and (n19859,n19860,n19861);
xor (n19860,n19858,n9643);
or (n19861,n19862,n19864);
and (n19862,n19863,n9400);
xor (n19863,n19779,n19780);
and (n19864,n19865,n19866);
xor (n19865,n19863,n9400);
or (n19866,n19867,n19869);
and (n19867,n19868,n8946);
xor (n19868,n19785,n19786);
and (n19869,n19870,n19871);
xor (n19870,n19868,n8946);
or (n19871,n19872,n19875);
and (n19872,n19873,n19874);
xor (n19873,n19791,n19792);
and (n19874,n7251,n7036);
and (n19875,n19876,n19877);
xor (n19876,n19873,n19874);
or (n19877,n19878,n19881);
and (n19878,n19879,n19880);
xor (n19879,n19797,n19798);
and (n19880,n7289,n7036);
and (n19881,n19882,n19883);
xor (n19882,n19879,n19880);
or (n19883,n19884,n19886);
and (n19884,n19885,n7892);
xor (n19885,n19803,n19804);
and (n19886,n19887,n19888);
xor (n19887,n19885,n7892);
or (n19888,n19889,n19891);
and (n19889,n19890,n7056);
xor (n19890,n19809,n19810);
and (n19891,n19892,n19893);
xor (n19892,n19890,n7056);
or (n19893,n19894,n19896);
and (n19894,n19895,n7037);
xor (n19895,n19815,n19816);
and (n19896,n19897,n19898);
xor (n19897,n19895,n7037);
and (n19898,n19899,n19900);
xor (n19899,n19821,n19822);
and (n19900,n7366,n7036);
and (n19901,n7745,n7758);
and (n19902,n19903,n19904);
xor (n19903,n18820,n19901);
or (n19904,n19905,n19908);
and (n19905,n19906,n19907);
xor (n19906,n19826,n19827);
and (n19907,n7383,n7758);
and (n19908,n19909,n19910);
xor (n19909,n19906,n19907);
or (n19910,n19911,n19914);
and (n19911,n19912,n19913);
xor (n19912,n19832,n19833);
and (n19913,n7391,n7758);
and (n19914,n19915,n19916);
xor (n19915,n19912,n19913);
or (n19916,n19917,n19920);
and (n19917,n19918,n19919);
xor (n19918,n19838,n19839);
and (n19919,n7558,n7758);
and (n19920,n19921,n19922);
xor (n19921,n19918,n19919);
or (n19922,n19923,n19926);
and (n19923,n19924,n19925);
xor (n19924,n19844,n19845);
and (n19925,n7173,n7758);
and (n19926,n19927,n19928);
xor (n19927,n19924,n19925);
or (n19928,n19929,n19932);
and (n19929,n19930,n19931);
xor (n19930,n19849,n19850);
and (n19931,n7194,n7758);
and (n19932,n19933,n19934);
xor (n19933,n19930,n19931);
or (n19934,n19935,n19938);
and (n19935,n19936,n19937);
xor (n19936,n19855,n19856);
and (n19937,n7223,n7758);
and (n19938,n19939,n19940);
xor (n19939,n19936,n19937);
or (n19940,n19941,n19944);
and (n19941,n19942,n19943);
xor (n19942,n19860,n19861);
and (n19943,n7204,n7758);
and (n19944,n19945,n19946);
xor (n19945,n19942,n19943);
or (n19946,n19947,n19950);
and (n19947,n19948,n19949);
xor (n19948,n19865,n19866);
and (n19949,n7270,n7758);
and (n19950,n19951,n19952);
xor (n19951,n19948,n19949);
or (n19952,n19953,n19956);
and (n19953,n19954,n19955);
xor (n19954,n19870,n19871);
and (n19955,n7251,n7758);
and (n19956,n19957,n19958);
xor (n19957,n19954,n19955);
or (n19958,n19959,n19962);
and (n19959,n19960,n19961);
xor (n19960,n19876,n19877);
and (n19961,n7289,n7758);
and (n19962,n19963,n19964);
xor (n19963,n19960,n19961);
or (n19964,n19965,n19968);
and (n19965,n19966,n19967);
xor (n19966,n19882,n19883);
and (n19967,n7339,n7758);
and (n19968,n19969,n19970);
xor (n19969,n19966,n19967);
or (n19970,n19971,n19974);
and (n19971,n19972,n19973);
xor (n19972,n19887,n19888);
and (n19973,n7055,n7758);
and (n19974,n19975,n19976);
xor (n19975,n19972,n19973);
or (n19976,n19977,n19980);
and (n19977,n19978,n19979);
xor (n19978,n19892,n19893);
and (n19979,n7034,n7758);
and (n19980,n19981,n19982);
xor (n19981,n19978,n19979);
and (n19982,n19983,n7849);
xor (n19983,n19897,n19898);
and (n19984,n7745,n7853);
and (n19985,n19986,n19987);
xor (n19986,n18817,n19984);
or (n19987,n19988,n19990);
and (n19988,n19989,n10287);
xor (n19989,n19903,n19904);
and (n19990,n19991,n19992);
xor (n19991,n19989,n10287);
or (n19992,n19993,n19996);
and (n19993,n19994,n19995);
xor (n19994,n19909,n19910);
and (n19995,n7391,n7853);
and (n19996,n19997,n19998);
xor (n19997,n19994,n19995);
or (n19998,n19999,n20002);
and (n19999,n20000,n20001);
xor (n20000,n19915,n19916);
and (n20001,n7558,n7853);
and (n20002,n20003,n20004);
xor (n20003,n20000,n20001);
or (n20004,n20005,n20008);
and (n20005,n20006,n20007);
xor (n20006,n19921,n19922);
and (n20007,n7173,n7853);
and (n20008,n20009,n20010);
xor (n20009,n20006,n20007);
or (n20010,n20011,n20014);
and (n20011,n20012,n20013);
xor (n20012,n19927,n19928);
and (n20013,n7194,n7853);
and (n20014,n20015,n20016);
xor (n20015,n20012,n20013);
or (n20016,n20017,n20020);
and (n20017,n20018,n20019);
xor (n20018,n19933,n19934);
and (n20019,n7223,n7853);
and (n20020,n20021,n20022);
xor (n20021,n20018,n20019);
or (n20022,n20023,n20026);
and (n20023,n20024,n20025);
xor (n20024,n19939,n19940);
and (n20025,n7204,n7853);
and (n20026,n20027,n20028);
xor (n20027,n20024,n20025);
or (n20028,n20029,n20032);
and (n20029,n20030,n20031);
xor (n20030,n19945,n19946);
and (n20031,n7270,n7853);
and (n20032,n20033,n20034);
xor (n20033,n20030,n20031);
or (n20034,n20035,n20037);
and (n20035,n20036,n9264);
xor (n20036,n19951,n19952);
and (n20037,n20038,n20039);
xor (n20038,n20036,n9264);
or (n20039,n20040,n20042);
and (n20040,n20041,n9004);
xor (n20041,n19957,n19958);
and (n20042,n20043,n20044);
xor (n20043,n20041,n9004);
or (n20044,n20045,n20048);
and (n20045,n20046,n20047);
xor (n20046,n19963,n19964);
and (n20047,n7339,n7853);
and (n20048,n20049,n20050);
xor (n20049,n20046,n20047);
or (n20050,n20051,n20054);
and (n20051,n20052,n20053);
xor (n20052,n19969,n19970);
and (n20053,n7055,n7853);
and (n20054,n20055,n20056);
xor (n20055,n20052,n20053);
or (n20056,n20057,n20060);
and (n20057,n20058,n20059);
xor (n20058,n19975,n19976);
and (n20059,n7034,n7853);
and (n20060,n20061,n20062);
xor (n20061,n20058,n20059);
and (n20062,n20063,n7977);
xor (n20063,n19981,n19982);
and (n20064,n20065,n20066);
xor (n20065,n18814,n19984);
or (n20066,n20067,n20069);
and (n20067,n20068,n10287);
xor (n20068,n19986,n19987);
and (n20069,n20070,n20071);
xor (n20070,n20068,n10287);
or (n20071,n20072,n20074);
and (n20072,n20073,n19995);
xor (n20073,n19991,n19992);
and (n20074,n20075,n20076);
xor (n20075,n20073,n19995);
or (n20076,n20077,n20079);
and (n20077,n20078,n20001);
xor (n20078,n19997,n19998);
and (n20079,n20080,n20081);
xor (n20080,n20078,n20001);
or (n20081,n20082,n20084);
and (n20082,n20083,n20007);
xor (n20083,n20003,n20004);
and (n20084,n20085,n20086);
xor (n20085,n20083,n20007);
or (n20086,n20087,n20089);
and (n20087,n20088,n20013);
xor (n20088,n20009,n20010);
and (n20089,n20090,n20091);
xor (n20090,n20088,n20013);
or (n20091,n20092,n20094);
and (n20092,n20093,n20019);
xor (n20093,n20015,n20016);
and (n20094,n20095,n20096);
xor (n20095,n20093,n20019);
or (n20096,n20097,n20099);
and (n20097,n20098,n20025);
xor (n20098,n20021,n20022);
and (n20099,n20100,n20101);
xor (n20100,n20098,n20025);
or (n20101,n20102,n20104);
and (n20102,n20103,n20031);
xor (n20103,n20027,n20028);
and (n20104,n20105,n20106);
xor (n20105,n20103,n20031);
or (n20106,n20107,n20109);
and (n20107,n20108,n9264);
xor (n20108,n20033,n20034);
and (n20109,n20110,n20111);
xor (n20110,n20108,n9264);
or (n20111,n20112,n20114);
and (n20112,n20113,n9004);
xor (n20113,n20038,n20039);
and (n20114,n20115,n20116);
xor (n20115,n20113,n9004);
or (n20116,n20117,n20119);
and (n20117,n20118,n20047);
xor (n20118,n20043,n20044);
and (n20119,n20120,n20121);
xor (n20120,n20118,n20047);
or (n20121,n20122,n20124);
and (n20122,n20123,n20053);
xor (n20123,n20049,n20050);
and (n20124,n20125,n20126);
xor (n20125,n20123,n20053);
or (n20126,n20127,n20129);
and (n20127,n20128,n20059);
xor (n20128,n20055,n20056);
and (n20129,n20130,n20131);
xor (n20130,n20128,n20059);
and (n20131,n20132,n7977);
xor (n20132,n20061,n20062);
or (n20133,n20134,n20136);
and (n20134,n20135,n10287);
xor (n20135,n20065,n20066);
and (n20136,n20137,n20138);
xor (n20137,n20135,n10287);
or (n20138,n20139,n20141);
and (n20139,n20140,n19995);
xor (n20140,n20070,n20071);
and (n20141,n20142,n20143);
xor (n20142,n20140,n19995);
or (n20143,n20144,n20146);
and (n20144,n20145,n20001);
xor (n20145,n20075,n20076);
and (n20146,n20147,n20148);
xor (n20147,n20145,n20001);
or (n20148,n20149,n20151);
and (n20149,n20150,n20007);
xor (n20150,n20080,n20081);
and (n20151,n20152,n20153);
xor (n20152,n20150,n20007);
or (n20153,n20154,n20156);
and (n20154,n20155,n20013);
xor (n20155,n20085,n20086);
and (n20156,n20157,n20158);
xor (n20157,n20155,n20013);
or (n20158,n20159,n20161);
and (n20159,n20160,n20019);
xor (n20160,n20090,n20091);
and (n20161,n20162,n20163);
xor (n20162,n20160,n20019);
or (n20163,n20164,n20166);
and (n20164,n20165,n20025);
xor (n20165,n20095,n20096);
and (n20166,n20167,n20168);
xor (n20167,n20165,n20025);
or (n20168,n20169,n20171);
and (n20169,n20170,n20031);
xor (n20170,n20100,n20101);
and (n20171,n20172,n20173);
xor (n20172,n20170,n20031);
or (n20173,n20174,n20176);
and (n20174,n20175,n9264);
xor (n20175,n20105,n20106);
and (n20176,n20177,n20178);
xor (n20177,n20175,n9264);
or (n20178,n20179,n20181);
and (n20179,n20180,n9004);
xor (n20180,n20110,n20111);
and (n20181,n20182,n20183);
xor (n20182,n20180,n9004);
or (n20183,n20184,n20186);
and (n20184,n20185,n20047);
xor (n20185,n20115,n20116);
and (n20186,n20187,n20188);
xor (n20187,n20185,n20047);
or (n20188,n20189,n20191);
and (n20189,n20190,n20053);
xor (n20190,n20120,n20121);
and (n20191,n20192,n20193);
xor (n20192,n20190,n20053);
or (n20193,n20194,n20196);
and (n20194,n20195,n20059);
xor (n20195,n20125,n20126);
and (n20196,n20197,n20198);
xor (n20197,n20195,n20059);
and (n20198,n20199,n7977);
xor (n20199,n20130,n20131);
or (n20200,n20201,n20203);
and (n20201,n20202,n19995);
xor (n20202,n20137,n20138);
and (n20203,n20204,n20205);
xor (n20204,n20202,n19995);
or (n20205,n20206,n20208);
and (n20206,n20207,n20001);
xor (n20207,n20142,n20143);
and (n20208,n20209,n20210);
xor (n20209,n20207,n20001);
or (n20210,n20211,n20213);
and (n20211,n20212,n20007);
xor (n20212,n20147,n20148);
and (n20213,n20214,n20215);
xor (n20214,n20212,n20007);
or (n20215,n20216,n20218);
and (n20216,n20217,n20013);
xor (n20217,n20152,n20153);
and (n20218,n20219,n20220);
xor (n20219,n20217,n20013);
or (n20220,n20221,n20223);
and (n20221,n20222,n20019);
xor (n20222,n20157,n20158);
and (n20223,n20224,n20225);
xor (n20224,n20222,n20019);
or (n20225,n20226,n20228);
and (n20226,n20227,n20025);
xor (n20227,n20162,n20163);
and (n20228,n20229,n20230);
xor (n20229,n20227,n20025);
or (n20230,n20231,n20233);
and (n20231,n20232,n20031);
xor (n20232,n20167,n20168);
and (n20233,n20234,n20235);
xor (n20234,n20232,n20031);
or (n20235,n20236,n20238);
and (n20236,n20237,n9264);
xor (n20237,n20172,n20173);
and (n20238,n20239,n20240);
xor (n20239,n20237,n9264);
or (n20240,n20241,n20243);
and (n20241,n20242,n9004);
xor (n20242,n20177,n20178);
and (n20243,n20244,n20245);
xor (n20244,n20242,n9004);
or (n20245,n20246,n20248);
and (n20246,n20247,n20047);
xor (n20247,n20182,n20183);
and (n20248,n20249,n20250);
xor (n20249,n20247,n20047);
or (n20250,n20251,n20253);
and (n20251,n20252,n20053);
xor (n20252,n20187,n20188);
and (n20253,n20254,n20255);
xor (n20254,n20252,n20053);
or (n20255,n20256,n20258);
and (n20256,n20257,n20059);
xor (n20257,n20192,n20193);
and (n20258,n20259,n20260);
xor (n20259,n20257,n20059);
and (n20260,n20261,n7977);
xor (n20261,n20197,n20198);
or (n20262,n20263,n20265);
and (n20263,n20264,n20001);
xor (n20264,n20204,n20205);
and (n20265,n20266,n20267);
xor (n20266,n20264,n20001);
or (n20267,n20268,n20270);
and (n20268,n20269,n20007);
xor (n20269,n20209,n20210);
and (n20270,n20271,n20272);
xor (n20271,n20269,n20007);
or (n20272,n20273,n20275);
and (n20273,n20274,n20013);
xor (n20274,n20214,n20215);
and (n20275,n20276,n20277);
xor (n20276,n20274,n20013);
or (n20277,n20278,n20280);
and (n20278,n20279,n20019);
xor (n20279,n20219,n20220);
and (n20280,n20281,n20282);
xor (n20281,n20279,n20019);
or (n20282,n20283,n20285);
and (n20283,n20284,n20025);
xor (n20284,n20224,n20225);
and (n20285,n20286,n20287);
xor (n20286,n20284,n20025);
or (n20287,n20288,n20290);
and (n20288,n20289,n20031);
xor (n20289,n20229,n20230);
and (n20290,n20291,n20292);
xor (n20291,n20289,n20031);
or (n20292,n20293,n20295);
and (n20293,n20294,n9264);
xor (n20294,n20234,n20235);
and (n20295,n20296,n20297);
xor (n20296,n20294,n9264);
or (n20297,n20298,n20300);
and (n20298,n20299,n9004);
xor (n20299,n20239,n20240);
and (n20300,n20301,n20302);
xor (n20301,n20299,n9004);
or (n20302,n20303,n20305);
and (n20303,n20304,n20047);
xor (n20304,n20244,n20245);
and (n20305,n20306,n20307);
xor (n20306,n20304,n20047);
or (n20307,n20308,n20310);
and (n20308,n20309,n20053);
xor (n20309,n20249,n20250);
and (n20310,n20311,n20312);
xor (n20311,n20309,n20053);
or (n20312,n20313,n20315);
and (n20313,n20314,n20059);
xor (n20314,n20254,n20255);
and (n20315,n20316,n20317);
xor (n20316,n20314,n20059);
and (n20317,n20318,n7977);
xor (n20318,n20259,n20260);
or (n20319,n20320,n20322);
and (n20320,n20321,n20007);
xor (n20321,n20266,n20267);
and (n20322,n20323,n20324);
xor (n20323,n20321,n20007);
or (n20324,n20325,n20327);
and (n20325,n20326,n20013);
xor (n20326,n20271,n20272);
and (n20327,n20328,n20329);
xor (n20328,n20326,n20013);
or (n20329,n20330,n20332);
and (n20330,n20331,n20019);
xor (n20331,n20276,n20277);
and (n20332,n20333,n20334);
xor (n20333,n20331,n20019);
or (n20334,n20335,n20337);
and (n20335,n20336,n20025);
xor (n20336,n20281,n20282);
and (n20337,n20338,n20339);
xor (n20338,n20336,n20025);
or (n20339,n20340,n20342);
and (n20340,n20341,n20031);
xor (n20341,n20286,n20287);
and (n20342,n20343,n20344);
xor (n20343,n20341,n20031);
or (n20344,n20345,n20347);
and (n20345,n20346,n9264);
xor (n20346,n20291,n20292);
and (n20347,n20348,n20349);
xor (n20348,n20346,n9264);
or (n20349,n20350,n20352);
and (n20350,n20351,n9004);
xor (n20351,n20296,n20297);
and (n20352,n20353,n20354);
xor (n20353,n20351,n9004);
or (n20354,n20355,n20357);
and (n20355,n20356,n20047);
xor (n20356,n20301,n20302);
and (n20357,n20358,n20359);
xor (n20358,n20356,n20047);
or (n20359,n20360,n20362);
and (n20360,n20361,n20053);
xor (n20361,n20306,n20307);
and (n20362,n20363,n20364);
xor (n20363,n20361,n20053);
or (n20364,n20365,n20367);
and (n20365,n20366,n20059);
xor (n20366,n20311,n20312);
and (n20367,n20368,n20369);
xor (n20368,n20366,n20059);
and (n20369,n20370,n7977);
xor (n20370,n20316,n20317);
or (n20371,n20372,n20374);
and (n20372,n20373,n20013);
xor (n20373,n20323,n20324);
and (n20374,n20375,n20376);
xor (n20375,n20373,n20013);
or (n20376,n20377,n20379);
and (n20377,n20378,n20019);
xor (n20378,n20328,n20329);
and (n20379,n20380,n20381);
xor (n20380,n20378,n20019);
or (n20381,n20382,n20384);
and (n20382,n20383,n20025);
xor (n20383,n20333,n20334);
and (n20384,n20385,n20386);
xor (n20385,n20383,n20025);
or (n20386,n20387,n20389);
and (n20387,n20388,n20031);
xor (n20388,n20338,n20339);
and (n20389,n20390,n20391);
xor (n20390,n20388,n20031);
or (n20391,n20392,n20394);
and (n20392,n20393,n9264);
xor (n20393,n20343,n20344);
and (n20394,n20395,n20396);
xor (n20395,n20393,n9264);
or (n20396,n20397,n20399);
and (n20397,n20398,n9004);
xor (n20398,n20348,n20349);
and (n20399,n20400,n20401);
xor (n20400,n20398,n9004);
or (n20401,n20402,n20404);
and (n20402,n20403,n20047);
xor (n20403,n20353,n20354);
and (n20404,n20405,n20406);
xor (n20405,n20403,n20047);
or (n20406,n20407,n20409);
and (n20407,n20408,n20053);
xor (n20408,n20358,n20359);
and (n20409,n20410,n20411);
xor (n20410,n20408,n20053);
or (n20411,n20412,n20414);
and (n20412,n20413,n20059);
xor (n20413,n20363,n20364);
and (n20414,n20415,n20416);
xor (n20415,n20413,n20059);
and (n20416,n20417,n7977);
xor (n20417,n20368,n20369);
or (n20418,n20419,n20421);
and (n20419,n20420,n20019);
xor (n20420,n20375,n20376);
and (n20421,n20422,n20423);
xor (n20422,n20420,n20019);
or (n20423,n20424,n20426);
and (n20424,n20425,n20025);
xor (n20425,n20380,n20381);
and (n20426,n20427,n20428);
xor (n20427,n20425,n20025);
or (n20428,n20429,n20431);
and (n20429,n20430,n20031);
xor (n20430,n20385,n20386);
and (n20431,n20432,n20433);
xor (n20432,n20430,n20031);
or (n20433,n20434,n20436);
and (n20434,n20435,n9264);
xor (n20435,n20390,n20391);
and (n20436,n20437,n20438);
xor (n20437,n20435,n9264);
or (n20438,n20439,n20441);
and (n20439,n20440,n9004);
xor (n20440,n20395,n20396);
and (n20441,n20442,n20443);
xor (n20442,n20440,n9004);
or (n20443,n20444,n20446);
and (n20444,n20445,n20047);
xor (n20445,n20400,n20401);
and (n20446,n20447,n20448);
xor (n20447,n20445,n20047);
or (n20448,n20449,n20451);
and (n20449,n20450,n20053);
xor (n20450,n20405,n20406);
and (n20451,n20452,n20453);
xor (n20452,n20450,n20053);
or (n20453,n20454,n20456);
and (n20454,n20455,n20059);
xor (n20455,n20410,n20411);
and (n20456,n20457,n20458);
xor (n20457,n20455,n20059);
and (n20458,n20459,n7977);
xor (n20459,n20415,n20416);
or (n20460,n20461,n20463);
and (n20461,n20462,n20025);
xor (n20462,n20422,n20423);
and (n20463,n20464,n20465);
xor (n20464,n20462,n20025);
or (n20465,n20466,n20468);
and (n20466,n20467,n20031);
xor (n20467,n20427,n20428);
and (n20468,n20469,n20470);
xor (n20469,n20467,n20031);
or (n20470,n20471,n20473);
and (n20471,n20472,n9264);
xor (n20472,n20432,n20433);
and (n20473,n20474,n20475);
xor (n20474,n20472,n9264);
or (n20475,n20476,n20478);
and (n20476,n20477,n9004);
xor (n20477,n20437,n20438);
and (n20478,n20479,n20480);
xor (n20479,n20477,n9004);
or (n20480,n20481,n20483);
and (n20481,n20482,n20047);
xor (n20482,n20442,n20443);
and (n20483,n20484,n20485);
xor (n20484,n20482,n20047);
or (n20485,n20486,n20488);
and (n20486,n20487,n20053);
xor (n20487,n20447,n20448);
and (n20488,n20489,n20490);
xor (n20489,n20487,n20053);
or (n20490,n20491,n20493);
and (n20491,n20492,n20059);
xor (n20492,n20452,n20453);
and (n20493,n20494,n20495);
xor (n20494,n20492,n20059);
and (n20495,n20496,n7977);
xor (n20496,n20457,n20458);
or (n20497,n20498,n20500);
and (n20498,n20499,n20031);
xor (n20499,n20464,n20465);
and (n20500,n20501,n20502);
xor (n20501,n20499,n20031);
or (n20502,n20503,n20505);
and (n20503,n20504,n9264);
xor (n20504,n20469,n20470);
and (n20505,n20506,n20507);
xor (n20506,n20504,n9264);
or (n20507,n20508,n20510);
and (n20508,n20509,n9004);
xor (n20509,n20474,n20475);
and (n20510,n20511,n20512);
xor (n20511,n20509,n9004);
or (n20512,n20513,n20515);
and (n20513,n20514,n20047);
xor (n20514,n20479,n20480);
and (n20515,n20516,n20517);
xor (n20516,n20514,n20047);
or (n20517,n20518,n20520);
and (n20518,n20519,n20053);
xor (n20519,n20484,n20485);
and (n20520,n20521,n20522);
xor (n20521,n20519,n20053);
or (n20522,n20523,n20525);
and (n20523,n20524,n20059);
xor (n20524,n20489,n20490);
and (n20525,n20526,n20527);
xor (n20526,n20524,n20059);
and (n20527,n20528,n7977);
xor (n20528,n20494,n20495);
or (n20529,n20530,n20532);
and (n20530,n20531,n9264);
xor (n20531,n20501,n20502);
and (n20532,n20533,n20534);
xor (n20533,n20531,n9264);
or (n20534,n20535,n20537);
and (n20535,n20536,n9004);
xor (n20536,n20506,n20507);
and (n20537,n20538,n20539);
xor (n20538,n20536,n9004);
or (n20539,n20540,n20542);
and (n20540,n20541,n20047);
xor (n20541,n20511,n20512);
and (n20542,n20543,n20544);
xor (n20543,n20541,n20047);
or (n20544,n20545,n20547);
and (n20545,n20546,n20053);
xor (n20546,n20516,n20517);
and (n20547,n20548,n20549);
xor (n20548,n20546,n20053);
or (n20549,n20550,n20552);
and (n20550,n20551,n20059);
xor (n20551,n20521,n20522);
and (n20552,n20553,n20554);
xor (n20553,n20551,n20059);
and (n20554,n20555,n7977);
xor (n20555,n20526,n20527);
or (n20556,n20557,n20559);
and (n20557,n20558,n9004);
xor (n20558,n20533,n20534);
and (n20559,n20560,n20561);
xor (n20560,n20558,n9004);
or (n20561,n20562,n20564);
and (n20562,n20563,n20047);
xor (n20563,n20538,n20539);
and (n20564,n20565,n20566);
xor (n20565,n20563,n20047);
or (n20566,n20567,n20569);
and (n20567,n20568,n20053);
xor (n20568,n20543,n20544);
and (n20569,n20570,n20571);
xor (n20570,n20568,n20053);
or (n20571,n20572,n20574);
and (n20572,n20573,n20059);
xor (n20573,n20548,n20549);
and (n20574,n20575,n20576);
xor (n20575,n20573,n20059);
and (n20576,n20577,n7977);
xor (n20577,n20553,n20554);
or (n20578,n20579,n20581);
and (n20579,n20580,n20047);
xor (n20580,n20560,n20561);
and (n20581,n20582,n20583);
xor (n20582,n20580,n20047);
or (n20583,n20584,n20586);
and (n20584,n20585,n20053);
xor (n20585,n20565,n20566);
and (n20586,n20587,n20588);
xor (n20587,n20585,n20053);
or (n20588,n20589,n20591);
and (n20589,n20590,n20059);
xor (n20590,n20570,n20571);
and (n20591,n20592,n20593);
xor (n20592,n20590,n20059);
and (n20593,n20594,n7977);
xor (n20594,n20575,n20576);
or (n20595,n20596,n20598);
and (n20596,n20597,n20053);
xor (n20597,n20582,n20583);
and (n20598,n20599,n20600);
xor (n20599,n20597,n20053);
or (n20600,n20601,n20603);
and (n20601,n20602,n20059);
xor (n20602,n20587,n20588);
and (n20603,n20604,n20605);
xor (n20604,n20602,n20059);
and (n20605,n20606,n7977);
xor (n20606,n20592,n20593);
or (n20607,n20608,n20610);
and (n20608,n20609,n20059);
xor (n20609,n20599,n20600);
and (n20610,n20611,n20612);
xor (n20611,n20609,n20059);
and (n20612,n20613,n7977);
xor (n20613,n20604,n20605);
and (n20614,n20615,n7977);
xor (n20615,n20611,n20612);
not (n20616,n20617);
xor (n20617,n20618,n8005);
xor (n20618,n20619,n22485);
xor (n20619,n20620,n8008);
xor (n20620,n20621,n22478);
xor (n20621,n20622,n9092);
xor (n20622,n20623,n22466);
xor (n20623,n20624,n21920);
xor (n20624,n20625,n22449);
xor (n20625,n20626,n9270);
xor (n20626,n20627,n22427);
xor (n20627,n20628,n21909);
xor (n20628,n20629,n22400);
xor (n20629,n20630,n21903);
xor (n20630,n20631,n22368);
xor (n20631,n20632,n21897);
xor (n20632,n20633,n22331);
xor (n20633,n20634,n9907);
xor (n20634,n20635,n22289);
xor (n20635,n20636,n10010);
xor (n20636,n20637,n22242);
xor (n20637,n20638,n10083);
xor (n20638,n20639,n22190);
xor (n20639,n20640,n10161);
xor (n20640,n20641,n22133);
xor (n20641,n20642,n10220);
xor (n20642,n20643,n22071);
xor (n20643,n20644,n10295);
xor (n20644,n20645,n22004);
xor (n20645,n20646,n10347);
xor (n20646,n20647,n20705);
xor (n20647,n20648,n10380);
xor (n20648,n20649,n20704);
xor (n20649,n20650,n10380);
xor (n20650,n20651,n20703);
xor (n20651,n20652,n20702);
xor (n20652,n20653,n20701);
xor (n20653,n20654,n10306);
xor (n20654,n20655,n20700);
xor (n20655,n20656,n20699);
xor (n20656,n20657,n20698);
xor (n20657,n20658,n10181);
xor (n20658,n20659,n20697);
xor (n20659,n20660,n20696);
xor (n20660,n20661,n20695);
xor (n20661,n20662,n20694);
xor (n20662,n20663,n20693);
xor (n20663,n20664,n20692);
xor (n20664,n20665,n20691);
xor (n20665,n20666,n20690);
xor (n20666,n20667,n20689);
xor (n20667,n20668,n20688);
xor (n20668,n20669,n20687);
xor (n20669,n20670,n20686);
xor (n20670,n20671,n20685);
xor (n20671,n20672,n20684);
xor (n20672,n20673,n20683);
xor (n20673,n20674,n20682);
xor (n20674,n20675,n20681);
xor (n20675,n20676,n20680);
xor (n20676,n20677,n20679);
xor (n20677,n20678,n7916);
and (n20678,n7917,n7237);
and (n20679,n20678,n7916);
and (n20680,n7917,n7124);
and (n20681,n20676,n20680);
and (n20682,n7917,n7120);
and (n20683,n20674,n20682);
and (n20684,n7917,n7154);
and (n20685,n20672,n20684);
and (n20686,n7917,n7147);
and (n20687,n20670,n20686);
and (n20688,n7917,n7479);
and (n20689,n20668,n20688);
and (n20690,n7917,n7483);
and (n20691,n20666,n20690);
and (n20692,n7917,n7527);
and (n20693,n20664,n20692);
and (n20694,n7917,n7078);
and (n20695,n20662,n20694);
and (n20696,n7917,n7072);
and (n20697,n20660,n20696);
and (n20698,n20658,n10181);
and (n20699,n7917,n7091);
and (n20700,n20656,n20699);
and (n20701,n20654,n10306);
and (n20702,n7917,n7753);
and (n20703,n20652,n20702);
and (n20704,n20650,n10380);
or (n20705,n20706,n21935);
and (n20706,n20707,n10347);
xor (n20707,n20649,n20708);
or (n20708,n20709,n21862);
and (n20709,n20710,n10347);
xor (n20710,n20651,n20711);
or (n20711,n20712,n21779);
and (n20712,n20713,n21778);
xor (n20713,n20653,n20714);
or (n20714,n20715,n21706);
and (n20715,n20716,n10255);
xor (n20716,n20655,n20717);
or (n20717,n20718,n21623);
and (n20718,n20719,n21622);
xor (n20719,n20657,n20720);
or (n20720,n20721,n21546);
and (n20721,n20722,n10105);
xor (n20722,n20659,n20723);
or (n20723,n20724,n21463);
and (n20724,n20725,n21462);
xor (n20725,n20661,n20726);
or (n20726,n20727,n21386);
and (n20727,n20728,n9936);
xor (n20728,n20663,n20729);
or (n20729,n20730,n21303);
and (n20730,n20731,n21302);
xor (n20731,n20665,n20732);
or (n20732,n20733,n21227);
and (n20733,n20734,n9627);
xor (n20734,n20667,n20735);
or (n20735,n20736,n21144);
and (n20736,n20737,n21143);
xor (n20737,n20669,n20738);
or (n20738,n20739,n21069);
and (n20739,n20740,n21068);
xor (n20740,n20671,n20741);
or (n20741,n20742,n20985);
and (n20742,n20743,n20984);
xor (n20743,n20673,n20744);
or (n20744,n20745,n20910);
and (n20745,n20746,n9113);
xor (n20746,n20675,n20747);
or (n20747,n20748,n20827);
and (n20748,n20749,n20826);
xor (n20749,n20677,n20750);
or (n20750,n20751,n20752);
and (n20751,n20678,n7241);
and (n20752,n20753,n20754);
xor (n20753,n20678,n7241);
or (n20754,n20755,n20758);
and (n20755,n20756,n20757);
and (n20756,n7242,n7237);
and (n20757,n7232,n7123);
and (n20758,n20759,n20760);
xor (n20759,n20756,n20757);
or (n20760,n20761,n20763);
and (n20761,n20762,n7281);
and (n20762,n7232,n7237);
and (n20763,n20764,n20765);
xor (n20764,n20762,n7281);
or (n20765,n20766,n20768);
and (n20766,n20767,n7429);
and (n20767,n7134,n7237);
and (n20768,n20769,n20770);
xor (n20769,n20767,n7429);
or (n20770,n20771,n20774);
and (n20771,n20772,n20773);
and (n20772,n7129,n7237);
and (n20773,n7165,n7123);
and (n20774,n20775,n20776);
xor (n20775,n20772,n20773);
or (n20776,n20777,n20779);
and (n20777,n20778,n8171);
and (n20778,n7165,n7237);
and (n20779,n20780,n20781);
xor (n20780,n20778,n8171);
or (n20781,n20782,n20785);
and (n20782,n20783,n20784);
and (n20783,n7146,n7237);
and (n20784,n7308,n7123);
and (n20785,n20786,n20787);
xor (n20786,n20783,n20784);
or (n20787,n20788,n20791);
and (n20788,n20789,n20790);
and (n20789,n7308,n7237);
and (n20790,n7471,n7123);
and (n20791,n20792,n20793);
xor (n20792,n20789,n20790);
or (n20793,n20794,n20796);
and (n20794,n20795,n8529);
and (n20795,n7471,n7237);
and (n20796,n20797,n20798);
xor (n20797,n20795,n8529);
or (n20798,n20799,n20802);
and (n20799,n20800,n20801);
and (n20800,n7463,n7237);
and (n20801,n7497,n7123);
and (n20802,n20803,n20804);
xor (n20803,n20800,n20801);
or (n20804,n20805,n20807);
and (n20805,n20806,n8660);
and (n20806,n7497,n7237);
and (n20807,n20808,n20809);
xor (n20808,n20806,n8660);
or (n20809,n20810,n20812);
and (n20810,n20811,n8706);
and (n20811,n7084,n7237);
and (n20812,n20813,n20814);
xor (n20813,n20811,n8706);
or (n20814,n20815,n20817);
and (n20815,n20816,n8775);
and (n20816,n7064,n7237);
and (n20817,n20818,n20819);
xor (n20818,n20816,n8775);
or (n20819,n20820,n20822);
and (n20820,n20821,n8823);
and (n20821,n7109,n7237);
and (n20822,n20823,n20824);
xor (n20823,n20821,n8823);
and (n20824,n20825,n8840);
and (n20825,n7102,n7237);
and (n20826,n7242,n7124);
and (n20827,n20828,n20829);
xor (n20828,n20749,n20826);
or (n20829,n20830,n20833);
and (n20830,n20831,n20832);
xor (n20831,n20753,n20754);
and (n20832,n7232,n7124);
and (n20833,n20834,n20835);
xor (n20834,n20831,n20832);
or (n20835,n20836,n20839);
and (n20836,n20837,n20838);
xor (n20837,n20759,n20760);
and (n20838,n7134,n7124);
and (n20839,n20840,n20841);
xor (n20840,n20837,n20838);
or (n20841,n20842,n20845);
and (n20842,n20843,n20844);
xor (n20843,n20764,n20765);
and (n20844,n7129,n7124);
and (n20845,n20846,n20847);
xor (n20846,n20843,n20844);
or (n20847,n20848,n20851);
and (n20848,n20849,n20850);
xor (n20849,n20769,n20770);
and (n20850,n7165,n7124);
and (n20851,n20852,n20853);
xor (n20852,n20849,n20850);
or (n20853,n20854,n20857);
and (n20854,n20855,n20856);
xor (n20855,n20775,n20776);
and (n20856,n7146,n7124);
and (n20857,n20858,n20859);
xor (n20858,n20855,n20856);
or (n20859,n20860,n20863);
and (n20860,n20861,n20862);
xor (n20861,n20780,n20781);
and (n20862,n7308,n7124);
and (n20863,n20864,n20865);
xor (n20864,n20861,n20862);
or (n20865,n20866,n20869);
and (n20866,n20867,n20868);
xor (n20867,n20786,n20787);
and (n20868,n7471,n7124);
and (n20869,n20870,n20871);
xor (n20870,n20867,n20868);
or (n20871,n20872,n20875);
and (n20872,n20873,n20874);
xor (n20873,n20792,n20793);
and (n20874,n7463,n7124);
and (n20875,n20876,n20877);
xor (n20876,n20873,n20874);
or (n20877,n20878,n20881);
and (n20878,n20879,n20880);
xor (n20879,n20797,n20798);
and (n20880,n7497,n7124);
and (n20881,n20882,n20883);
xor (n20882,n20879,n20880);
or (n20883,n20884,n20887);
and (n20884,n20885,n20886);
xor (n20885,n20803,n20804);
and (n20886,n7084,n7124);
and (n20887,n20888,n20889);
xor (n20888,n20885,n20886);
or (n20889,n20890,n20893);
and (n20890,n20891,n20892);
xor (n20891,n20808,n20809);
and (n20892,n7064,n7124);
and (n20893,n20894,n20895);
xor (n20894,n20891,n20892);
or (n20895,n20896,n20899);
and (n20896,n20897,n20898);
xor (n20897,n20813,n20814);
and (n20898,n7109,n7124);
and (n20899,n20900,n20901);
xor (n20900,n20897,n20898);
or (n20901,n20902,n20905);
and (n20902,n20903,n20904);
xor (n20903,n20818,n20819);
and (n20904,n7102,n7124);
and (n20905,n20906,n20907);
xor (n20906,n20903,n20904);
and (n20907,n20908,n20909);
xor (n20908,n20823,n20824);
and (n20909,n7355,n7124);
and (n20910,n20911,n20912);
xor (n20911,n20746,n9113);
or (n20912,n20913,n20915);
and (n20913,n20914,n7926);
xor (n20914,n20828,n20829);
and (n20915,n20916,n20917);
xor (n20916,n20914,n7926);
or (n20917,n20918,n20921);
and (n20918,n20919,n20920);
xor (n20919,n20834,n20835);
not (n20920,n7135);
and (n20921,n20922,n20923);
xor (n20922,n20919,n20920);
or (n20923,n20924,n20927);
and (n20924,n20925,n20926);
xor (n20925,n20840,n20841);
not (n20926,n7130);
and (n20927,n20928,n20929);
xor (n20928,n20925,n20926);
or (n20929,n20930,n20933);
and (n20930,n20931,n20932);
xor (n20931,n20846,n20847);
not (n20932,n7297);
and (n20933,n20934,n20935);
xor (n20934,n20931,n20932);
or (n20935,n20936,n20939);
and (n20936,n20937,n20938);
xor (n20937,n20852,n20853);
not (n20938,n7436);
and (n20939,n20940,n20941);
xor (n20940,n20937,n20938);
or (n20941,n20942,n20944);
and (n20942,n20943,n7441);
xor (n20943,n20858,n20859);
and (n20944,n20945,n20946);
xor (n20945,n20943,n7441);
or (n20946,n20947,n20950);
and (n20947,n20948,n20949);
xor (n20948,n20864,n20865);
not (n20949,n8081);
and (n20950,n20951,n20952);
xor (n20951,n20948,n20949);
or (n20952,n20953,n20955);
and (n20953,n20954,n8262);
xor (n20954,n20870,n20871);
and (n20955,n20956,n20957);
xor (n20956,n20954,n8262);
or (n20957,n20958,n20960);
and (n20958,n20959,n8353);
xor (n20959,n20876,n20877);
and (n20960,n20961,n20962);
xor (n20961,n20959,n8353);
or (n20962,n20963,n20965);
and (n20963,n20964,n8535);
xor (n20964,n20882,n20883);
and (n20965,n20966,n20967);
xor (n20966,n20964,n8535);
or (n20967,n20968,n20970);
and (n20968,n20969,n8581);
xor (n20969,n20888,n20889);
and (n20970,n20971,n20972);
xor (n20971,n20969,n8581);
or (n20972,n20973,n20975);
and (n20973,n20974,n8617);
xor (n20974,n20894,n20895);
and (n20975,n20976,n20977);
xor (n20976,n20974,n8617);
or (n20977,n20978,n20980);
and (n20978,n20979,n8733);
xor (n20979,n20900,n20901);
and (n20980,n20981,n20982);
xor (n20981,n20979,n8733);
and (n20982,n20983,n8781);
xor (n20983,n20906,n20907);
and (n20984,n7242,n7154);
and (n20985,n20986,n20987);
xor (n20986,n20743,n20984);
or (n20987,n20988,n20991);
and (n20988,n20989,n20990);
xor (n20989,n20911,n20912);
and (n20990,n7232,n7154);
and (n20991,n20992,n20993);
xor (n20992,n20989,n20990);
or (n20993,n20994,n20997);
and (n20994,n20995,n20996);
xor (n20995,n20916,n20917);
and (n20996,n7134,n7154);
and (n20997,n20998,n20999);
xor (n20998,n20995,n20996);
or (n20999,n21000,n21003);
and (n21000,n21001,n21002);
xor (n21001,n20922,n20923);
and (n21002,n7129,n7154);
and (n21003,n21004,n21005);
xor (n21004,n21001,n21002);
or (n21005,n21006,n21009);
and (n21006,n21007,n21008);
xor (n21007,n20928,n20929);
and (n21008,n7165,n7154);
and (n21009,n21010,n21011);
xor (n21010,n21007,n21008);
or (n21011,n21012,n21015);
and (n21012,n21013,n21014);
xor (n21013,n20934,n20935);
and (n21014,n7146,n7154);
and (n21015,n21016,n21017);
xor (n21016,n21013,n21014);
or (n21017,n21018,n21021);
and (n21018,n21019,n21020);
xor (n21019,n20940,n20941);
and (n21020,n7308,n7154);
and (n21021,n21022,n21023);
xor (n21022,n21019,n21020);
or (n21023,n21024,n21027);
and (n21024,n21025,n21026);
xor (n21025,n20945,n20946);
and (n21026,n7471,n7154);
and (n21027,n21028,n21029);
xor (n21028,n21025,n21026);
or (n21029,n21030,n21033);
and (n21030,n21031,n21032);
xor (n21031,n20951,n20952);
and (n21032,n7463,n7154);
and (n21033,n21034,n21035);
xor (n21034,n21031,n21032);
or (n21035,n21036,n21039);
and (n21036,n21037,n21038);
xor (n21037,n20956,n20957);
and (n21038,n7497,n7154);
and (n21039,n21040,n21041);
xor (n21040,n21037,n21038);
or (n21041,n21042,n21045);
and (n21042,n21043,n21044);
xor (n21043,n20961,n20962);
and (n21044,n7084,n7154);
and (n21045,n21046,n21047);
xor (n21046,n21043,n21044);
or (n21047,n21048,n21051);
and (n21048,n21049,n21050);
xor (n21049,n20966,n20967);
and (n21050,n7064,n7154);
and (n21051,n21052,n21053);
xor (n21052,n21049,n21050);
or (n21053,n21054,n21057);
and (n21054,n21055,n21056);
xor (n21055,n20971,n20972);
and (n21056,n7109,n7154);
and (n21057,n21058,n21059);
xor (n21058,n21055,n21056);
or (n21059,n21060,n21063);
and (n21060,n21061,n21062);
xor (n21061,n20976,n20977);
and (n21062,n7102,n7154);
and (n21063,n21064,n21065);
xor (n21064,n21061,n21062);
and (n21065,n21066,n21067);
xor (n21066,n20981,n20982);
and (n21067,n7355,n7154);
and (n21068,n7242,n7147);
and (n21069,n21070,n21071);
xor (n21070,n20740,n21068);
or (n21071,n21072,n21075);
and (n21072,n21073,n21074);
xor (n21073,n20986,n20987);
and (n21074,n7232,n7147);
and (n21075,n21076,n21077);
xor (n21076,n21073,n21074);
or (n21077,n21078,n21080);
and (n21078,n21079,n9127);
xor (n21079,n20992,n20993);
and (n21080,n21081,n21082);
xor (n21081,n21079,n9127);
or (n21082,n21083,n21086);
and (n21083,n21084,n21085);
xor (n21084,n20998,n20999);
not (n21085,n8030);
and (n21086,n21087,n21088);
xor (n21087,n21084,n21085);
or (n21088,n21089,n21091);
and (n21089,n21090,n7166);
xor (n21090,n21004,n21005);
and (n21091,n21092,n21093);
xor (n21092,n21090,n7166);
or (n21093,n21094,n21097);
and (n21094,n21095,n21096);
xor (n21095,n21010,n21011);
and (n21096,n7146,n7147);
and (n21097,n21098,n21099);
xor (n21098,n21095,n21096);
or (n21099,n21100,n21102);
and (n21100,n21101,n7307);
xor (n21101,n21016,n21017);
and (n21102,n21103,n21104);
xor (n21103,n21101,n7307);
or (n21104,n21105,n21107);
and (n21105,n21106,n7472);
xor (n21106,n21022,n21023);
and (n21107,n21108,n21109);
xor (n21108,n21106,n7472);
or (n21109,n21110,n21112);
and (n21110,n21111,n7462);
xor (n21111,n21028,n21029);
and (n21112,n21113,n21114);
xor (n21113,n21111,n7462);
or (n21114,n21115,n21118);
and (n21115,n21116,n21117);
xor (n21116,n21034,n21035);
and (n21117,n7497,n7147);
and (n21118,n21119,n21120);
xor (n21119,n21116,n21117);
or (n21120,n21121,n21123);
and (n21121,n21122,n8267);
xor (n21122,n21040,n21041);
and (n21123,n21124,n21125);
xor (n21124,n21122,n8267);
or (n21125,n21126,n21129);
and (n21126,n21127,n21128);
xor (n21127,n21046,n21047);
and (n21128,n7064,n7147);
and (n21129,n21130,n21131);
xor (n21130,n21127,n21128);
or (n21131,n21132,n21134);
and (n21132,n21133,n8461);
xor (n21133,n21052,n21053);
and (n21134,n21135,n21136);
xor (n21135,n21133,n8461);
or (n21136,n21137,n21139);
and (n21137,n21138,n8628);
xor (n21138,n21058,n21059);
and (n21139,n21140,n21141);
xor (n21140,n21138,n8628);
and (n21141,n21142,n8624);
xor (n21142,n21064,n21065);
and (n21143,n7242,n7479);
and (n21144,n21145,n21146);
xor (n21145,n20737,n21143);
or (n21146,n21147,n21150);
and (n21147,n21148,n21149);
xor (n21148,n21070,n21071);
and (n21149,n7232,n7479);
and (n21150,n21151,n21152);
xor (n21151,n21148,n21149);
or (n21152,n21153,n21156);
and (n21153,n21154,n21155);
xor (n21154,n21076,n21077);
and (n21155,n7134,n7479);
and (n21156,n21157,n21158);
xor (n21157,n21154,n21155);
or (n21158,n21159,n21162);
and (n21159,n21160,n21161);
xor (n21160,n21081,n21082);
and (n21161,n7129,n7479);
and (n21162,n21163,n21164);
xor (n21163,n21160,n21161);
or (n21164,n21165,n21168);
and (n21165,n21166,n21167);
xor (n21166,n21087,n21088);
and (n21167,n7165,n7479);
and (n21168,n21169,n21170);
xor (n21169,n21166,n21167);
or (n21170,n21171,n21174);
and (n21171,n21172,n21173);
xor (n21172,n21092,n21093);
and (n21173,n7146,n7479);
and (n21174,n21175,n21176);
xor (n21175,n21172,n21173);
or (n21176,n21177,n21180);
and (n21177,n21178,n21179);
xor (n21178,n21098,n21099);
and (n21179,n7308,n7479);
and (n21180,n21181,n21182);
xor (n21181,n21178,n21179);
or (n21182,n21183,n21186);
and (n21183,n21184,n21185);
xor (n21184,n21103,n21104);
and (n21185,n7471,n7479);
and (n21186,n21187,n21188);
xor (n21187,n21184,n21185);
or (n21188,n21189,n21192);
and (n21189,n21190,n21191);
xor (n21190,n21108,n21109);
and (n21191,n7463,n7479);
and (n21192,n21193,n21194);
xor (n21193,n21190,n21191);
or (n21194,n21195,n21198);
and (n21195,n21196,n21197);
xor (n21196,n21113,n21114);
and (n21197,n7497,n7479);
and (n21198,n21199,n21200);
xor (n21199,n21196,n21197);
or (n21200,n21201,n21204);
and (n21201,n21202,n21203);
xor (n21202,n21119,n21120);
and (n21203,n7084,n7479);
and (n21204,n21205,n21206);
xor (n21205,n21202,n21203);
or (n21206,n21207,n21210);
and (n21207,n21208,n21209);
xor (n21208,n21124,n21125);
and (n21209,n7064,n7479);
and (n21210,n21211,n21212);
xor (n21211,n21208,n21209);
or (n21212,n21213,n21216);
and (n21213,n21214,n21215);
xor (n21214,n21130,n21131);
and (n21215,n7109,n7479);
and (n21216,n21217,n21218);
xor (n21217,n21214,n21215);
or (n21218,n21219,n21222);
and (n21219,n21220,n21221);
xor (n21220,n21135,n21136);
and (n21221,n7102,n7479);
and (n21222,n21223,n21224);
xor (n21223,n21220,n21221);
and (n21224,n21225,n21226);
xor (n21225,n21140,n21141);
and (n21226,n7355,n7479);
and (n21227,n21228,n21229);
xor (n21228,n20734,n9627);
or (n21229,n21230,n21233);
and (n21230,n21231,n21232);
xor (n21231,n21145,n21146);
and (n21232,n7232,n7483);
and (n21233,n21234,n21235);
xor (n21234,n21231,n21232);
or (n21235,n21236,n21239);
and (n21236,n21237,n21238);
xor (n21237,n21151,n21152);
and (n21238,n7134,n7483);
and (n21239,n21240,n21241);
xor (n21240,n21237,n21238);
or (n21241,n21242,n21244);
and (n21242,n21243,n8972);
xor (n21243,n21157,n21158);
and (n21244,n21245,n21246);
xor (n21245,n21243,n8972);
or (n21246,n21247,n21249);
and (n21247,n21248,n9155);
xor (n21248,n21163,n21164);
and (n21249,n21250,n21251);
xor (n21250,n21248,n9155);
or (n21251,n21252,n21255);
and (n21252,n21253,n21254);
xor (n21253,n21169,n21170);
not (n21254,n7885);
and (n21255,n21256,n21257);
xor (n21256,n21253,n21254);
or (n21257,n21258,n21261);
and (n21258,n21259,n21260);
xor (n21259,n21175,n21176);
and (n21260,n7308,n7483);
and (n21261,n21262,n21263);
xor (n21262,n21259,n21260);
or (n21263,n21264,n21266);
and (n21264,n21265,n7690);
xor (n21265,n21181,n21182);
and (n21266,n21267,n21268);
xor (n21267,n21265,n7690);
or (n21268,n21269,n21271);
and (n21269,n21270,n7654);
xor (n21270,n21187,n21188);
and (n21271,n21272,n21273);
xor (n21272,n21270,n7654);
or (n21273,n21274,n21277);
and (n21274,n21275,n21276);
xor (n21275,n21193,n21194);
and (n21276,n7497,n7483);
and (n21277,n21278,n21279);
xor (n21278,n21275,n21276);
or (n21279,n21280,n21282);
and (n21280,n21281,n7490);
xor (n21281,n21199,n21200);
and (n21282,n21283,n21284);
xor (n21283,n21281,n7490);
or (n21284,n21285,n21287);
and (n21285,n21286,n8110);
xor (n21286,n21205,n21206);
and (n21287,n21288,n21289);
xor (n21288,n21286,n8110);
or (n21289,n21290,n21293);
and (n21290,n21291,n21292);
xor (n21291,n21211,n21212);
not (n21292,n8216);
and (n21293,n21294,n21295);
xor (n21294,n21291,n21292);
or (n21295,n21296,n21298);
and (n21296,n21297,n8397);
xor (n21297,n21217,n21218);
and (n21298,n21299,n21300);
xor (n21299,n21297,n8397);
and (n21300,n21301,n8470);
xor (n21301,n21223,n21224);
and (n21302,n7242,n7527);
and (n21303,n21304,n21305);
xor (n21304,n20731,n21302);
or (n21305,n21306,n21309);
and (n21306,n21307,n21308);
xor (n21307,n21228,n21229);
and (n21308,n7232,n7527);
and (n21309,n21310,n21311);
xor (n21310,n21307,n21308);
or (n21311,n21312,n21315);
and (n21312,n21313,n21314);
xor (n21313,n21234,n21235);
and (n21314,n7134,n7527);
and (n21315,n21316,n21317);
xor (n21316,n21313,n21314);
or (n21317,n21318,n21321);
and (n21318,n21319,n21320);
xor (n21319,n21240,n21241);
and (n21320,n7129,n7527);
and (n21321,n21322,n21323);
xor (n21322,n21319,n21320);
or (n21323,n21324,n21327);
and (n21324,n21325,n21326);
xor (n21325,n21245,n21246);
and (n21326,n7165,n7527);
and (n21327,n21328,n21329);
xor (n21328,n21325,n21326);
or (n21329,n21330,n21333);
and (n21330,n21331,n21332);
xor (n21331,n21250,n21251);
and (n21332,n7146,n7527);
and (n21333,n21334,n21335);
xor (n21334,n21331,n21332);
or (n21335,n21336,n21339);
and (n21336,n21337,n21338);
xor (n21337,n21256,n21257);
and (n21338,n7308,n7527);
and (n21339,n21340,n21341);
xor (n21340,n21337,n21338);
or (n21341,n21342,n21345);
and (n21342,n21343,n21344);
xor (n21343,n21262,n21263);
and (n21344,n7471,n7527);
and (n21345,n21346,n21347);
xor (n21346,n21343,n21344);
or (n21347,n21348,n21351);
and (n21348,n21349,n21350);
xor (n21349,n21267,n21268);
and (n21350,n7463,n7527);
and (n21351,n21352,n21353);
xor (n21352,n21349,n21350);
or (n21353,n21354,n21357);
and (n21354,n21355,n21356);
xor (n21355,n21272,n21273);
and (n21356,n7497,n7527);
and (n21357,n21358,n21359);
xor (n21358,n21355,n21356);
or (n21359,n21360,n21363);
and (n21360,n21361,n21362);
xor (n21361,n21278,n21279);
and (n21362,n7084,n7527);
and (n21363,n21364,n21365);
xor (n21364,n21361,n21362);
or (n21365,n21366,n21369);
and (n21366,n21367,n21368);
xor (n21367,n21283,n21284);
and (n21368,n7064,n7527);
and (n21369,n21370,n21371);
xor (n21370,n21367,n21368);
or (n21371,n21372,n21375);
and (n21372,n21373,n21374);
xor (n21373,n21288,n21289);
and (n21374,n7109,n7527);
and (n21375,n21376,n21377);
xor (n21376,n21373,n21374);
or (n21377,n21378,n21381);
and (n21378,n21379,n21380);
xor (n21379,n21294,n21295);
and (n21380,n7102,n7527);
and (n21381,n21382,n21383);
xor (n21382,n21379,n21380);
and (n21383,n21384,n21385);
xor (n21384,n21299,n21300);
and (n21385,n7355,n7527);
and (n21386,n21387,n21388);
xor (n21387,n20728,n9936);
or (n21388,n21389,n21391);
and (n21389,n21390,n9741);
xor (n21390,n21304,n21305);
and (n21391,n21392,n21393);
xor (n21392,n21390,n9741);
or (n21393,n21394,n21396);
and (n21394,n21395,n9633);
xor (n21395,n21310,n21311);
and (n21396,n21397,n21398);
xor (n21397,n21395,n9633);
or (n21398,n21399,n21401);
and (n21399,n21400,n9392);
xor (n21400,n21316,n21317);
and (n21401,n21402,n21403);
xor (n21402,n21400,n9392);
or (n21403,n21404,n21406);
and (n21404,n21405,n8985);
xor (n21405,n21322,n21323);
and (n21406,n21407,n21408);
xor (n21407,n21405,n8985);
or (n21408,n21409,n21412);
and (n21409,n21410,n21411);
xor (n21410,n21328,n21329);
not (n21411,n8990);
and (n21412,n21413,n21414);
xor (n21413,n21410,n21411);
or (n21414,n21415,n21417);
and (n21415,n21416,n9161);
xor (n21416,n21334,n21335);
and (n21417,n21418,n21419);
xor (n21418,n21416,n9161);
or (n21419,n21420,n21423);
and (n21420,n21421,n21422);
xor (n21421,n21340,n21341);
and (n21422,n7471,n7078);
and (n21423,n21424,n21425);
xor (n21424,n21421,n21422);
or (n21425,n21426,n21428);
and (n21426,n21427,n7705);
xor (n21427,n21346,n21347);
and (n21428,n21429,n21430);
xor (n21429,n21427,n7705);
or (n21430,n21431,n21434);
and (n21431,n21432,n21433);
xor (n21432,n21352,n21353);
and (n21433,n7497,n7078);
and (n21434,n21435,n21436);
xor (n21435,n21432,n21433);
or (n21436,n21437,n21440);
and (n21437,n21438,n21439);
xor (n21438,n21358,n21359);
and (n21439,n7084,n7078);
and (n21440,n21441,n21442);
xor (n21441,n21438,n21439);
or (n21442,n21443,n21446);
and (n21443,n21444,n21445);
xor (n21444,n21364,n21365);
not (n21445,n7535);
and (n21446,n21447,n21448);
xor (n21447,n21444,n21445);
or (n21448,n21449,n21452);
and (n21449,n21450,n21451);
xor (n21450,n21370,n21371);
and (n21451,n7109,n7078);
and (n21452,n21453,n21454);
xor (n21453,n21450,n21451);
or (n21454,n21455,n21458);
and (n21455,n21456,n21457);
xor (n21456,n21376,n21377);
and (n21457,n7102,n7078);
and (n21458,n21459,n21460);
xor (n21459,n21456,n21457);
and (n21460,n21461,n8222);
xor (n21461,n21382,n21383);
and (n21462,n7242,n7072);
and (n21463,n21464,n21465);
xor (n21464,n20725,n21462);
or (n21465,n21466,n21469);
and (n21466,n21467,n21468);
xor (n21467,n21387,n21388);
and (n21468,n7232,n7072);
and (n21469,n21470,n21471);
xor (n21470,n21467,n21468);
or (n21471,n21472,n21475);
and (n21472,n21473,n21474);
xor (n21473,n21392,n21393);
and (n21474,n7134,n7072);
and (n21475,n21476,n21477);
xor (n21476,n21473,n21474);
or (n21477,n21478,n21481);
and (n21478,n21479,n21480);
xor (n21479,n21397,n21398);
and (n21480,n7129,n7072);
and (n21481,n21482,n21483);
xor (n21482,n21479,n21480);
or (n21483,n21484,n21487);
and (n21484,n21485,n21486);
xor (n21485,n21402,n21403);
and (n21486,n7165,n7072);
and (n21487,n21488,n21489);
xor (n21488,n21485,n21486);
or (n21489,n21490,n21493);
and (n21490,n21491,n21492);
xor (n21491,n21407,n21408);
and (n21492,n7146,n7072);
and (n21493,n21494,n21495);
xor (n21494,n21491,n21492);
or (n21495,n21496,n21499);
and (n21496,n21497,n21498);
xor (n21497,n21413,n21414);
and (n21498,n7308,n7072);
and (n21499,n21500,n21501);
xor (n21500,n21497,n21498);
or (n21501,n21502,n21505);
and (n21502,n21503,n21504);
xor (n21503,n21418,n21419);
and (n21504,n7471,n7072);
and (n21505,n21506,n21507);
xor (n21506,n21503,n21504);
or (n21507,n21508,n21511);
and (n21508,n21509,n21510);
xor (n21509,n21424,n21425);
and (n21510,n7463,n7072);
and (n21511,n21512,n21513);
xor (n21512,n21509,n21510);
or (n21513,n21514,n21517);
and (n21514,n21515,n21516);
xor (n21515,n21429,n21430);
and (n21516,n7497,n7072);
and (n21517,n21518,n21519);
xor (n21518,n21515,n21516);
or (n21519,n21520,n21523);
and (n21520,n21521,n21522);
xor (n21521,n21435,n21436);
and (n21522,n7084,n7072);
and (n21523,n21524,n21525);
xor (n21524,n21521,n21522);
or (n21525,n21526,n21529);
and (n21526,n21527,n21528);
xor (n21527,n21441,n21442);
and (n21528,n7064,n7072);
and (n21529,n21530,n21531);
xor (n21530,n21527,n21528);
or (n21531,n21532,n21535);
and (n21532,n21533,n21534);
xor (n21533,n21447,n21448);
and (n21534,n7109,n7072);
and (n21535,n21536,n21537);
xor (n21536,n21533,n21534);
or (n21537,n21538,n21541);
and (n21538,n21539,n21540);
xor (n21539,n21453,n21454);
and (n21540,n7102,n7072);
and (n21541,n21542,n21543);
xor (n21542,n21539,n21540);
and (n21543,n21544,n21545);
xor (n21544,n21459,n21460);
and (n21545,n7355,n7072);
and (n21546,n21547,n21548);
xor (n21547,n20722,n10105);
or (n21548,n21549,n21551);
and (n21549,n21550,n10031);
xor (n21550,n21464,n21465);
and (n21551,n21552,n21553);
xor (n21552,n21550,n10031);
or (n21553,n21554,n21556);
and (n21554,n21555,n9884);
xor (n21555,n21470,n21471);
and (n21556,n21557,n21558);
xor (n21557,n21555,n9884);
or (n21558,n21559,n21561);
and (n21559,n21560,n9769);
xor (n21560,n21476,n21477);
and (n21561,n21562,n21563);
xor (n21562,n21560,n9769);
or (n21563,n21564,n21567);
and (n21564,n21565,n21566);
xor (n21565,n21482,n21483);
and (n21566,n7165,n7065);
and (n21567,n21568,n21569);
xor (n21568,n21565,n21566);
or (n21569,n21570,n21572);
and (n21570,n21571,n9362);
xor (n21571,n21488,n21489);
and (n21572,n21573,n21574);
xor (n21573,n21571,n9362);
or (n21574,n21575,n21578);
and (n21575,n21576,n21577);
xor (n21576,n21494,n21495);
not (n21577,n8956);
and (n21578,n21579,n21580);
xor (n21579,n21576,n21577);
or (n21580,n21581,n21584);
and (n21581,n21582,n21583);
xor (n21582,n21500,n21501);
and (n21583,n7471,n7065);
and (n21584,n21585,n21586);
xor (n21585,n21582,n21583);
or (n21586,n21587,n21590);
and (n21587,n21588,n21589);
xor (n21588,n21506,n21507);
and (n21589,n7463,n7065);
and (n21590,n21591,n21592);
xor (n21591,n21588,n21589);
or (n21592,n21593,n21595);
and (n21593,n21594,n7842);
xor (n21594,n21512,n21513);
and (n21595,n21596,n21597);
xor (n21596,n21594,n7842);
or (n21597,n21598,n21601);
and (n21598,n21599,n21600);
xor (n21599,n21518,n21519);
and (n21600,n7084,n7065);
and (n21601,n21602,n21603);
xor (n21602,n21599,n21600);
or (n21603,n21604,n21607);
and (n21604,n21605,n21606);
xor (n21605,n21524,n21525);
and (n21606,n7064,n7065);
and (n21607,n21608,n21609);
xor (n21608,n21605,n21606);
or (n21609,n21610,n21612);
and (n21610,n21611,n7347);
xor (n21611,n21530,n21531);
and (n21612,n21613,n21614);
xor (n21613,n21611,n7347);
or (n21614,n21615,n21618);
and (n21615,n21616,n21617);
xor (n21616,n21536,n21537);
and (n21617,n7102,n7065);
and (n21618,n21619,n21620);
xor (n21619,n21616,n21617);
and (n21620,n21621,n7543);
xor (n21621,n21542,n21543);
and (n21622,n7242,n7091);
and (n21623,n21624,n21625);
xor (n21624,n20719,n21622);
or (n21625,n21626,n21629);
and (n21626,n21627,n21628);
xor (n21627,n21547,n21548);
and (n21628,n7232,n7091);
and (n21629,n21630,n21631);
xor (n21630,n21627,n21628);
or (n21631,n21632,n21635);
and (n21632,n21633,n21634);
xor (n21633,n21552,n21553);
and (n21634,n7134,n7091);
and (n21635,n21636,n21637);
xor (n21636,n21633,n21634);
or (n21637,n21638,n21641);
and (n21638,n21639,n21640);
xor (n21639,n21557,n21558);
and (n21640,n7129,n7091);
and (n21641,n21642,n21643);
xor (n21642,n21639,n21640);
or (n21643,n21644,n21647);
and (n21644,n21645,n21646);
xor (n21645,n21562,n21563);
and (n21646,n7165,n7091);
and (n21647,n21648,n21649);
xor (n21648,n21645,n21646);
or (n21649,n21650,n21653);
and (n21650,n21651,n21652);
xor (n21651,n21568,n21569);
and (n21652,n7146,n7091);
and (n21653,n21654,n21655);
xor (n21654,n21651,n21652);
or (n21655,n21656,n21659);
and (n21656,n21657,n21658);
xor (n21657,n21573,n21574);
and (n21658,n7308,n7091);
and (n21659,n21660,n21661);
xor (n21660,n21657,n21658);
or (n21661,n21662,n21665);
and (n21662,n21663,n21664);
xor (n21663,n21579,n21580);
and (n21664,n7471,n7091);
and (n21665,n21666,n21667);
xor (n21666,n21663,n21664);
or (n21667,n21668,n21671);
and (n21668,n21669,n21670);
xor (n21669,n21585,n21586);
and (n21670,n7463,n7091);
and (n21671,n21672,n21673);
xor (n21672,n21669,n21670);
or (n21673,n21674,n21677);
and (n21674,n21675,n21676);
xor (n21675,n21591,n21592);
and (n21676,n7497,n7091);
and (n21677,n21678,n21679);
xor (n21678,n21675,n21676);
or (n21679,n21680,n21683);
and (n21680,n21681,n21682);
xor (n21681,n21596,n21597);
and (n21682,n7084,n7091);
and (n21683,n21684,n21685);
xor (n21684,n21681,n21682);
or (n21685,n21686,n21689);
and (n21686,n21687,n21688);
xor (n21687,n21602,n21603);
and (n21688,n7064,n7091);
and (n21689,n21690,n21691);
xor (n21690,n21687,n21688);
or (n21691,n21692,n21695);
and (n21692,n21693,n21694);
xor (n21693,n21608,n21609);
and (n21694,n7109,n7091);
and (n21695,n21696,n21697);
xor (n21696,n21693,n21694);
or (n21697,n21698,n21701);
and (n21698,n21699,n21700);
xor (n21699,n21613,n21614);
and (n21700,n7102,n7091);
and (n21701,n21702,n21703);
xor (n21702,n21699,n21700);
and (n21703,n21704,n21705);
xor (n21704,n21619,n21620);
and (n21705,n7355,n7091);
and (n21706,n21707,n21708);
xor (n21707,n20716,n10255);
or (n21708,n21709,n21712);
and (n21709,n21710,n21711);
xor (n21710,n21624,n21625);
and (n21711,n7232,n7093);
and (n21712,n21713,n21714);
xor (n21713,n21710,n21711);
or (n21714,n21715,n21717);
and (n21715,n21716,n10121);
xor (n21716,n21630,n21631);
and (n21717,n21718,n21719);
xor (n21718,n21716,n10121);
or (n21719,n21720,n21722);
and (n21720,n21721,n10037);
xor (n21721,n21636,n21637);
and (n21722,n21723,n21724);
xor (n21723,n21721,n10037);
or (n21724,n21725,n21727);
and (n21725,n21726,n9891);
xor (n21726,n21642,n21643);
and (n21727,n21728,n21729);
xor (n21728,n21726,n9891);
or (n21729,n21730,n21732);
and (n21730,n21731,n9775);
xor (n21731,n21648,n21649);
and (n21732,n21733,n21734);
xor (n21733,n21731,n9775);
or (n21734,n21735,n21737);
and (n21735,n21736,n9657);
xor (n21736,n21654,n21655);
and (n21737,n21738,n21739);
xor (n21738,n21736,n9657);
or (n21739,n21740,n21743);
and (n21740,n21741,n21742);
xor (n21741,n21660,n21661);
and (n21742,n7471,n7093);
and (n21743,n21744,n21745);
xor (n21744,n21741,n21742);
or (n21745,n21746,n21749);
and (n21746,n21747,n21748);
xor (n21747,n21666,n21667);
and (n21748,n7463,n7093);
and (n21749,n21750,n21751);
xor (n21750,n21747,n21748);
or (n21751,n21752,n21754);
and (n21752,n21753,n9040);
xor (n21753,n21672,n21673);
and (n21754,n21755,n21756);
xor (n21755,n21753,n9040);
or (n21756,n21757,n21759);
and (n21757,n21758,n9035);
xor (n21758,n21678,n21679);
and (n21759,n21760,n21761);
xor (n21760,n21758,n9035);
or (n21761,n21762,n21764);
and (n21762,n21763,n7993);
xor (n21763,n21684,n21685);
and (n21764,n21765,n21766);
xor (n21765,n21763,n7993);
or (n21766,n21767,n21769);
and (n21767,n21768,n7108);
xor (n21768,n21690,n21691);
and (n21769,n21770,n21771);
xor (n21770,n21768,n7108);
or (n21771,n21772,n21774);
and (n21772,n21773,n7103);
xor (n21773,n21696,n21697);
and (n21774,n21775,n21776);
xor (n21775,n21773,n7103);
and (n21776,n21777,n7357);
xor (n21777,n21702,n21703);
and (n21778,n7242,n7753);
and (n21779,n21780,n21781);
xor (n21780,n20713,n21778);
or (n21781,n21782,n21785);
and (n21782,n21783,n21784);
xor (n21783,n21707,n21708);
and (n21784,n7232,n7753);
and (n21785,n21786,n21787);
xor (n21786,n21783,n21784);
or (n21787,n21788,n21791);
and (n21788,n21789,n21790);
xor (n21789,n21713,n21714);
and (n21790,n7134,n7753);
and (n21791,n21792,n21793);
xor (n21792,n21789,n21790);
or (n21793,n21794,n21797);
and (n21794,n21795,n21796);
xor (n21795,n21718,n21719);
and (n21796,n7129,n7753);
and (n21797,n21798,n21799);
xor (n21798,n21795,n21796);
or (n21799,n21800,n21803);
and (n21800,n21801,n21802);
xor (n21801,n21723,n21724);
and (n21802,n7165,n7753);
and (n21803,n21804,n21805);
xor (n21804,n21801,n21802);
or (n21805,n21806,n21809);
and (n21806,n21807,n21808);
xor (n21807,n21728,n21729);
and (n21808,n7146,n7753);
and (n21809,n21810,n21811);
xor (n21810,n21807,n21808);
or (n21811,n21812,n21815);
and (n21812,n21813,n21814);
xor (n21813,n21733,n21734);
and (n21814,n7308,n7753);
and (n21815,n21816,n21817);
xor (n21816,n21813,n21814);
or (n21817,n21818,n21821);
and (n21818,n21819,n21820);
xor (n21819,n21738,n21739);
and (n21820,n7471,n7753);
and (n21821,n21822,n21823);
xor (n21822,n21819,n21820);
or (n21823,n21824,n21827);
and (n21824,n21825,n21826);
xor (n21825,n21744,n21745);
and (n21826,n7463,n7753);
and (n21827,n21828,n21829);
xor (n21828,n21825,n21826);
or (n21829,n21830,n21833);
and (n21830,n21831,n21832);
xor (n21831,n21750,n21751);
and (n21832,n7497,n7753);
and (n21833,n21834,n21835);
xor (n21834,n21831,n21832);
or (n21835,n21836,n21839);
and (n21836,n21837,n21838);
xor (n21837,n21755,n21756);
and (n21838,n7084,n7753);
and (n21839,n21840,n21841);
xor (n21840,n21837,n21838);
or (n21841,n21842,n21845);
and (n21842,n21843,n21844);
xor (n21843,n21760,n21761);
and (n21844,n7064,n7753);
and (n21845,n21846,n21847);
xor (n21846,n21843,n21844);
or (n21847,n21848,n21851);
and (n21848,n21849,n21850);
xor (n21849,n21765,n21766);
and (n21850,n7109,n7753);
and (n21851,n21852,n21853);
xor (n21852,n21849,n21850);
or (n21853,n21854,n21857);
and (n21854,n21855,n21856);
xor (n21855,n21770,n21771);
and (n21856,n7102,n7753);
and (n21857,n21858,n21859);
xor (n21858,n21855,n21856);
and (n21859,n21860,n21861);
xor (n21860,n21775,n21776);
and (n21861,n7355,n7753);
and (n21862,n21863,n21864);
xor (n21863,n20710,n10347);
or (n21864,n21865,n21867);
and (n21865,n21866,n10295);
xor (n21866,n21780,n21781);
and (n21867,n21868,n21869);
xor (n21868,n21866,n10295);
or (n21869,n21870,n21872);
and (n21870,n21871,n10220);
xor (n21871,n21786,n21787);
and (n21872,n21873,n21874);
xor (n21873,n21871,n10220);
or (n21874,n21875,n21877);
and (n21875,n21876,n10161);
xor (n21876,n21792,n21793);
and (n21877,n21878,n21879);
xor (n21878,n21876,n10161);
or (n21879,n21880,n21882);
and (n21880,n21881,n10083);
xor (n21881,n21798,n21799);
and (n21882,n21883,n21884);
xor (n21883,n21881,n10083);
or (n21884,n21885,n21887);
and (n21885,n21886,n10010);
xor (n21886,n21804,n21805);
and (n21887,n21888,n21889);
xor (n21888,n21886,n10010);
or (n21889,n21890,n21892);
and (n21890,n21891,n9907);
xor (n21891,n21810,n21811);
and (n21892,n21893,n21894);
xor (n21893,n21891,n9907);
or (n21894,n21895,n21898);
and (n21895,n21896,n21897);
xor (n21896,n21816,n21817);
and (n21897,n7471,n7859);
and (n21898,n21899,n21900);
xor (n21899,n21896,n21897);
or (n21900,n21901,n21904);
and (n21901,n21902,n21903);
xor (n21902,n21822,n21823);
and (n21903,n7463,n7859);
and (n21904,n21905,n21906);
xor (n21905,n21902,n21903);
or (n21906,n21907,n21910);
and (n21907,n21908,n21909);
xor (n21908,n21828,n21829);
and (n21909,n7497,n7859);
and (n21910,n21911,n21912);
xor (n21911,n21908,n21909);
or (n21912,n21913,n21915);
and (n21913,n21914,n9270);
xor (n21914,n21834,n21835);
and (n21915,n21916,n21917);
xor (n21916,n21914,n9270);
or (n21917,n21918,n21921);
and (n21918,n21919,n21920);
xor (n21919,n21840,n21841);
and (n21920,n7064,n7859);
and (n21921,n21922,n21923);
xor (n21922,n21919,n21920);
or (n21923,n21924,n21926);
and (n21924,n21925,n9092);
xor (n21925,n21846,n21847);
and (n21926,n21927,n21928);
xor (n21927,n21925,n9092);
or (n21928,n21929,n21931);
and (n21929,n21930,n8008);
xor (n21930,n21852,n21853);
and (n21931,n21932,n21933);
xor (n21932,n21930,n8008);
and (n21933,n21934,n8005);
xor (n21934,n21858,n21859);
and (n21935,n21936,n21937);
xor (n21936,n20707,n10347);
or (n21937,n21938,n21940);
and (n21938,n21939,n10295);
xor (n21939,n21863,n21864);
and (n21940,n21941,n21942);
xor (n21941,n21939,n10295);
or (n21942,n21943,n21945);
and (n21943,n21944,n10220);
xor (n21944,n21868,n21869);
and (n21945,n21946,n21947);
xor (n21946,n21944,n10220);
or (n21947,n21948,n21950);
and (n21948,n21949,n10161);
xor (n21949,n21873,n21874);
and (n21950,n21951,n21952);
xor (n21951,n21949,n10161);
or (n21952,n21953,n21955);
and (n21953,n21954,n10083);
xor (n21954,n21878,n21879);
and (n21955,n21956,n21957);
xor (n21956,n21954,n10083);
or (n21957,n21958,n21960);
and (n21958,n21959,n10010);
xor (n21959,n21883,n21884);
and (n21960,n21961,n21962);
xor (n21961,n21959,n10010);
or (n21962,n21963,n21965);
and (n21963,n21964,n9907);
xor (n21964,n21888,n21889);
and (n21965,n21966,n21967);
xor (n21966,n21964,n9907);
or (n21967,n21968,n21970);
and (n21968,n21969,n21897);
xor (n21969,n21893,n21894);
and (n21970,n21971,n21972);
xor (n21971,n21969,n21897);
or (n21972,n21973,n21975);
and (n21973,n21974,n21903);
xor (n21974,n21899,n21900);
and (n21975,n21976,n21977);
xor (n21976,n21974,n21903);
or (n21977,n21978,n21980);
and (n21978,n21979,n21909);
xor (n21979,n21905,n21906);
and (n21980,n21981,n21982);
xor (n21981,n21979,n21909);
or (n21982,n21983,n21985);
and (n21983,n21984,n9270);
xor (n21984,n21911,n21912);
and (n21985,n21986,n21987);
xor (n21986,n21984,n9270);
or (n21987,n21988,n21990);
and (n21988,n21989,n21920);
xor (n21989,n21916,n21917);
and (n21990,n21991,n21992);
xor (n21991,n21989,n21920);
or (n21992,n21993,n21995);
and (n21993,n21994,n9092);
xor (n21994,n21922,n21923);
and (n21995,n21996,n21997);
xor (n21996,n21994,n9092);
or (n21997,n21998,n22000);
and (n21998,n21999,n8008);
xor (n21999,n21927,n21928);
and (n22000,n22001,n22002);
xor (n22001,n21999,n8008);
and (n22002,n22003,n8005);
xor (n22003,n21932,n21933);
or (n22004,n22005,n22007);
and (n22005,n22006,n10295);
xor (n22006,n21936,n21937);
and (n22007,n22008,n22009);
xor (n22008,n22006,n10295);
or (n22009,n22010,n22012);
and (n22010,n22011,n10220);
xor (n22011,n21941,n21942);
and (n22012,n22013,n22014);
xor (n22013,n22011,n10220);
or (n22014,n22015,n22017);
and (n22015,n22016,n10161);
xor (n22016,n21946,n21947);
and (n22017,n22018,n22019);
xor (n22018,n22016,n10161);
or (n22019,n22020,n22022);
and (n22020,n22021,n10083);
xor (n22021,n21951,n21952);
and (n22022,n22023,n22024);
xor (n22023,n22021,n10083);
or (n22024,n22025,n22027);
and (n22025,n22026,n10010);
xor (n22026,n21956,n21957);
and (n22027,n22028,n22029);
xor (n22028,n22026,n10010);
or (n22029,n22030,n22032);
and (n22030,n22031,n9907);
xor (n22031,n21961,n21962);
and (n22032,n22033,n22034);
xor (n22033,n22031,n9907);
or (n22034,n22035,n22037);
and (n22035,n22036,n21897);
xor (n22036,n21966,n21967);
and (n22037,n22038,n22039);
xor (n22038,n22036,n21897);
or (n22039,n22040,n22042);
and (n22040,n22041,n21903);
xor (n22041,n21971,n21972);
and (n22042,n22043,n22044);
xor (n22043,n22041,n21903);
or (n22044,n22045,n22047);
and (n22045,n22046,n21909);
xor (n22046,n21976,n21977);
and (n22047,n22048,n22049);
xor (n22048,n22046,n21909);
or (n22049,n22050,n22052);
and (n22050,n22051,n9270);
xor (n22051,n21981,n21982);
and (n22052,n22053,n22054);
xor (n22053,n22051,n9270);
or (n22054,n22055,n22057);
and (n22055,n22056,n21920);
xor (n22056,n21986,n21987);
and (n22057,n22058,n22059);
xor (n22058,n22056,n21920);
or (n22059,n22060,n22062);
and (n22060,n22061,n9092);
xor (n22061,n21991,n21992);
and (n22062,n22063,n22064);
xor (n22063,n22061,n9092);
or (n22064,n22065,n22067);
and (n22065,n22066,n8008);
xor (n22066,n21996,n21997);
and (n22067,n22068,n22069);
xor (n22068,n22066,n8008);
and (n22069,n22070,n8005);
xor (n22070,n22001,n22002);
or (n22071,n22072,n22074);
and (n22072,n22073,n10220);
xor (n22073,n22008,n22009);
and (n22074,n22075,n22076);
xor (n22075,n22073,n10220);
or (n22076,n22077,n22079);
and (n22077,n22078,n10161);
xor (n22078,n22013,n22014);
and (n22079,n22080,n22081);
xor (n22080,n22078,n10161);
or (n22081,n22082,n22084);
and (n22082,n22083,n10083);
xor (n22083,n22018,n22019);
and (n22084,n22085,n22086);
xor (n22085,n22083,n10083);
or (n22086,n22087,n22089);
and (n22087,n22088,n10010);
xor (n22088,n22023,n22024);
and (n22089,n22090,n22091);
xor (n22090,n22088,n10010);
or (n22091,n22092,n22094);
and (n22092,n22093,n9907);
xor (n22093,n22028,n22029);
and (n22094,n22095,n22096);
xor (n22095,n22093,n9907);
or (n22096,n22097,n22099);
and (n22097,n22098,n21897);
xor (n22098,n22033,n22034);
and (n22099,n22100,n22101);
xor (n22100,n22098,n21897);
or (n22101,n22102,n22104);
and (n22102,n22103,n21903);
xor (n22103,n22038,n22039);
and (n22104,n22105,n22106);
xor (n22105,n22103,n21903);
or (n22106,n22107,n22109);
and (n22107,n22108,n21909);
xor (n22108,n22043,n22044);
and (n22109,n22110,n22111);
xor (n22110,n22108,n21909);
or (n22111,n22112,n22114);
and (n22112,n22113,n9270);
xor (n22113,n22048,n22049);
and (n22114,n22115,n22116);
xor (n22115,n22113,n9270);
or (n22116,n22117,n22119);
and (n22117,n22118,n21920);
xor (n22118,n22053,n22054);
and (n22119,n22120,n22121);
xor (n22120,n22118,n21920);
or (n22121,n22122,n22124);
and (n22122,n22123,n9092);
xor (n22123,n22058,n22059);
and (n22124,n22125,n22126);
xor (n22125,n22123,n9092);
or (n22126,n22127,n22129);
and (n22127,n22128,n8008);
xor (n22128,n22063,n22064);
and (n22129,n22130,n22131);
xor (n22130,n22128,n8008);
and (n22131,n22132,n8005);
xor (n22132,n22068,n22069);
or (n22133,n22134,n22136);
and (n22134,n22135,n10161);
xor (n22135,n22075,n22076);
and (n22136,n22137,n22138);
xor (n22137,n22135,n10161);
or (n22138,n22139,n22141);
and (n22139,n22140,n10083);
xor (n22140,n22080,n22081);
and (n22141,n22142,n22143);
xor (n22142,n22140,n10083);
or (n22143,n22144,n22146);
and (n22144,n22145,n10010);
xor (n22145,n22085,n22086);
and (n22146,n22147,n22148);
xor (n22147,n22145,n10010);
or (n22148,n22149,n22151);
and (n22149,n22150,n9907);
xor (n22150,n22090,n22091);
and (n22151,n22152,n22153);
xor (n22152,n22150,n9907);
or (n22153,n22154,n22156);
and (n22154,n22155,n21897);
xor (n22155,n22095,n22096);
and (n22156,n22157,n22158);
xor (n22157,n22155,n21897);
or (n22158,n22159,n22161);
and (n22159,n22160,n21903);
xor (n22160,n22100,n22101);
and (n22161,n22162,n22163);
xor (n22162,n22160,n21903);
or (n22163,n22164,n22166);
and (n22164,n22165,n21909);
xor (n22165,n22105,n22106);
and (n22166,n22167,n22168);
xor (n22167,n22165,n21909);
or (n22168,n22169,n22171);
and (n22169,n22170,n9270);
xor (n22170,n22110,n22111);
and (n22171,n22172,n22173);
xor (n22172,n22170,n9270);
or (n22173,n22174,n22176);
and (n22174,n22175,n21920);
xor (n22175,n22115,n22116);
and (n22176,n22177,n22178);
xor (n22177,n22175,n21920);
or (n22178,n22179,n22181);
and (n22179,n22180,n9092);
xor (n22180,n22120,n22121);
and (n22181,n22182,n22183);
xor (n22182,n22180,n9092);
or (n22183,n22184,n22186);
and (n22184,n22185,n8008);
xor (n22185,n22125,n22126);
and (n22186,n22187,n22188);
xor (n22187,n22185,n8008);
and (n22188,n22189,n8005);
xor (n22189,n22130,n22131);
or (n22190,n22191,n22193);
and (n22191,n22192,n10083);
xor (n22192,n22137,n22138);
and (n22193,n22194,n22195);
xor (n22194,n22192,n10083);
or (n22195,n22196,n22198);
and (n22196,n22197,n10010);
xor (n22197,n22142,n22143);
and (n22198,n22199,n22200);
xor (n22199,n22197,n10010);
or (n22200,n22201,n22203);
and (n22201,n22202,n9907);
xor (n22202,n22147,n22148);
and (n22203,n22204,n22205);
xor (n22204,n22202,n9907);
or (n22205,n22206,n22208);
and (n22206,n22207,n21897);
xor (n22207,n22152,n22153);
and (n22208,n22209,n22210);
xor (n22209,n22207,n21897);
or (n22210,n22211,n22213);
and (n22211,n22212,n21903);
xor (n22212,n22157,n22158);
and (n22213,n22214,n22215);
xor (n22214,n22212,n21903);
or (n22215,n22216,n22218);
and (n22216,n22217,n21909);
xor (n22217,n22162,n22163);
and (n22218,n22219,n22220);
xor (n22219,n22217,n21909);
or (n22220,n22221,n22223);
and (n22221,n22222,n9270);
xor (n22222,n22167,n22168);
and (n22223,n22224,n22225);
xor (n22224,n22222,n9270);
or (n22225,n22226,n22228);
and (n22226,n22227,n21920);
xor (n22227,n22172,n22173);
and (n22228,n22229,n22230);
xor (n22229,n22227,n21920);
or (n22230,n22231,n22233);
and (n22231,n22232,n9092);
xor (n22232,n22177,n22178);
and (n22233,n22234,n22235);
xor (n22234,n22232,n9092);
or (n22235,n22236,n22238);
and (n22236,n22237,n8008);
xor (n22237,n22182,n22183);
and (n22238,n22239,n22240);
xor (n22239,n22237,n8008);
and (n22240,n22241,n8005);
xor (n22241,n22187,n22188);
or (n22242,n22243,n22245);
and (n22243,n22244,n10010);
xor (n22244,n22194,n22195);
and (n22245,n22246,n22247);
xor (n22246,n22244,n10010);
or (n22247,n22248,n22250);
and (n22248,n22249,n9907);
xor (n22249,n22199,n22200);
and (n22250,n22251,n22252);
xor (n22251,n22249,n9907);
or (n22252,n22253,n22255);
and (n22253,n22254,n21897);
xor (n22254,n22204,n22205);
and (n22255,n22256,n22257);
xor (n22256,n22254,n21897);
or (n22257,n22258,n22260);
and (n22258,n22259,n21903);
xor (n22259,n22209,n22210);
and (n22260,n22261,n22262);
xor (n22261,n22259,n21903);
or (n22262,n22263,n22265);
and (n22263,n22264,n21909);
xor (n22264,n22214,n22215);
and (n22265,n22266,n22267);
xor (n22266,n22264,n21909);
or (n22267,n22268,n22270);
and (n22268,n22269,n9270);
xor (n22269,n22219,n22220);
and (n22270,n22271,n22272);
xor (n22271,n22269,n9270);
or (n22272,n22273,n22275);
and (n22273,n22274,n21920);
xor (n22274,n22224,n22225);
and (n22275,n22276,n22277);
xor (n22276,n22274,n21920);
or (n22277,n22278,n22280);
and (n22278,n22279,n9092);
xor (n22279,n22229,n22230);
and (n22280,n22281,n22282);
xor (n22281,n22279,n9092);
or (n22282,n22283,n22285);
and (n22283,n22284,n8008);
xor (n22284,n22234,n22235);
and (n22285,n22286,n22287);
xor (n22286,n22284,n8008);
and (n22287,n22288,n8005);
xor (n22288,n22239,n22240);
or (n22289,n22290,n22292);
and (n22290,n22291,n9907);
xor (n22291,n22246,n22247);
and (n22292,n22293,n22294);
xor (n22293,n22291,n9907);
or (n22294,n22295,n22297);
and (n22295,n22296,n21897);
xor (n22296,n22251,n22252);
and (n22297,n22298,n22299);
xor (n22298,n22296,n21897);
or (n22299,n22300,n22302);
and (n22300,n22301,n21903);
xor (n22301,n22256,n22257);
and (n22302,n22303,n22304);
xor (n22303,n22301,n21903);
or (n22304,n22305,n22307);
and (n22305,n22306,n21909);
xor (n22306,n22261,n22262);
and (n22307,n22308,n22309);
xor (n22308,n22306,n21909);
or (n22309,n22310,n22312);
and (n22310,n22311,n9270);
xor (n22311,n22266,n22267);
and (n22312,n22313,n22314);
xor (n22313,n22311,n9270);
or (n22314,n22315,n22317);
and (n22315,n22316,n21920);
xor (n22316,n22271,n22272);
and (n22317,n22318,n22319);
xor (n22318,n22316,n21920);
or (n22319,n22320,n22322);
and (n22320,n22321,n9092);
xor (n22321,n22276,n22277);
and (n22322,n22323,n22324);
xor (n22323,n22321,n9092);
or (n22324,n22325,n22327);
and (n22325,n22326,n8008);
xor (n22326,n22281,n22282);
and (n22327,n22328,n22329);
xor (n22328,n22326,n8008);
and (n22329,n22330,n8005);
xor (n22330,n22286,n22287);
or (n22331,n22332,n22334);
and (n22332,n22333,n21897);
xor (n22333,n22293,n22294);
and (n22334,n22335,n22336);
xor (n22335,n22333,n21897);
or (n22336,n22337,n22339);
and (n22337,n22338,n21903);
xor (n22338,n22298,n22299);
and (n22339,n22340,n22341);
xor (n22340,n22338,n21903);
or (n22341,n22342,n22344);
and (n22342,n22343,n21909);
xor (n22343,n22303,n22304);
and (n22344,n22345,n22346);
xor (n22345,n22343,n21909);
or (n22346,n22347,n22349);
and (n22347,n22348,n9270);
xor (n22348,n22308,n22309);
and (n22349,n22350,n22351);
xor (n22350,n22348,n9270);
or (n22351,n22352,n22354);
and (n22352,n22353,n21920);
xor (n22353,n22313,n22314);
and (n22354,n22355,n22356);
xor (n22355,n22353,n21920);
or (n22356,n22357,n22359);
and (n22357,n22358,n9092);
xor (n22358,n22318,n22319);
and (n22359,n22360,n22361);
xor (n22360,n22358,n9092);
or (n22361,n22362,n22364);
and (n22362,n22363,n8008);
xor (n22363,n22323,n22324);
and (n22364,n22365,n22366);
xor (n22365,n22363,n8008);
and (n22366,n22367,n8005);
xor (n22367,n22328,n22329);
or (n22368,n22369,n22371);
and (n22369,n22370,n21903);
xor (n22370,n22335,n22336);
and (n22371,n22372,n22373);
xor (n22372,n22370,n21903);
or (n22373,n22374,n22376);
and (n22374,n22375,n21909);
xor (n22375,n22340,n22341);
and (n22376,n22377,n22378);
xor (n22377,n22375,n21909);
or (n22378,n22379,n22381);
and (n22379,n22380,n9270);
xor (n22380,n22345,n22346);
and (n22381,n22382,n22383);
xor (n22382,n22380,n9270);
or (n22383,n22384,n22386);
and (n22384,n22385,n21920);
xor (n22385,n22350,n22351);
and (n22386,n22387,n22388);
xor (n22387,n22385,n21920);
or (n22388,n22389,n22391);
and (n22389,n22390,n9092);
xor (n22390,n22355,n22356);
and (n22391,n22392,n22393);
xor (n22392,n22390,n9092);
or (n22393,n22394,n22396);
and (n22394,n22395,n8008);
xor (n22395,n22360,n22361);
and (n22396,n22397,n22398);
xor (n22397,n22395,n8008);
and (n22398,n22399,n8005);
xor (n22399,n22365,n22366);
or (n22400,n22401,n22403);
and (n22401,n22402,n21909);
xor (n22402,n22372,n22373);
and (n22403,n22404,n22405);
xor (n22404,n22402,n21909);
or (n22405,n22406,n22408);
and (n22406,n22407,n9270);
xor (n22407,n22377,n22378);
and (n22408,n22409,n22410);
xor (n22409,n22407,n9270);
or (n22410,n22411,n22413);
and (n22411,n22412,n21920);
xor (n22412,n22382,n22383);
and (n22413,n22414,n22415);
xor (n22414,n22412,n21920);
or (n22415,n22416,n22418);
and (n22416,n22417,n9092);
xor (n22417,n22387,n22388);
and (n22418,n22419,n22420);
xor (n22419,n22417,n9092);
or (n22420,n22421,n22423);
and (n22421,n22422,n8008);
xor (n22422,n22392,n22393);
and (n22423,n22424,n22425);
xor (n22424,n22422,n8008);
and (n22425,n22426,n8005);
xor (n22426,n22397,n22398);
or (n22427,n22428,n22430);
and (n22428,n22429,n9270);
xor (n22429,n22404,n22405);
and (n22430,n22431,n22432);
xor (n22431,n22429,n9270);
or (n22432,n22433,n22435);
and (n22433,n22434,n21920);
xor (n22434,n22409,n22410);
and (n22435,n22436,n22437);
xor (n22436,n22434,n21920);
or (n22437,n22438,n22440);
and (n22438,n22439,n9092);
xor (n22439,n22414,n22415);
and (n22440,n22441,n22442);
xor (n22441,n22439,n9092);
or (n22442,n22443,n22445);
and (n22443,n22444,n8008);
xor (n22444,n22419,n22420);
and (n22445,n22446,n22447);
xor (n22446,n22444,n8008);
and (n22447,n22448,n8005);
xor (n22448,n22424,n22425);
or (n22449,n22450,n22452);
and (n22450,n22451,n21920);
xor (n22451,n22431,n22432);
and (n22452,n22453,n22454);
xor (n22453,n22451,n21920);
or (n22454,n22455,n22457);
and (n22455,n22456,n9092);
xor (n22456,n22436,n22437);
and (n22457,n22458,n22459);
xor (n22458,n22456,n9092);
or (n22459,n22460,n22462);
and (n22460,n22461,n8008);
xor (n22461,n22441,n22442);
and (n22462,n22463,n22464);
xor (n22463,n22461,n8008);
and (n22464,n22465,n8005);
xor (n22465,n22446,n22447);
or (n22466,n22467,n22469);
and (n22467,n22468,n9092);
xor (n22468,n22453,n22454);
and (n22469,n22470,n22471);
xor (n22470,n22468,n9092);
or (n22471,n22472,n22474);
and (n22472,n22473,n8008);
xor (n22473,n22458,n22459);
and (n22474,n22475,n22476);
xor (n22475,n22473,n8008);
and (n22476,n22477,n8005);
xor (n22477,n22463,n22464);
or (n22478,n22479,n22481);
and (n22479,n22480,n8008);
xor (n22480,n22470,n22471);
and (n22481,n22482,n22483);
xor (n22482,n22480,n8008);
and (n22483,n22484,n8005);
xor (n22484,n22475,n22476);
and (n22485,n22486,n8005);
xor (n22486,n22482,n22483);
or (n22487,n22488,n22492,n22699);
and (n22488,n22489,n22490);
xor (n22489,n20615,n7977);
not (n22490,n22491);
xor (n22491,n22486,n8005);
and (n22492,n22490,n22493);
or (n22493,n22494,n22498,n22698);
and (n22494,n22495,n22496);
xor (n22495,n20613,n7977);
not (n22496,n22497);
xor (n22497,n22484,n8005);
and (n22498,n22496,n22499);
or (n22499,n22500,n22504,n22697);
and (n22500,n22501,n22502);
xor (n22501,n20606,n7977);
not (n22502,n22503);
xor (n22503,n22477,n8005);
and (n22504,n22502,n22505);
or (n22505,n22506,n22510,n22696);
and (n22506,n22507,n22508);
xor (n22507,n20594,n7977);
not (n22508,n22509);
xor (n22509,n22465,n8005);
and (n22510,n22508,n22511);
or (n22511,n22512,n22516,n22695);
and (n22512,n22513,n22514);
xor (n22513,n20577,n7977);
not (n22514,n22515);
xor (n22515,n22448,n8005);
and (n22516,n22514,n22517);
or (n22517,n22518,n22522,n22694);
and (n22518,n22519,n22520);
xor (n22519,n20555,n7977);
not (n22520,n22521);
xor (n22521,n22426,n8005);
and (n22522,n22520,n22523);
or (n22523,n22524,n22528,n22693);
and (n22524,n22525,n22526);
xor (n22525,n20528,n7977);
not (n22526,n22527);
xor (n22527,n22399,n8005);
and (n22528,n22526,n22529);
or (n22529,n22530,n22534,n22692);
and (n22530,n22531,n22532);
xor (n22531,n20496,n7977);
not (n22532,n22533);
xor (n22533,n22367,n8005);
and (n22534,n22532,n22535);
or (n22535,n22536,n22540,n22691);
and (n22536,n22537,n22538);
xor (n22537,n20459,n7977);
not (n22538,n22539);
xor (n22539,n22330,n8005);
and (n22540,n22538,n22541);
or (n22541,n22542,n22546,n22690);
and (n22542,n22543,n22544);
xor (n22543,n20417,n7977);
not (n22544,n22545);
xor (n22545,n22288,n8005);
and (n22546,n22544,n22547);
or (n22547,n22548,n22552,n22689);
and (n22548,n22549,n22550);
xor (n22549,n20370,n7977);
not (n22550,n22551);
xor (n22551,n22241,n8005);
and (n22552,n22550,n22553);
or (n22553,n22554,n22558,n22688);
and (n22554,n22555,n22556);
xor (n22555,n20318,n7977);
not (n22556,n22557);
xor (n22557,n22189,n8005);
and (n22558,n22556,n22559);
or (n22559,n22560,n22564,n22687);
and (n22560,n22561,n22562);
xor (n22561,n20261,n7977);
not (n22562,n22563);
xor (n22563,n22132,n8005);
and (n22564,n22562,n22565);
or (n22565,n22566,n22570,n22686);
and (n22566,n22567,n22568);
xor (n22567,n20199,n7977);
not (n22568,n22569);
xor (n22569,n22070,n8005);
and (n22570,n22568,n22571);
or (n22571,n22572,n22576,n22685);
and (n22572,n22573,n22574);
xor (n22573,n20132,n7977);
not (n22574,n22575);
xor (n22575,n22003,n8005);
and (n22576,n22574,n22577);
or (n22577,n22578,n22582,n22684);
and (n22578,n22579,n22580);
xor (n22579,n20063,n7977);
not (n22580,n22581);
xor (n22581,n21934,n8005);
and (n22582,n22580,n22583);
or (n22583,n22584,n22588,n22683);
and (n22584,n22585,n22586);
xor (n22585,n19983,n7849);
not (n22586,n22587);
xor (n22587,n21860,n21861);
and (n22588,n22586,n22589);
or (n22589,n22590,n22594,n22682);
and (n22590,n22591,n22592);
xor (n22591,n19899,n19900);
not (n22592,n22593);
xor (n22593,n21777,n7357);
and (n22594,n22592,n22595);
or (n22595,n22596,n22600,n22681);
and (n22596,n22597,n22598);
xor (n22597,n19823,n7365);
not (n22598,n22599);
xor (n22599,n21704,n21705);
and (n22600,n22598,n22601);
or (n22601,n22602,n22606,n22680);
and (n22602,n22603,n22604);
xor (n22603,n19739,n19740);
not (n22604,n22605);
xor (n22605,n21621,n7543);
and (n22606,n22604,n22607);
or (n22607,n22608,n22612,n22679);
and (n22608,n22609,n22610);
xor (n22609,n19663,n7577);
not (n22610,n22611);
xor (n22611,n21544,n21545);
and (n22612,n22610,n22613);
or (n22613,n22614,n22618,n22678);
and (n22614,n22615,n22616);
xor (n22615,n19580,n8209);
not (n22616,n22617);
xor (n22617,n21461,n8222);
and (n22618,n22616,n22619);
or (n22619,n22620,n22624,n22677);
and (n22620,n22621,n22622);
xor (n22621,n19504,n8232);
not (n22622,n22623);
xor (n22623,n21384,n21385);
and (n22624,n22622,n22625);
or (n22625,n22626,n22630,n22676);
and (n22626,n22627,n22628);
xor (n22627,n19420,n19421);
not (n22628,n22629);
xor (n22629,n21301,n8470);
and (n22630,n22628,n22631);
or (n22631,n22632,n22636,n22675);
and (n22632,n22633,n22634);
xor (n22633,n19342,n8439);
not (n22634,n22635);
xor (n22635,n21225,n21226);
and (n22636,n22634,n22637);
or (n22637,n22638,n22642,n22674);
and (n22638,n22639,n22640);
xor (n22639,n19258,n19259);
not (n22640,n22641);
xor (n22641,n21142,n8624);
and (n22642,n22640,n22643);
or (n22643,n22644,n22648,n22673);
and (n22644,n22645,n22646);
xor (n22645,n19179,n8670);
not (n22646,n22647);
xor (n22647,n21066,n21067);
and (n22648,n22646,n22649);
or (n22649,n22650,n22654,n22672);
and (n22650,n22651,n22652);
xor (n22651,n19095,n19096);
not (n22652,n22653);
xor (n22653,n20983,n8781);
and (n22654,n22652,n22655);
or (n22655,n22656,n22660,n22671);
and (n22656,n22657,n22658);
xor (n22657,n19019,n8745);
not (n22658,n22659);
xor (n22659,n20908,n20909);
and (n22660,n22658,n22661);
or (n22661,n22662,n22666,n22670);
and (n22662,n22663,n22664);
xor (n22663,n18935,n18936);
not (n22664,n22665);
xor (n22665,n20825,n8840);
and (n22666,n22664,n22667);
or (n22667,n8832,n22668);
not (n22668,n22669);
and (n22669,n7355,n7237);
and (n22670,n22663,n22667);
and (n22671,n22657,n22661);
and (n22672,n22651,n22655);
and (n22673,n22645,n22649);
and (n22674,n22639,n22643);
and (n22675,n22633,n22637);
and (n22676,n22627,n22631);
and (n22677,n22621,n22625);
and (n22678,n22615,n22619);
and (n22679,n22609,n22613);
and (n22680,n22603,n22607);
and (n22681,n22597,n22601);
and (n22682,n22591,n22595);
and (n22683,n22585,n22589);
and (n22684,n22579,n22583);
and (n22685,n22573,n22577);
and (n22686,n22567,n22571);
and (n22687,n22561,n22565);
and (n22688,n22555,n22559);
and (n22689,n22549,n22553);
and (n22690,n22543,n22547);
and (n22691,n22537,n22541);
and (n22692,n22531,n22535);
and (n22693,n22525,n22529);
and (n22694,n22519,n22523);
and (n22695,n22513,n22517);
and (n22696,n22507,n22511);
and (n22697,n22501,n22505);
and (n22698,n22495,n22499);
and (n22699,n22489,n22493);
and (n22700,n10717,n22701);
not (n22701,n10713);
endmodule
