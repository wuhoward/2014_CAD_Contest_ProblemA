module top (out,n21,n26,n27,n28,n30,n31,n42,n45,n48
        ,n51,n54,n57,n60,n63,n66,n69,n72,n75,n78
        ,n81,n84,n87,n90,n93,n95,n98,n101,n111,n121
        ,n128,n133,n168,n173,n176,n179,n182,n185,n188,n191
        ,n194,n197,n200,n203,n206,n209,n212,n215,n218,n227
        ,n495,n546);
output out;
input n21;
input n26;
input n27;
input n28;
input n30;
input n31;
input n42;
input n45;
input n48;
input n51;
input n54;
input n57;
input n60;
input n63;
input n66;
input n69;
input n72;
input n75;
input n78;
input n81;
input n84;
input n87;
input n90;
input n93;
input n95;
input n98;
input n101;
input n111;
input n121;
input n128;
input n133;
input n168;
input n173;
input n176;
input n179;
input n182;
input n185;
input n188;
input n191;
input n194;
input n197;
input n200;
input n203;
input n206;
input n209;
input n212;
input n215;
input n218;
input n227;
input n495;
input n546;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n29;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n46;
wire n47;
wire n49;
wire n50;
wire n52;
wire n53;
wire n55;
wire n56;
wire n58;
wire n59;
wire n61;
wire n62;
wire n64;
wire n65;
wire n67;
wire n68;
wire n70;
wire n71;
wire n73;
wire n74;
wire n76;
wire n77;
wire n79;
wire n80;
wire n82;
wire n83;
wire n85;
wire n86;
wire n88;
wire n89;
wire n91;
wire n92;
wire n94;
wire n96;
wire n97;
wire n99;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n177;
wire n178;
wire n180;
wire n181;
wire n183;
wire n184;
wire n186;
wire n187;
wire n189;
wire n190;
wire n192;
wire n193;
wire n195;
wire n196;
wire n198;
wire n199;
wire n201;
wire n202;
wire n204;
wire n205;
wire n207;
wire n208;
wire n210;
wire n211;
wire n213;
wire n214;
wire n216;
wire n217;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
xor (out,n0,n1776);
nand (n0,n1,n1775);
or (n1,n2,n896);
not (n2,n3);
nor (n3,n4,n895);
nor (n4,n5,n832);
not (n5,n6);
xor (n6,n7,n747);
xor (n7,n8,n558);
xor (n8,n9,n476);
xor (n9,n10,n339);
xor (n10,n11,n233);
xor (n11,n12,n136);
nand (n12,n13,n123);
or (n13,n14,n117);
nand (n14,n15,n107);
nor (n15,n16,n105);
and (n16,n17,n99);
not (n17,n18);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n96);
and (s0n18,notn18,n19);
and (s1n18,n96,n38);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,1'b0);
and (s1n19,n22,n21);
or (n22,n23,n34);
or (n23,n24,n32);
nor (n24,n25,n27,n28,n29,n31);
not (n25,n26);
not (n29,n30);
nor (n32,n26,n33,n28,n29,n31);
not (n33,n27);
or (n34,n35,n37);
and (n35,n25,n27,n28,n29,n36);
not (n36,n31);
nor (n37,n25,n33,n28,n29,n31);
xor (n38,n39,n40);
not (n39,n21);
and (n40,n41,n43);
not (n41,n42);
and (n43,n44,n46);
not (n44,n45);
and (n46,n47,n49);
not (n47,n48);
and (n49,n50,n52);
not (n50,n51);
and (n52,n53,n55);
not (n53,n54);
and (n55,n56,n58);
not (n56,n57);
and (n58,n59,n61);
not (n59,n60);
and (n61,n62,n64);
not (n62,n63);
and (n64,n65,n67);
not (n65,n66);
and (n67,n68,n70);
not (n68,n69);
and (n70,n71,n73);
not (n71,n72);
and (n73,n74,n76);
not (n74,n75);
and (n76,n77,n79);
not (n77,n78);
and (n79,n80,n82);
not (n80,n81);
and (n82,n83,n85);
not (n83,n84);
and (n85,n86,n88);
not (n86,n87);
and (n88,n89,n91);
not (n89,n90);
and (n91,n92,n94);
not (n92,n93);
not (n94,n95);
and (n96,n97,n98);
or (n97,n24,n35);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n96);
and (s0n99,notn99,n100);
and (s1n99,n96,n102);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n22);
and (s0n100,notn100,1'b0);
and (s1n100,n22,n101);
xor (n102,n103,n104);
not (n103,n101);
and (n104,n39,n40);
and (n105,n18,n106);
not (n106,n99);
nand (n107,n108,n115);
or (n108,n106,n109);
wire s0n109,s1n109,notn109;
or (n109,s0n109,s1n109);
not(notn109,n96);
and (s0n109,notn109,n110);
and (s1n109,n96,n112);
wire s0n110,s1n110,notn110;
or (n110,s0n110,s1n110);
not(notn110,n22);
and (s0n110,notn110,1'b0);
and (s1n110,n22,n111);
xor (n112,n113,n114);
not (n113,n111);
and (n114,n103,n104);
or (n115,n99,n116);
not (n116,n109);
nor (n117,n118,n122);
and (n118,n109,n119);
not (n119,n120);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n22);
and (s0n120,notn120,1'b0);
and (s1n120,n22,n121);
and (n122,n116,n120);
or (n123,n15,n124);
nor (n124,n125,n134);
and (n125,n126,n116);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n132);
and (s0n126,notn126,n127);
and (s1n126,n132,n129);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n22);
and (s0n127,notn127,1'b0);
and (s1n127,n22,n128);
xor (n129,n130,n131);
not (n130,n128);
not (n131,n121);
and (n132,n97,n133);
and (n134,n135,n109);
not (n135,n126);
xor (n136,n137,n143);
nor (n137,n138,n116);
nor (n138,n139,n142);
and (n139,n140,n17);
not (n140,n141);
and (n141,n120,n99);
and (n142,n106,n119);
nand (n143,n144,n222);
or (n144,n145,n164);
nand (n145,n146,n157);
nor (n146,n147,n155);
and (n147,n148,n152);
not (n148,n149);
wire s0n149,s1n149,notn149;
or (n149,s0n149,s1n149);
not(notn149,n96);
and (s0n149,notn149,n150);
and (s1n149,n96,n151);
wire s0n150,s1n150,notn150;
or (n150,s0n150,s1n150);
not(notn150,n22);
and (s0n150,notn150,1'b0);
and (s1n150,n22,n93);
xor (n151,n92,n94);
wire s0n152,s1n152,notn152;
or (n152,s0n152,s1n152);
not(notn152,n96);
and (s0n152,notn152,n153);
and (s1n152,n96,n154);
wire s0n153,s1n153,notn153;
or (n153,s0n153,s1n153);
not(notn153,n22);
and (s0n153,notn153,1'b0);
and (s1n153,n22,n90);
xor (n154,n89,n91);
and (n155,n149,n156);
not (n156,n152);
nand (n157,n158,n163);
or (n158,n159,n152);
not (n159,n160);
wire s0n160,s1n160,notn160;
or (n160,s0n160,s1n160);
not(notn160,n96);
and (s0n160,notn160,n161);
and (s1n160,n96,n162);
wire s0n161,s1n161,notn161;
or (n161,s0n161,s1n161);
not(notn161,n22);
and (s0n161,notn161,1'b0);
and (s1n161,n22,n87);
xor (n162,n86,n88);
nand (n163,n159,n152);
nor (n164,n165,n220);
and (n165,n166,n159);
wire s0n166,s1n166,notn166;
or (n166,s0n166,s1n166);
not(notn166,n132);
and (s0n166,notn166,n167);
and (s1n166,n132,n169);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n22);
and (s0n167,notn167,1'b0);
and (s1n167,n22,n168);
xor (n169,n170,n171);
not (n170,n168);
and (n171,n172,n174);
not (n172,n173);
and (n174,n175,n177);
not (n175,n176);
and (n177,n178,n180);
not (n178,n179);
and (n180,n181,n183);
not (n181,n182);
and (n183,n184,n186);
not (n184,n185);
and (n186,n187,n189);
not (n187,n188);
and (n189,n190,n192);
not (n190,n191);
and (n192,n193,n195);
not (n193,n194);
and (n195,n196,n198);
not (n196,n197);
and (n198,n199,n201);
not (n199,n200);
and (n201,n202,n204);
not (n202,n203);
and (n204,n205,n207);
not (n205,n206);
and (n207,n208,n210);
not (n208,n209);
and (n210,n211,n213);
not (n211,n212);
and (n213,n214,n216);
not (n214,n215);
and (n216,n217,n219);
not (n217,n218);
and (n219,n130,n131);
and (n220,n221,n160);
not (n221,n166);
or (n222,n146,n223);
nor (n223,n224,n231);
and (n224,n225,n159);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n132);
and (s0n225,notn225,n226);
and (s1n225,n132,n228);
wire s0n226,s1n226,notn226;
or (n226,s0n226,s1n226);
not(notn226,n22);
and (s0n226,notn226,1'b0);
and (s1n226,n22,n227);
xor (n228,n229,n230);
not (n229,n227);
and (n230,n170,n171);
and (n231,n232,n160);
not (n232,n225);
or (n233,n234,n338);
and (n234,n235,n306);
xor (n235,n236,n273);
nand (n236,n237,n265);
or (n237,n238,n258);
nand (n238,n239,n250);
nor (n239,n240,n247);
and (n240,n241,n244);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n96);
and (s0n241,notn241,n242);
and (s1n241,n96,n243);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n22);
and (s0n242,notn242,1'b0);
and (s1n242,n22,n72);
xor (n243,n71,n73);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n96);
and (s0n244,notn244,n245);
and (s1n244,n96,n246);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n22);
and (s0n245,notn245,1'b0);
and (s1n245,n22,n69);
xor (n246,n68,n70);
and (n247,n248,n249);
not (n248,n241);
not (n249,n244);
not (n250,n251);
nor (n251,n252,n256);
and (n252,n253,n241);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n96);
and (s0n253,notn253,n254);
and (s1n253,n96,n255);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n22);
and (s0n254,notn254,1'b0);
and (s1n254,n22,n75);
xor (n255,n74,n76);
and (n256,n257,n248);
not (n257,n253);
nor (n258,n259,n263);
and (n259,n249,n260);
wire s0n260,s1n260,notn260;
or (n260,s0n260,s1n260);
not(notn260,n132);
and (s0n260,notn260,n261);
and (s1n260,n132,n262);
wire s0n261,s1n261,notn261;
or (n261,s0n261,s1n261);
not(notn261,n22);
and (s0n261,notn261,1'b0);
and (s1n261,n22,n191);
xor (n262,n190,n192);
and (n263,n244,n264);
not (n264,n260);
or (n265,n266,n250);
nor (n266,n267,n271);
and (n267,n249,n268);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n132);
and (s0n268,notn268,n269);
and (s1n268,n132,n270);
wire s0n269,s1n269,notn269;
or (n269,s0n269,s1n269);
not(notn269,n22);
and (s0n269,notn269,1'b0);
and (s1n269,n22,n188);
xor (n270,n187,n189);
and (n271,n244,n272);
not (n272,n268);
nand (n273,n274,n298);
or (n274,n275,n291);
nand (n275,n276,n283);
not (n276,n277);
nand (n277,n278,n282);
or (n278,n159,n279);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n96);
and (s0n279,notn279,n280);
and (s1n279,n96,n281);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n22);
and (s0n280,notn280,1'b0);
and (s1n280,n22,n84);
xor (n281,n83,n85);
nand (n282,n279,n159);
nor (n283,n284,n290);
and (n284,n285,n289);
not (n285,n286);
wire s0n286,s1n286,notn286;
or (n286,s0n286,s1n286);
not(notn286,n96);
and (s0n286,notn286,n287);
and (s1n286,n96,n288);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n22);
and (s0n287,notn287,1'b0);
and (s1n287,n22,n81);
xor (n288,n80,n82);
not (n289,n279);
and (n290,n286,n279);
nor (n291,n292,n296);
and (n292,n293,n285);
wire s0n293,s1n293,notn293;
or (n293,s0n293,s1n293);
not(notn293,n132);
and (s0n293,notn293,n294);
and (s1n293,n132,n295);
wire s0n294,s1n294,notn294;
or (n294,s0n294,s1n294);
not(notn294,n22);
and (s0n294,notn294,1'b0);
and (s1n294,n22,n179);
xor (n295,n178,n180);
and (n296,n297,n286);
not (n297,n293);
or (n298,n276,n299);
nor (n299,n300,n304);
and (n300,n301,n285);
wire s0n301,s1n301,notn301;
or (n301,s0n301,s1n301);
not(notn301,n132);
and (s0n301,notn301,n302);
and (s1n301,n132,n303);
wire s0n302,s1n302,notn302;
or (n302,s0n302,s1n302);
not(notn302,n22);
and (s0n302,notn302,1'b0);
and (s1n302,n22,n176);
xor (n303,n175,n177);
and (n304,n305,n286);
not (n305,n301);
nand (n306,n307,n330);
or (n307,n308,n323);
nand (n308,n309,n316);
or (n309,n310,n314);
and (n310,n311,n244);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n96);
and (s0n311,notn311,n312);
and (s1n311,n96,n313);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n22);
and (s0n312,notn312,1'b0);
and (s1n312,n22,n66);
xor (n313,n65,n67);
and (n314,n315,n249);
not (n315,n311);
nand (n316,n317,n321);
or (n317,n315,n318);
wire s0n318,s1n318,notn318;
or (n318,s0n318,s1n318);
not(notn318,n96);
and (s0n318,notn318,n319);
and (s1n318,n96,n320);
wire s0n319,s1n319,notn319;
or (n319,s0n319,s1n319);
not(notn319,n22);
and (s0n319,notn319,1'b0);
and (s1n319,n22,n63);
xor (n320,n62,n64);
or (n321,n322,n311);
not (n322,n318);
nor (n323,n324,n328);
and (n324,n322,n325);
wire s0n325,s1n325,notn325;
or (n325,s0n325,s1n325);
not(notn325,n132);
and (s0n325,notn325,n326);
and (s1n325,n132,n327);
wire s0n326,s1n326,notn326;
or (n326,s0n326,s1n326);
not(notn326,n22);
and (s0n326,notn326,1'b0);
and (s1n326,n22,n197);
xor (n327,n196,n198);
and (n328,n318,n329);
not (n329,n325);
or (n330,n309,n331);
nor (n331,n332,n336);
and (n332,n322,n333);
wire s0n333,s1n333,notn333;
or (n333,s0n333,s1n333);
not(notn333,n132);
and (s0n333,notn333,n334);
and (s1n333,n132,n335);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n22);
and (s0n334,notn334,1'b0);
and (s1n334,n22,n194);
xor (n335,n193,n195);
and (n336,n318,n337);
not (n337,n333);
and (n338,n236,n273);
or (n339,n340,n475);
and (n340,n341,n474);
xor (n341,n342,n441);
or (n342,n343,n440);
and (n343,n344,n407);
xor (n344,n345,n369);
nand (n345,n346,n361);
or (n346,n347,n358);
nand (n347,n348,n355);
or (n348,n349,n353);
and (n349,n286,n350);
wire s0n350,s1n350,notn350;
or (n350,s0n350,s1n350);
not(notn350,n96);
and (s0n350,notn350,n351);
and (s1n350,n96,n352);
wire s0n351,s1n351,notn351;
or (n351,s0n351,s1n351);
not(notn351,n22);
and (s0n351,notn351,1'b0);
and (s1n351,n22,n78);
xor (n352,n77,n79);
and (n353,n285,n354);
not (n354,n350);
nor (n355,n356,n357);
and (n356,n253,n350);
and (n357,n257,n354);
nor (n358,n359,n360);
and (n359,n268,n257);
and (n360,n272,n253);
or (n361,n348,n362);
nor (n362,n363,n367);
and (n363,n364,n257);
wire s0n364,s1n364,notn364;
or (n364,s0n364,s1n364);
not(notn364,n132);
and (s0n364,notn364,n365);
and (s1n364,n132,n366);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n22);
and (s0n365,notn365,1'b0);
and (s1n365,n22,n185);
xor (n366,n184,n186);
and (n367,n368,n253);
not (n368,n364);
nand (n369,n370,n398);
or (n370,n371,n391);
not (n371,n372);
nor (n372,n373,n383);
nand (n373,n374,n382);
or (n374,n375,n379);
not (n375,n376);
wire s0n376,s1n376,notn376;
or (n376,s0n376,s1n376);
not(notn376,n96);
and (s0n376,notn376,n377);
and (s1n376,n96,n378);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n22);
and (s0n377,notn377,1'b0);
and (s1n377,n22,n57);
xor (n378,n56,n58);
wire s0n379,s1n379,notn379;
or (n379,s0n379,s1n379);
not(notn379,n96);
and (s0n379,notn379,n380);
and (s1n379,n96,n381);
wire s0n380,s1n380,notn380;
or (n380,s0n380,s1n380);
not(notn380,n22);
and (s0n380,notn380,1'b0);
and (s1n380,n22,n54);
xor (n381,n53,n55);
nand (n382,n375,n379);
nor (n383,n384,n389);
and (n384,n385,n379);
not (n385,n386);
wire s0n386,s1n386,notn386;
or (n386,s0n386,s1n386);
not(notn386,n96);
and (s0n386,notn386,n387);
and (s1n386,n96,n388);
wire s0n387,s1n387,notn387;
or (n387,s0n387,s1n387);
not(notn387,n22);
and (s0n387,notn387,1'b0);
and (s1n387,n22,n51);
xor (n388,n50,n52);
and (n389,n390,n386);
not (n390,n379);
nor (n391,n392,n396);
and (n392,n385,n393);
wire s0n393,s1n393,notn393;
or (n393,s0n393,s1n393);
not(notn393,n132);
and (s0n393,notn393,n394);
and (s1n393,n132,n395);
wire s0n394,s1n394,notn394;
or (n394,s0n394,s1n394);
not(notn394,n22);
and (s0n394,notn394,1'b0);
and (s1n394,n22,n212);
xor (n395,n211,n213);
and (n396,n397,n386);
not (n397,n393);
or (n398,n399,n400);
not (n399,n373);
nor (n400,n401,n405);
and (n401,n402,n385);
wire s0n402,s1n402,notn402;
or (n402,s0n402,s1n402);
not(notn402,n132);
and (s0n402,notn402,n403);
and (s1n402,n132,n404);
wire s0n403,s1n403,notn403;
or (n403,s0n403,s1n403);
not(notn403,n22);
and (s0n403,notn403,1'b0);
and (s1n403,n22,n209);
xor (n404,n208,n210);
and (n405,n406,n386);
not (n406,n402);
nand (n407,n408,n432);
or (n408,n409,n425);
not (n409,n410);
and (n410,n411,n418);
nor (n411,n412,n417);
and (n412,n386,n413);
not (n413,n414);
wire s0n414,s1n414,notn414;
or (n414,s0n414,s1n414);
not(notn414,n96);
and (s0n414,notn414,n415);
and (s1n414,n96,n416);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n22);
and (s0n415,notn415,1'b0);
and (s1n415,n22,n48);
xor (n416,n47,n49);
and (n417,n385,n414);
nand (n418,n419,n423);
or (n419,n413,n420);
wire s0n420,s1n420,notn420;
or (n420,s0n420,s1n420);
not(notn420,n96);
and (s0n420,notn420,n421);
and (s1n420,n96,n422);
wire s0n421,s1n421,notn421;
or (n421,s0n421,s1n421);
not(notn421,n22);
and (s0n421,notn421,1'b0);
and (s1n421,n22,n45);
xor (n422,n44,n46);
or (n423,n424,n414);
not (n424,n420);
nor (n425,n426,n430);
and (n426,n427,n424);
wire s0n427,s1n427,notn427;
or (n427,s0n427,s1n427);
not(notn427,n132);
and (s0n427,notn427,n428);
and (s1n427,n132,n429);
wire s0n428,s1n428,notn428;
or (n428,s0n428,s1n428);
not(notn428,n22);
and (s0n428,notn428,1'b0);
and (s1n428,n22,n218);
xor (n429,n217,n219);
and (n430,n431,n420);
not (n431,n427);
or (n432,n433,n411);
nor (n433,n434,n438);
and (n434,n435,n424);
wire s0n435,s1n435,notn435;
or (n435,s0n435,s1n435);
not(notn435,n132);
and (s0n435,notn435,n436);
and (s1n435,n132,n437);
wire s0n436,s1n436,notn436;
or (n436,s0n436,s1n436);
not(notn436,n22);
and (s0n436,notn436,1'b0);
and (s1n436,n22,n215);
xor (n437,n214,n216);
and (n438,n439,n420);
not (n439,n435);
and (n440,n345,n369);
or (n441,n442,n473);
and (n442,n443,n463);
xor (n443,n444,n457);
nand (n444,n445,n449);
or (n445,n145,n446);
nor (n446,n447,n448);
and (n447,n159,n301);
and (n448,n305,n160);
or (n449,n450,n146);
nor (n450,n451,n455);
and (n451,n452,n159);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n132);
and (s0n452,notn452,n453);
and (s1n452,n132,n454);
wire s0n453,s1n453,notn453;
or (n453,s0n453,s1n453);
not(notn453,n22);
and (s0n453,notn453,1'b0);
and (s1n453,n22,n173);
xor (n454,n172,n174);
and (n455,n456,n160);
not (n456,n452);
nand (n457,n458,n462);
or (n458,n238,n459);
nor (n459,n460,n461);
and (n460,n249,n333);
and (n461,n244,n337);
or (n462,n258,n250);
nand (n463,n464,n472);
or (n464,n275,n465);
nor (n465,n466,n470);
and (n466,n467,n285);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n132);
and (s0n467,notn467,n468);
and (s1n467,n132,n469);
wire s0n468,s1n468,notn468;
or (n468,s0n468,s1n468);
not(notn468,n22);
and (s0n468,notn468,1'b0);
and (s1n468,n22,n182);
xor (n469,n181,n183);
and (n470,n471,n286);
not (n471,n467);
or (n472,n276,n291);
and (n473,n444,n457);
xor (n474,n235,n306);
and (n475,n342,n441);
xor (n476,n477,n531);
xor (n477,n478,n508);
or (n478,n479,n507);
and (n479,n480,n501);
xor (n480,n481,n482);
nor (n481,n15,n119);
nand (n482,n483,n490);
or (n483,n484,n487);
nor (n484,n485,n486);
and (n485,n225,n148);
and (n486,n232,n149);
nand (n487,n149,n488);
not (n488,n489);
wire s0n489,s1n489,notn489;
or (n489,s0n489,s1n489);
not(notn489,n22);
and (s0n489,notn489,1'b0);
and (s1n489,n22,n95);
or (n490,n491,n488);
nor (n491,n492,n499);
and (n492,n493,n148);
wire s0n493,s1n493,notn493;
or (n493,s0n493,s1n493);
not(notn493,n132);
and (s0n493,notn493,n494);
and (s1n493,n132,n496);
wire s0n494,s1n494,notn494;
or (n494,s0n494,s1n494);
not(notn494,n22);
and (s0n494,notn494,1'b0);
and (s1n494,n22,n495);
xor (n496,n497,n498);
not (n497,n495);
and (n498,n229,n230);
and (n499,n500,n149);
not (n500,n493);
nand (n501,n502,n503);
or (n502,n347,n362);
or (n503,n348,n504);
nor (n504,n505,n506);
and (n505,n467,n257);
and (n506,n471,n253);
and (n507,n481,n482);
or (n508,n509,n530);
and (n509,n510,n527);
xor (n510,n511,n521);
nand (n511,n512,n513);
or (n512,n371,n400);
or (n513,n514,n399);
nor (n514,n515,n519);
and (n515,n385,n516);
wire s0n516,s1n516,notn516;
or (n516,s0n516,s1n516);
not(notn516,n132);
and (s0n516,notn516,n517);
and (s1n516,n132,n518);
wire s0n517,s1n517,notn517;
or (n517,s0n517,s1n517);
not(notn517,n22);
and (s0n517,notn517,1'b0);
and (s1n517,n22,n206);
xor (n518,n205,n207);
and (n519,n386,n520);
not (n520,n516);
nand (n521,n522,n523);
or (n522,n409,n433);
or (n523,n524,n411);
nor (n524,n525,n526);
and (n525,n424,n393);
and (n526,n420,n397);
nand (n527,n528,n529);
or (n528,n145,n450);
or (n529,n146,n164);
and (n530,n511,n521);
xor (n531,n532,n552);
xor (n532,n533,n539);
nand (n533,n534,n535);
or (n534,n238,n266);
or (n535,n536,n250);
nor (n536,n537,n538);
and (n537,n249,n364);
and (n538,n244,n368);
nand (n539,n540,n541);
or (n540,n491,n487);
or (n541,n542,n488);
nor (n542,n543,n550);
and (n543,n544,n148);
wire s0n544,s1n544,notn544;
or (n544,s0n544,s1n544);
not(notn544,n132);
and (s0n544,notn544,n545);
and (s1n544,n132,n547);
wire s0n545,s1n545,notn545;
or (n545,s0n545,s1n545);
not(notn545,n22);
and (s0n545,notn545,1'b0);
and (s1n545,n22,n546);
xor (n547,n548,n549);
not (n548,n546);
and (n549,n497,n498);
and (n550,n551,n149);
not (n551,n544);
nand (n552,n553,n554);
or (n553,n275,n299);
or (n554,n555,n276);
nor (n555,n556,n557);
and (n556,n452,n285);
and (n557,n456,n286);
xor (n558,n559,n697);
xor (n559,n560,n626);
or (n560,n561,n625);
and (n561,n562,n565);
xor (n562,n563,n564);
xor (n563,n480,n501);
xor (n564,n510,n527);
or (n565,n566,n624);
and (n566,n567,n603);
xor (n567,n568,n578);
nand (n568,n569,n577);
or (n569,n308,n570);
nor (n570,n571,n575);
and (n571,n322,n572);
wire s0n572,s1n572,notn572;
or (n572,s0n572,s1n572);
not(notn572,n132);
and (s0n572,notn572,n573);
and (s1n572,n132,n574);
wire s0n573,s1n573,notn573;
or (n573,s0n573,s1n573);
not(notn573,n22);
and (s0n573,notn573,1'b0);
and (s1n573,n22,n200);
xor (n574,n199,n201);
and (n575,n318,n576);
not (n576,n572);
or (n577,n309,n323);
nand (n578,n579,n594);
or (n579,n580,n591);
or (n580,n581,n588);
nor (n581,n582,n586);
and (n582,n375,n583);
wire s0n583,s1n583,notn583;
or (n583,s0n583,s1n583);
not(notn583,n96);
and (s0n583,notn583,n584);
and (s1n583,n96,n585);
wire s0n584,s1n584,notn584;
or (n584,s0n584,s1n584);
not(notn584,n22);
and (s0n584,notn584,1'b0);
and (s1n584,n22,n60);
xor (n585,n59,n61);
and (n586,n587,n376);
not (n587,n583);
nor (n588,n589,n590);
and (n589,n583,n318);
and (n590,n587,n322);
nor (n591,n592,n593);
and (n592,n375,n516);
and (n593,n376,n520);
or (n594,n595,n602);
nor (n595,n596,n600);
and (n596,n375,n597);
wire s0n597,s1n597,notn597;
or (n597,s0n597,s1n597);
not(notn597,n132);
and (s0n597,notn597,n598);
and (s1n597,n132,n599);
wire s0n598,s1n598,notn598;
or (n598,s0n598,s1n598);
not(notn598,n22);
and (s0n598,notn598,1'b0);
and (s1n598,n22,n203);
xor (n599,n202,n204);
and (n600,n376,n601);
not (n601,n597);
not (n602,n588);
nand (n603,n604,n619);
or (n604,n605,n616);
or (n605,n606,n613);
nor (n606,n607,n611);
and (n607,n608,n420);
wire s0n608,s1n608,notn608;
or (n608,s0n608,s1n608);
not(notn608,n96);
and (s0n608,notn608,n609);
and (s1n608,n96,n610);
wire s0n609,s1n609,notn609;
or (n609,s0n609,s1n609);
not(notn609,n22);
and (s0n609,notn609,1'b0);
and (s1n609,n22,n42);
xor (n610,n41,n43);
and (n611,n612,n424);
not (n612,n608);
nor (n613,n614,n615);
and (n614,n608,n17);
and (n615,n612,n18);
nor (n616,n617,n618);
and (n617,n18,n119);
and (n618,n17,n120);
or (n619,n620,n621);
not (n620,n606);
nor (n621,n622,n623);
and (n622,n126,n17);
and (n623,n135,n18);
and (n624,n568,n578);
and (n625,n563,n564);
xor (n626,n627,n674);
xor (n627,n628,n648);
xor (n628,n629,n642);
xor (n629,n630,n636);
nand (n630,n631,n632);
or (n631,n347,n504);
or (n632,n348,n633);
nor (n633,n634,n635);
and (n634,n293,n257);
and (n635,n297,n253);
nand (n636,n637,n638);
or (n637,n371,n514);
or (n638,n639,n399);
nor (n639,n640,n641);
and (n640,n385,n597);
and (n641,n386,n601);
nand (n642,n643,n644);
or (n643,n409,n524);
or (n644,n645,n411);
nor (n645,n646,n647);
and (n646,n424,n402);
and (n647,n420,n406);
xor (n648,n649,n665);
xor (n649,n650,n656);
nand (n650,n651,n652);
or (n651,n308,n331);
or (n652,n309,n653);
nor (n653,n654,n655);
and (n654,n322,n260);
and (n655,n318,n264);
nand (n656,n657,n661);
or (n657,n580,n658);
nor (n658,n659,n660);
and (n659,n375,n572);
and (n660,n376,n576);
or (n661,n602,n662);
nor (n662,n663,n664);
and (n663,n375,n325);
and (n664,n376,n329);
nand (n665,n666,n670);
or (n666,n605,n667);
nor (n667,n668,n669);
and (n668,n427,n17);
and (n669,n431,n18);
or (n670,n620,n671);
nor (n671,n672,n673);
and (n672,n435,n17);
and (n673,n439,n18);
or (n674,n675,n696);
and (n675,n676,n683);
xor (n676,n677,n680);
nand (n677,n678,n679);
or (n678,n580,n595);
or (n679,n602,n658);
nand (n680,n681,n682);
or (n681,n605,n621);
or (n682,n620,n667);
and (n683,n684,n690);
nor (n684,n685,n17);
nor (n685,n686,n689);
and (n686,n687,n424);
not (n687,n688);
and (n688,n120,n608);
and (n689,n612,n119);
nand (n690,n691,n695);
or (n691,n692,n487);
nor (n692,n693,n694);
and (n693,n166,n148);
and (n694,n221,n149);
or (n695,n484,n488);
and (n696,n677,n680);
or (n697,n698,n746);
and (n698,n699,n745);
xor (n699,n700,n701);
xor (n700,n676,n683);
or (n701,n702,n744);
and (n702,n703,n722);
xor (n703,n704,n705);
xor (n704,n684,n690);
or (n705,n706,n721);
and (n706,n707,n715);
xor (n707,n708,n709);
nor (n708,n620,n119);
nand (n709,n710,n714);
or (n710,n711,n487);
nor (n711,n712,n713);
and (n712,n452,n148);
and (n713,n456,n149);
or (n714,n692,n488);
nand (n715,n716,n717);
or (n716,n358,n348);
or (n717,n347,n718);
nor (n718,n719,n720);
and (n719,n260,n257);
and (n720,n264,n253);
and (n721,n708,n709);
or (n722,n723,n743);
and (n723,n724,n737);
xor (n724,n725,n731);
nand (n725,n726,n730);
or (n726,n371,n727);
nor (n727,n728,n729);
and (n728,n435,n385);
and (n729,n439,n386);
or (n730,n391,n399);
nand (n731,n732,n736);
or (n732,n409,n733);
nor (n733,n734,n735);
and (n734,n126,n424);
and (n735,n135,n420);
or (n736,n425,n411);
nand (n737,n738,n742);
or (n738,n145,n739);
nor (n739,n740,n741);
and (n740,n159,n293);
and (n741,n297,n160);
or (n742,n146,n446);
and (n743,n725,n731);
and (n744,n704,n705);
xor (n745,n341,n474);
and (n746,n700,n701);
or (n747,n748,n831);
and (n748,n749,n779);
xor (n749,n750,n778);
or (n750,n751,n777);
and (n751,n752,n776);
xor (n752,n753,n775);
or (n753,n754,n774);
and (n754,n755,n768);
xor (n755,n756,n762);
nand (n756,n757,n761);
or (n757,n238,n758);
nor (n758,n759,n760);
and (n759,n249,n325);
and (n760,n244,n329);
or (n761,n459,n250);
nand (n762,n763,n767);
or (n763,n275,n764);
nor (n764,n765,n766);
and (n765,n364,n285);
and (n766,n368,n286);
or (n767,n276,n465);
nand (n768,n769,n773);
or (n769,n308,n770);
nor (n770,n771,n772);
and (n771,n322,n597);
and (n772,n318,n601);
or (n773,n309,n570);
and (n774,n756,n762);
xor (n775,n443,n463);
xor (n776,n344,n407);
and (n777,n753,n775);
xor (n778,n562,n565);
or (n779,n780,n830);
and (n780,n781,n829);
xor (n781,n782,n783);
xor (n782,n567,n603);
or (n783,n784,n828);
and (n784,n785,n805);
xor (n785,n786,n792);
nand (n786,n787,n791);
or (n787,n580,n788);
nor (n788,n789,n790);
and (n789,n375,n402);
and (n790,n376,n406);
or (n791,n591,n602);
and (n792,n793,n799);
nor (n793,n794,n424);
nor (n794,n795,n798);
and (n795,n385,n796);
not (n796,n797);
and (n797,n120,n414);
and (n798,n413,n119);
nand (n799,n800,n804);
or (n800,n801,n487);
nor (n801,n802,n803);
and (n802,n301,n148);
and (n803,n305,n149);
or (n804,n711,n488);
or (n805,n806,n827);
and (n806,n807,n820);
xor (n807,n808,n814);
nand (n808,n809,n813);
or (n809,n347,n810);
nor (n810,n811,n812);
and (n811,n333,n257);
and (n812,n337,n253);
or (n813,n718,n348);
nand (n814,n815,n819);
or (n815,n371,n816);
nor (n816,n817,n818);
and (n817,n427,n385);
and (n818,n431,n386);
or (n819,n399,n727);
nand (n820,n821,n826);
or (n821,n822,n409);
not (n822,n823);
nand (n823,n824,n825);
or (n824,n424,n120);
or (n825,n420,n119);
or (n826,n733,n411);
and (n827,n808,n814);
and (n828,n786,n792);
xor (n829,n703,n722);
and (n830,n782,n783);
and (n831,n750,n778);
not (n832,n833);
or (n833,n834,n894);
and (n834,n835,n893);
xor (n835,n836,n837);
xor (n836,n699,n745);
or (n837,n838,n892);
and (n838,n839,n869);
xor (n839,n840,n868);
or (n840,n841,n867);
and (n841,n842,n866);
xor (n842,n843,n865);
or (n843,n844,n864);
and (n844,n845,n858);
xor (n845,n846,n852);
nand (n846,n847,n851);
or (n847,n145,n848);
nor (n848,n849,n850);
and (n849,n159,n467);
and (n850,n471,n160);
or (n851,n146,n739);
nand (n852,n853,n857);
or (n853,n238,n854);
nor (n854,n855,n856);
and (n855,n249,n572);
and (n856,n244,n576);
or (n857,n758,n250);
nand (n858,n859,n863);
or (n859,n860,n275);
nor (n860,n861,n862);
and (n861,n268,n285);
and (n862,n272,n286);
or (n863,n276,n764);
and (n864,n846,n852);
xor (n865,n755,n768);
xor (n866,n707,n715);
and (n867,n843,n865);
xor (n868,n752,n776);
or (n869,n870,n891);
and (n870,n871,n890);
xor (n871,n872,n873);
xor (n872,n724,n737);
or (n873,n874,n889);
and (n874,n875,n888);
xor (n875,n876,n882);
nand (n876,n877,n881);
or (n877,n308,n878);
nor (n878,n879,n880);
and (n879,n322,n516);
and (n880,n318,n520);
or (n881,n770,n309);
nand (n882,n883,n887);
or (n883,n580,n884);
nor (n884,n885,n886);
and (n885,n375,n393);
and (n886,n397,n376);
or (n887,n602,n788);
xor (n888,n793,n799);
and (n889,n876,n882);
xor (n890,n785,n805);
and (n891,n872,n873);
and (n892,n840,n868);
xor (n893,n749,n779);
and (n894,n836,n837);
and (n895,n5,n832);
not (n896,n897);
and (n897,n898,n1774);
nand (n898,n899,n1769);
not (n899,n900);
nor (n900,n901,n1758);
nor (n901,n902,n1727);
nand (n902,n903,n1634);
or (n903,n904,n1633);
and (n904,n905,n1223);
xor (n905,n906,n1137);
or (n906,n907,n1136);
and (n907,n908,n1085);
xor (n908,n909,n992);
xor (n909,n910,n961);
xor (n910,n911,n932);
xor (n911,n912,n923);
xor (n912,n913,n914);
nor (n913,n399,n119);
nand (n914,n915,n919);
or (n915,n916,n487);
nor (n916,n917,n918);
and (n917,n148,n364);
and (n918,n368,n149);
or (n919,n920,n488);
nor (n920,n921,n922);
and (n921,n467,n148);
and (n922,n471,n149);
nand (n923,n924,n928);
or (n924,n145,n925);
nor (n925,n926,n927);
and (n926,n159,n260);
and (n927,n264,n160);
or (n928,n146,n929);
nor (n929,n930,n931);
and (n930,n268,n159);
and (n931,n272,n160);
or (n932,n933,n960);
and (n933,n934,n950);
xor (n934,n935,n941);
nand (n935,n936,n940);
or (n936,n145,n937);
nor (n937,n938,n939);
and (n938,n159,n333);
and (n939,n337,n160);
or (n940,n146,n925);
nand (n941,n942,n946);
or (n942,n347,n943);
nor (n943,n944,n945);
and (n944,n516,n257);
and (n945,n520,n253);
or (n946,n348,n947);
nor (n947,n948,n949);
and (n948,n597,n257);
and (n949,n601,n253);
nand (n950,n951,n956);
or (n951,n952,n238);
not (n952,n953);
nand (n953,n954,n955);
or (n954,n244,n397);
or (n955,n249,n393);
or (n956,n957,n250);
nor (n957,n958,n959);
and (n958,n249,n402);
and (n959,n244,n406);
and (n960,n935,n941);
or (n961,n962,n991);
and (n962,n963,n982);
xor (n963,n964,n973);
nand (n964,n965,n969);
or (n965,n275,n966);
nor (n966,n967,n968);
and (n967,n572,n285);
and (n968,n576,n286);
or (n969,n970,n276);
nor (n970,n971,n972);
and (n971,n325,n285);
and (n972,n329,n286);
nand (n973,n974,n978);
or (n974,n308,n975);
nor (n975,n976,n977);
and (n976,n427,n322);
and (n977,n431,n318);
or (n978,n979,n309);
nor (n979,n980,n981);
and (n980,n435,n322);
and (n981,n439,n318);
nand (n982,n983,n987);
or (n983,n602,n984);
nor (n984,n985,n986);
and (n985,n126,n375);
and (n986,n135,n376);
or (n987,n580,n988);
nor (n988,n989,n990);
and (n989,n376,n119);
and (n990,n375,n120);
and (n991,n964,n973);
xor (n992,n993,n1041);
xor (n993,n994,n1021);
xor (n994,n995,n1008);
xor (n995,n996,n1002);
nand (n996,n997,n998);
or (n997,n308,n979);
or (n998,n999,n309);
nor (n999,n1000,n1001);
and (n1000,n322,n393);
and (n1001,n318,n397);
nand (n1002,n1003,n1004);
or (n1003,n580,n984);
or (n1004,n1005,n602);
nor (n1005,n1006,n1007);
and (n1006,n427,n375);
and (n1007,n431,n376);
and (n1008,n1009,n1015);
nand (n1009,n1010,n1014);
or (n1010,n1011,n487);
nor (n1011,n1012,n1013);
and (n1012,n148,n268);
and (n1013,n272,n149);
or (n1014,n916,n488);
nor (n1015,n1016,n375);
nor (n1016,n1017,n1020);
and (n1017,n322,n1018);
not (n1018,n1019);
and (n1019,n120,n583);
and (n1020,n587,n119);
xor (n1021,n1022,n1035);
xor (n1022,n1023,n1029);
nand (n1023,n1024,n1025);
or (n1024,n347,n947);
or (n1025,n1026,n348);
nor (n1026,n1027,n1028);
and (n1027,n572,n257);
and (n1028,n576,n253);
nand (n1029,n1030,n1031);
or (n1030,n238,n957);
or (n1031,n1032,n250);
nor (n1032,n1033,n1034);
and (n1033,n249,n516);
and (n1034,n244,n520);
nand (n1035,n1036,n1040);
or (n1036,n276,n1037);
nor (n1037,n1038,n1039);
and (n1038,n333,n285);
and (n1039,n337,n286);
or (n1040,n275,n970);
or (n1041,n1042,n1084);
and (n1042,n1043,n1062);
xor (n1043,n1044,n1045);
xor (n1044,n1009,n1015);
or (n1045,n1046,n1061);
and (n1046,n1047,n1055);
xor (n1047,n1048,n1049);
nor (n1048,n602,n119);
nand (n1049,n1050,n1054);
or (n1050,n1051,n487);
nor (n1051,n1052,n1053);
and (n1052,n148,n260);
and (n1053,n264,n149);
or (n1054,n1011,n488);
nand (n1055,n1056,n1057);
or (n1056,n146,n937);
or (n1057,n145,n1058);
nor (n1058,n1059,n1060);
and (n1059,n325,n159);
and (n1060,n329,n160);
and (n1061,n1048,n1049);
or (n1062,n1063,n1083);
and (n1063,n1064,n1077);
xor (n1064,n1065,n1071);
nand (n1065,n1066,n1070);
or (n1066,n347,n1067);
nor (n1067,n1068,n1069);
and (n1068,n402,n257);
and (n1069,n406,n253);
or (n1070,n943,n348);
nand (n1071,n1072,n1073);
or (n1072,n250,n952);
or (n1073,n238,n1074);
nor (n1074,n1075,n1076);
and (n1075,n249,n435);
and (n1076,n244,n439);
nand (n1077,n1078,n1079);
or (n1078,n309,n975);
or (n1079,n308,n1080);
nor (n1080,n1081,n1082);
and (n1081,n126,n322);
and (n1082,n135,n318);
and (n1083,n1065,n1071);
and (n1084,n1044,n1045);
or (n1085,n1086,n1135);
and (n1086,n1087,n1090);
xor (n1087,n1088,n1089);
xor (n1088,n963,n982);
xor (n1089,n934,n950);
or (n1090,n1091,n1134);
and (n1091,n1092,n1112);
xor (n1092,n1093,n1099);
nand (n1093,n1094,n1098);
or (n1094,n275,n1095);
nor (n1095,n1096,n1097);
and (n1096,n597,n285);
and (n1097,n601,n286);
or (n1098,n276,n966);
and (n1099,n1100,n1106);
nand (n1100,n1101,n1105);
or (n1101,n1102,n487);
nor (n1102,n1103,n1104);
and (n1103,n333,n148);
and (n1104,n337,n149);
or (n1105,n1051,n488);
nor (n1106,n1107,n322);
nor (n1107,n1108,n1111);
and (n1108,n249,n1109);
not (n1109,n1110);
and (n1110,n120,n311);
and (n1111,n315,n119);
or (n1112,n1113,n1133);
and (n1113,n1114,n1127);
xor (n1114,n1115,n1121);
nand (n1115,n1116,n1120);
or (n1116,n145,n1117);
nor (n1117,n1118,n1119);
and (n1118,n572,n159);
and (n1119,n576,n160);
or (n1120,n146,n1058);
nand (n1121,n1122,n1126);
or (n1122,n347,n1123);
nor (n1123,n1124,n1125);
and (n1124,n393,n257);
and (n1125,n397,n253);
or (n1126,n1067,n348);
nand (n1127,n1128,n1132);
or (n1128,n238,n1129);
nor (n1129,n1130,n1131);
and (n1130,n427,n249);
and (n1131,n431,n244);
or (n1132,n1074,n250);
and (n1133,n1115,n1121);
and (n1134,n1093,n1099);
and (n1135,n1088,n1089);
and (n1136,n909,n992);
xor (n1137,n1138,n1171);
xor (n1138,n1139,n1168);
xor (n1139,n1140,n1147);
xor (n1140,n1141,n1144);
or (n1141,n1142,n1143);
and (n1142,n1022,n1035);
and (n1143,n1023,n1029);
or (n1144,n1145,n1146);
and (n1145,n995,n1008);
and (n1146,n996,n1002);
xor (n1147,n1148,n1161);
xor (n1148,n1149,n1155);
nand (n1149,n1150,n1151);
or (n1150,n238,n1032);
or (n1151,n1152,n250);
nor (n1152,n1153,n1154);
and (n1153,n249,n597);
and (n1154,n244,n601);
nand (n1155,n1156,n1157);
or (n1156,n275,n1037);
or (n1157,n276,n1158);
nor (n1158,n1159,n1160);
and (n1159,n260,n285);
and (n1160,n264,n286);
nand (n1161,n1162,n1167);
or (n1162,n309,n1163);
not (n1163,n1164);
nand (n1164,n1165,n1166);
or (n1165,n406,n318);
or (n1166,n322,n402);
or (n1167,n308,n999);
or (n1168,n1169,n1170);
and (n1169,n993,n1041);
and (n1170,n994,n1021);
xor (n1171,n1172,n1199);
xor (n1172,n1173,n1196);
xor (n1173,n1174,n1190);
xor (n1174,n1175,n1181);
nand (n1175,n1176,n1177);
or (n1176,n145,n929);
or (n1177,n146,n1178);
nor (n1178,n1179,n1180);
and (n1179,n159,n364);
and (n1180,n368,n160);
nand (n1181,n1182,n1186);
or (n1182,n371,n1183);
nor (n1183,n1184,n1185);
and (n1184,n386,n119);
and (n1185,n385,n120);
or (n1186,n1187,n399);
nor (n1187,n1188,n1189);
and (n1188,n126,n385);
and (n1189,n135,n386);
nand (n1190,n1191,n1195);
or (n1191,n1192,n348);
nor (n1192,n1193,n1194);
and (n1193,n325,n257);
and (n1194,n329,n253);
or (n1195,n347,n1026);
or (n1196,n1197,n1198);
and (n1197,n910,n961);
and (n1198,n911,n932);
xor (n1199,n1200,n1220);
xor (n1200,n1201,n1207);
nand (n1201,n1202,n1203);
or (n1202,n580,n1005);
or (n1203,n1204,n602);
nor (n1204,n1205,n1206);
and (n1205,n435,n375);
and (n1206,n439,n376);
xor (n1207,n1208,n1214);
nand (n1208,n1209,n1210);
or (n1209,n920,n487);
or (n1210,n1211,n488);
nor (n1211,n1212,n1213);
and (n1212,n293,n148);
and (n1213,n297,n149);
nor (n1214,n1215,n385);
nor (n1215,n1216,n1219);
and (n1216,n375,n1217);
not (n1217,n1218);
and (n1218,n120,n379);
and (n1219,n390,n119);
or (n1220,n1221,n1222);
and (n1221,n912,n923);
and (n1222,n913,n914);
or (n1223,n1224,n1632);
and (n1224,n1225,n1256);
xor (n1225,n1226,n1255);
or (n1226,n1227,n1254);
and (n1227,n1228,n1253);
xor (n1228,n1229,n1252);
or (n1229,n1230,n1251);
and (n1230,n1231,n1234);
xor (n1231,n1232,n1233);
xor (n1232,n1047,n1055);
xor (n1233,n1064,n1077);
or (n1234,n1235,n1250);
and (n1235,n1236,n1249);
xor (n1236,n1237,n1243);
nand (n1237,n1238,n1242);
or (n1238,n308,n1239);
nor (n1239,n1240,n1241);
and (n1240,n318,n119);
and (n1241,n322,n120);
or (n1242,n1080,n309);
nand (n1243,n1244,n1248);
or (n1244,n275,n1245);
nor (n1245,n1246,n1247);
and (n1246,n516,n285);
and (n1247,n520,n286);
or (n1248,n1095,n276);
xor (n1249,n1100,n1106);
and (n1250,n1237,n1243);
and (n1251,n1232,n1233);
xor (n1252,n1043,n1062);
xor (n1253,n1087,n1090);
and (n1254,n1229,n1252);
xor (n1255,n908,n1085);
nand (n1256,n1257,n1629,n1631);
or (n1257,n1258,n1624);
nand (n1258,n1259,n1613);
or (n1259,n1260,n1612);
and (n1260,n1261,n1382);
xor (n1261,n1262,n1367);
or (n1262,n1263,n1366);
and (n1263,n1264,n1332);
xor (n1264,n1265,n1287);
xor (n1265,n1266,n1281);
xor (n1266,n1267,n1274);
nand (n1267,n1268,n1273);
or (n1268,n347,n1269);
not (n1269,n1270);
nor (n1270,n1271,n1272);
and (n1271,n257,n439);
and (n1272,n435,n253);
or (n1273,n1123,n348);
nand (n1274,n1275,n1280);
or (n1275,n1276,n238);
not (n1276,n1277);
nand (n1277,n1278,n1279);
or (n1278,n135,n244);
or (n1279,n126,n249);
or (n1280,n1129,n250);
nand (n1281,n1282,n1286);
or (n1282,n275,n1283);
nor (n1283,n1284,n1285);
and (n1284,n402,n285);
and (n1285,n406,n286);
or (n1286,n276,n1245);
or (n1287,n1288,n1331);
and (n1288,n1289,n1311);
xor (n1289,n1290,n1296);
nand (n1290,n1291,n1295);
or (n1291,n275,n1292);
nor (n1292,n1293,n1294);
and (n1293,n393,n285);
and (n1294,n397,n286);
or (n1295,n1283,n276);
xor (n1296,n1297,n1303);
nor (n1297,n1298,n249);
nor (n1298,n1299,n1302);
and (n1299,n1300,n257);
not (n1300,n1301);
and (n1301,n120,n241);
and (n1302,n248,n119);
nand (n1303,n1304,n1307);
or (n1304,n487,n1305);
not (n1305,n1306);
xnor (n1306,n572,n148);
or (n1307,n1308,n488);
nor (n1308,n1309,n1310);
and (n1309,n148,n325);
and (n1310,n329,n149);
or (n1311,n1312,n1330);
and (n1312,n1313,n1321);
xor (n1313,n1314,n1315);
nor (n1314,n250,n119);
nand (n1315,n1316,n1317);
or (n1316,n488,n1305);
or (n1317,n1318,n487);
nor (n1318,n1319,n1320);
and (n1319,n148,n597);
and (n1320,n601,n149);
nand (n1321,n1322,n1326);
or (n1322,n347,n1323);
nor (n1323,n1324,n1325);
and (n1324,n126,n257);
and (n1325,n135,n253);
or (n1326,n1327,n348);
nor (n1327,n1328,n1329);
and (n1328,n427,n257);
and (n1329,n431,n253);
and (n1330,n1314,n1315);
and (n1331,n1290,n1296);
xor (n1332,n1333,n1347);
xor (n1333,n1334,n1335);
and (n1334,n1297,n1303);
xor (n1335,n1336,n1341);
xor (n1336,n1337,n1338);
nor (n1337,n309,n119);
nand (n1338,n1339,n1340);
or (n1339,n1308,n487);
or (n1340,n1102,n488);
nand (n1341,n1342,n1346);
or (n1342,n145,n1343);
nor (n1343,n1344,n1345);
and (n1344,n597,n159);
and (n1345,n601,n160);
or (n1346,n146,n1117);
or (n1347,n1348,n1365);
and (n1348,n1349,n1359);
xor (n1349,n1350,n1356);
nand (n1350,n1351,n1355);
or (n1351,n145,n1352);
nor (n1352,n1353,n1354);
and (n1353,n159,n516);
and (n1354,n520,n160);
or (n1355,n1343,n146);
nand (n1356,n1357,n1358);
or (n1357,n348,n1269);
or (n1358,n1327,n347);
nand (n1359,n1360,n1361);
or (n1360,n250,n1276);
or (n1361,n238,n1362);
nor (n1362,n1363,n1364);
and (n1363,n244,n119);
and (n1364,n249,n120);
and (n1365,n1350,n1356);
and (n1366,n1265,n1287);
xor (n1367,n1368,n1373);
xor (n1368,n1369,n1370);
xor (n1369,n1114,n1127);
or (n1370,n1371,n1372);
and (n1371,n1333,n1347);
and (n1372,n1334,n1335);
xor (n1373,n1374,n1381);
xor (n1374,n1375,n1378);
or (n1375,n1376,n1377);
and (n1376,n1336,n1341);
and (n1377,n1337,n1338);
or (n1378,n1379,n1380);
and (n1379,n1266,n1281);
and (n1380,n1267,n1274);
xor (n1381,n1236,n1249);
or (n1382,n1383,n1611);
and (n1383,n1384,n1421);
xor (n1384,n1385,n1420);
or (n1385,n1386,n1419);
and (n1386,n1387,n1418);
xor (n1387,n1388,n1417);
or (n1388,n1389,n1416);
and (n1389,n1390,n1403);
xor (n1390,n1391,n1397);
nand (n1391,n1392,n1396);
or (n1392,n145,n1393);
nor (n1393,n1394,n1395);
and (n1394,n402,n159);
and (n1395,n160,n406);
or (n1396,n1352,n146);
nand (n1397,n1398,n1402);
or (n1398,n275,n1399);
nor (n1399,n1400,n1401);
and (n1400,n435,n285);
and (n1401,n439,n286);
or (n1402,n1292,n276);
and (n1403,n1404,n1410);
nor (n1404,n1405,n257);
nor (n1405,n1406,n1409);
and (n1406,n1407,n285);
not (n1407,n1408);
and (n1408,n120,n350);
and (n1409,n354,n119);
nand (n1410,n1411,n1415);
or (n1411,n1412,n487);
nor (n1412,n1413,n1414);
and (n1413,n148,n516);
and (n1414,n520,n149);
or (n1415,n1318,n488);
and (n1416,n1391,n1397);
xor (n1417,n1349,n1359);
xor (n1418,n1289,n1311);
and (n1419,n1388,n1417);
xor (n1420,n1264,n1332);
nand (n1421,n1422,n1608,n1610);
or (n1422,n1423,n1481);
nand (n1423,n1424,n1476);
not (n1424,n1425);
nor (n1425,n1426,n1452);
xor (n1426,n1427,n1451);
xor (n1427,n1428,n1450);
or (n1428,n1429,n1449);
and (n1429,n1430,n1443);
xor (n1430,n1431,n1437);
nand (n1431,n1432,n1436);
or (n1432,n347,n1433);
nor (n1433,n1434,n1435);
and (n1434,n253,n119);
and (n1435,n257,n120);
or (n1436,n1323,n348);
nand (n1437,n1438,n1442);
or (n1438,n1439,n145);
nor (n1439,n1440,n1441);
and (n1440,n160,n397);
and (n1441,n159,n393);
or (n1442,n1393,n146);
nand (n1443,n1444,n1448);
or (n1444,n275,n1445);
nor (n1445,n1446,n1447);
and (n1446,n427,n285);
and (n1447,n431,n286);
or (n1448,n1399,n276);
and (n1449,n1431,n1437);
xor (n1450,n1313,n1321);
xor (n1451,n1390,n1403);
or (n1452,n1453,n1475);
and (n1453,n1454,n1474);
xor (n1454,n1455,n1456);
xor (n1455,n1404,n1410);
or (n1456,n1457,n1473);
and (n1457,n1458,n1467);
xor (n1458,n1459,n1460);
nor (n1459,n348,n119);
nand (n1460,n1461,n1466);
or (n1461,n1462,n487);
not (n1462,n1463);
nand (n1463,n1464,n1465);
or (n1464,n149,n406);
nand (n1465,n406,n149);
or (n1466,n1412,n488);
nand (n1467,n1468,n1472);
or (n1468,n145,n1469);
nor (n1469,n1470,n1471);
and (n1470,n159,n435);
and (n1471,n160,n439);
or (n1472,n1439,n146);
and (n1473,n1459,n1460);
xor (n1474,n1430,n1443);
and (n1475,n1455,n1456);
or (n1476,n1477,n1478);
xor (n1477,n1387,n1418);
or (n1478,n1479,n1480);
and (n1479,n1427,n1451);
and (n1480,n1428,n1450);
nor (n1481,n1482,n1607);
and (n1482,n1483,n1602);
or (n1483,n1484,n1601);
and (n1484,n1485,n1526);
xor (n1485,n1486,n1519);
or (n1486,n1487,n1518);
and (n1487,n1488,n1504);
xor (n1488,n1489,n1495);
nand (n1489,n1490,n1494);
or (n1490,n145,n1491);
nor (n1491,n1492,n1493);
and (n1492,n160,n431);
and (n1493,n159,n427);
or (n1494,n1469,n146);
or (n1495,n1496,n1500);
nor (n1496,n1497,n276);
nor (n1497,n1498,n1499);
and (n1498,n285,n126);
and (n1499,n286,n135);
nor (n1500,n275,n1501);
nor (n1501,n1502,n1503);
and (n1502,n286,n119);
and (n1503,n285,n120);
xor (n1504,n1505,n1511);
nor (n1505,n1506,n285);
nor (n1506,n1507,n1510);
and (n1507,n1508,n159);
not (n1508,n1509);
and (n1509,n120,n279);
and (n1510,n289,n119);
nand (n1511,n1512,n1517);
or (n1512,n487,n1513);
not (n1513,n1514);
nand (n1514,n1515,n1516);
or (n1515,n148,n393);
nand (n1516,n393,n148);
nand (n1517,n1463,n489);
and (n1518,n1489,n1495);
xor (n1519,n1520,n1525);
xor (n1520,n1521,n1524);
nand (n1521,n1522,n1523);
or (n1522,n275,n1497);
or (n1523,n1445,n276);
and (n1524,n1505,n1511);
xor (n1525,n1458,n1467);
or (n1526,n1527,n1600);
and (n1527,n1528,n1548);
xor (n1528,n1529,n1547);
or (n1529,n1530,n1546);
and (n1530,n1531,n1540);
xor (n1531,n1532,n1533);
and (n1532,n277,n120);
nand (n1533,n1534,n1539);
or (n1534,n487,n1535);
not (n1535,n1536);
nand (n1536,n1537,n1538);
or (n1537,n149,n439);
nand (n1538,n439,n149);
nand (n1539,n1514,n489);
nand (n1540,n1541,n1545);
or (n1541,n145,n1542);
nor (n1542,n1543,n1544);
and (n1543,n159,n126);
and (n1544,n160,n135);
or (n1545,n1491,n146);
and (n1546,n1532,n1533);
xor (n1547,n1488,n1504);
or (n1548,n1549,n1599);
and (n1549,n1550,n1567);
xor (n1550,n1551,n1566);
and (n1551,n1552,n1558);
and (n1552,n1553,n160);
nand (n1553,n1554,n1557);
nand (n1554,n1555,n148);
not (n1555,n1556);
and (n1556,n120,n152);
nand (n1557,n156,n119);
nand (n1558,n1559,n1560);
or (n1559,n488,n1535);
nand (n1560,n1561,n1565);
not (n1561,n1562);
nor (n1562,n1563,n1564);
and (n1563,n431,n149);
and (n1564,n427,n148);
not (n1565,n487);
xor (n1566,n1531,n1540);
or (n1567,n1568,n1598);
and (n1568,n1569,n1577);
xor (n1569,n1570,n1576);
nand (n1570,n1571,n1575);
or (n1571,n145,n1572);
nor (n1572,n1573,n1574);
and (n1573,n160,n119);
and (n1574,n159,n120);
or (n1575,n1542,n146);
xor (n1576,n1552,n1558);
or (n1577,n1578,n1597);
and (n1578,n1579,n1587);
xor (n1579,n1580,n1581);
nor (n1580,n146,n119);
nand (n1581,n1582,n1586);
or (n1582,n1583,n487);
or (n1583,n1584,n1585);
and (n1584,n148,n135);
and (n1585,n126,n149);
or (n1586,n1562,n488);
nor (n1587,n1588,n1595);
nor (n1588,n1589,n1591);
and (n1589,n1590,n489);
not (n1590,n1583);
and (n1591,n1592,n1565);
nand (n1592,n1593,n1594);
or (n1593,n148,n120);
or (n1594,n149,n119);
or (n1595,n148,n1596);
and (n1596,n120,n489);
and (n1597,n1580,n1581);
and (n1598,n1570,n1576);
and (n1599,n1551,n1566);
and (n1600,n1529,n1547);
and (n1601,n1486,n1519);
or (n1602,n1603,n1604);
xor (n1603,n1454,n1474);
or (n1604,n1605,n1606);
and (n1605,n1520,n1525);
and (n1606,n1521,n1524);
and (n1607,n1603,n1604);
nand (n1608,n1476,n1609);
and (n1609,n1426,n1452);
nand (n1610,n1477,n1478);
and (n1611,n1385,n1420);
and (n1612,n1262,n1367);
or (n1613,n1614,n1621);
xor (n1614,n1615,n1620);
xor (n1615,n1616,n1617);
xor (n1616,n1092,n1112);
or (n1617,n1618,n1619);
and (n1618,n1374,n1381);
and (n1619,n1375,n1378);
xor (n1620,n1231,n1234);
or (n1621,n1622,n1623);
and (n1622,n1368,n1373);
and (n1623,n1369,n1370);
nor (n1624,n1625,n1626);
xor (n1625,n1228,n1253);
or (n1626,n1627,n1628);
and (n1627,n1615,n1620);
and (n1628,n1616,n1617);
or (n1629,n1624,n1630);
nand (n1630,n1614,n1621);
nand (n1631,n1625,n1626);
and (n1632,n1226,n1255);
and (n1633,n906,n1137);
nor (n1634,n1635,n1722);
nor (n1635,n1636,n1713);
xor (n1636,n1637,n1668);
xor (n1637,n1638,n1643);
xor (n1638,n1639,n1642);
xor (n1639,n1640,n1641);
xor (n1640,n807,n820);
xor (n1641,n845,n858);
xor (n1642,n875,n888);
or (n1643,n1644,n1667);
and (n1644,n1645,n1652);
xor (n1645,n1646,n1649);
or (n1646,n1647,n1648);
and (n1647,n1200,n1220);
and (n1648,n1201,n1207);
or (n1649,n1650,n1651);
and (n1650,n1140,n1147);
and (n1651,n1141,n1144);
xor (n1652,n1653,n1664);
xor (n1653,n1654,n1655);
and (n1654,n1208,n1214);
xor (n1655,n1656,n1661);
xor (n1656,n1657,n1658);
nor (n1657,n411,n119);
nand (n1658,n1659,n1660);
or (n1659,n1211,n487);
or (n1660,n801,n488);
nand (n1661,n1662,n1663);
or (n1662,n145,n1178);
or (n1663,n146,n848);
or (n1664,n1665,n1666);
and (n1665,n1174,n1190);
and (n1666,n1175,n1181);
and (n1667,n1646,n1649);
xor (n1668,n1669,n1704);
xor (n1669,n1670,n1673);
or (n1670,n1671,n1672);
and (n1671,n1653,n1664);
and (n1672,n1654,n1655);
xor (n1673,n1674,n1691);
xor (n1674,n1675,n1678);
or (n1675,n1676,n1677);
and (n1676,n1656,n1661);
and (n1677,n1657,n1658);
or (n1678,n1679,n1690);
and (n1679,n1680,n1687);
xor (n1680,n1681,n1684);
nand (n1681,n1682,n1683);
or (n1682,n275,n1158);
or (n1683,n276,n860);
nand (n1684,n1685,n1686);
or (n1685,n1163,n308);
or (n1686,n878,n309);
nand (n1687,n1688,n1689);
or (n1688,n580,n1204);
or (n1689,n884,n602);
and (n1690,n1681,n1684);
or (n1691,n1692,n1703);
and (n1692,n1693,n1700);
xor (n1693,n1694,n1697);
nand (n1694,n1695,n1696);
or (n1695,n371,n1187);
or (n1696,n816,n399);
nand (n1697,n1698,n1699);
or (n1698,n347,n1192);
or (n1699,n810,n348);
nand (n1700,n1701,n1702);
or (n1701,n238,n1152);
or (n1702,n854,n250);
and (n1703,n1694,n1697);
or (n1704,n1705,n1712);
and (n1705,n1706,n1711);
xor (n1706,n1707,n1710);
or (n1707,n1708,n1709);
and (n1708,n1148,n1161);
and (n1709,n1149,n1155);
xor (n1710,n1680,n1687);
xor (n1711,n1693,n1700);
and (n1712,n1707,n1710);
or (n1713,n1714,n1721);
and (n1714,n1715,n1720);
xor (n1715,n1716,n1717);
xor (n1716,n1706,n1711);
or (n1717,n1718,n1719);
and (n1718,n1172,n1199);
and (n1719,n1173,n1196);
xor (n1720,n1645,n1652);
and (n1721,n1716,n1717);
nor (n1722,n1723,n1724);
xor (n1723,n1715,n1720);
or (n1724,n1725,n1726);
and (n1725,n1138,n1171);
and (n1726,n1139,n1168);
or (n1727,n1728,n1753);
nor (n1728,n1729,n1744);
xor (n1729,n1730,n1743);
xor (n1730,n1731,n1732);
xor (n1731,n781,n829);
or (n1732,n1733,n1742);
and (n1733,n1734,n1741);
xor (n1734,n1735,n1738);
or (n1735,n1736,n1737);
and (n1736,n1674,n1691);
and (n1737,n1675,n1678);
or (n1738,n1739,n1740);
and (n1739,n1639,n1642);
and (n1740,n1640,n1641);
xor (n1741,n842,n866);
and (n1742,n1735,n1738);
xor (n1743,n839,n869);
or (n1744,n1745,n1752);
and (n1745,n1746,n1751);
xor (n1746,n1747,n1748);
xor (n1747,n871,n890);
or (n1748,n1749,n1750);
and (n1749,n1669,n1704);
and (n1750,n1670,n1673);
xor (n1751,n1734,n1741);
and (n1752,n1747,n1748);
nor (n1753,n1754,n1757);
or (n1754,n1755,n1756);
and (n1755,n1637,n1668);
and (n1756,n1638,n1643);
xor (n1757,n1746,n1751);
nand (n1758,n1759,n1768);
or (n1759,n1760,n1728);
nor (n1760,n1761,n1767);
and (n1761,n1762,n1766);
nand (n1762,n1763,n1765);
or (n1763,n1635,n1764);
nand (n1764,n1723,n1724);
nand (n1765,n1636,n1713);
not (n1766,n1753);
and (n1767,n1754,n1757);
nand (n1768,n1729,n1744);
or (n1769,n1770,n1771);
xor (n1770,n835,n893);
or (n1771,n1772,n1773);
and (n1772,n1730,n1743);
and (n1773,n1731,n1732);
nand (n1774,n1770,n1771);
or (n1775,n897,n3);
xor (n1776,n1777,n3026);
xor (n1777,n1778,n3024);
xor (n1778,n1779,n3023);
xor (n1779,n1780,n3014);
xor (n1780,n1781,n3013);
xor (n1781,n1782,n2999);
xor (n1782,n1783,n2998);
xor (n1783,n1784,n2977);
xor (n1784,n1785,n2976);
xor (n1785,n1786,n2950);
xor (n1786,n1787,n2949);
xor (n1787,n1788,n2916);
xor (n1788,n1789,n2915);
xor (n1789,n1790,n2877);
xor (n1790,n1791,n2876);
xor (n1791,n1792,n2831);
xor (n1792,n1793,n2830);
xor (n1793,n1794,n2780);
xor (n1794,n1795,n2779);
xor (n1795,n1796,n2722);
xor (n1796,n1797,n2721);
xor (n1797,n1798,n2659);
xor (n1798,n1799,n2658);
xor (n1799,n1800,n2589);
xor (n1800,n1801,n2588);
xor (n1801,n1802,n2514);
xor (n1802,n1803,n2513);
xor (n1803,n1804,n2433);
xor (n1804,n1805,n2432);
xor (n1805,n1806,n2346);
xor (n1806,n1807,n2345);
xor (n1807,n1808,n2252);
xor (n1808,n1809,n2251);
xor (n1809,n1810,n2153);
xor (n1810,n1811,n2152);
xor (n1811,n1812,n2047);
xor (n1812,n1813,n2046);
xor (n1813,n1814,n1936);
xor (n1814,n1815,n1935);
xor (n1815,n1816,n1819);
xor (n1816,n1817,n1818);
and (n1817,n544,n489);
and (n1818,n493,n149);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
and (n1821,n493,n489);
and (n1822,n225,n149);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
and (n1827,n225,n489);
and (n1828,n166,n149);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
or (n1831,n1832,n1835);
and (n1832,n1833,n1834);
and (n1833,n166,n489);
and (n1834,n452,n149);
and (n1835,n1836,n1837);
xor (n1836,n1833,n1834);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
and (n1839,n452,n489);
and (n1840,n301,n149);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
or (n1843,n1844,n1847);
and (n1844,n1845,n1846);
and (n1845,n301,n489);
and (n1846,n293,n149);
and (n1847,n1848,n1849);
xor (n1848,n1845,n1846);
or (n1849,n1850,n1853);
and (n1850,n1851,n1852);
and (n1851,n293,n489);
and (n1852,n467,n149);
and (n1853,n1854,n1855);
xor (n1854,n1851,n1852);
or (n1855,n1856,n1859);
and (n1856,n1857,n1858);
and (n1857,n467,n489);
and (n1858,n364,n149);
and (n1859,n1860,n1861);
xor (n1860,n1857,n1858);
or (n1861,n1862,n1865);
and (n1862,n1863,n1864);
and (n1863,n364,n489);
and (n1864,n268,n149);
and (n1865,n1866,n1867);
xor (n1866,n1863,n1864);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
and (n1869,n268,n489);
and (n1870,n260,n149);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
or (n1873,n1874,n1877);
and (n1874,n1875,n1876);
and (n1875,n260,n489);
and (n1876,n333,n149);
and (n1877,n1878,n1879);
xor (n1878,n1875,n1876);
or (n1879,n1880,n1883);
and (n1880,n1881,n1882);
and (n1881,n333,n489);
and (n1882,n325,n149);
and (n1883,n1884,n1885);
xor (n1884,n1881,n1882);
or (n1885,n1886,n1889);
and (n1886,n1887,n1888);
and (n1887,n325,n489);
and (n1888,n572,n149);
and (n1889,n1890,n1891);
xor (n1890,n1887,n1888);
or (n1891,n1892,n1895);
and (n1892,n1893,n1894);
and (n1893,n572,n489);
and (n1894,n597,n149);
and (n1895,n1896,n1897);
xor (n1896,n1893,n1894);
or (n1897,n1898,n1901);
and (n1898,n1899,n1900);
and (n1899,n597,n489);
and (n1900,n516,n149);
and (n1901,n1902,n1903);
xor (n1902,n1899,n1900);
or (n1903,n1904,n1907);
and (n1904,n1905,n1906);
and (n1905,n516,n489);
and (n1906,n402,n149);
and (n1907,n1908,n1909);
xor (n1908,n1905,n1906);
or (n1909,n1910,n1913);
and (n1910,n1911,n1912);
and (n1911,n402,n489);
and (n1912,n393,n149);
and (n1913,n1914,n1915);
xor (n1914,n1911,n1912);
or (n1915,n1916,n1919);
and (n1916,n1917,n1918);
and (n1917,n393,n489);
and (n1918,n435,n149);
and (n1919,n1920,n1921);
xor (n1920,n1917,n1918);
or (n1921,n1922,n1925);
and (n1922,n1923,n1924);
and (n1923,n435,n489);
and (n1924,n427,n149);
and (n1925,n1926,n1927);
xor (n1926,n1923,n1924);
or (n1927,n1928,n1930);
and (n1928,n1929,n1585);
and (n1929,n427,n489);
and (n1930,n1931,n1932);
xor (n1931,n1929,n1585);
and (n1932,n1933,n1934);
and (n1933,n126,n489);
and (n1934,n120,n149);
and (n1935,n225,n152);
or (n1936,n1937,n1940);
and (n1937,n1938,n1939);
xor (n1938,n1824,n1825);
and (n1939,n166,n152);
and (n1940,n1941,n1942);
xor (n1941,n1938,n1939);
or (n1942,n1943,n1946);
and (n1943,n1944,n1945);
xor (n1944,n1830,n1831);
and (n1945,n452,n152);
and (n1946,n1947,n1948);
xor (n1947,n1944,n1945);
or (n1948,n1949,n1952);
and (n1949,n1950,n1951);
xor (n1950,n1836,n1837);
and (n1951,n301,n152);
and (n1952,n1953,n1954);
xor (n1953,n1950,n1951);
or (n1954,n1955,n1958);
and (n1955,n1956,n1957);
xor (n1956,n1842,n1843);
and (n1957,n293,n152);
and (n1958,n1959,n1960);
xor (n1959,n1956,n1957);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
xor (n1962,n1848,n1849);
and (n1963,n467,n152);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
xor (n1968,n1854,n1855);
and (n1969,n364,n152);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
xor (n1974,n1860,n1861);
and (n1975,n268,n152);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
xor (n1980,n1866,n1867);
and (n1981,n260,n152);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
xor (n1986,n1872,n1873);
and (n1987,n333,n152);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
or (n1990,n1991,n1994);
and (n1991,n1992,n1993);
xor (n1992,n1878,n1879);
and (n1993,n325,n152);
and (n1994,n1995,n1996);
xor (n1995,n1992,n1993);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
xor (n1998,n1884,n1885);
and (n1999,n572,n152);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2006);
and (n2003,n2004,n2005);
xor (n2004,n1890,n1891);
and (n2005,n597,n152);
and (n2006,n2007,n2008);
xor (n2007,n2004,n2005);
or (n2008,n2009,n2012);
and (n2009,n2010,n2011);
xor (n2010,n1896,n1897);
and (n2011,n516,n152);
and (n2012,n2013,n2014);
xor (n2013,n2010,n2011);
or (n2014,n2015,n2018);
and (n2015,n2016,n2017);
xor (n2016,n1902,n1903);
and (n2017,n402,n152);
and (n2018,n2019,n2020);
xor (n2019,n2016,n2017);
or (n2020,n2021,n2024);
and (n2021,n2022,n2023);
xor (n2022,n1908,n1909);
and (n2023,n393,n152);
and (n2024,n2025,n2026);
xor (n2025,n2022,n2023);
or (n2026,n2027,n2030);
and (n2027,n2028,n2029);
xor (n2028,n1914,n1915);
and (n2029,n435,n152);
and (n2030,n2031,n2032);
xor (n2031,n2028,n2029);
or (n2032,n2033,n2036);
and (n2033,n2034,n2035);
xor (n2034,n1920,n1921);
and (n2035,n427,n152);
and (n2036,n2037,n2038);
xor (n2037,n2034,n2035);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
xor (n2040,n1926,n1927);
and (n2041,n126,n152);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
and (n2044,n2045,n1556);
xor (n2045,n1931,n1932);
and (n2046,n166,n160);
or (n2047,n2048,n2051);
and (n2048,n2049,n2050);
xor (n2049,n1941,n1942);
and (n2050,n452,n160);
and (n2051,n2052,n2053);
xor (n2052,n2049,n2050);
or (n2053,n2054,n2057);
and (n2054,n2055,n2056);
xor (n2055,n1947,n1948);
and (n2056,n301,n160);
and (n2057,n2058,n2059);
xor (n2058,n2055,n2056);
or (n2059,n2060,n2063);
and (n2060,n2061,n2062);
xor (n2061,n1953,n1954);
and (n2062,n293,n160);
and (n2063,n2064,n2065);
xor (n2064,n2061,n2062);
or (n2065,n2066,n2069);
and (n2066,n2067,n2068);
xor (n2067,n1959,n1960);
and (n2068,n467,n160);
and (n2069,n2070,n2071);
xor (n2070,n2067,n2068);
or (n2071,n2072,n2075);
and (n2072,n2073,n2074);
xor (n2073,n1965,n1966);
and (n2074,n364,n160);
and (n2075,n2076,n2077);
xor (n2076,n2073,n2074);
or (n2077,n2078,n2081);
and (n2078,n2079,n2080);
xor (n2079,n1971,n1972);
and (n2080,n268,n160);
and (n2081,n2082,n2083);
xor (n2082,n2079,n2080);
or (n2083,n2084,n2087);
and (n2084,n2085,n2086);
xor (n2085,n1977,n1978);
and (n2086,n260,n160);
and (n2087,n2088,n2089);
xor (n2088,n2085,n2086);
or (n2089,n2090,n2093);
and (n2090,n2091,n2092);
xor (n2091,n1983,n1984);
and (n2092,n333,n160);
and (n2093,n2094,n2095);
xor (n2094,n2091,n2092);
or (n2095,n2096,n2099);
and (n2096,n2097,n2098);
xor (n2097,n1989,n1990);
and (n2098,n325,n160);
and (n2099,n2100,n2101);
xor (n2100,n2097,n2098);
or (n2101,n2102,n2105);
and (n2102,n2103,n2104);
xor (n2103,n1995,n1996);
and (n2104,n572,n160);
and (n2105,n2106,n2107);
xor (n2106,n2103,n2104);
or (n2107,n2108,n2111);
and (n2108,n2109,n2110);
xor (n2109,n2001,n2002);
and (n2110,n597,n160);
and (n2111,n2112,n2113);
xor (n2112,n2109,n2110);
or (n2113,n2114,n2117);
and (n2114,n2115,n2116);
xor (n2115,n2007,n2008);
and (n2116,n516,n160);
and (n2117,n2118,n2119);
xor (n2118,n2115,n2116);
or (n2119,n2120,n2123);
and (n2120,n2121,n2122);
xor (n2121,n2013,n2014);
and (n2122,n402,n160);
and (n2123,n2124,n2125);
xor (n2124,n2121,n2122);
or (n2125,n2126,n2129);
and (n2126,n2127,n2128);
xor (n2127,n2019,n2020);
and (n2128,n393,n160);
and (n2129,n2130,n2131);
xor (n2130,n2127,n2128);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2025,n2026);
and (n2134,n435,n160);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2031,n2032);
and (n2140,n427,n160);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2037,n2038);
and (n2146,n126,n160);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
and (n2149,n2150,n2151);
xor (n2150,n2043,n2044);
and (n2151,n120,n160);
and (n2152,n452,n279);
or (n2153,n2154,n2157);
and (n2154,n2155,n2156);
xor (n2155,n2052,n2053);
and (n2156,n301,n279);
and (n2157,n2158,n2159);
xor (n2158,n2155,n2156);
or (n2159,n2160,n2163);
and (n2160,n2161,n2162);
xor (n2161,n2058,n2059);
and (n2162,n293,n279);
and (n2163,n2164,n2165);
xor (n2164,n2161,n2162);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2064,n2065);
and (n2168,n467,n279);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2070,n2071);
and (n2174,n364,n279);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
or (n2177,n2178,n2181);
and (n2178,n2179,n2180);
xor (n2179,n2076,n2077);
and (n2180,n268,n279);
and (n2181,n2182,n2183);
xor (n2182,n2179,n2180);
or (n2183,n2184,n2187);
and (n2184,n2185,n2186);
xor (n2185,n2082,n2083);
and (n2186,n260,n279);
and (n2187,n2188,n2189);
xor (n2188,n2185,n2186);
or (n2189,n2190,n2193);
and (n2190,n2191,n2192);
xor (n2191,n2088,n2089);
and (n2192,n333,n279);
and (n2193,n2194,n2195);
xor (n2194,n2191,n2192);
or (n2195,n2196,n2199);
and (n2196,n2197,n2198);
xor (n2197,n2094,n2095);
and (n2198,n325,n279);
and (n2199,n2200,n2201);
xor (n2200,n2197,n2198);
or (n2201,n2202,n2205);
and (n2202,n2203,n2204);
xor (n2203,n2100,n2101);
and (n2204,n572,n279);
and (n2205,n2206,n2207);
xor (n2206,n2203,n2204);
or (n2207,n2208,n2211);
and (n2208,n2209,n2210);
xor (n2209,n2106,n2107);
and (n2210,n597,n279);
and (n2211,n2212,n2213);
xor (n2212,n2209,n2210);
or (n2213,n2214,n2217);
and (n2214,n2215,n2216);
xor (n2215,n2112,n2113);
and (n2216,n516,n279);
and (n2217,n2218,n2219);
xor (n2218,n2215,n2216);
or (n2219,n2220,n2223);
and (n2220,n2221,n2222);
xor (n2221,n2118,n2119);
and (n2222,n402,n279);
and (n2223,n2224,n2225);
xor (n2224,n2221,n2222);
or (n2225,n2226,n2229);
and (n2226,n2227,n2228);
xor (n2227,n2124,n2125);
and (n2228,n393,n279);
and (n2229,n2230,n2231);
xor (n2230,n2227,n2228);
or (n2231,n2232,n2235);
and (n2232,n2233,n2234);
xor (n2233,n2130,n2131);
and (n2234,n435,n279);
and (n2235,n2236,n2237);
xor (n2236,n2233,n2234);
or (n2237,n2238,n2241);
and (n2238,n2239,n2240);
xor (n2239,n2136,n2137);
and (n2240,n427,n279);
and (n2241,n2242,n2243);
xor (n2242,n2239,n2240);
or (n2243,n2244,n2247);
and (n2244,n2245,n2246);
xor (n2245,n2142,n2143);
and (n2246,n126,n279);
and (n2247,n2248,n2249);
xor (n2248,n2245,n2246);
and (n2249,n2250,n1509);
xor (n2250,n2148,n2149);
and (n2251,n301,n286);
or (n2252,n2253,n2256);
and (n2253,n2254,n2255);
xor (n2254,n2158,n2159);
and (n2255,n293,n286);
and (n2256,n2257,n2258);
xor (n2257,n2254,n2255);
or (n2258,n2259,n2262);
and (n2259,n2260,n2261);
xor (n2260,n2164,n2165);
and (n2261,n467,n286);
and (n2262,n2263,n2264);
xor (n2263,n2260,n2261);
or (n2264,n2265,n2268);
and (n2265,n2266,n2267);
xor (n2266,n2170,n2171);
and (n2267,n364,n286);
and (n2268,n2269,n2270);
xor (n2269,n2266,n2267);
or (n2270,n2271,n2274);
and (n2271,n2272,n2273);
xor (n2272,n2176,n2177);
and (n2273,n268,n286);
and (n2274,n2275,n2276);
xor (n2275,n2272,n2273);
or (n2276,n2277,n2280);
and (n2277,n2278,n2279);
xor (n2278,n2182,n2183);
and (n2279,n260,n286);
and (n2280,n2281,n2282);
xor (n2281,n2278,n2279);
or (n2282,n2283,n2286);
and (n2283,n2284,n2285);
xor (n2284,n2188,n2189);
and (n2285,n333,n286);
and (n2286,n2287,n2288);
xor (n2287,n2284,n2285);
or (n2288,n2289,n2292);
and (n2289,n2290,n2291);
xor (n2290,n2194,n2195);
and (n2291,n325,n286);
and (n2292,n2293,n2294);
xor (n2293,n2290,n2291);
or (n2294,n2295,n2298);
and (n2295,n2296,n2297);
xor (n2296,n2200,n2201);
and (n2297,n572,n286);
and (n2298,n2299,n2300);
xor (n2299,n2296,n2297);
or (n2300,n2301,n2304);
and (n2301,n2302,n2303);
xor (n2302,n2206,n2207);
and (n2303,n597,n286);
and (n2304,n2305,n2306);
xor (n2305,n2302,n2303);
or (n2306,n2307,n2310);
and (n2307,n2308,n2309);
xor (n2308,n2212,n2213);
and (n2309,n516,n286);
and (n2310,n2311,n2312);
xor (n2311,n2308,n2309);
or (n2312,n2313,n2316);
and (n2313,n2314,n2315);
xor (n2314,n2218,n2219);
and (n2315,n402,n286);
and (n2316,n2317,n2318);
xor (n2317,n2314,n2315);
or (n2318,n2319,n2322);
and (n2319,n2320,n2321);
xor (n2320,n2224,n2225);
and (n2321,n393,n286);
and (n2322,n2323,n2324);
xor (n2323,n2320,n2321);
or (n2324,n2325,n2328);
and (n2325,n2326,n2327);
xor (n2326,n2230,n2231);
and (n2327,n435,n286);
and (n2328,n2329,n2330);
xor (n2329,n2326,n2327);
or (n2330,n2331,n2334);
and (n2331,n2332,n2333);
xor (n2332,n2236,n2237);
and (n2333,n427,n286);
and (n2334,n2335,n2336);
xor (n2335,n2332,n2333);
or (n2336,n2337,n2340);
and (n2337,n2338,n2339);
xor (n2338,n2242,n2243);
and (n2339,n126,n286);
and (n2340,n2341,n2342);
xor (n2341,n2338,n2339);
and (n2342,n2343,n2344);
xor (n2343,n2248,n2249);
and (n2344,n120,n286);
and (n2345,n293,n350);
or (n2346,n2347,n2350);
and (n2347,n2348,n2349);
xor (n2348,n2257,n2258);
and (n2349,n467,n350);
and (n2350,n2351,n2352);
xor (n2351,n2348,n2349);
or (n2352,n2353,n2356);
and (n2353,n2354,n2355);
xor (n2354,n2263,n2264);
and (n2355,n364,n350);
and (n2356,n2357,n2358);
xor (n2357,n2354,n2355);
or (n2358,n2359,n2362);
and (n2359,n2360,n2361);
xor (n2360,n2269,n2270);
and (n2361,n268,n350);
and (n2362,n2363,n2364);
xor (n2363,n2360,n2361);
or (n2364,n2365,n2368);
and (n2365,n2366,n2367);
xor (n2366,n2275,n2276);
and (n2367,n260,n350);
and (n2368,n2369,n2370);
xor (n2369,n2366,n2367);
or (n2370,n2371,n2374);
and (n2371,n2372,n2373);
xor (n2372,n2281,n2282);
and (n2373,n333,n350);
and (n2374,n2375,n2376);
xor (n2375,n2372,n2373);
or (n2376,n2377,n2380);
and (n2377,n2378,n2379);
xor (n2378,n2287,n2288);
and (n2379,n325,n350);
and (n2380,n2381,n2382);
xor (n2381,n2378,n2379);
or (n2382,n2383,n2386);
and (n2383,n2384,n2385);
xor (n2384,n2293,n2294);
and (n2385,n572,n350);
and (n2386,n2387,n2388);
xor (n2387,n2384,n2385);
or (n2388,n2389,n2392);
and (n2389,n2390,n2391);
xor (n2390,n2299,n2300);
and (n2391,n597,n350);
and (n2392,n2393,n2394);
xor (n2393,n2390,n2391);
or (n2394,n2395,n2398);
and (n2395,n2396,n2397);
xor (n2396,n2305,n2306);
and (n2397,n516,n350);
and (n2398,n2399,n2400);
xor (n2399,n2396,n2397);
or (n2400,n2401,n2404);
and (n2401,n2402,n2403);
xor (n2402,n2311,n2312);
and (n2403,n402,n350);
and (n2404,n2405,n2406);
xor (n2405,n2402,n2403);
or (n2406,n2407,n2410);
and (n2407,n2408,n2409);
xor (n2408,n2317,n2318);
and (n2409,n393,n350);
and (n2410,n2411,n2412);
xor (n2411,n2408,n2409);
or (n2412,n2413,n2416);
and (n2413,n2414,n2415);
xor (n2414,n2323,n2324);
and (n2415,n435,n350);
and (n2416,n2417,n2418);
xor (n2417,n2414,n2415);
or (n2418,n2419,n2422);
and (n2419,n2420,n2421);
xor (n2420,n2329,n2330);
and (n2421,n427,n350);
and (n2422,n2423,n2424);
xor (n2423,n2420,n2421);
or (n2424,n2425,n2428);
and (n2425,n2426,n2427);
xor (n2426,n2335,n2336);
and (n2427,n126,n350);
and (n2428,n2429,n2430);
xor (n2429,n2426,n2427);
and (n2430,n2431,n1408);
xor (n2431,n2341,n2342);
and (n2432,n467,n253);
or (n2433,n2434,n2437);
and (n2434,n2435,n2436);
xor (n2435,n2351,n2352);
and (n2436,n364,n253);
and (n2437,n2438,n2439);
xor (n2438,n2435,n2436);
or (n2439,n2440,n2443);
and (n2440,n2441,n2442);
xor (n2441,n2357,n2358);
and (n2442,n268,n253);
and (n2443,n2444,n2445);
xor (n2444,n2441,n2442);
or (n2445,n2446,n2449);
and (n2446,n2447,n2448);
xor (n2447,n2363,n2364);
and (n2448,n260,n253);
and (n2449,n2450,n2451);
xor (n2450,n2447,n2448);
or (n2451,n2452,n2455);
and (n2452,n2453,n2454);
xor (n2453,n2369,n2370);
and (n2454,n333,n253);
and (n2455,n2456,n2457);
xor (n2456,n2453,n2454);
or (n2457,n2458,n2461);
and (n2458,n2459,n2460);
xor (n2459,n2375,n2376);
and (n2460,n325,n253);
and (n2461,n2462,n2463);
xor (n2462,n2459,n2460);
or (n2463,n2464,n2467);
and (n2464,n2465,n2466);
xor (n2465,n2381,n2382);
and (n2466,n572,n253);
and (n2467,n2468,n2469);
xor (n2468,n2465,n2466);
or (n2469,n2470,n2473);
and (n2470,n2471,n2472);
xor (n2471,n2387,n2388);
and (n2472,n597,n253);
and (n2473,n2474,n2475);
xor (n2474,n2471,n2472);
or (n2475,n2476,n2479);
and (n2476,n2477,n2478);
xor (n2477,n2393,n2394);
and (n2478,n516,n253);
and (n2479,n2480,n2481);
xor (n2480,n2477,n2478);
or (n2481,n2482,n2485);
and (n2482,n2483,n2484);
xor (n2483,n2399,n2400);
and (n2484,n402,n253);
and (n2485,n2486,n2487);
xor (n2486,n2483,n2484);
or (n2487,n2488,n2491);
and (n2488,n2489,n2490);
xor (n2489,n2405,n2406);
and (n2490,n393,n253);
and (n2491,n2492,n2493);
xor (n2492,n2489,n2490);
or (n2493,n2494,n2496);
and (n2494,n2495,n1272);
xor (n2495,n2411,n2412);
and (n2496,n2497,n2498);
xor (n2497,n2495,n1272);
or (n2498,n2499,n2502);
and (n2499,n2500,n2501);
xor (n2500,n2417,n2418);
and (n2501,n427,n253);
and (n2502,n2503,n2504);
xor (n2503,n2500,n2501);
or (n2504,n2505,n2508);
and (n2505,n2506,n2507);
xor (n2506,n2423,n2424);
and (n2507,n126,n253);
and (n2508,n2509,n2510);
xor (n2509,n2506,n2507);
and (n2510,n2511,n2512);
xor (n2511,n2429,n2430);
and (n2512,n120,n253);
and (n2513,n364,n241);
or (n2514,n2515,n2518);
and (n2515,n2516,n2517);
xor (n2516,n2438,n2439);
and (n2517,n268,n241);
and (n2518,n2519,n2520);
xor (n2519,n2516,n2517);
or (n2520,n2521,n2524);
and (n2521,n2522,n2523);
xor (n2522,n2444,n2445);
and (n2523,n260,n241);
and (n2524,n2525,n2526);
xor (n2525,n2522,n2523);
or (n2526,n2527,n2530);
and (n2527,n2528,n2529);
xor (n2528,n2450,n2451);
and (n2529,n333,n241);
and (n2530,n2531,n2532);
xor (n2531,n2528,n2529);
or (n2532,n2533,n2536);
and (n2533,n2534,n2535);
xor (n2534,n2456,n2457);
and (n2535,n325,n241);
and (n2536,n2537,n2538);
xor (n2537,n2534,n2535);
or (n2538,n2539,n2542);
and (n2539,n2540,n2541);
xor (n2540,n2462,n2463);
and (n2541,n572,n241);
and (n2542,n2543,n2544);
xor (n2543,n2540,n2541);
or (n2544,n2545,n2548);
and (n2545,n2546,n2547);
xor (n2546,n2468,n2469);
and (n2547,n597,n241);
and (n2548,n2549,n2550);
xor (n2549,n2546,n2547);
or (n2550,n2551,n2554);
and (n2551,n2552,n2553);
xor (n2552,n2474,n2475);
and (n2553,n516,n241);
and (n2554,n2555,n2556);
xor (n2555,n2552,n2553);
or (n2556,n2557,n2560);
and (n2557,n2558,n2559);
xor (n2558,n2480,n2481);
and (n2559,n402,n241);
and (n2560,n2561,n2562);
xor (n2561,n2558,n2559);
or (n2562,n2563,n2566);
and (n2563,n2564,n2565);
xor (n2564,n2486,n2487);
and (n2565,n393,n241);
and (n2566,n2567,n2568);
xor (n2567,n2564,n2565);
or (n2568,n2569,n2572);
and (n2569,n2570,n2571);
xor (n2570,n2492,n2493);
and (n2571,n435,n241);
and (n2572,n2573,n2574);
xor (n2573,n2570,n2571);
or (n2574,n2575,n2578);
and (n2575,n2576,n2577);
xor (n2576,n2497,n2498);
and (n2577,n427,n241);
and (n2578,n2579,n2580);
xor (n2579,n2576,n2577);
or (n2580,n2581,n2584);
and (n2581,n2582,n2583);
xor (n2582,n2503,n2504);
and (n2583,n126,n241);
and (n2584,n2585,n2586);
xor (n2585,n2582,n2583);
and (n2586,n2587,n1301);
xor (n2587,n2509,n2510);
and (n2588,n268,n244);
or (n2589,n2590,n2593);
and (n2590,n2591,n2592);
xor (n2591,n2519,n2520);
and (n2592,n260,n244);
and (n2593,n2594,n2595);
xor (n2594,n2591,n2592);
or (n2595,n2596,n2599);
and (n2596,n2597,n2598);
xor (n2597,n2525,n2526);
and (n2598,n333,n244);
and (n2599,n2600,n2601);
xor (n2600,n2597,n2598);
or (n2601,n2602,n2605);
and (n2602,n2603,n2604);
xor (n2603,n2531,n2532);
and (n2604,n325,n244);
and (n2605,n2606,n2607);
xor (n2606,n2603,n2604);
or (n2607,n2608,n2611);
and (n2608,n2609,n2610);
xor (n2609,n2537,n2538);
and (n2610,n572,n244);
and (n2611,n2612,n2613);
xor (n2612,n2609,n2610);
or (n2613,n2614,n2617);
and (n2614,n2615,n2616);
xor (n2615,n2543,n2544);
and (n2616,n597,n244);
and (n2617,n2618,n2619);
xor (n2618,n2615,n2616);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
xor (n2621,n2549,n2550);
and (n2622,n516,n244);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
xor (n2627,n2555,n2556);
and (n2628,n402,n244);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
xor (n2633,n2561,n2562);
and (n2634,n393,n244);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
xor (n2639,n2567,n2568);
and (n2640,n435,n244);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
or (n2643,n2644,n2647);
and (n2644,n2645,n2646);
xor (n2645,n2573,n2574);
and (n2646,n427,n244);
and (n2647,n2648,n2649);
xor (n2648,n2645,n2646);
or (n2649,n2650,n2653);
and (n2650,n2651,n2652);
xor (n2651,n2579,n2580);
and (n2652,n126,n244);
and (n2653,n2654,n2655);
xor (n2654,n2651,n2652);
and (n2655,n2656,n2657);
xor (n2656,n2585,n2586);
and (n2657,n120,n244);
and (n2658,n260,n311);
or (n2659,n2660,n2663);
and (n2660,n2661,n2662);
xor (n2661,n2594,n2595);
and (n2662,n333,n311);
and (n2663,n2664,n2665);
xor (n2664,n2661,n2662);
or (n2665,n2666,n2669);
and (n2666,n2667,n2668);
xor (n2667,n2600,n2601);
and (n2668,n325,n311);
and (n2669,n2670,n2671);
xor (n2670,n2667,n2668);
or (n2671,n2672,n2675);
and (n2672,n2673,n2674);
xor (n2673,n2606,n2607);
and (n2674,n572,n311);
and (n2675,n2676,n2677);
xor (n2676,n2673,n2674);
or (n2677,n2678,n2681);
and (n2678,n2679,n2680);
xor (n2679,n2612,n2613);
and (n2680,n597,n311);
and (n2681,n2682,n2683);
xor (n2682,n2679,n2680);
or (n2683,n2684,n2687);
and (n2684,n2685,n2686);
xor (n2685,n2618,n2619);
and (n2686,n516,n311);
and (n2687,n2688,n2689);
xor (n2688,n2685,n2686);
or (n2689,n2690,n2693);
and (n2690,n2691,n2692);
xor (n2691,n2624,n2625);
and (n2692,n402,n311);
and (n2693,n2694,n2695);
xor (n2694,n2691,n2692);
or (n2695,n2696,n2699);
and (n2696,n2697,n2698);
xor (n2697,n2630,n2631);
and (n2698,n393,n311);
and (n2699,n2700,n2701);
xor (n2700,n2697,n2698);
or (n2701,n2702,n2705);
and (n2702,n2703,n2704);
xor (n2703,n2636,n2637);
and (n2704,n435,n311);
and (n2705,n2706,n2707);
xor (n2706,n2703,n2704);
or (n2707,n2708,n2711);
and (n2708,n2709,n2710);
xor (n2709,n2642,n2643);
and (n2710,n427,n311);
and (n2711,n2712,n2713);
xor (n2712,n2709,n2710);
or (n2713,n2714,n2717);
and (n2714,n2715,n2716);
xor (n2715,n2648,n2649);
and (n2716,n126,n311);
and (n2717,n2718,n2719);
xor (n2718,n2715,n2716);
and (n2719,n2720,n1110);
xor (n2720,n2654,n2655);
and (n2721,n333,n318);
or (n2722,n2723,n2726);
and (n2723,n2724,n2725);
xor (n2724,n2664,n2665);
and (n2725,n325,n318);
and (n2726,n2727,n2728);
xor (n2727,n2724,n2725);
or (n2728,n2729,n2732);
and (n2729,n2730,n2731);
xor (n2730,n2670,n2671);
and (n2731,n572,n318);
and (n2732,n2733,n2734);
xor (n2733,n2730,n2731);
or (n2734,n2735,n2738);
and (n2735,n2736,n2737);
xor (n2736,n2676,n2677);
and (n2737,n597,n318);
and (n2738,n2739,n2740);
xor (n2739,n2736,n2737);
or (n2740,n2741,n2744);
and (n2741,n2742,n2743);
xor (n2742,n2682,n2683);
and (n2743,n516,n318);
and (n2744,n2745,n2746);
xor (n2745,n2742,n2743);
or (n2746,n2747,n2750);
and (n2747,n2748,n2749);
xor (n2748,n2688,n2689);
and (n2749,n402,n318);
and (n2750,n2751,n2752);
xor (n2751,n2748,n2749);
or (n2752,n2753,n2756);
and (n2753,n2754,n2755);
xor (n2754,n2694,n2695);
and (n2755,n393,n318);
and (n2756,n2757,n2758);
xor (n2757,n2754,n2755);
or (n2758,n2759,n2762);
and (n2759,n2760,n2761);
xor (n2760,n2700,n2701);
and (n2761,n435,n318);
and (n2762,n2763,n2764);
xor (n2763,n2760,n2761);
or (n2764,n2765,n2768);
and (n2765,n2766,n2767);
xor (n2766,n2706,n2707);
and (n2767,n427,n318);
and (n2768,n2769,n2770);
xor (n2769,n2766,n2767);
or (n2770,n2771,n2774);
and (n2771,n2772,n2773);
xor (n2772,n2712,n2713);
and (n2773,n126,n318);
and (n2774,n2775,n2776);
xor (n2775,n2772,n2773);
and (n2776,n2777,n2778);
xor (n2777,n2718,n2719);
and (n2778,n120,n318);
and (n2779,n325,n583);
or (n2780,n2781,n2784);
and (n2781,n2782,n2783);
xor (n2782,n2727,n2728);
and (n2783,n572,n583);
and (n2784,n2785,n2786);
xor (n2785,n2782,n2783);
or (n2786,n2787,n2790);
and (n2787,n2788,n2789);
xor (n2788,n2733,n2734);
and (n2789,n597,n583);
and (n2790,n2791,n2792);
xor (n2791,n2788,n2789);
or (n2792,n2793,n2796);
and (n2793,n2794,n2795);
xor (n2794,n2739,n2740);
and (n2795,n516,n583);
and (n2796,n2797,n2798);
xor (n2797,n2794,n2795);
or (n2798,n2799,n2802);
and (n2799,n2800,n2801);
xor (n2800,n2745,n2746);
and (n2801,n402,n583);
and (n2802,n2803,n2804);
xor (n2803,n2800,n2801);
or (n2804,n2805,n2808);
and (n2805,n2806,n2807);
xor (n2806,n2751,n2752);
and (n2807,n393,n583);
and (n2808,n2809,n2810);
xor (n2809,n2806,n2807);
or (n2810,n2811,n2814);
and (n2811,n2812,n2813);
xor (n2812,n2757,n2758);
and (n2813,n435,n583);
and (n2814,n2815,n2816);
xor (n2815,n2812,n2813);
or (n2816,n2817,n2820);
and (n2817,n2818,n2819);
xor (n2818,n2763,n2764);
and (n2819,n427,n583);
and (n2820,n2821,n2822);
xor (n2821,n2818,n2819);
or (n2822,n2823,n2826);
and (n2823,n2824,n2825);
xor (n2824,n2769,n2770);
and (n2825,n126,n583);
and (n2826,n2827,n2828);
xor (n2827,n2824,n2825);
and (n2828,n2829,n1019);
xor (n2829,n2775,n2776);
and (n2830,n572,n376);
or (n2831,n2832,n2835);
and (n2832,n2833,n2834);
xor (n2833,n2785,n2786);
and (n2834,n597,n376);
and (n2835,n2836,n2837);
xor (n2836,n2833,n2834);
or (n2837,n2838,n2841);
and (n2838,n2839,n2840);
xor (n2839,n2791,n2792);
and (n2840,n516,n376);
and (n2841,n2842,n2843);
xor (n2842,n2839,n2840);
or (n2843,n2844,n2847);
and (n2844,n2845,n2846);
xor (n2845,n2797,n2798);
and (n2846,n402,n376);
and (n2847,n2848,n2849);
xor (n2848,n2845,n2846);
or (n2849,n2850,n2853);
and (n2850,n2851,n2852);
xor (n2851,n2803,n2804);
and (n2852,n393,n376);
and (n2853,n2854,n2855);
xor (n2854,n2851,n2852);
or (n2855,n2856,n2859);
and (n2856,n2857,n2858);
xor (n2857,n2809,n2810);
and (n2858,n435,n376);
and (n2859,n2860,n2861);
xor (n2860,n2857,n2858);
or (n2861,n2862,n2865);
and (n2862,n2863,n2864);
xor (n2863,n2815,n2816);
and (n2864,n427,n376);
and (n2865,n2866,n2867);
xor (n2866,n2863,n2864);
or (n2867,n2868,n2871);
and (n2868,n2869,n2870);
xor (n2869,n2821,n2822);
and (n2870,n126,n376);
and (n2871,n2872,n2873);
xor (n2872,n2869,n2870);
and (n2873,n2874,n2875);
xor (n2874,n2827,n2828);
and (n2875,n120,n376);
and (n2876,n597,n379);
or (n2877,n2878,n2881);
and (n2878,n2879,n2880);
xor (n2879,n2836,n2837);
and (n2880,n516,n379);
and (n2881,n2882,n2883);
xor (n2882,n2879,n2880);
or (n2883,n2884,n2887);
and (n2884,n2885,n2886);
xor (n2885,n2842,n2843);
and (n2886,n402,n379);
and (n2887,n2888,n2889);
xor (n2888,n2885,n2886);
or (n2889,n2890,n2893);
and (n2890,n2891,n2892);
xor (n2891,n2848,n2849);
and (n2892,n393,n379);
and (n2893,n2894,n2895);
xor (n2894,n2891,n2892);
or (n2895,n2896,n2899);
and (n2896,n2897,n2898);
xor (n2897,n2854,n2855);
and (n2898,n435,n379);
and (n2899,n2900,n2901);
xor (n2900,n2897,n2898);
or (n2901,n2902,n2905);
and (n2902,n2903,n2904);
xor (n2903,n2860,n2861);
and (n2904,n427,n379);
and (n2905,n2906,n2907);
xor (n2906,n2903,n2904);
or (n2907,n2908,n2911);
and (n2908,n2909,n2910);
xor (n2909,n2866,n2867);
and (n2910,n126,n379);
and (n2911,n2912,n2913);
xor (n2912,n2909,n2910);
and (n2913,n2914,n1218);
xor (n2914,n2872,n2873);
and (n2915,n516,n386);
or (n2916,n2917,n2920);
and (n2917,n2918,n2919);
xor (n2918,n2882,n2883);
and (n2919,n402,n386);
and (n2920,n2921,n2922);
xor (n2921,n2918,n2919);
or (n2922,n2923,n2926);
and (n2923,n2924,n2925);
xor (n2924,n2888,n2889);
and (n2925,n393,n386);
and (n2926,n2927,n2928);
xor (n2927,n2924,n2925);
or (n2928,n2929,n2932);
and (n2929,n2930,n2931);
xor (n2930,n2894,n2895);
and (n2931,n435,n386);
and (n2932,n2933,n2934);
xor (n2933,n2930,n2931);
or (n2934,n2935,n2938);
and (n2935,n2936,n2937);
xor (n2936,n2900,n2901);
and (n2937,n427,n386);
and (n2938,n2939,n2940);
xor (n2939,n2936,n2937);
or (n2940,n2941,n2944);
and (n2941,n2942,n2943);
xor (n2942,n2906,n2907);
and (n2943,n126,n386);
and (n2944,n2945,n2946);
xor (n2945,n2942,n2943);
and (n2946,n2947,n2948);
xor (n2947,n2912,n2913);
and (n2948,n120,n386);
and (n2949,n402,n414);
or (n2950,n2951,n2954);
and (n2951,n2952,n2953);
xor (n2952,n2921,n2922);
and (n2953,n393,n414);
and (n2954,n2955,n2956);
xor (n2955,n2952,n2953);
or (n2956,n2957,n2960);
and (n2957,n2958,n2959);
xor (n2958,n2927,n2928);
and (n2959,n435,n414);
and (n2960,n2961,n2962);
xor (n2961,n2958,n2959);
or (n2962,n2963,n2966);
and (n2963,n2964,n2965);
xor (n2964,n2933,n2934);
and (n2965,n427,n414);
and (n2966,n2967,n2968);
xor (n2967,n2964,n2965);
or (n2968,n2969,n2972);
and (n2969,n2970,n2971);
xor (n2970,n2939,n2940);
and (n2971,n126,n414);
and (n2972,n2973,n2974);
xor (n2973,n2970,n2971);
and (n2974,n2975,n797);
xor (n2975,n2945,n2946);
and (n2976,n393,n420);
or (n2977,n2978,n2981);
and (n2978,n2979,n2980);
xor (n2979,n2955,n2956);
and (n2980,n435,n420);
and (n2981,n2982,n2983);
xor (n2982,n2979,n2980);
or (n2983,n2984,n2987);
and (n2984,n2985,n2986);
xor (n2985,n2961,n2962);
and (n2986,n427,n420);
and (n2987,n2988,n2989);
xor (n2988,n2985,n2986);
or (n2989,n2990,n2993);
and (n2990,n2991,n2992);
xor (n2991,n2967,n2968);
and (n2992,n126,n420);
and (n2993,n2994,n2995);
xor (n2994,n2991,n2992);
and (n2995,n2996,n2997);
xor (n2996,n2973,n2974);
and (n2997,n120,n420);
and (n2998,n435,n608);
or (n2999,n3000,n3003);
and (n3000,n3001,n3002);
xor (n3001,n2982,n2983);
and (n3002,n427,n608);
and (n3003,n3004,n3005);
xor (n3004,n3001,n3002);
or (n3005,n3006,n3009);
and (n3006,n3007,n3008);
xor (n3007,n2988,n2989);
and (n3008,n126,n608);
and (n3009,n3010,n3011);
xor (n3010,n3007,n3008);
and (n3011,n3012,n688);
xor (n3012,n2994,n2995);
and (n3013,n427,n18);
or (n3014,n3015,n3018);
and (n3015,n3016,n3017);
xor (n3016,n3004,n3005);
and (n3017,n126,n18);
and (n3018,n3019,n3020);
xor (n3019,n3016,n3017);
and (n3020,n3021,n3022);
xor (n3021,n3010,n3011);
and (n3022,n120,n18);
and (n3023,n126,n99);
and (n3024,n3025,n141);
xor (n3025,n3019,n3020);
and (n3026,n120,n109);
endmodule
