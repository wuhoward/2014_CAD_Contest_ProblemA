module top (out,n8,n21,n24,n25,n33,n34,n40,n41,n46
        ,n54,n56,n57,n66,n67,n77,n92,n93,n96,n102
        ,n124,n125,n132,n243,n246,n247,n257,n266,n274,n280
        ,n290,n296,n303,n309,n668,n746,n758,n773,n779,n783
        ,n788,n793,n799,n805,n810,n832,n843,n858,n869);
output out;
input n8;
input n21;
input n24;
input n25;
input n33;
input n34;
input n40;
input n41;
input n46;
input n54;
input n56;
input n57;
input n66;
input n67;
input n77;
input n92;
input n93;
input n96;
input n102;
input n124;
input n125;
input n132;
input n243;
input n246;
input n247;
input n257;
input n266;
input n274;
input n280;
input n290;
input n296;
input n303;
input n309;
input n668;
input n746;
input n758;
input n773;
input n779;
input n783;
input n788;
input n793;
input n799;
input n805;
input n810;
input n832;
input n843;
input n858;
input n869;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n244;
wire n245;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n780;
wire n781;
wire n782;
wire n784;
wire n785;
wire n786;
wire n787;
wire n789;
wire n790;
wire n791;
wire n792;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n806;
wire n807;
wire n808;
wire n809;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
xor (out,n0,n887);
nand (n0,n1,n886);
or (n1,n2,n670);
not (n2,n3);
and (n3,n4,n669);
or (n4,n5,n668);
nand (n5,n6,n228);
or (n6,n7,n9);
not (n7,n8);
not (n9,n10);
xor (n10,n11,n144);
xor (n11,n12,n107);
or (n12,n13,n106);
and (n13,n14,n80);
xor (n14,n15,n49);
nand (n15,n16,n43);
or (n16,n17,n27);
not (n17,n18);
nor (n18,n19,n26);
and (n19,n20,n22);
not (n20,n21);
not (n22,n23);
wire s0n23,s1n23,notn23;
or (n23,s0n23,s1n23);
not(notn23,n8);
and (s0n23,notn23,n24);
and (s1n23,n8,n25);
and (n26,n21,n23);
not (n27,n28);
and (n28,n29,n36);
nand (n29,n30,n35);
or (n30,n31,n23);
not (n31,n32);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n8);
and (s0n32,notn32,n33);
and (s1n32,n8,n34);
nand (n35,n23,n31);
not (n36,n37);
nand (n37,n38,n42);
or (n38,n31,n39);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n8);
and (s0n39,notn39,n40);
and (s1n39,n8,n41);
nand (n42,n39,n31);
nand (n43,n37,n44);
nor (n44,n45,n47);
and (n45,n46,n23);
and (n47,n22,n48);
not (n48,n46);
nand (n49,n50,n69);
or (n50,n51,n61);
not (n51,n52);
nor (n52,n53,n58);
and (n53,n54,n55);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n8);
and (s0n55,notn55,n56);
and (s1n55,n8,n57);
and (n58,n59,n60);
not (n59,n54);
not (n60,n55);
not (n61,n62);
nand (n62,n63,n68);
or (n63,n64,n23);
not (n64,n65);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n8);
and (s0n65,notn65,n66);
and (s1n65,n8,n67);
nand (n68,n23,n64);
nand (n69,n70,n75);
not (n70,n71);
nand (n71,n61,n72);
nand (n72,n73,n74);
or (n73,n64,n55);
nand (n74,n55,n64);
nand (n75,n76,n78);
or (n76,n60,n77);
or (n78,n55,n79);
not (n79,n77);
xor (n80,n81,n86);
and (n81,n82,n55);
nand (n82,n83,n85);
or (n83,n23,n84);
and (n84,n77,n65);
or (n85,n65,n77);
nand (n86,n87,n99);
or (n87,n88,n94);
not (n88,n89);
nor (n89,n90,n91);
not (n90,n39);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n8);
and (s0n91,notn91,n92);
and (s1n91,n8,n93);
nor (n94,n95,n97);
and (n95,n90,n96);
and (n97,n39,n98);
not (n98,n96);
or (n99,n100,n105);
nor (n100,n101,n103);
and (n101,n102,n90);
and (n103,n104,n39);
not (n104,n102);
not (n105,n91);
and (n106,n15,n49);
xor (n107,n108,n116);
xor (n108,n109,n115);
nand (n109,n110,n111);
or (n110,n51,n71);
or (n111,n61,n112);
nor (n112,n113,n114);
and (n113,n60,n21);
and (n114,n55,n20);
and (n115,n81,n86);
xor (n116,n117,n137);
xor (n117,n118,n127);
and (n118,n119,n77);
not (n119,n120);
nor (n120,n121,n126);
and (n121,n122,n55);
not (n122,n123);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n8);
and (s0n123,notn123,n124);
and (s1n123,n8,n125);
and (n126,n123,n60);
nand (n127,n128,n135);
or (n128,n105,n129);
not (n129,n130);
nor (n130,n131,n133);
and (n131,n132,n39);
and (n133,n134,n90);
not (n134,n132);
nand (n135,n136,n89);
not (n136,n100);
nand (n137,n138,n140);
or (n138,n139,n27);
not (n139,n44);
nand (n140,n37,n141);
nand (n141,n142,n143);
or (n142,n23,n98);
or (n143,n22,n96);
or (n144,n145,n227);
and (n145,n146,n167);
xor (n146,n147,n166);
or (n147,n148,n165);
and (n148,n149,n158);
xor (n149,n150,n151);
and (n150,n62,n77);
nand (n151,n152,n157);
or (n152,n153,n27);
not (n153,n154);
nor (n154,n155,n156);
and (n155,n54,n23);
and (n156,n59,n22);
nand (n157,n18,n37);
nand (n158,n159,n164);
or (n159,n88,n160);
not (n160,n161);
nor (n161,n162,n163);
and (n162,n48,n90);
and (n163,n46,n39);
or (n164,n94,n105);
and (n165,n150,n151);
xor (n166,n14,n80);
or (n167,n168,n226);
and (n168,n169,n225);
xor (n169,n170,n184);
nor (n170,n171,n179);
not (n171,n172);
nand (n172,n173,n178);
or (n173,n174,n88);
not (n174,n175);
nand (n175,n176,n177);
or (n176,n20,n39);
nand (n177,n39,n20);
nand (n178,n161,n91);
nand (n179,n180,n23);
nand (n180,n181,n183);
or (n181,n39,n182);
and (n182,n77,n32);
or (n183,n32,n77);
nand (n184,n185,n223);
or (n185,n186,n209);
not (n186,n187);
nand (n187,n188,n208);
or (n188,n189,n198);
nor (n189,n190,n197);
nand (n190,n191,n196);
or (n191,n192,n88);
not (n192,n193);
nand (n193,n194,n195);
or (n194,n59,n39);
nand (n195,n39,n59);
nand (n196,n175,n91);
nor (n197,n36,n79);
nand (n198,n199,n206);
nand (n199,n200,n205);
or (n200,n201,n88);
not (n201,n202);
nand (n202,n203,n204);
or (n203,n90,n77);
or (n204,n39,n79);
nand (n205,n193,n91);
nor (n206,n207,n90);
and (n207,n77,n91);
nand (n208,n190,n197);
not (n209,n210);
nand (n210,n211,n219);
not (n211,n212);
nand (n212,n213,n218);
or (n213,n214,n27);
not (n214,n215);
nand (n215,n216,n217);
or (n216,n22,n77);
or (n217,n23,n79);
nand (n218,n37,n154);
nor (n219,n220,n222);
and (n220,n171,n221);
not (n221,n179);
and (n222,n172,n179);
nand (n223,n224,n212);
not (n224,n219);
xor (n225,n149,n158);
and (n226,n170,n184);
and (n227,n147,n166);
nand (n228,n229,n7);
nand (n229,n230,n667);
or (n230,n231,n432);
not (n231,n232);
nand (n232,n233,n431);
nand (n233,n234,n385);
not (n234,n235);
xor (n235,n236,n345);
xor (n236,n237,n283);
xor (n237,n238,n270);
xor (n238,n239,n260);
nand (n239,n240,n254);
or (n240,n241,n250);
nor (n241,n242,n248);
and (n242,n243,n244);
not (n244,n245);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n8);
and (s0n245,notn245,n246);
and (s1n245,n8,n247);
and (n248,n249,n245);
not (n249,n243);
nand (n250,n120,n251);
nand (n251,n252,n253);
or (n252,n122,n245);
nand (n253,n245,n122);
nand (n254,n119,n255);
nor (n255,n256,n258);
and (n256,n257,n245);
and (n258,n259,n244);
not (n259,n257);
nor (n260,n261,n267);
nand (n261,n245,n262);
not (n262,n263);
wire s0n263,s1n263,notn263;
or (n263,s0n263,s1n263);
not(notn263,n8);
and (s0n263,notn263,1'b0);
and (s1n263,n8,n265);
and (n265,n266,n247);
nor (n267,n268,n269);
and (n268,n263,n134);
and (n269,n262,n132);
nand (n270,n271,n277);
or (n271,n71,n272);
nor (n272,n273,n275);
and (n273,n60,n274);
and (n275,n55,n276);
not (n276,n274);
or (n277,n61,n278);
nor (n278,n279,n281);
and (n279,n60,n280);
and (n281,n55,n282);
not (n282,n280);
xor (n283,n284,n325);
xor (n284,n285,n312);
xor (n285,n286,n299);
nand (n286,n287,n293);
or (n287,n88,n288);
nor (n288,n289,n291);
and (n289,n90,n290);
and (n291,n39,n292);
not (n292,n290);
or (n293,n294,n105);
nor (n294,n295,n297);
and (n295,n90,n296);
and (n297,n39,n298);
not (n298,n296);
nand (n299,n300,n306);
or (n300,n27,n301);
nor (n301,n302,n304);
and (n302,n22,n303);
and (n304,n23,n305);
not (n305,n303);
or (n306,n36,n307);
nor (n307,n308,n310);
and (n308,n22,n309);
and (n310,n23,n311);
not (n311,n309);
and (n312,n313,n319);
nand (n313,n314,n318);
or (n314,n88,n315);
nor (n315,n316,n317);
and (n316,n90,n309);
and (n317,n39,n311);
or (n318,n288,n105);
nand (n319,n320,n324);
or (n320,n27,n321);
nor (n321,n322,n323);
and (n322,n22,n280);
and (n323,n23,n282);
or (n324,n301,n36);
or (n325,n326,n344);
and (n326,n327,n338);
xor (n327,n328,n334);
nand (n328,n329,n333);
or (n329,n250,n330);
nor (n330,n331,n332);
and (n331,n244,n132);
and (n332,n245,n134);
or (n333,n120,n241);
nor (n334,n261,n335);
nor (n335,n336,n337);
and (n336,n263,n104);
and (n337,n262,n102);
nand (n338,n339,n340);
or (n339,n272,n61);
or (n340,n71,n341);
nor (n341,n342,n343);
and (n342,n60,n257);
and (n343,n55,n259);
and (n344,n328,n334);
or (n345,n346,n384);
and (n346,n347,n362);
xor (n347,n348,n349);
xor (n348,n313,n319);
and (n349,n350,n356);
nand (n350,n351,n355);
or (n351,n88,n352);
nor (n352,n353,n354);
and (n353,n90,n303);
and (n354,n39,n305);
or (n355,n315,n105);
nand (n356,n357,n361);
or (n357,n27,n358);
nor (n358,n359,n360);
and (n359,n22,n274);
and (n360,n23,n276);
or (n361,n321,n36);
or (n362,n363,n383);
and (n363,n364,n377);
xor (n364,n365,n373);
nand (n365,n366,n371);
or (n366,n367,n250);
not (n367,n368);
nor (n368,n369,n370);
and (n369,n102,n245);
and (n370,n104,n244);
nand (n371,n372,n119);
not (n372,n330);
nor (n373,n261,n374);
nor (n374,n375,n376);
and (n375,n263,n98);
and (n376,n262,n96);
nand (n377,n378,n382);
or (n378,n71,n379);
nor (n379,n380,n381);
and (n380,n60,n243);
and (n381,n55,n249);
or (n382,n61,n341);
and (n383,n365,n373);
and (n384,n348,n349);
not (n385,n386);
or (n386,n387,n430);
and (n387,n388,n391);
xor (n388,n389,n390);
xor (n389,n327,n338);
xor (n390,n347,n362);
or (n391,n392,n429);
and (n392,n393,n408);
xor (n393,n394,n395);
xor (n394,n350,n356);
and (n395,n396,n402);
nand (n396,n397,n401);
or (n397,n88,n398);
nor (n398,n399,n400);
and (n399,n90,n280);
and (n400,n39,n282);
or (n401,n352,n105);
nand (n402,n403,n407);
or (n403,n27,n404);
nor (n404,n405,n406);
and (n405,n22,n257);
and (n406,n23,n259);
or (n407,n36,n358);
or (n408,n409,n428);
and (n409,n410,n422);
xor (n410,n411,n418);
nand (n411,n412,n417);
or (n412,n413,n250);
not (n413,n414);
nor (n414,n415,n416);
and (n415,n96,n245);
and (n416,n98,n244);
nand (n417,n119,n368);
nor (n418,n261,n419);
nor (n419,n420,n421);
and (n420,n263,n48);
and (n421,n262,n46);
nand (n422,n423,n427);
or (n423,n71,n424);
nor (n424,n425,n426);
and (n425,n60,n132);
and (n426,n55,n134);
or (n427,n61,n379);
and (n428,n411,n418);
and (n429,n394,n395);
and (n430,n389,n390);
nand (n431,n235,n386);
not (n432,n433);
nand (n433,n434,n662);
or (n434,n435,n516);
nand (n435,n436,n484);
not (n436,n437);
nor (n437,n438,n439);
xor (n438,n388,n391);
or (n439,n440,n483);
and (n440,n441,n444);
xor (n441,n442,n443);
xor (n442,n364,n377);
xor (n443,n393,n408);
or (n444,n445,n482);
and (n445,n446,n461);
xor (n446,n447,n448);
xor (n447,n396,n402);
and (n448,n449,n455);
nand (n449,n450,n454);
or (n450,n88,n451);
nor (n451,n452,n453);
and (n452,n90,n274);
and (n453,n39,n276);
or (n454,n398,n105);
nand (n455,n456,n460);
or (n456,n27,n457);
nor (n457,n458,n459);
and (n458,n22,n243);
and (n459,n23,n249);
or (n460,n404,n36);
or (n461,n462,n481);
and (n462,n463,n475);
xor (n463,n464,n471);
nand (n464,n465,n470);
or (n465,n466,n250);
not (n466,n467);
nor (n467,n468,n469);
and (n468,n46,n245);
and (n469,n48,n244);
nand (n470,n119,n414);
nor (n471,n261,n472);
nor (n472,n473,n474);
and (n473,n263,n20);
and (n474,n262,n21);
nand (n475,n476,n480);
or (n476,n71,n477);
nor (n477,n478,n479);
and (n478,n60,n102);
and (n479,n55,n104);
or (n480,n61,n424);
and (n481,n464,n471);
and (n482,n447,n448);
and (n483,n442,n443);
nand (n484,n485,n487);
not (n485,n486);
xor (n486,n441,n444);
not (n487,n488);
or (n488,n489,n515);
and (n489,n490,n493);
xor (n490,n491,n492);
xor (n491,n410,n422);
xor (n492,n446,n461);
and (n493,n494,n495);
xor (n494,n449,n455);
or (n495,n496,n514);
and (n496,n497,n508);
xor (n497,n498,n504);
nand (n498,n499,n503);
or (n499,n500,n250);
nor (n500,n501,n502);
and (n501,n21,n244);
and (n502,n20,n245);
nand (n503,n467,n119);
nor (n504,n261,n505);
nor (n505,n506,n507);
and (n506,n263,n59);
and (n507,n262,n54);
nand (n508,n509,n513);
or (n509,n88,n510);
nor (n510,n511,n512);
and (n511,n90,n257);
and (n512,n39,n259);
or (n513,n451,n105);
and (n514,n498,n504);
and (n515,n491,n492);
not (n516,n517);
nand (n517,n518,n643,n661);
nand (n518,n519,n636);
nand (n519,n520,n635);
or (n520,n521,n624);
nor (n521,n522,n623);
and (n522,n523,n611);
not (n523,n524);
nor (n524,n525,n594);
or (n525,n526,n593);
and (n526,n527,n568);
xor (n527,n528,n555);
or (n528,n529,n554);
and (n529,n530,n548);
xor (n530,n531,n541);
nand (n531,n532,n537);
or (n532,n533,n250);
not (n533,n534);
nand (n534,n535,n536);
or (n535,n244,n77);
or (n536,n245,n79);
or (n537,n120,n538);
nor (n538,n539,n540);
and (n539,n54,n244);
and (n540,n59,n245);
nand (n541,n542,n544);
or (n542,n543,n27);
not (n543,n141);
nand (n544,n37,n545);
nor (n545,n546,n547);
and (n546,n102,n23);
and (n547,n104,n22);
nand (n548,n549,n550);
or (n549,n71,n112);
or (n550,n61,n551);
nor (n551,n552,n553);
and (n552,n60,n46);
and (n553,n55,n48);
and (n554,n531,n541);
xor (n555,n556,n565);
xor (n556,n557,n559);
and (n557,n558,n77);
not (n558,n261);
nand (n559,n560,n564);
or (n560,n88,n561);
nor (n561,n562,n563);
and (n562,n249,n39);
and (n563,n243,n90);
or (n564,n510,n105);
nand (n565,n566,n567);
or (n566,n250,n538);
or (n567,n120,n500);
xor (n568,n569,n583);
xor (n569,n570,n577);
nand (n570,n571,n573);
or (n571,n27,n572);
not (n572,n545);
or (n573,n36,n574);
nor (n574,n575,n576);
and (n575,n22,n132);
and (n576,n23,n134);
nand (n577,n578,n579);
or (n578,n71,n551);
or (n579,n61,n580);
nor (n580,n581,n582);
and (n581,n60,n96);
and (n582,n55,n98);
and (n583,n584,n589);
nor (n584,n585,n244);
nor (n585,n586,n588);
and (n586,n60,n587);
nand (n587,n123,n77);
and (n588,n122,n79);
nand (n589,n590,n591);
or (n590,n129,n88);
nand (n591,n592,n91);
not (n592,n561);
and (n593,n528,n555);
xor (n594,n595,n600);
xor (n595,n596,n597);
xor (n596,n497,n508);
or (n597,n598,n599);
and (n598,n569,n583);
and (n599,n570,n577);
xor (n600,n601,n608);
xor (n601,n602,n605);
nand (n602,n603,n604);
or (n603,n71,n580);
or (n604,n61,n477);
nand (n605,n606,n607);
or (n606,n27,n574);
or (n607,n457,n36);
or (n608,n609,n610);
and (n609,n556,n565);
and (n610,n557,n559);
not (n611,n612);
nand (n612,n613,n614);
xor (n613,n527,n568);
or (n614,n615,n622);
and (n615,n616,n621);
xor (n616,n617,n618);
xor (n617,n584,n589);
or (n618,n619,n620);
and (n619,n117,n137);
and (n620,n118,n127);
xor (n621,n530,n548);
and (n622,n617,n618);
and (n623,n525,n594);
nor (n624,n625,n632);
xor (n625,n626,n629);
xor (n626,n627,n628);
xor (n627,n463,n475);
xor (n628,n494,n495);
or (n629,n630,n631);
and (n630,n601,n608);
and (n631,n602,n605);
or (n632,n633,n634);
and (n633,n595,n600);
and (n634,n596,n597);
nand (n635,n625,n632);
nand (n636,n637,n639);
not (n637,n638);
xor (n638,n490,n493);
not (n639,n640);
or (n640,n641,n642);
and (n641,n626,n629);
and (n642,n627,n628);
nand (n643,n636,n644,n660);
nor (n644,n645,n657);
nor (n645,n646,n655);
and (n646,n647,n650);
or (n647,n648,n649);
and (n648,n11,n144);
and (n649,n12,n107);
or (n650,n651,n652);
xor (n651,n616,n621);
or (n652,n653,n654);
and (n653,n108,n116);
and (n654,n109,n115);
not (n655,n656);
nand (n656,n651,n652);
nand (n657,n658,n523);
not (n658,n659);
nor (n659,n613,n614);
not (n660,n624);
nand (n661,n638,n640);
not (n662,n663);
nand (n663,n664,n666);
or (n664,n437,n665);
nand (n665,n486,n488);
nand (n666,n438,n439);
or (n667,n433,n232);
nand (n669,n5,n668);
not (n670,n671);
nor (n671,n672,n870,n882);
and (n672,n673,n759);
nor (n673,n674,n747);
nor (n674,n675,n746);
nand (n675,n676,n736);
or (n676,n7,n677);
not (n677,n678);
xor (n678,n679,n735);
xor (n679,n680,n733);
xor (n680,n681,n732);
xor (n681,n682,n724);
xor (n682,n683,n26);
xor (n683,n684,n710);
xor (n684,n685,n709);
xor (n685,n686,n689);
xor (n686,n687,n688);
and (n687,n102,n91);
and (n688,n96,n39);
or (n689,n690,n692);
and (n690,n691,n163);
and (n691,n96,n91);
and (n692,n693,n694);
xor (n693,n691,n163);
or (n694,n695,n698);
and (n695,n696,n697);
and (n696,n46,n91);
and (n697,n21,n39);
and (n698,n699,n700);
xor (n699,n696,n697);
or (n700,n701,n704);
and (n701,n702,n703);
and (n702,n21,n91);
and (n703,n54,n39);
and (n704,n705,n706);
xor (n705,n702,n703);
and (n706,n707,n708);
and (n707,n54,n91);
and (n708,n77,n39);
and (n709,n46,n32);
or (n710,n711,n714);
and (n711,n712,n713);
xor (n712,n693,n694);
and (n713,n21,n32);
and (n714,n715,n716);
xor (n715,n712,n713);
or (n716,n717,n720);
and (n717,n718,n719);
xor (n718,n699,n700);
and (n719,n54,n32);
and (n720,n721,n722);
xor (n721,n718,n719);
and (n722,n723,n182);
xor (n723,n705,n706);
or (n724,n725,n727);
and (n725,n726,n155);
xor (n726,n715,n716);
and (n727,n728,n729);
xor (n728,n726,n155);
and (n729,n730,n731);
xor (n730,n721,n722);
and (n731,n77,n23);
and (n732,n54,n65);
and (n733,n734,n84);
xor (n734,n728,n729);
and (n735,n77,n55);
nand (n736,n737,n7);
nand (n737,n738,n745);
or (n738,n739,n741);
not (n739,n740);
nand (n740,n436,n666);
not (n741,n742);
nand (n742,n743,n665);
or (n743,n744,n516);
not (n744,n484);
or (n745,n742,n740);
nor (n747,n748,n758);
nand (n748,n749,n752);
or (n749,n7,n750);
not (n750,n751);
xor (n751,n734,n84);
nand (n752,n753,n7);
nand (n753,n754,n757);
or (n754,n755,n516);
not (n755,n756);
nand (n756,n484,n665);
or (n757,n517,n756);
not (n759,n760);
nand (n760,n761,n819,n844);
not (n761,n762);
not (n762,n763);
or (n763,n764,n774,n818);
not (n764,n765);
nand (n765,n766,n773);
and (n766,n767,n7);
nand (n767,n768,n772);
or (n768,n769,n770);
not (n769,n647);
not (n770,n771);
nand (n771,n650,n656);
or (n772,n771,n647);
and (n774,n766,n775);
or (n775,n776,n780,n817);
not (n776,n777);
nand (n777,n778,n779);
and (n778,n10,n7);
and (n780,n778,n781);
or (n781,n782,n785,n816);
and (n782,n783,n784);
wire s0n784,s1n784,notn784;
or (n784,s0n784,s1n784);
not(notn784,n8);
and (s0n784,notn784,n678);
and (s1n784,n8,1'b0);
and (n785,n784,n786);
or (n786,n787,n790,n815);
and (n787,n788,n789);
wire s0n789,s1n789,notn789;
or (n789,s0n789,s1n789);
not(notn789,n8);
and (s0n789,notn789,n751);
and (s1n789,n8,1'b0);
and (n790,n789,n791);
or (n791,n792,n796,n814);
and (n792,n793,n794);
wire s0n794,s1n794,notn794;
or (n794,s0n794,s1n794);
not(notn794,n8);
and (s0n794,notn794,n795);
and (s1n794,n8,1'b0);
xor (n795,n730,n731);
and (n796,n794,n797);
or (n797,n798,n802,n813);
and (n798,n799,n800);
wire s0n800,s1n800,notn800;
or (n800,s0n800,s1n800);
not(notn800,n8);
and (s0n800,notn800,n801);
and (s1n800,n8,1'b0);
xor (n801,n723,n182);
and (n802,n800,n803);
or (n803,n804,n808,n812);
and (n804,n805,n806);
wire s0n806,s1n806,notn806;
or (n806,s0n806,s1n806);
not(notn806,n8);
and (s0n806,notn806,n807);
and (s1n806,n8,1'b0);
xor (n807,n707,n708);
and (n808,n806,n809);
and (n809,n810,n811);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n8);
and (s0n811,notn811,n207);
and (s1n811,n8,1'b0);
and (n812,n805,n809);
and (n813,n799,n803);
and (n814,n793,n797);
and (n815,n788,n791);
and (n816,n783,n786);
and (n817,n779,n781);
and (n818,n773,n775);
nor (n819,n820,n833);
nor (n820,n821,n832);
nand (n821,n822,n824);
or (n822,n7,n823);
not (n823,n795);
nand (n824,n825,n7);
xnor (n825,n826,n827);
nand (n826,n636,n661);
nand (n827,n828,n635);
or (n828,n624,n829);
not (n829,n830);
nand (n830,n831,n521);
not (n831,n644);
nor (n833,n834,n843);
nand (n834,n835,n837);
or (n835,n7,n836);
not (n836,n801);
nand (n837,n838,n7);
nand (n838,n839,n842);
or (n839,n840,n829);
not (n840,n841);
nand (n841,n660,n635);
or (n842,n830,n841);
nor (n844,n845,n859);
nor (n845,n846,n858);
nand (n846,n847,n849);
or (n847,n7,n848);
not (n848,n807);
nand (n849,n850,n7);
nand (n850,n851,n857);
or (n851,n852,n854);
not (n852,n853);
or (n853,n623,n524);
not (n854,n855);
nand (n855,n856,n612);
or (n856,n645,n659);
or (n857,n855,n853);
nor (n859,n860,n869);
or (n860,n861,n862);
and (n861,n8,n207);
and (n862,n7,n863);
nand (n863,n864,n868);
or (n864,n865,n866);
not (n865,n645);
not (n866,n867);
nor (n867,n611,n659);
or (n868,n867,n645);
and (n870,n673,n871);
not (n871,n872);
nor (n872,n873,n878);
and (n873,n819,n874);
nand (n874,n875,n877);
or (n875,n845,n876);
nand (n876,n860,n869);
nand (n877,n846,n858);
nand (n878,n879,n881);
or (n879,n820,n880);
nand (n880,n834,n843);
nand (n881,n821,n832);
nand (n882,n883,n885);
or (n883,n674,n884);
nand (n884,n748,n758);
nand (n885,n675,n746);
or (n886,n671,n3);
xor (n887,n888,n1349);
xor (n888,n668,n889);
wire s0n889,s1n889,notn889;
or (n889,s0n889,s1n889);
not(notn889,n8);
and (s0n889,notn889,n890);
and (s1n889,n8,n10);
xor (n890,n891,n1288);
xor (n891,n892,n1347);
xor (n892,n893,n1283);
xor (n893,n894,n1340);
xor (n894,n895,n1277);
xor (n895,n896,n1328);
xor (n896,n897,n1271);
xor (n897,n898,n1311);
xor (n898,n899,n1265);
xor (n899,n900,n1289);
xor (n900,n901,n1259);
xor (n901,n902,n1256);
xor (n902,n903,n1255);
xor (n903,n904,n1219);
xor (n904,n905,n1218);
xor (n905,n906,n1173);
xor (n906,n907,n1172);
xor (n907,n908,n1124);
xor (n908,n909,n1123);
xor (n909,n910,n1072);
xor (n910,n911,n1071);
xor (n911,n912,n1022);
xor (n912,n913,n1021);
xor (n913,n914,n970);
xor (n914,n915,n969);
xor (n915,n916,n919);
xor (n916,n917,n918);
and (n917,n296,n91);
and (n918,n290,n39);
or (n919,n920,n923);
and (n920,n921,n922);
and (n921,n290,n91);
and (n922,n309,n39);
and (n923,n924,n925);
xor (n924,n921,n922);
or (n925,n926,n929);
and (n926,n927,n928);
and (n927,n309,n91);
and (n928,n303,n39);
and (n929,n930,n931);
xor (n930,n927,n928);
or (n931,n932,n935);
and (n932,n933,n934);
and (n933,n303,n91);
and (n934,n280,n39);
and (n935,n936,n937);
xor (n936,n933,n934);
or (n937,n938,n941);
and (n938,n939,n940);
and (n939,n280,n91);
and (n940,n274,n39);
and (n941,n942,n943);
xor (n942,n939,n940);
or (n943,n944,n947);
and (n944,n945,n946);
and (n945,n274,n91);
and (n946,n257,n39);
and (n947,n948,n949);
xor (n948,n945,n946);
or (n949,n950,n953);
and (n950,n951,n952);
and (n951,n257,n91);
and (n952,n243,n39);
and (n953,n954,n955);
xor (n954,n951,n952);
or (n955,n956,n958);
and (n956,n957,n131);
and (n957,n243,n91);
and (n958,n959,n960);
xor (n959,n957,n131);
or (n960,n961,n964);
and (n961,n962,n963);
and (n962,n132,n91);
and (n963,n102,n39);
and (n964,n965,n966);
xor (n965,n962,n963);
or (n966,n967,n968);
and (n967,n687,n688);
and (n968,n686,n689);
and (n969,n309,n32);
or (n970,n971,n974);
and (n971,n972,n973);
xor (n972,n924,n925);
and (n973,n303,n32);
and (n974,n975,n976);
xor (n975,n972,n973);
or (n976,n977,n980);
and (n977,n978,n979);
xor (n978,n930,n931);
and (n979,n280,n32);
and (n980,n981,n982);
xor (n981,n978,n979);
or (n982,n983,n986);
and (n983,n984,n985);
xor (n984,n936,n937);
and (n985,n274,n32);
and (n986,n987,n988);
xor (n987,n984,n985);
or (n988,n989,n992);
and (n989,n990,n991);
xor (n990,n942,n943);
and (n991,n257,n32);
and (n992,n993,n994);
xor (n993,n990,n991);
or (n994,n995,n998);
and (n995,n996,n997);
xor (n996,n948,n949);
and (n997,n243,n32);
and (n998,n999,n1000);
xor (n999,n996,n997);
or (n1000,n1001,n1004);
and (n1001,n1002,n1003);
xor (n1002,n954,n955);
and (n1003,n132,n32);
and (n1004,n1005,n1006);
xor (n1005,n1002,n1003);
or (n1006,n1007,n1010);
and (n1007,n1008,n1009);
xor (n1008,n959,n960);
and (n1009,n102,n32);
and (n1010,n1011,n1012);
xor (n1011,n1008,n1009);
or (n1012,n1013,n1016);
and (n1013,n1014,n1015);
xor (n1014,n965,n966);
and (n1015,n96,n32);
and (n1016,n1017,n1018);
xor (n1017,n1014,n1015);
or (n1018,n1019,n1020);
and (n1019,n685,n709);
and (n1020,n684,n710);
and (n1021,n303,n23);
or (n1022,n1023,n1026);
and (n1023,n1024,n1025);
xor (n1024,n975,n976);
and (n1025,n280,n23);
and (n1026,n1027,n1028);
xor (n1027,n1024,n1025);
or (n1028,n1029,n1032);
and (n1029,n1030,n1031);
xor (n1030,n981,n982);
and (n1031,n274,n23);
and (n1032,n1033,n1034);
xor (n1033,n1030,n1031);
or (n1034,n1035,n1038);
and (n1035,n1036,n1037);
xor (n1036,n987,n988);
and (n1037,n257,n23);
and (n1038,n1039,n1040);
xor (n1039,n1036,n1037);
or (n1040,n1041,n1044);
and (n1041,n1042,n1043);
xor (n1042,n993,n994);
and (n1043,n243,n23);
and (n1044,n1045,n1046);
xor (n1045,n1042,n1043);
or (n1046,n1047,n1050);
and (n1047,n1048,n1049);
xor (n1048,n999,n1000);
and (n1049,n132,n23);
and (n1050,n1051,n1052);
xor (n1051,n1048,n1049);
or (n1052,n1053,n1055);
and (n1053,n1054,n546);
xor (n1054,n1005,n1006);
and (n1055,n1056,n1057);
xor (n1056,n1054,n546);
or (n1057,n1058,n1061);
and (n1058,n1059,n1060);
xor (n1059,n1011,n1012);
and (n1060,n96,n23);
and (n1061,n1062,n1063);
xor (n1062,n1059,n1060);
or (n1063,n1064,n1066);
and (n1064,n1065,n45);
xor (n1065,n1017,n1018);
and (n1066,n1067,n1068);
xor (n1067,n1065,n45);
or (n1068,n1069,n1070);
and (n1069,n683,n26);
and (n1070,n682,n724);
and (n1071,n280,n65);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1027,n1028);
and (n1075,n274,n65);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1033,n1034);
and (n1081,n257,n65);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
xor (n1086,n1039,n1040);
and (n1087,n243,n65);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
xor (n1092,n1045,n1046);
and (n1093,n132,n65);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
or (n1096,n1097,n1100);
and (n1097,n1098,n1099);
xor (n1098,n1051,n1052);
and (n1099,n102,n65);
and (n1100,n1101,n1102);
xor (n1101,n1098,n1099);
or (n1102,n1103,n1106);
and (n1103,n1104,n1105);
xor (n1104,n1056,n1057);
and (n1105,n96,n65);
and (n1106,n1107,n1108);
xor (n1107,n1104,n1105);
or (n1108,n1109,n1112);
and (n1109,n1110,n1111);
xor (n1110,n1062,n1063);
and (n1111,n46,n65);
and (n1112,n1113,n1114);
xor (n1113,n1110,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
xor (n1116,n1067,n1068);
and (n1117,n21,n65);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1122);
and (n1121,n681,n732);
and (n1122,n680,n733);
and (n1123,n274,n55);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1077,n1078);
and (n1127,n257,n55);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1083,n1084);
and (n1133,n243,n55);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1089,n1090);
and (n1139,n132,n55);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1095,n1096);
and (n1145,n102,n55);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1101,n1102);
and (n1151,n96,n55);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1107,n1108);
and (n1157,n46,n55);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1113,n1114);
and (n1163,n21,n55);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1169);
and (n1167,n1168,n53);
xor (n1168,n1119,n1120);
and (n1169,n1170,n1171);
xor (n1170,n1168,n53);
and (n1171,n679,n735);
and (n1172,n257,n123);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1129,n1130);
and (n1176,n243,n123);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1135,n1136);
and (n1182,n132,n123);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1141,n1142);
and (n1188,n102,n123);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1147,n1148);
and (n1194,n96,n123);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1153,n1154);
and (n1200,n46,n123);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1159,n1160);
and (n1206,n21,n123);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1165,n1166);
and (n1212,n54,n123);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
and (n1215,n1216,n1217);
xor (n1216,n1170,n1171);
not (n1217,n587);
and (n1218,n243,n245);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1178,n1179);
and (n1222,n132,n245);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1228);
and (n1226,n1227,n369);
xor (n1227,n1184,n1185);
and (n1228,n1229,n1230);
xor (n1229,n1227,n369);
or (n1230,n1231,n1233);
and (n1231,n1232,n415);
xor (n1232,n1190,n1191);
and (n1233,n1234,n1235);
xor (n1234,n1232,n415);
or (n1235,n1236,n1238);
and (n1236,n1237,n468);
xor (n1237,n1196,n1197);
and (n1238,n1239,n1240);
xor (n1239,n1237,n468);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1202,n1203);
and (n1243,n21,n245);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1208,n1209);
and (n1249,n54,n245);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
and (n1252,n1253,n1254);
xor (n1253,n1214,n1215);
and (n1254,n77,n245);
and (n1255,n132,n263);
or (n1256,n1257,n1260);
and (n1257,n1258,n1259);
xor (n1258,n1224,n1225);
and (n1259,n102,n263);
and (n1260,n1261,n1262);
xor (n1261,n1258,n1259);
or (n1262,n1263,n1266);
and (n1263,n1264,n1265);
xor (n1264,n1229,n1230);
and (n1265,n96,n263);
and (n1266,n1267,n1268);
xor (n1267,n1264,n1265);
or (n1268,n1269,n1272);
and (n1269,n1270,n1271);
xor (n1270,n1234,n1235);
and (n1271,n46,n263);
and (n1272,n1273,n1274);
xor (n1273,n1270,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1239,n1240);
and (n1277,n21,n263);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1245,n1246);
and (n1283,n54,n263);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
and (n1286,n1287,n1288);
xor (n1287,n1251,n1252);
and (n1288,n77,n263);
or (n1289,n1290,n1292);
and (n1290,n1291,n1265);
xor (n1291,n1261,n1262);
and (n1292,n1293,n1294);
xor (n1293,n1291,n1265);
or (n1294,n1295,n1297);
and (n1295,n1296,n1271);
xor (n1296,n1267,n1268);
and (n1297,n1298,n1299);
xor (n1298,n1296,n1271);
or (n1299,n1300,n1302);
and (n1300,n1301,n1277);
xor (n1301,n1273,n1274);
and (n1302,n1303,n1304);
xor (n1303,n1301,n1277);
or (n1304,n1305,n1307);
and (n1305,n1306,n1283);
xor (n1306,n1279,n1280);
and (n1307,n1308,n1309);
xor (n1308,n1306,n1283);
and (n1309,n1310,n1288);
xor (n1310,n1285,n1286);
or (n1311,n1312,n1314);
and (n1312,n1313,n1271);
xor (n1313,n1293,n1294);
and (n1314,n1315,n1316);
xor (n1315,n1313,n1271);
or (n1316,n1317,n1319);
and (n1317,n1318,n1277);
xor (n1318,n1298,n1299);
and (n1319,n1320,n1321);
xor (n1320,n1318,n1277);
or (n1321,n1322,n1324);
and (n1322,n1323,n1283);
xor (n1323,n1303,n1304);
and (n1324,n1325,n1326);
xor (n1325,n1323,n1283);
and (n1326,n1327,n1288);
xor (n1327,n1308,n1309);
or (n1328,n1329,n1331);
and (n1329,n1330,n1277);
xor (n1330,n1315,n1316);
and (n1331,n1332,n1333);
xor (n1332,n1330,n1277);
or (n1333,n1334,n1336);
and (n1334,n1335,n1283);
xor (n1335,n1320,n1321);
and (n1336,n1337,n1338);
xor (n1337,n1335,n1283);
and (n1338,n1339,n1288);
xor (n1339,n1325,n1326);
or (n1340,n1341,n1343);
and (n1341,n1342,n1283);
xor (n1342,n1332,n1333);
and (n1343,n1344,n1345);
xor (n1344,n1342,n1283);
and (n1345,n1346,n1288);
xor (n1346,n1337,n1338);
and (n1347,n1348,n1288);
xor (n1348,n1344,n1345);
or (n1349,n1350,n1353,n1384);
and (n1350,n746,n1351);
wire s0n1351,s1n1351,notn1351;
or (n1351,s0n1351,s1n1351);
not(notn1351,n8);
and (s0n1351,notn1351,n1352);
and (s1n1351,n8,n678);
xor (n1352,n1348,n1288);
and (n1353,n1351,n1354);
or (n1354,n1355,n1358,n1383);
and (n1355,n758,n1356);
wire s0n1356,s1n1356,notn1356;
or (n1356,s0n1356,s1n1356);
not(notn1356,n8);
and (s0n1356,notn1356,n1357);
and (s1n1356,n8,n751);
xor (n1357,n1346,n1288);
and (n1358,n1356,n1359);
or (n1359,n1360,n1363,n1382);
and (n1360,n832,n1361);
wire s0n1361,s1n1361,notn1361;
or (n1361,s0n1361,s1n1361);
not(notn1361,n8);
and (s0n1361,notn1361,n1362);
and (s1n1361,n8,n795);
xor (n1362,n1339,n1288);
and (n1363,n1361,n1364);
or (n1364,n1365,n1368,n1381);
and (n1365,n843,n1366);
wire s0n1366,s1n1366,notn1366;
or (n1366,s0n1366,s1n1366);
not(notn1366,n8);
and (s0n1366,notn1366,n1367);
and (s1n1366,n8,n801);
xor (n1367,n1327,n1288);
and (n1368,n1366,n1369);
or (n1369,n1370,n1373,n1380);
and (n1370,n858,n1371);
wire s0n1371,s1n1371,notn1371;
or (n1371,s0n1371,s1n1371);
not(notn1371,n8);
and (s0n1371,notn1371,n1372);
and (s1n1371,n8,n807);
xor (n1372,n1310,n1288);
and (n1373,n1371,n1374);
or (n1374,n1375,n1378,n1379);
and (n1375,n869,n1376);
wire s0n1376,s1n1376,notn1376;
or (n1376,s0n1376,s1n1376);
not(notn1376,n8);
and (s0n1376,notn1376,n1377);
and (s1n1376,n8,n207);
xor (n1377,n1287,n1288);
and (n1378,n1376,n763);
and (n1379,n869,n763);
and (n1380,n858,n1374);
and (n1381,n843,n1369);
and (n1382,n832,n1364);
and (n1383,n758,n1359);
and (n1384,n746,n1354);
endmodule
