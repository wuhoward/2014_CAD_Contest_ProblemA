module top (out,n4,n20,n22,n23,n32,n33,n35,n36,n46
        ,n55,n59,n69,n70,n72,n73,n80,n86,n98,n99
        ,n101,n102,n105,n111,n123,n124,n133,n138,n166,n205
        ,n284,n290,n299,n309,n315,n1024);
output out;
input n4;
input n20;
input n22;
input n23;
input n32;
input n33;
input n35;
input n36;
input n46;
input n55;
input n59;
input n69;
input n70;
input n72;
input n73;
input n80;
input n86;
input n98;
input n99;
input n101;
input n102;
input n105;
input n111;
input n123;
input n124;
input n133;
input n138;
input n166;
input n205;
input n284;
input n290;
input n299;
input n309;
input n315;
input n1024;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n71;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
xnor (out,n0,n1025);
nand (n0,n1,n1024);
nand (n1,n2,n765);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
xor (n6,n7,n263);
and (n7,n8,n261);
not (n8,n9);
nor (n9,n10,n216);
or (n10,n11,n215);
and (n11,n12,n175);
xor (n12,n13,n89);
xor (n13,n14,n61);
xor (n14,n15,n49);
nand (n15,n16,n42);
or (n16,n17,n27);
not (n17,n18);
nor (n18,n19,n24);
and (n19,n20,n21);
wire s0n21,s1n21,notn21;
or (n21,s0n21,s1n21);
not(notn21,n4);
and (s0n21,notn21,n22);
and (s1n21,n4,n23);
and (n24,n25,n26);
not (n25,n20);
not (n26,n21);
nand (n27,n28,n39);
nor (n28,n29,n37);
and (n29,n30,n34);
not (n30,n31);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n4);
and (s0n31,notn31,n32);
and (s1n31,n4,n33);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n4);
and (s0n34,notn34,n35);
and (s1n34,n4,n36);
and (n37,n31,n38);
not (n38,n34);
nand (n39,n40,n41);
or (n40,n30,n21);
nand (n41,n21,n30);
nand (n42,n43,n44);
not (n43,n28);
nor (n44,n45,n47);
and (n45,n46,n21);
and (n47,n48,n26);
not (n48,n46);
nor (n49,n50,n56);
nand (n50,n21,n51);
not (n51,n52);
wire s0n52,s1n52,notn52;
or (n52,s0n52,s1n52);
not(notn52,n4);
and (s0n52,notn52,1'b0);
and (s1n52,n4,n54);
and (n54,n55,n23);
nor (n56,n57,n60);
and (n57,n52,n58);
not (n58,n59);
and (n60,n51,n59);
nand (n61,n62,n83);
or (n62,n63,n78);
nand (n63,n64,n75);
not (n64,n65);
nand (n65,n66,n74);
or (n66,n67,n71);
not (n67,n68);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n4);
and (s0n68,notn68,n69);
and (s1n68,n4,n70);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n4);
and (s0n71,notn71,n72);
and (s1n71,n4,n73);
nand (n74,n71,n67);
nand (n75,n76,n77);
or (n76,n67,n34);
nand (n77,n34,n67);
nor (n78,n79,n81);
and (n79,n38,n80);
and (n81,n34,n82);
not (n82,n80);
or (n83,n64,n84);
nor (n84,n85,n87);
and (n85,n38,n86);
and (n87,n34,n88);
not (n88,n86);
xor (n89,n90,n153);
xor (n90,n91,n139);
xor (n91,n92,n115);
nand (n92,n93,n108);
or (n93,n94,n103);
not (n94,n95);
nor (n95,n96,n100);
not (n96,n97);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n4);
and (s0n97,notn97,n98);
and (s1n97,n4,n99);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n4);
and (s0n100,notn100,n101);
and (s1n100,n4,n102);
nor (n103,n104,n106);
and (n104,n96,n105);
and (n106,n97,n107);
not (n107,n105);
or (n108,n109,n114);
nor (n109,n110,n112);
and (n110,n96,n111);
and (n112,n97,n113);
not (n113,n111);
not (n114,n100);
nand (n115,n116,n136);
or (n116,n117,n130);
not (n117,n118);
and (n118,n119,n126);
nand (n119,n120,n125);
or (n120,n121,n71);
not (n121,n122);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n4);
and (s0n122,notn122,n123);
and (s1n122,n4,n124);
nand (n125,n71,n121);
not (n126,n127);
nand (n127,n128,n129);
or (n128,n121,n97);
nand (n129,n97,n121);
nor (n130,n131,n134);
and (n131,n132,n133);
not (n132,n71);
and (n134,n71,n135);
not (n135,n133);
or (n136,n137,n126);
xor (n137,n138,n132);
and (n139,n140,n147);
nand (n140,n141,n146);
or (n141,n94,n142);
nor (n142,n143,n144);
and (n143,n96,n138);
and (n144,n97,n145);
not (n145,n138);
or (n146,n103,n114);
nand (n147,n148,n152);
or (n148,n117,n149);
nor (n149,n150,n151);
and (n150,n132,n86);
and (n151,n71,n88);
or (n152,n126,n130);
or (n153,n154,n174);
and (n154,n155,n168);
xor (n155,n156,n162);
nand (n156,n157,n161);
or (n157,n158,n27);
nor (n158,n159,n160);
and (n159,n59,n26);
and (n160,n58,n21);
nand (n161,n43,n18);
nor (n162,n50,n163);
nor (n163,n164,n167);
and (n164,n52,n165);
not (n165,n166);
and (n167,n51,n166);
nand (n168,n169,n173);
or (n169,n63,n170);
nor (n170,n171,n172);
and (n171,n38,n46);
and (n172,n34,n48);
or (n173,n64,n78);
and (n174,n156,n162);
or (n175,n176,n214);
and (n176,n177,n192);
xor (n177,n178,n179);
xor (n178,n140,n147);
and (n179,n180,n186);
nand (n180,n181,n185);
or (n181,n94,n182);
nor (n182,n183,n184);
and (n183,n96,n133);
and (n184,n97,n135);
or (n185,n142,n114);
nand (n186,n187,n191);
or (n187,n117,n188);
nor (n188,n189,n190);
and (n189,n132,n80);
and (n190,n71,n82);
or (n191,n149,n126);
or (n192,n193,n213);
and (n193,n194,n207);
xor (n194,n195,n201);
nand (n195,n196,n200);
or (n196,n27,n197);
nor (n197,n198,n199);
and (n198,n26,n166);
and (n199,n21,n165);
or (n200,n28,n158);
nor (n201,n50,n202);
nor (n202,n203,n206);
and (n203,n52,n204);
not (n204,n205);
and (n206,n51,n205);
nand (n207,n208,n209);
or (n208,n170,n64);
or (n209,n63,n210);
nor (n210,n211,n212);
and (n211,n38,n20);
and (n212,n34,n25);
and (n213,n195,n201);
and (n214,n178,n179);
and (n215,n13,n89);
xor (n216,n217,n258);
xor (n217,n218,n237);
xor (n218,n219,n231);
xor (n219,n220,n227);
nand (n220,n221,n223);
or (n221,n222,n27);
not (n222,n44);
or (n223,n28,n224);
nor (n224,n225,n226);
and (n225,n26,n80);
and (n226,n21,n82);
nor (n227,n50,n228);
nor (n228,n229,n230);
and (n229,n52,n25);
and (n230,n51,n20);
nand (n231,n232,n233);
or (n232,n63,n84);
or (n233,n64,n234);
nor (n234,n235,n236);
and (n235,n38,n133);
and (n236,n34,n135);
xor (n237,n238,n255);
xor (n238,n239,n254);
xor (n239,n240,n248);
nand (n240,n241,n242);
or (n241,n94,n109);
or (n242,n243,n114);
nor (n243,n244,n246);
and (n244,n96,n245);
and (n245,n55,n111);
and (n246,n97,n247);
not (n247,n245);
nand (n248,n249,n250);
or (n249,n137,n117);
nand (n250,n127,n251);
nand (n251,n252,n253);
or (n252,n71,n107);
or (n253,n132,n105);
and (n254,n92,n115);
or (n255,n256,n257);
and (n256,n14,n61);
and (n257,n15,n49);
or (n258,n259,n260);
and (n259,n90,n153);
and (n260,n91,n139);
not (n261,n262);
and (n262,n10,n216);
nand (n263,n264,n754,n764);
nand (n264,n265,n675);
nand (n265,n266,n530,n674);
nand (n266,n267,n483);
nand (n267,n268,n482);
or (n268,n269,n437);
nor (n269,n270,n436);
and (n270,n271,n408);
not (n271,n272);
nor (n272,n273,n368);
or (n273,n274,n367);
and (n274,n275,n338);
xor (n275,n276,n319);
or (n276,n277,n318);
and (n277,n278,n305);
xor (n278,n279,n293);
nand (n279,n280,n287);
or (n280,n281,n27);
not (n281,n282);
nand (n282,n283,n285);
or (n283,n26,n284);
or (n285,n21,n286);
not (n286,n284);
or (n287,n28,n288);
nor (n288,n289,n291);
and (n289,n290,n26);
and (n291,n292,n21);
not (n292,n290);
nand (n293,n294,n301);
or (n294,n295,n117);
not (n295,n296);
nand (n296,n297,n300);
or (n297,n71,n298);
not (n298,n299);
or (n300,n132,n299);
nand (n301,n127,n302);
nor (n302,n303,n304);
and (n303,n205,n71);
and (n304,n204,n132);
nand (n305,n306,n312);
or (n306,n63,n307);
nor (n307,n308,n310);
and (n308,n38,n309);
and (n310,n34,n311);
not (n311,n309);
or (n312,n64,n313);
nor (n313,n314,n316);
and (n314,n38,n315);
and (n316,n34,n317);
not (n317,n315);
and (n318,n279,n293);
xor (n319,n320,n332);
xor (n320,n321,n323);
and (n321,n322,n284);
not (n322,n50);
nand (n323,n324,n328);
or (n324,n94,n325);
nor (n325,n326,n327);
and (n326,n58,n97);
and (n327,n59,n96);
or (n328,n329,n114);
nor (n329,n330,n331);
and (n330,n96,n20);
and (n331,n97,n25);
nand (n332,n333,n334);
or (n333,n27,n288);
or (n334,n28,n335);
nor (n335,n336,n337);
and (n336,n309,n26);
and (n337,n311,n21);
xor (n338,n339,n353);
xor (n339,n340,n347);
nand (n340,n341,n343);
or (n341,n117,n342);
not (n342,n302);
or (n343,n126,n344);
nor (n344,n345,n346);
and (n345,n132,n166);
and (n346,n71,n165);
nand (n347,n348,n349);
or (n348,n63,n313);
or (n349,n64,n350);
nor (n350,n351,n352);
and (n351,n38,n299);
and (n352,n34,n298);
and (n353,n354,n359);
nor (n354,n355,n26);
nor (n355,n356,n358);
and (n356,n38,n357);
nand (n357,n31,n284);
and (n358,n30,n286);
nand (n359,n360,n365);
or (n360,n361,n94);
not (n361,n362);
nor (n362,n363,n364);
and (n363,n166,n97);
and (n364,n165,n96);
nand (n365,n366,n100);
not (n366,n325);
and (n367,n276,n319);
xor (n368,n369,n391);
xor (n369,n370,n388);
xor (n370,n371,n382);
xor (n371,n372,n378);
nand (n372,n373,n374);
or (n373,n335,n27);
nand (n374,n375,n43);
nor (n375,n376,n377);
and (n376,n315,n21);
and (n377,n317,n26);
nor (n378,n50,n379);
nor (n379,n380,n381);
and (n380,n52,n292);
and (n381,n51,n290);
nand (n382,n383,n384);
or (n383,n94,n329);
or (n384,n385,n114);
nor (n385,n386,n387);
and (n386,n96,n46);
and (n387,n97,n48);
or (n388,n389,n390);
and (n389,n339,n353);
and (n390,n340,n347);
xor (n391,n392,n405);
xor (n392,n393,n399);
nand (n393,n394,n395);
or (n394,n63,n350);
or (n395,n64,n396);
nor (n396,n397,n398);
and (n397,n38,n205);
and (n398,n34,n204);
nand (n399,n400,n401);
or (n400,n117,n344);
or (n401,n402,n126);
nor (n402,n403,n404);
and (n403,n132,n59);
and (n404,n71,n58);
or (n405,n406,n407);
and (n406,n320,n332);
and (n407,n321,n323);
not (n408,n409);
nand (n409,n410,n411);
xor (n410,n275,n338);
or (n411,n412,n435);
and (n412,n413,n434);
xor (n413,n414,n415);
xor (n414,n354,n359);
or (n415,n416,n433);
and (n416,n417,n426);
xor (n417,n418,n419);
and (n418,n43,n284);
nand (n419,n420,n421);
or (n420,n114,n361);
nand (n421,n422,n95);
not (n422,n423);
nor (n423,n424,n425);
and (n424,n205,n96);
and (n425,n204,n97);
nand (n426,n427,n432);
or (n427,n428,n117);
not (n428,n429);
nor (n429,n430,n431);
and (n430,n315,n71);
and (n431,n132,n317);
nand (n432,n127,n296);
and (n433,n418,n419);
xor (n434,n278,n305);
and (n435,n414,n415);
and (n436,n273,n368);
nor (n437,n438,n479);
xor (n438,n439,n476);
xor (n439,n440,n459);
xor (n440,n441,n453);
xor (n441,n442,n449);
nand (n442,n443,n445);
or (n443,n444,n27);
not (n444,n375);
nand (n445,n43,n446);
nor (n446,n447,n448);
and (n447,n299,n21);
and (n448,n298,n26);
nor (n449,n50,n450);
nor (n450,n451,n452);
and (n451,n52,n311);
and (n452,n51,n309);
nand (n453,n454,n455);
or (n454,n63,n396);
or (n455,n64,n456);
nor (n456,n457,n458);
and (n457,n38,n166);
and (n458,n34,n165);
xor (n459,n460,n473);
xor (n460,n461,n467);
nand (n461,n462,n463);
or (n462,n94,n385);
or (n463,n464,n114);
nor (n464,n465,n466);
and (n465,n96,n80);
and (n466,n97,n82);
nand (n467,n468,n469);
or (n468,n117,n402);
or (n469,n470,n126);
nor (n470,n471,n472);
and (n471,n132,n20);
and (n472,n71,n25);
or (n473,n474,n475);
and (n474,n371,n382);
and (n475,n372,n378);
or (n476,n477,n478);
and (n477,n392,n405);
and (n478,n393,n399);
or (n479,n480,n481);
and (n480,n369,n391);
and (n481,n370,n388);
nand (n482,n438,n479);
nand (n483,n484,n526);
not (n484,n485);
xor (n485,n486,n525);
xor (n486,n487,n506);
xor (n487,n488,n500);
xor (n488,n489,n496);
nand (n489,n490,n492);
or (n490,n491,n27);
not (n491,n446);
nand (n492,n43,n493);
nor (n493,n494,n495);
and (n494,n205,n21);
and (n495,n204,n26);
nor (n496,n50,n497);
nor (n497,n498,n499);
and (n498,n52,n317);
and (n499,n51,n315);
nand (n500,n501,n502);
or (n501,n63,n456);
or (n502,n64,n503);
nor (n503,n504,n505);
and (n504,n38,n59);
and (n505,n34,n58);
xor (n506,n507,n522);
xor (n507,n508,n521);
xor (n508,n509,n515);
nand (n509,n510,n511);
or (n510,n94,n464);
or (n511,n512,n114);
nor (n512,n513,n514);
and (n513,n96,n86);
and (n514,n97,n88);
nand (n515,n516,n517);
or (n516,n117,n470);
or (n517,n126,n518);
nor (n518,n519,n520);
and (n519,n132,n46);
and (n520,n71,n48);
and (n521,n461,n467);
or (n522,n523,n524);
and (n523,n441,n453);
and (n524,n442,n449);
and (n525,n460,n473);
not (n526,n527);
or (n527,n528,n529);
and (n528,n439,n476);
and (n529,n440,n459);
nand (n530,n483,n531,n673);
nor (n531,n532,n670);
nor (n532,n533,n668);
and (n533,n534,n663);
or (n534,n535,n662);
and (n535,n536,n578);
xor (n536,n537,n571);
or (n537,n538,n570);
and (n538,n539,n558);
xor (n539,n540,n547);
nand (n540,n541,n546);
or (n541,n542,n117);
not (n542,n543);
nor (n543,n544,n545);
and (n544,n311,n132);
and (n545,n309,n71);
nand (n546,n127,n429);
nand (n547,n548,n553);
or (n548,n549,n64);
not (n549,n550);
nor (n550,n551,n552);
and (n551,n290,n34);
and (n552,n292,n38);
nand (n553,n554,n555);
not (n554,n63);
nand (n555,n556,n557);
or (n556,n38,n284);
or (n557,n34,n286);
xor (n558,n559,n564);
and (n559,n560,n34);
nand (n560,n561,n563);
or (n561,n71,n562);
and (n562,n284,n68);
or (n563,n68,n284);
nand (n564,n565,n569);
or (n565,n94,n566);
nor (n566,n567,n568);
and (n567,n96,n299);
and (n568,n97,n298);
or (n569,n423,n114);
and (n570,n540,n547);
xor (n571,n572,n577);
xor (n572,n573,n576);
nand (n573,n574,n575);
or (n574,n549,n63);
or (n575,n64,n307);
and (n576,n559,n564);
xor (n577,n417,n426);
or (n578,n579,n661);
and (n579,n580,n601);
xor (n580,n581,n600);
or (n581,n582,n599);
and (n582,n583,n592);
xor (n583,n584,n585);
and (n584,n65,n284);
nand (n585,n586,n591);
or (n586,n587,n117);
not (n587,n588);
nor (n588,n589,n590);
and (n589,n290,n71);
and (n590,n292,n132);
nand (n591,n543,n127);
nand (n592,n593,n598);
or (n593,n94,n594);
not (n594,n595);
nor (n595,n596,n597);
and (n596,n317,n96);
and (n597,n315,n97);
or (n598,n566,n114);
and (n599,n584,n585);
xor (n600,n539,n558);
or (n601,n602,n660);
and (n602,n603,n659);
xor (n603,n604,n618);
nor (n604,n605,n613);
not (n605,n606);
nand (n606,n607,n612);
or (n607,n608,n94);
not (n608,n609);
nand (n609,n610,n611);
or (n610,n311,n97);
nand (n611,n97,n311);
nand (n612,n595,n100);
nand (n613,n614,n71);
nand (n614,n615,n617);
or (n615,n97,n616);
and (n616,n284,n122);
or (n617,n122,n284);
nand (n618,n619,n657);
or (n619,n620,n643);
not (n620,n621);
nand (n621,n622,n642);
or (n622,n623,n632);
nor (n623,n624,n631);
nand (n624,n625,n630);
or (n625,n626,n94);
not (n626,n627);
nand (n627,n628,n629);
or (n628,n292,n97);
nand (n629,n97,n292);
nand (n630,n609,n100);
nor (n631,n126,n286);
nand (n632,n633,n640);
nand (n633,n634,n639);
or (n634,n635,n94);
not (n635,n636);
nand (n636,n637,n638);
or (n637,n96,n284);
or (n638,n97,n286);
nand (n639,n627,n100);
nor (n640,n641,n96);
and (n641,n284,n100);
nand (n642,n624,n631);
not (n643,n644);
nand (n644,n645,n653);
not (n645,n646);
nand (n646,n647,n652);
or (n647,n648,n117);
not (n648,n649);
nand (n649,n650,n651);
or (n650,n132,n284);
or (n651,n71,n286);
nand (n652,n127,n588);
nor (n653,n654,n656);
and (n654,n605,n655);
not (n655,n613);
and (n656,n606,n613);
nand (n657,n658,n646);
not (n658,n653);
xor (n659,n583,n592);
and (n660,n604,n618);
and (n661,n581,n600);
and (n662,n537,n571);
or (n663,n664,n665);
xor (n664,n413,n434);
or (n665,n666,n667);
and (n666,n572,n577);
and (n667,n573,n576);
not (n668,n669);
nand (n669,n664,n665);
nand (n670,n671,n271);
not (n671,n672);
nor (n672,n410,n411);
not (n673,n437);
nand (n674,n485,n527);
nor (n675,n676,n733);
nand (n676,n677,n726);
not (n677,n678);
nor (n678,n679,n717);
xor (n679,n680,n708);
xor (n680,n681,n682);
xor (n681,n194,n207);
xor (n682,n683,n692);
xor (n683,n684,n685);
xor (n684,n180,n186);
and (n685,n686,n689);
nand (n686,n687,n688);
or (n687,n94,n512);
or (n688,n182,n114);
nand (n689,n690,n691);
or (n690,n117,n518);
or (n691,n188,n126);
or (n692,n693,n707);
and (n693,n694,n704);
xor (n694,n695,n700);
nand (n695,n696,n698);
or (n696,n697,n27);
not (n697,n493);
nand (n698,n699,n43);
not (n699,n197);
nor (n700,n50,n701);
nor (n701,n702,n703);
and (n702,n52,n298);
and (n703,n51,n299);
nand (n704,n705,n706);
or (n705,n63,n503);
or (n706,n64,n210);
and (n707,n695,n700);
or (n708,n709,n716);
and (n709,n710,n713);
xor (n710,n711,n712);
xor (n711,n686,n689);
and (n712,n509,n515);
or (n713,n714,n715);
and (n714,n488,n500);
and (n715,n489,n496);
and (n716,n711,n712);
or (n717,n718,n725);
and (n718,n719,n722);
xor (n719,n720,n721);
xor (n720,n694,n704);
xor (n721,n710,n713);
or (n722,n723,n724);
and (n723,n507,n522);
and (n724,n508,n521);
and (n725,n720,n721);
nand (n726,n727,n729);
not (n727,n728);
xor (n728,n719,n722);
not (n729,n730);
or (n730,n731,n732);
and (n731,n486,n525);
and (n732,n487,n506);
nand (n733,n734,n747);
nand (n734,n735,n743);
not (n735,n736);
xor (n736,n737,n740);
xor (n737,n738,n739);
xor (n738,n155,n168);
xor (n739,n177,n192);
or (n740,n741,n742);
and (n741,n683,n692);
and (n742,n684,n685);
not (n743,n744);
or (n744,n745,n746);
and (n745,n680,n708);
and (n746,n681,n682);
nand (n747,n748,n750);
not (n748,n749);
xor (n749,n12,n175);
not (n750,n751);
or (n751,n752,n753);
and (n752,n737,n740);
and (n753,n738,n739);
nand (n754,n755,n747);
nand (n755,n756,n763);
or (n756,n757,n758);
not (n757,n734);
not (n758,n759);
nand (n759,n760,n762);
or (n760,n678,n761);
nand (n761,n728,n730);
nand (n762,n679,n717);
nand (n763,n736,n744);
nand (n764,n751,n749);
not (n765,n766);
and (n766,n767,n3,n55);
nand (n767,n768,n1023);
or (n768,n769,n822);
not (n769,n770);
nor (n770,n771,n821);
and (n771,n772,n810);
not (n772,n773);
or (n773,n774,n809);
and (n774,n775,n790);
xor (n775,n776,n786);
nand (n776,n777,n782);
or (n777,n778,n28);
not (n778,n779);
nand (n779,n780,n781);
or (n780,n21,n247);
or (n781,n26,n245);
or (n782,n27,n783);
nor (n783,n784,n785);
and (n784,n26,n111);
and (n785,n21,n113);
nand (n786,n787,n788,n322);
or (n787,n52,n105);
not (n788,n789);
and (n789,n105,n52);
or (n790,n791,n808);
and (n791,n792,n804);
xor (n792,n793,n798);
nand (n793,n794,n795);
or (n794,n554,n65);
nand (n795,n796,n797);
or (n796,n34,n247);
or (n797,n38,n245);
nand (n798,n799,n803);
or (n799,n27,n800);
nor (n800,n801,n802);
and (n801,n26,n105);
and (n802,n21,n107);
or (n803,n28,n783);
nor (n804,n50,n805);
nor (n805,n806,n807);
and (n806,n52,n145);
and (n807,n51,n138);
and (n808,n793,n798);
and (n809,n776,n786);
not (n810,n811);
xor (n811,n812,n820);
xor (n812,n813,n816);
nand (n813,n814,n779);
or (n814,n815,n43);
not (n815,n27);
nor (n816,n50,n817);
nor (n817,n818,n819);
and (n818,n52,n113);
and (n819,n51,n111);
not (n820,n786);
and (n821,n773,n811);
nand (n822,n823,n1000,n1022);
nand (n823,n263,n824);
and (n824,n825,n956,n995);
and (n825,n826,n878,n950);
nor (n826,n9,n827);
not (n827,n828);
nand (n828,n829,n874);
not (n829,n830);
xor (n830,n831,n850);
xor (n831,n832,n847);
xor (n832,n833,n841);
xor (n833,n834,n838);
nor (n834,n50,n835);
nor (n835,n836,n837);
and (n836,n52,n48);
and (n837,n51,n46);
nand (n838,n839,n840);
or (n839,n100,n95);
not (n840,n243);
nand (n841,n842,n846);
or (n842,n843,n64);
nor (n843,n844,n845);
and (n844,n138,n38);
and (n845,n145,n34);
or (n846,n63,n234);
or (n847,n848,n849);
and (n848,n238,n255);
and (n849,n239,n254);
xor (n850,n851,n856);
xor (n851,n852,n853);
and (n852,n240,n248);
or (n853,n854,n855);
and (n854,n219,n231);
and (n855,n220,n227);
nand (n856,n857,n873);
or (n857,n858,n866);
not (n858,n859);
nand (n859,n860,n862);
or (n860,n117,n861);
not (n861,n251);
or (n862,n126,n863);
nor (n863,n864,n865);
and (n864,n132,n111);
and (n865,n71,n113);
not (n866,n867);
nand (n867,n868,n869);
or (n868,n27,n224);
or (n869,n28,n870);
nor (n870,n871,n872);
and (n871,n26,n86);
and (n872,n21,n88);
or (n873,n867,n859);
not (n874,n875);
or (n875,n876,n877);
and (n876,n217,n258);
and (n877,n218,n237);
nand (n878,n879,n940);
not (n879,n880);
xor (n880,n881,n932);
xor (n881,n882,n902);
xor (n882,n883,n898);
xor (n883,n884,n889);
nand (n884,n885,n886);
or (n885,n118,n127);
nand (n886,n887,n888);
or (n887,n71,n247);
or (n888,n132,n245);
nand (n889,n890,n894);
or (n890,n63,n891);
nor (n891,n892,n893);
and (n892,n38,n105);
and (n893,n34,n107);
or (n894,n64,n895);
nor (n895,n896,n897);
and (n896,n38,n111);
and (n897,n34,n113);
nor (n898,n50,n899);
nor (n899,n900,n901);
and (n900,n52,n88);
and (n901,n51,n86);
xor (n902,n903,n918);
xor (n903,n904,n913);
nand (n904,n905,n909);
or (n905,n27,n906);
nor (n906,n907,n908);
and (n907,n26,n133);
and (n908,n21,n135);
or (n909,n28,n910);
nor (n910,n911,n912);
and (n911,n26,n138);
and (n912,n21,n145);
nand (n913,n914,n916);
or (n914,n915,n126);
not (n915,n886);
nand (n916,n917,n118);
not (n917,n863);
or (n918,n919,n931);
and (n919,n920,n928);
xor (n920,n921,n925);
nor (n921,n50,n922);
nor (n922,n923,n924);
and (n923,n52,n82);
and (n924,n51,n80);
nand (n925,n926,n927);
or (n926,n63,n843);
or (n927,n64,n891);
nand (n928,n929,n930);
or (n929,n27,n870);
or (n930,n28,n906);
and (n931,n921,n925);
or (n932,n933,n939);
and (n933,n934,n936);
xor (n934,n935,n873);
not (n935,n913);
or (n936,n937,n938);
and (n937,n833,n841);
and (n938,n834,n838);
and (n939,n935,n873);
not (n940,n941);
or (n941,n942,n949);
and (n942,n943,n946);
xor (n943,n944,n945);
xor (n944,n920,n928);
xor (n945,n934,n936);
or (n946,n947,n948);
and (n947,n851,n856);
and (n948,n852,n853);
and (n949,n944,n945);
not (n950,n951);
nor (n951,n952,n953);
xor (n952,n943,n946);
or (n953,n954,n955);
and (n954,n831,n850);
and (n955,n832,n847);
nor (n956,n957,n982);
nor (n957,n958,n961);
or (n958,n959,n960);
and (n959,n881,n932);
and (n960,n882,n902);
xor (n961,n962,n979);
xor (n962,n963,n966);
or (n963,n964,n965);
and (n964,n883,n898);
and (n965,n884,n889);
xor (n966,n967,n975);
xor (n967,n968,n971);
nand (n968,n969,n970);
or (n969,n27,n910);
or (n970,n28,n800);
nor (n971,n50,n972);
nor (n972,n973,n974);
and (n973,n52,n135);
and (n974,n51,n133);
nor (n975,n976,n978);
and (n976,n554,n977);
not (n977,n895);
and (n978,n65,n795);
or (n979,n980,n981);
and (n980,n903,n918);
and (n981,n904,n913);
and (n982,n983,n987);
not (n983,n984);
or (n984,n985,n986);
and (n985,n962,n979);
and (n986,n963,n966);
not (n987,n988);
xor (n988,n989,n992);
xor (n989,n990,n991);
not (n990,n975);
xor (n991,n792,n804);
or (n992,n993,n994);
and (n993,n967,n975);
and (n994,n968,n971);
or (n995,n996,n999);
or (n996,n997,n998);
and (n997,n989,n992);
and (n998,n990,n991);
xor (n999,n775,n790);
nand (n1000,n1001,n995);
nand (n1001,n1002,n1016);
or (n1002,n1003,n1004);
not (n1003,n956);
not (n1004,n1005);
nand (n1005,n1006,n1015);
or (n1006,n1007,n1008);
not (n1007,n878);
not (n1008,n1009);
nand (n1009,n1010,n1014);
or (n1010,n1011,n951);
nor (n1011,n1012,n1013);
and (n1012,n262,n828);
nor (n1013,n829,n874);
nand (n1014,n952,n953);
or (n1015,n879,n940);
nor (n1016,n1017,n1021);
and (n1017,n1018,n1020);
not (n1018,n1019);
nand (n1019,n958,n961);
not (n1020,n982);
nor (n1021,n983,n987);
nand (n1022,n996,n999);
nand (n1023,n769,n822);
and (n1025,n1024,n1026);
wire s0n1026,s1n1026,notn1026;
or (n1026,s0n1026,s1n1026);
not(notn1026,n4);
and (s0n1026,notn1026,n1027);
and (s1n1026,n4,n2327);
and (n1027,n55,n1028);
xor (n1028,n1029,n1843);
xor (n1029,n1030,n2325);
xor (n1030,n1031,n1838);
xor (n1031,n1032,n2318);
xor (n1032,n1033,n1832);
xor (n1033,n1034,n2306);
xor (n1034,n1035,n1826);
xor (n1035,n1036,n2289);
xor (n1036,n1037,n1820);
xor (n1037,n1038,n2267);
xor (n1038,n1039,n1814);
xor (n1039,n1040,n2240);
xor (n1040,n1041,n1808);
xor (n1041,n1042,n2208);
xor (n1042,n1043,n1802);
xor (n1043,n1044,n2171);
xor (n1044,n1045,n1796);
xor (n1045,n1046,n2129);
xor (n1046,n1047,n1790);
xor (n1047,n1048,n2082);
xor (n1048,n1049,n1784);
xor (n1049,n1050,n2030);
xor (n1050,n1051,n1778);
xor (n1051,n1052,n1973);
xor (n1052,n1053,n1772);
xor (n1053,n1054,n1911);
xor (n1054,n1055,n1766);
xor (n1055,n1056,n1844);
xor (n1056,n1057,n789);
xor (n1057,n1058,n1758);
xor (n1058,n1059,n1757);
xor (n1059,n1060,n1669);
xor (n1060,n1061,n1668);
xor (n1061,n1062,n1570);
xor (n1062,n1063,n1569);
xor (n1063,n1064,n1467);
xor (n1064,n1065,n1466);
xor (n1065,n1066,n1359);
xor (n1066,n1067,n1358);
xor (n1067,n1068,n1079);
xor (n1068,n1069,n1078);
xor (n1069,n1070,n1077);
xor (n1070,n1071,n1076);
xor (n1071,n1072,n1075);
xor (n1072,n1073,n1074);
and (n1073,n245,n100);
and (n1074,n245,n97);
and (n1075,n1073,n1074);
and (n1076,n245,n122);
and (n1077,n1071,n1076);
and (n1078,n245,n71);
or (n1079,n1080,n1081);
and (n1080,n1069,n1078);
and (n1081,n1068,n1082);
or (n1082,n1080,n1083);
and (n1083,n1068,n1084);
or (n1084,n1080,n1085);
and (n1085,n1068,n1086);
or (n1086,n1080,n1087);
and (n1087,n1068,n1088);
or (n1088,n1089,n1273);
and (n1089,n1090,n1272);
xor (n1090,n1070,n1091);
or (n1091,n1092,n1184);
and (n1092,n1093,n1183);
xor (n1093,n1072,n1094);
or (n1094,n1075,n1095);
and (n1095,n1096,n1098);
xor (n1096,n1073,n1097);
and (n1097,n111,n97);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
and (n1100,n111,n100);
and (n1101,n105,n97);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
and (n1106,n105,n100);
and (n1107,n138,n97);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1114);
and (n1111,n1112,n1113);
and (n1112,n138,n100);
and (n1113,n133,n97);
and (n1114,n1115,n1116);
xor (n1115,n1112,n1113);
or (n1116,n1117,n1120);
and (n1117,n1118,n1119);
and (n1118,n133,n100);
and (n1119,n86,n97);
and (n1120,n1121,n1122);
xor (n1121,n1118,n1119);
or (n1122,n1123,n1126);
and (n1123,n1124,n1125);
and (n1124,n86,n100);
and (n1125,n80,n97);
and (n1126,n1127,n1128);
xor (n1127,n1124,n1125);
or (n1128,n1129,n1132);
and (n1129,n1130,n1131);
and (n1130,n80,n100);
and (n1131,n46,n97);
and (n1132,n1133,n1134);
xor (n1133,n1130,n1131);
or (n1134,n1135,n1138);
and (n1135,n1136,n1137);
and (n1136,n46,n100);
and (n1137,n20,n97);
and (n1138,n1139,n1140);
xor (n1139,n1136,n1137);
or (n1140,n1141,n1144);
and (n1141,n1142,n1143);
and (n1142,n20,n100);
and (n1143,n59,n97);
and (n1144,n1145,n1146);
xor (n1145,n1142,n1143);
or (n1146,n1147,n1149);
and (n1147,n1148,n363);
and (n1148,n59,n100);
and (n1149,n1150,n1151);
xor (n1150,n1148,n363);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
and (n1153,n166,n100);
and (n1154,n205,n97);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
and (n1159,n205,n100);
and (n1160,n299,n97);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1166);
and (n1164,n1165,n597);
and (n1165,n299,n100);
and (n1166,n1167,n1168);
xor (n1167,n1165,n597);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
and (n1170,n315,n100);
and (n1171,n309,n97);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
and (n1176,n309,n100);
and (n1177,n290,n97);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
and (n1180,n1181,n1182);
and (n1181,n290,n100);
and (n1182,n284,n97);
and (n1183,n111,n122);
and (n1184,n1185,n1186);
xor (n1185,n1093,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1096,n1098);
and (n1189,n105,n122);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1196);
and (n1193,n1194,n1195);
xor (n1194,n1103,n1104);
and (n1195,n138,n122);
and (n1196,n1197,n1198);
xor (n1197,n1194,n1195);
or (n1198,n1199,n1202);
and (n1199,n1200,n1201);
xor (n1200,n1109,n1110);
and (n1201,n133,n122);
and (n1202,n1203,n1204);
xor (n1203,n1200,n1201);
or (n1204,n1205,n1208);
and (n1205,n1206,n1207);
xor (n1206,n1115,n1116);
and (n1207,n86,n122);
and (n1208,n1209,n1210);
xor (n1209,n1206,n1207);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1121,n1122);
and (n1213,n80,n122);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1220);
and (n1217,n1218,n1219);
xor (n1218,n1127,n1128);
and (n1219,n46,n122);
and (n1220,n1221,n1222);
xor (n1221,n1218,n1219);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1133,n1134);
and (n1225,n20,n122);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1139,n1140);
and (n1231,n59,n122);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1145,n1146);
and (n1237,n166,n122);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1150,n1151);
and (n1243,n205,n122);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1156,n1157);
and (n1249,n299,n122);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1162,n1163);
and (n1255,n315,n122);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1167,n1168);
and (n1261,n309,n122);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1173,n1174);
and (n1267,n290,n122);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
and (n1270,n1271,n616);
xor (n1271,n1179,n1180);
and (n1272,n111,n71);
and (n1273,n1274,n1275);
xor (n1274,n1090,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1185,n1186);
and (n1278,n105,n71);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1191,n1192);
and (n1284,n138,n71);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1197,n1198);
and (n1290,n133,n71);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1203,n1204);
and (n1296,n86,n71);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1209,n1210);
and (n1302,n80,n71);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1215,n1216);
and (n1308,n46,n71);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1221,n1222);
and (n1314,n20,n71);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1227,n1228);
and (n1320,n59,n71);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1233,n1234);
and (n1326,n166,n71);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1332);
and (n1330,n1331,n303);
xor (n1331,n1239,n1240);
and (n1332,n1333,n1334);
xor (n1333,n1331,n303);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1245,n1246);
and (n1337,n299,n71);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
or (n1340,n1341,n1343);
and (n1341,n1342,n430);
xor (n1342,n1251,n1252);
and (n1343,n1344,n1345);
xor (n1344,n1342,n430);
or (n1345,n1346,n1348);
and (n1346,n1347,n545);
xor (n1347,n1257,n1258);
and (n1348,n1349,n1350);
xor (n1349,n1347,n545);
or (n1350,n1351,n1353);
and (n1351,n1352,n589);
xor (n1352,n1263,n1264);
and (n1353,n1354,n1355);
xor (n1354,n1352,n589);
and (n1355,n1356,n1357);
xor (n1356,n1269,n1270);
and (n1357,n284,n71);
and (n1358,n245,n68);
or (n1359,n1360,n1362);
and (n1360,n1361,n1358);
xor (n1361,n1068,n1082);
and (n1362,n1363,n1364);
xor (n1363,n1361,n1358);
or (n1364,n1365,n1367);
and (n1365,n1366,n1358);
xor (n1366,n1068,n1084);
and (n1367,n1368,n1369);
xor (n1368,n1366,n1358);
or (n1369,n1370,n1372);
and (n1370,n1371,n1358);
xor (n1371,n1068,n1086);
and (n1372,n1373,n1374);
xor (n1373,n1371,n1358);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1068,n1088);
and (n1377,n111,n68);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1274,n1275);
and (n1383,n105,n68);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1280,n1281);
and (n1389,n138,n68);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
or (n1392,n1393,n1396);
and (n1393,n1394,n1395);
xor (n1394,n1286,n1287);
and (n1395,n133,n68);
and (n1396,n1397,n1398);
xor (n1397,n1394,n1395);
or (n1398,n1399,n1402);
and (n1399,n1400,n1401);
xor (n1400,n1292,n1293);
and (n1401,n86,n68);
and (n1402,n1403,n1404);
xor (n1403,n1400,n1401);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1298,n1299);
and (n1407,n80,n68);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1414);
and (n1411,n1412,n1413);
xor (n1412,n1304,n1305);
and (n1413,n46,n68);
and (n1414,n1415,n1416);
xor (n1415,n1412,n1413);
or (n1416,n1417,n1420);
and (n1417,n1418,n1419);
xor (n1418,n1310,n1311);
and (n1419,n20,n68);
and (n1420,n1421,n1422);
xor (n1421,n1418,n1419);
or (n1422,n1423,n1426);
and (n1423,n1424,n1425);
xor (n1424,n1316,n1317);
and (n1425,n59,n68);
and (n1426,n1427,n1428);
xor (n1427,n1424,n1425);
or (n1428,n1429,n1432);
and (n1429,n1430,n1431);
xor (n1430,n1322,n1323);
and (n1431,n166,n68);
and (n1432,n1433,n1434);
xor (n1433,n1430,n1431);
or (n1434,n1435,n1438);
and (n1435,n1436,n1437);
xor (n1436,n1328,n1329);
and (n1437,n205,n68);
and (n1438,n1439,n1440);
xor (n1439,n1436,n1437);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1333,n1334);
and (n1443,n299,n68);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1339,n1340);
and (n1449,n315,n68);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1344,n1345);
and (n1455,n309,n68);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1349,n1350);
and (n1461,n290,n68);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
and (n1464,n1465,n562);
xor (n1465,n1354,n1355);
and (n1466,n245,n34);
or (n1467,n1468,n1470);
and (n1468,n1469,n1466);
xor (n1469,n1363,n1364);
and (n1470,n1471,n1472);
xor (n1471,n1469,n1466);
or (n1472,n1473,n1475);
and (n1473,n1474,n1466);
xor (n1474,n1368,n1369);
and (n1475,n1476,n1477);
xor (n1476,n1474,n1466);
or (n1477,n1478,n1481);
and (n1478,n1479,n1480);
xor (n1479,n1373,n1374);
and (n1480,n111,n34);
and (n1481,n1482,n1483);
xor (n1482,n1479,n1480);
or (n1483,n1484,n1487);
and (n1484,n1485,n1486);
xor (n1485,n1379,n1380);
and (n1486,n105,n34);
and (n1487,n1488,n1489);
xor (n1488,n1485,n1486);
or (n1489,n1490,n1493);
and (n1490,n1491,n1492);
xor (n1491,n1385,n1386);
and (n1492,n138,n34);
and (n1493,n1494,n1495);
xor (n1494,n1491,n1492);
or (n1495,n1496,n1499);
and (n1496,n1497,n1498);
xor (n1497,n1391,n1392);
and (n1498,n133,n34);
and (n1499,n1500,n1501);
xor (n1500,n1497,n1498);
or (n1501,n1502,n1505);
and (n1502,n1503,n1504);
xor (n1503,n1397,n1398);
and (n1504,n86,n34);
and (n1505,n1506,n1507);
xor (n1506,n1503,n1504);
or (n1507,n1508,n1511);
and (n1508,n1509,n1510);
xor (n1509,n1403,n1404);
and (n1510,n80,n34);
and (n1511,n1512,n1513);
xor (n1512,n1509,n1510);
or (n1513,n1514,n1517);
and (n1514,n1515,n1516);
xor (n1515,n1409,n1410);
and (n1516,n46,n34);
and (n1517,n1518,n1519);
xor (n1518,n1515,n1516);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1415,n1416);
and (n1522,n20,n34);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1421,n1422);
and (n1528,n59,n34);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1427,n1428);
and (n1534,n166,n34);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1433,n1434);
and (n1540,n205,n34);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1439,n1440);
and (n1546,n299,n34);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1445,n1446);
and (n1552,n315,n34);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1451,n1452);
and (n1558,n309,n34);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1564);
and (n1562,n1563,n551);
xor (n1563,n1457,n1458);
and (n1564,n1565,n1566);
xor (n1565,n1563,n551);
and (n1566,n1567,n1568);
xor (n1567,n1463,n1464);
and (n1568,n284,n34);
and (n1569,n245,n31);
or (n1570,n1571,n1573);
and (n1571,n1572,n1569);
xor (n1572,n1471,n1472);
and (n1573,n1574,n1575);
xor (n1574,n1572,n1569);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1476,n1477);
and (n1578,n111,n31);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1482,n1483);
and (n1584,n105,n31);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1591);
and (n1588,n1589,n1590);
xor (n1589,n1488,n1489);
and (n1590,n138,n31);
and (n1591,n1592,n1593);
xor (n1592,n1589,n1590);
or (n1593,n1594,n1597);
and (n1594,n1595,n1596);
xor (n1595,n1494,n1495);
and (n1596,n133,n31);
and (n1597,n1598,n1599);
xor (n1598,n1595,n1596);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
xor (n1601,n1500,n1501);
and (n1602,n86,n31);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1506,n1507);
and (n1608,n80,n31);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1512,n1513);
and (n1614,n46,n31);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1518,n1519);
and (n1620,n20,n31);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1524,n1525);
and (n1626,n59,n31);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1633);
and (n1630,n1631,n1632);
xor (n1631,n1530,n1531);
and (n1632,n166,n31);
and (n1633,n1634,n1635);
xor (n1634,n1631,n1632);
or (n1635,n1636,n1639);
and (n1636,n1637,n1638);
xor (n1637,n1536,n1537);
and (n1638,n205,n31);
and (n1639,n1640,n1641);
xor (n1640,n1637,n1638);
or (n1641,n1642,n1645);
and (n1642,n1643,n1644);
xor (n1643,n1542,n1543);
and (n1644,n299,n31);
and (n1645,n1646,n1647);
xor (n1646,n1643,n1644);
or (n1647,n1648,n1651);
and (n1648,n1649,n1650);
xor (n1649,n1548,n1549);
and (n1650,n315,n31);
and (n1651,n1652,n1653);
xor (n1652,n1649,n1650);
or (n1653,n1654,n1657);
and (n1654,n1655,n1656);
xor (n1655,n1554,n1555);
and (n1656,n309,n31);
and (n1657,n1658,n1659);
xor (n1658,n1655,n1656);
or (n1659,n1660,n1663);
and (n1660,n1661,n1662);
xor (n1661,n1560,n1561);
and (n1662,n290,n31);
and (n1663,n1664,n1665);
xor (n1664,n1661,n1662);
and (n1665,n1666,n1667);
xor (n1666,n1565,n1566);
not (n1667,n357);
and (n1668,n245,n21);
or (n1669,n1670,n1673);
and (n1670,n1671,n1672);
xor (n1671,n1574,n1575);
and (n1672,n111,n21);
and (n1673,n1674,n1675);
xor (n1674,n1671,n1672);
or (n1675,n1676,n1679);
and (n1676,n1677,n1678);
xor (n1677,n1580,n1581);
and (n1678,n105,n21);
and (n1679,n1680,n1681);
xor (n1680,n1677,n1678);
or (n1681,n1682,n1685);
and (n1682,n1683,n1684);
xor (n1683,n1586,n1587);
and (n1684,n138,n21);
and (n1685,n1686,n1687);
xor (n1686,n1683,n1684);
or (n1687,n1688,n1691);
and (n1688,n1689,n1690);
xor (n1689,n1592,n1593);
and (n1690,n133,n21);
and (n1691,n1692,n1693);
xor (n1692,n1689,n1690);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1598,n1599);
and (n1696,n86,n21);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1604,n1605);
and (n1702,n80,n21);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
or (n1705,n1706,n1708);
and (n1706,n1707,n45);
xor (n1707,n1610,n1611);
and (n1708,n1709,n1710);
xor (n1709,n1707,n45);
or (n1710,n1711,n1713);
and (n1711,n1712,n19);
xor (n1712,n1616,n1617);
and (n1713,n1714,n1715);
xor (n1714,n1712,n19);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1622,n1623);
and (n1718,n59,n21);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1628,n1629);
and (n1724,n166,n21);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1730);
and (n1728,n1729,n494);
xor (n1729,n1634,n1635);
and (n1730,n1731,n1732);
xor (n1731,n1729,n494);
or (n1732,n1733,n1735);
and (n1733,n1734,n447);
xor (n1734,n1640,n1641);
and (n1735,n1736,n1737);
xor (n1736,n1734,n447);
or (n1737,n1738,n1740);
and (n1738,n1739,n376);
xor (n1739,n1646,n1647);
and (n1740,n1741,n1742);
xor (n1741,n1739,n376);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1652,n1653);
and (n1745,n309,n21);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1658,n1659);
and (n1751,n290,n21);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
and (n1754,n1755,n1756);
xor (n1755,n1664,n1665);
and (n1756,n284,n21);
and (n1757,n111,n52);
or (n1758,n1759,n1761);
and (n1759,n1760,n789);
xor (n1760,n1674,n1675);
and (n1761,n1762,n1763);
xor (n1762,n1760,n789);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1680,n1681);
and (n1766,n138,n52);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1686,n1687);
and (n1772,n133,n52);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1692,n1693);
and (n1778,n86,n52);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1698,n1699);
and (n1784,n80,n52);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1704,n1705);
and (n1790,n46,n52);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1709,n1710);
and (n1796,n20,n52);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1714,n1715);
and (n1802,n59,n52);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1720,n1721);
and (n1808,n166,n52);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
or (n1811,n1812,n1815);
and (n1812,n1813,n1814);
xor (n1813,n1726,n1727);
and (n1814,n205,n52);
and (n1815,n1816,n1817);
xor (n1816,n1813,n1814);
or (n1817,n1818,n1821);
and (n1818,n1819,n1820);
xor (n1819,n1731,n1732);
and (n1820,n299,n52);
and (n1821,n1822,n1823);
xor (n1822,n1819,n1820);
or (n1823,n1824,n1827);
and (n1824,n1825,n1826);
xor (n1825,n1736,n1737);
and (n1826,n315,n52);
and (n1827,n1828,n1829);
xor (n1828,n1825,n1826);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1741,n1742);
and (n1832,n309,n52);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1747,n1748);
and (n1838,n290,n52);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
and (n1841,n1842,n1843);
xor (n1842,n1753,n1754);
and (n1843,n284,n52);
or (n1844,n1845,n1847);
and (n1845,n1846,n1766);
xor (n1846,n1762,n1763);
and (n1847,n1848,n1849);
xor (n1848,n1846,n1766);
or (n1849,n1850,n1852);
and (n1850,n1851,n1772);
xor (n1851,n1768,n1769);
and (n1852,n1853,n1854);
xor (n1853,n1851,n1772);
or (n1854,n1855,n1857);
and (n1855,n1856,n1778);
xor (n1856,n1774,n1775);
and (n1857,n1858,n1859);
xor (n1858,n1856,n1778);
or (n1859,n1860,n1862);
and (n1860,n1861,n1784);
xor (n1861,n1780,n1781);
and (n1862,n1863,n1864);
xor (n1863,n1861,n1784);
or (n1864,n1865,n1867);
and (n1865,n1866,n1790);
xor (n1866,n1786,n1787);
and (n1867,n1868,n1869);
xor (n1868,n1866,n1790);
or (n1869,n1870,n1872);
and (n1870,n1871,n1796);
xor (n1871,n1792,n1793);
and (n1872,n1873,n1874);
xor (n1873,n1871,n1796);
or (n1874,n1875,n1877);
and (n1875,n1876,n1802);
xor (n1876,n1798,n1799);
and (n1877,n1878,n1879);
xor (n1878,n1876,n1802);
or (n1879,n1880,n1882);
and (n1880,n1881,n1808);
xor (n1881,n1804,n1805);
and (n1882,n1883,n1884);
xor (n1883,n1881,n1808);
or (n1884,n1885,n1887);
and (n1885,n1886,n1814);
xor (n1886,n1810,n1811);
and (n1887,n1888,n1889);
xor (n1888,n1886,n1814);
or (n1889,n1890,n1892);
and (n1890,n1891,n1820);
xor (n1891,n1816,n1817);
and (n1892,n1893,n1894);
xor (n1893,n1891,n1820);
or (n1894,n1895,n1897);
and (n1895,n1896,n1826);
xor (n1896,n1822,n1823);
and (n1897,n1898,n1899);
xor (n1898,n1896,n1826);
or (n1899,n1900,n1902);
and (n1900,n1901,n1832);
xor (n1901,n1828,n1829);
and (n1902,n1903,n1904);
xor (n1903,n1901,n1832);
or (n1904,n1905,n1907);
and (n1905,n1906,n1838);
xor (n1906,n1834,n1835);
and (n1907,n1908,n1909);
xor (n1908,n1906,n1838);
and (n1909,n1910,n1843);
xor (n1910,n1840,n1841);
or (n1911,n1912,n1914);
and (n1912,n1913,n1772);
xor (n1913,n1848,n1849);
and (n1914,n1915,n1916);
xor (n1915,n1913,n1772);
or (n1916,n1917,n1919);
and (n1917,n1918,n1778);
xor (n1918,n1853,n1854);
and (n1919,n1920,n1921);
xor (n1920,n1918,n1778);
or (n1921,n1922,n1924);
and (n1922,n1923,n1784);
xor (n1923,n1858,n1859);
and (n1924,n1925,n1926);
xor (n1925,n1923,n1784);
or (n1926,n1927,n1929);
and (n1927,n1928,n1790);
xor (n1928,n1863,n1864);
and (n1929,n1930,n1931);
xor (n1930,n1928,n1790);
or (n1931,n1932,n1934);
and (n1932,n1933,n1796);
xor (n1933,n1868,n1869);
and (n1934,n1935,n1936);
xor (n1935,n1933,n1796);
or (n1936,n1937,n1939);
and (n1937,n1938,n1802);
xor (n1938,n1873,n1874);
and (n1939,n1940,n1941);
xor (n1940,n1938,n1802);
or (n1941,n1942,n1944);
and (n1942,n1943,n1808);
xor (n1943,n1878,n1879);
and (n1944,n1945,n1946);
xor (n1945,n1943,n1808);
or (n1946,n1947,n1949);
and (n1947,n1948,n1814);
xor (n1948,n1883,n1884);
and (n1949,n1950,n1951);
xor (n1950,n1948,n1814);
or (n1951,n1952,n1954);
and (n1952,n1953,n1820);
xor (n1953,n1888,n1889);
and (n1954,n1955,n1956);
xor (n1955,n1953,n1820);
or (n1956,n1957,n1959);
and (n1957,n1958,n1826);
xor (n1958,n1893,n1894);
and (n1959,n1960,n1961);
xor (n1960,n1958,n1826);
or (n1961,n1962,n1964);
and (n1962,n1963,n1832);
xor (n1963,n1898,n1899);
and (n1964,n1965,n1966);
xor (n1965,n1963,n1832);
or (n1966,n1967,n1969);
and (n1967,n1968,n1838);
xor (n1968,n1903,n1904);
and (n1969,n1970,n1971);
xor (n1970,n1968,n1838);
and (n1971,n1972,n1843);
xor (n1972,n1908,n1909);
or (n1973,n1974,n1976);
and (n1974,n1975,n1778);
xor (n1975,n1915,n1916);
and (n1976,n1977,n1978);
xor (n1977,n1975,n1778);
or (n1978,n1979,n1981);
and (n1979,n1980,n1784);
xor (n1980,n1920,n1921);
and (n1981,n1982,n1983);
xor (n1982,n1980,n1784);
or (n1983,n1984,n1986);
and (n1984,n1985,n1790);
xor (n1985,n1925,n1926);
and (n1986,n1987,n1988);
xor (n1987,n1985,n1790);
or (n1988,n1989,n1991);
and (n1989,n1990,n1796);
xor (n1990,n1930,n1931);
and (n1991,n1992,n1993);
xor (n1992,n1990,n1796);
or (n1993,n1994,n1996);
and (n1994,n1995,n1802);
xor (n1995,n1935,n1936);
and (n1996,n1997,n1998);
xor (n1997,n1995,n1802);
or (n1998,n1999,n2001);
and (n1999,n2000,n1808);
xor (n2000,n1940,n1941);
and (n2001,n2002,n2003);
xor (n2002,n2000,n1808);
or (n2003,n2004,n2006);
and (n2004,n2005,n1814);
xor (n2005,n1945,n1946);
and (n2006,n2007,n2008);
xor (n2007,n2005,n1814);
or (n2008,n2009,n2011);
and (n2009,n2010,n1820);
xor (n2010,n1950,n1951);
and (n2011,n2012,n2013);
xor (n2012,n2010,n1820);
or (n2013,n2014,n2016);
and (n2014,n2015,n1826);
xor (n2015,n1955,n1956);
and (n2016,n2017,n2018);
xor (n2017,n2015,n1826);
or (n2018,n2019,n2021);
and (n2019,n2020,n1832);
xor (n2020,n1960,n1961);
and (n2021,n2022,n2023);
xor (n2022,n2020,n1832);
or (n2023,n2024,n2026);
and (n2024,n2025,n1838);
xor (n2025,n1965,n1966);
and (n2026,n2027,n2028);
xor (n2027,n2025,n1838);
and (n2028,n2029,n1843);
xor (n2029,n1970,n1971);
or (n2030,n2031,n2033);
and (n2031,n2032,n1784);
xor (n2032,n1977,n1978);
and (n2033,n2034,n2035);
xor (n2034,n2032,n1784);
or (n2035,n2036,n2038);
and (n2036,n2037,n1790);
xor (n2037,n1982,n1983);
and (n2038,n2039,n2040);
xor (n2039,n2037,n1790);
or (n2040,n2041,n2043);
and (n2041,n2042,n1796);
xor (n2042,n1987,n1988);
and (n2043,n2044,n2045);
xor (n2044,n2042,n1796);
or (n2045,n2046,n2048);
and (n2046,n2047,n1802);
xor (n2047,n1992,n1993);
and (n2048,n2049,n2050);
xor (n2049,n2047,n1802);
or (n2050,n2051,n2053);
and (n2051,n2052,n1808);
xor (n2052,n1997,n1998);
and (n2053,n2054,n2055);
xor (n2054,n2052,n1808);
or (n2055,n2056,n2058);
and (n2056,n2057,n1814);
xor (n2057,n2002,n2003);
and (n2058,n2059,n2060);
xor (n2059,n2057,n1814);
or (n2060,n2061,n2063);
and (n2061,n2062,n1820);
xor (n2062,n2007,n2008);
and (n2063,n2064,n2065);
xor (n2064,n2062,n1820);
or (n2065,n2066,n2068);
and (n2066,n2067,n1826);
xor (n2067,n2012,n2013);
and (n2068,n2069,n2070);
xor (n2069,n2067,n1826);
or (n2070,n2071,n2073);
and (n2071,n2072,n1832);
xor (n2072,n2017,n2018);
and (n2073,n2074,n2075);
xor (n2074,n2072,n1832);
or (n2075,n2076,n2078);
and (n2076,n2077,n1838);
xor (n2077,n2022,n2023);
and (n2078,n2079,n2080);
xor (n2079,n2077,n1838);
and (n2080,n2081,n1843);
xor (n2081,n2027,n2028);
or (n2082,n2083,n2085);
and (n2083,n2084,n1790);
xor (n2084,n2034,n2035);
and (n2085,n2086,n2087);
xor (n2086,n2084,n1790);
or (n2087,n2088,n2090);
and (n2088,n2089,n1796);
xor (n2089,n2039,n2040);
and (n2090,n2091,n2092);
xor (n2091,n2089,n1796);
or (n2092,n2093,n2095);
and (n2093,n2094,n1802);
xor (n2094,n2044,n2045);
and (n2095,n2096,n2097);
xor (n2096,n2094,n1802);
or (n2097,n2098,n2100);
and (n2098,n2099,n1808);
xor (n2099,n2049,n2050);
and (n2100,n2101,n2102);
xor (n2101,n2099,n1808);
or (n2102,n2103,n2105);
and (n2103,n2104,n1814);
xor (n2104,n2054,n2055);
and (n2105,n2106,n2107);
xor (n2106,n2104,n1814);
or (n2107,n2108,n2110);
and (n2108,n2109,n1820);
xor (n2109,n2059,n2060);
and (n2110,n2111,n2112);
xor (n2111,n2109,n1820);
or (n2112,n2113,n2115);
and (n2113,n2114,n1826);
xor (n2114,n2064,n2065);
and (n2115,n2116,n2117);
xor (n2116,n2114,n1826);
or (n2117,n2118,n2120);
and (n2118,n2119,n1832);
xor (n2119,n2069,n2070);
and (n2120,n2121,n2122);
xor (n2121,n2119,n1832);
or (n2122,n2123,n2125);
and (n2123,n2124,n1838);
xor (n2124,n2074,n2075);
and (n2125,n2126,n2127);
xor (n2126,n2124,n1838);
and (n2127,n2128,n1843);
xor (n2128,n2079,n2080);
or (n2129,n2130,n2132);
and (n2130,n2131,n1796);
xor (n2131,n2086,n2087);
and (n2132,n2133,n2134);
xor (n2133,n2131,n1796);
or (n2134,n2135,n2137);
and (n2135,n2136,n1802);
xor (n2136,n2091,n2092);
and (n2137,n2138,n2139);
xor (n2138,n2136,n1802);
or (n2139,n2140,n2142);
and (n2140,n2141,n1808);
xor (n2141,n2096,n2097);
and (n2142,n2143,n2144);
xor (n2143,n2141,n1808);
or (n2144,n2145,n2147);
and (n2145,n2146,n1814);
xor (n2146,n2101,n2102);
and (n2147,n2148,n2149);
xor (n2148,n2146,n1814);
or (n2149,n2150,n2152);
and (n2150,n2151,n1820);
xor (n2151,n2106,n2107);
and (n2152,n2153,n2154);
xor (n2153,n2151,n1820);
or (n2154,n2155,n2157);
and (n2155,n2156,n1826);
xor (n2156,n2111,n2112);
and (n2157,n2158,n2159);
xor (n2158,n2156,n1826);
or (n2159,n2160,n2162);
and (n2160,n2161,n1832);
xor (n2161,n2116,n2117);
and (n2162,n2163,n2164);
xor (n2163,n2161,n1832);
or (n2164,n2165,n2167);
and (n2165,n2166,n1838);
xor (n2166,n2121,n2122);
and (n2167,n2168,n2169);
xor (n2168,n2166,n1838);
and (n2169,n2170,n1843);
xor (n2170,n2126,n2127);
or (n2171,n2172,n2174);
and (n2172,n2173,n1802);
xor (n2173,n2133,n2134);
and (n2174,n2175,n2176);
xor (n2175,n2173,n1802);
or (n2176,n2177,n2179);
and (n2177,n2178,n1808);
xor (n2178,n2138,n2139);
and (n2179,n2180,n2181);
xor (n2180,n2178,n1808);
or (n2181,n2182,n2184);
and (n2182,n2183,n1814);
xor (n2183,n2143,n2144);
and (n2184,n2185,n2186);
xor (n2185,n2183,n1814);
or (n2186,n2187,n2189);
and (n2187,n2188,n1820);
xor (n2188,n2148,n2149);
and (n2189,n2190,n2191);
xor (n2190,n2188,n1820);
or (n2191,n2192,n2194);
and (n2192,n2193,n1826);
xor (n2193,n2153,n2154);
and (n2194,n2195,n2196);
xor (n2195,n2193,n1826);
or (n2196,n2197,n2199);
and (n2197,n2198,n1832);
xor (n2198,n2158,n2159);
and (n2199,n2200,n2201);
xor (n2200,n2198,n1832);
or (n2201,n2202,n2204);
and (n2202,n2203,n1838);
xor (n2203,n2163,n2164);
and (n2204,n2205,n2206);
xor (n2205,n2203,n1838);
and (n2206,n2207,n1843);
xor (n2207,n2168,n2169);
or (n2208,n2209,n2211);
and (n2209,n2210,n1808);
xor (n2210,n2175,n2176);
and (n2211,n2212,n2213);
xor (n2212,n2210,n1808);
or (n2213,n2214,n2216);
and (n2214,n2215,n1814);
xor (n2215,n2180,n2181);
and (n2216,n2217,n2218);
xor (n2217,n2215,n1814);
or (n2218,n2219,n2221);
and (n2219,n2220,n1820);
xor (n2220,n2185,n2186);
and (n2221,n2222,n2223);
xor (n2222,n2220,n1820);
or (n2223,n2224,n2226);
and (n2224,n2225,n1826);
xor (n2225,n2190,n2191);
and (n2226,n2227,n2228);
xor (n2227,n2225,n1826);
or (n2228,n2229,n2231);
and (n2229,n2230,n1832);
xor (n2230,n2195,n2196);
and (n2231,n2232,n2233);
xor (n2232,n2230,n1832);
or (n2233,n2234,n2236);
and (n2234,n2235,n1838);
xor (n2235,n2200,n2201);
and (n2236,n2237,n2238);
xor (n2237,n2235,n1838);
and (n2238,n2239,n1843);
xor (n2239,n2205,n2206);
or (n2240,n2241,n2243);
and (n2241,n2242,n1814);
xor (n2242,n2212,n2213);
and (n2243,n2244,n2245);
xor (n2244,n2242,n1814);
or (n2245,n2246,n2248);
and (n2246,n2247,n1820);
xor (n2247,n2217,n2218);
and (n2248,n2249,n2250);
xor (n2249,n2247,n1820);
or (n2250,n2251,n2253);
and (n2251,n2252,n1826);
xor (n2252,n2222,n2223);
and (n2253,n2254,n2255);
xor (n2254,n2252,n1826);
or (n2255,n2256,n2258);
and (n2256,n2257,n1832);
xor (n2257,n2227,n2228);
and (n2258,n2259,n2260);
xor (n2259,n2257,n1832);
or (n2260,n2261,n2263);
and (n2261,n2262,n1838);
xor (n2262,n2232,n2233);
and (n2263,n2264,n2265);
xor (n2264,n2262,n1838);
and (n2265,n2266,n1843);
xor (n2266,n2237,n2238);
or (n2267,n2268,n2270);
and (n2268,n2269,n1820);
xor (n2269,n2244,n2245);
and (n2270,n2271,n2272);
xor (n2271,n2269,n1820);
or (n2272,n2273,n2275);
and (n2273,n2274,n1826);
xor (n2274,n2249,n2250);
and (n2275,n2276,n2277);
xor (n2276,n2274,n1826);
or (n2277,n2278,n2280);
and (n2278,n2279,n1832);
xor (n2279,n2254,n2255);
and (n2280,n2281,n2282);
xor (n2281,n2279,n1832);
or (n2282,n2283,n2285);
and (n2283,n2284,n1838);
xor (n2284,n2259,n2260);
and (n2285,n2286,n2287);
xor (n2286,n2284,n1838);
and (n2287,n2288,n1843);
xor (n2288,n2264,n2265);
or (n2289,n2290,n2292);
and (n2290,n2291,n1826);
xor (n2291,n2271,n2272);
and (n2292,n2293,n2294);
xor (n2293,n2291,n1826);
or (n2294,n2295,n2297);
and (n2295,n2296,n1832);
xor (n2296,n2276,n2277);
and (n2297,n2298,n2299);
xor (n2298,n2296,n1832);
or (n2299,n2300,n2302);
and (n2300,n2301,n1838);
xor (n2301,n2281,n2282);
and (n2302,n2303,n2304);
xor (n2303,n2301,n1838);
and (n2304,n2305,n1843);
xor (n2305,n2286,n2287);
or (n2306,n2307,n2309);
and (n2307,n2308,n1832);
xor (n2308,n2293,n2294);
and (n2309,n2310,n2311);
xor (n2310,n2308,n1832);
or (n2311,n2312,n2314);
and (n2312,n2313,n1838);
xor (n2313,n2298,n2299);
and (n2314,n2315,n2316);
xor (n2315,n2313,n1838);
and (n2316,n2317,n1843);
xor (n2317,n2303,n2304);
or (n2318,n2319,n2321);
and (n2319,n2320,n1838);
xor (n2320,n2310,n2311);
and (n2321,n2322,n2323);
xor (n2322,n2320,n1838);
and (n2323,n2324,n1843);
xor (n2324,n2315,n2316);
and (n2325,n2326,n1843);
xor (n2326,n2322,n2323);
xor (n2327,n2239,n1843);
endmodule
