module top (out,n6,n10,n12,n13,n15,n17,n18,n38,n39
        ,n47,n48,n50,n51,n68,n69,n71,n80,n81,n90
        ,n101,n102,n109,n115,n128,n137,n142,n160,n204,n398);
output out;
input n6;
input n10;
input n12;
input n13;
input n15;
input n17;
input n18;
input n38;
input n39;
input n47;
input n48;
input n50;
input n51;
input n68;
input n69;
input n71;
input n80;
input n81;
input n90;
input n101;
input n102;
input n109;
input n115;
input n128;
input n137;
input n142;
input n160;
input n204;
input n398;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n7;
wire n8;
wire n9;
wire n11;
wire n14;
wire n16;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n49;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
xnor (out,n0,n400);
nand (n0,n1,n399);
not (n1,n2);
nor (n2,n3,n398);
nand (n3,n4,n19);
or (n4,n5,n7);
not (n5,n6);
not (n7,n8);
xor (n8,n9,n14);
and (n9,n10,n11);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n6);
and (s0n11,notn11,n12);
and (s1n11,n6,n13);
and (n14,n15,n16);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n6);
and (s0n16,notn16,n17);
and (s1n16,n6,n18);
nand (n19,n20,n5);
nand (n20,n21,n397);
or (n21,n22,n228);
not (n22,n23);
or (n23,n24,n227);
and (n24,n25,n184);
or (n25,n26,n183);
and (n26,n27,n152);
xor (n27,n28,n119);
or (n28,n29,n118);
and (n29,n30,n93);
xor (n30,n31,n62);
nand (n31,n32,n57);
or (n32,n33,n42);
not (n33,n34);
nand (n34,n35,n40);
or (n35,n36,n15);
not (n36,n37);
wire s0n37,s1n37,notn37;
or (n37,s0n37,s1n37);
not(notn37,n6);
and (s0n37,notn37,n38);
and (s1n37,n6,n39);
or (n40,n37,n41);
not (n41,n15);
nand (n42,n43,n54);
nor (n43,n44,n52);
and (n44,n45,n49);
not (n45,n46);
wire s0n46,s1n46,notn46;
or (n46,s0n46,s1n46);
not(notn46,n6);
and (s0n46,notn46,n47);
and (s1n46,n6,n48);
wire s0n49,s1n49,notn49;
or (n49,s0n49,s1n49);
not(notn49,n6);
and (s0n49,notn49,n50);
and (s1n49,n6,n51);
and (n52,n46,n53);
not (n53,n49);
nand (n54,n55,n56);
or (n55,n45,n37);
nand (n56,n37,n45);
or (n57,n43,n58);
nor (n58,n59,n60);
and (n59,n10,n36);
and (n60,n61,n37);
not (n61,n10);
nand (n62,n63,n87);
or (n63,n64,n74);
not (n64,n65);
nand (n65,n66,n72);
or (n66,n67,n70);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n6);
and (s0n67,notn67,n68);
and (s1n67,n6,n69);
not (n70,n71);
or (n72,n73,n71);
not (n73,n67);
not (n74,n75);
and (n75,n76,n83);
nand (n76,n77,n82);
or (n77,n78,n67);
not (n78,n79);
wire s0n79,s1n79,notn79;
or (n79,s0n79,s1n79);
not(notn79,n6);
and (s0n79,notn79,n80);
and (s1n79,n6,n81);
nand (n82,n67,n78);
not (n83,n84);
nand (n84,n85,n86);
or (n85,n78,n16);
nand (n86,n16,n78);
nand (n87,n84,n88);
nor (n88,n89,n91);
and (n89,n90,n67);
and (n91,n92,n73);
not (n92,n90);
nand (n93,n94,n112);
or (n94,n95,n107);
nand (n95,n96,n104);
not (n96,n97);
nand (n97,n98,n103);
or (n98,n99,n67);
not (n99,n100);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n6);
and (s0n100,notn100,n101);
and (s1n100,n6,n102);
nand (n103,n67,n99);
nand (n104,n105,n106);
or (n105,n99,n49);
nand (n106,n49,n99);
nor (n107,n108,n110);
and (n108,n53,n109);
and (n110,n49,n111);
not (n111,n109);
or (n112,n96,n113);
nor (n113,n114,n116);
and (n114,n53,n115);
and (n116,n49,n117);
not (n117,n115);
and (n118,n31,n62);
xor (n119,n120,n146);
xor (n120,n121,n129);
and (n121,n122,n15);
not (n122,n123);
nand (n123,n37,n124);
not (n124,n125);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n6);
and (s0n125,notn125,1'b0);
and (s1n125,n6,n127);
and (n127,n128,n39);
nand (n129,n130,n139);
or (n130,n131,n134);
not (n131,n132);
nor (n132,n133,n11);
not (n133,n16);
nor (n134,n135,n138);
and (n135,n136,n16);
not (n136,n137);
and (n138,n137,n133);
or (n139,n140,n145);
nor (n140,n141,n143);
and (n141,n133,n142);
and (n143,n16,n144);
not (n144,n142);
not (n145,n11);
nand (n146,n147,n148);
or (n147,n42,n58);
or (n148,n43,n149);
nor (n149,n150,n151);
and (n150,n109,n36);
and (n151,n111,n37);
xor (n152,n153,n169);
xor (n153,n154,n163);
nand (n154,n155,n157);
or (n155,n74,n156);
not (n156,n88);
or (n157,n83,n158);
nor (n158,n159,n161);
and (n159,n73,n160);
and (n161,n67,n162);
not (n162,n160);
nand (n163,n164,n165);
or (n164,n95,n113);
or (n165,n96,n166);
nor (n166,n167,n168);
and (n167,n53,n71);
and (n168,n49,n70);
and (n169,n170,n175);
nor (n170,n171,n36);
nor (n171,n172,n174);
and (n172,n53,n173);
nand (n173,n46,n15);
and (n174,n45,n41);
nand (n175,n176,n181);
or (n176,n177,n131);
not (n177,n178);
nor (n178,n179,n180);
and (n179,n160,n16);
and (n180,n162,n133);
nand (n181,n182,n11);
not (n182,n134);
and (n183,n28,n119);
xor (n184,n185,n210);
xor (n185,n186,n207);
xor (n186,n187,n199);
xor (n187,n188,n195);
nand (n188,n189,n190);
or (n189,n149,n42);
nand (n190,n191,n194);
nor (n191,n192,n193);
and (n192,n115,n37);
and (n193,n117,n36);
not (n194,n43);
nor (n195,n123,n196);
nor (n196,n197,n198);
and (n197,n125,n61);
and (n198,n124,n10);
nand (n199,n200,n201);
or (n200,n131,n140);
or (n201,n202,n145);
nor (n202,n203,n205);
and (n203,n133,n204);
and (n205,n16,n206);
not (n206,n204);
or (n207,n208,n209);
and (n208,n153,n169);
and (n209,n154,n163);
xor (n210,n211,n224);
xor (n211,n212,n218);
nand (n212,n213,n214);
or (n213,n95,n166);
or (n214,n96,n215);
nor (n215,n216,n217);
and (n216,n53,n90);
and (n217,n49,n92);
nand (n218,n219,n220);
or (n219,n74,n158);
or (n220,n221,n83);
nor (n221,n222,n223);
and (n222,n73,n137);
and (n223,n67,n136);
or (n224,n225,n226);
and (n225,n120,n146);
and (n226,n121,n129);
nor (n227,n25,n184);
not (n228,n229);
nand (n229,n230,n396);
or (n230,n231,n391);
nor (n231,n232,n389);
and (n232,n233,n378);
or (n233,n234,n377);
and (n234,n235,n293);
xor (n235,n236,n276);
or (n236,n237,n275);
and (n237,n238,n260);
xor (n238,n239,n249);
nand (n239,n240,n245);
or (n240,n241,n74);
not (n241,n242);
nor (n242,n243,n244);
and (n243,n111,n73);
and (n244,n109,n67);
nand (n245,n84,n246);
nor (n246,n247,n248);
and (n247,n115,n67);
and (n248,n73,n117);
nand (n249,n250,n255);
or (n250,n251,n96);
not (n251,n252);
nor (n252,n253,n254);
and (n253,n10,n49);
and (n254,n61,n53);
nand (n255,n256,n257);
not (n256,n95);
nand (n257,n258,n259);
or (n258,n53,n15);
or (n259,n49,n41);
xor (n260,n261,n266);
and (n261,n262,n49);
nand (n262,n263,n265);
or (n263,n67,n264);
and (n264,n15,n100);
or (n265,n100,n15);
nand (n266,n267,n271);
or (n267,n131,n268);
nor (n268,n269,n270);
and (n269,n133,n71);
and (n270,n16,n70);
or (n271,n272,n145);
nor (n272,n273,n274);
and (n273,n90,n133);
and (n274,n92,n16);
and (n275,n239,n249);
xor (n276,n277,n282);
xor (n277,n278,n281);
nand (n278,n279,n280);
or (n279,n251,n95);
or (n280,n96,n107);
and (n281,n261,n266);
xor (n282,n283,n289);
xor (n283,n284,n285);
and (n284,n194,n15);
nand (n285,n286,n287);
or (n286,n145,n177);
nand (n287,n288,n132);
not (n288,n272);
nand (n289,n290,n292);
or (n290,n291,n74);
not (n291,n246);
nand (n292,n84,n65);
or (n293,n294,n376);
and (n294,n295,n316);
xor (n295,n296,n315);
or (n296,n297,n314);
and (n297,n298,n307);
xor (n298,n299,n300);
and (n299,n97,n15);
nand (n300,n301,n306);
or (n301,n302,n74);
not (n302,n303);
nor (n303,n304,n305);
and (n304,n10,n67);
and (n305,n61,n73);
nand (n306,n242,n84);
nand (n307,n308,n313);
or (n308,n131,n309);
not (n309,n310);
nor (n310,n311,n312);
and (n311,n117,n133);
and (n312,n115,n16);
or (n313,n268,n145);
and (n314,n299,n300);
xor (n315,n238,n260);
or (n316,n317,n375);
and (n317,n318,n374);
xor (n318,n319,n333);
nor (n319,n320,n328);
not (n320,n321);
nand (n321,n322,n327);
or (n322,n323,n131);
not (n323,n324);
nand (n324,n325,n326);
or (n325,n111,n16);
nand (n326,n16,n111);
nand (n327,n310,n11);
nand (n328,n329,n67);
nand (n329,n330,n332);
or (n330,n16,n331);
and (n331,n15,n79);
or (n332,n79,n15);
nand (n333,n334,n372);
or (n334,n335,n358);
not (n335,n336);
nand (n336,n337,n357);
or (n337,n338,n347);
nor (n338,n339,n346);
nand (n339,n340,n345);
or (n340,n341,n131);
not (n341,n342);
nand (n342,n343,n344);
or (n343,n61,n16);
nand (n344,n16,n61);
nand (n345,n324,n11);
nor (n346,n83,n41);
nand (n347,n348,n355);
nand (n348,n349,n354);
or (n349,n350,n131);
not (n350,n351);
nand (n351,n352,n353);
or (n352,n133,n15);
or (n353,n16,n41);
nand (n354,n342,n11);
nor (n355,n356,n133);
and (n356,n15,n11);
nand (n357,n339,n346);
not (n358,n359);
nand (n359,n360,n368);
not (n360,n361);
nand (n361,n362,n367);
or (n362,n363,n74);
not (n363,n364);
nand (n364,n365,n366);
or (n365,n73,n15);
or (n366,n67,n41);
nand (n367,n84,n303);
nor (n368,n369,n371);
and (n369,n320,n370);
not (n370,n328);
and (n371,n321,n328);
nand (n372,n373,n361);
not (n373,n368);
xor (n374,n298,n307);
and (n375,n319,n333);
and (n376,n296,n315);
and (n377,n236,n276);
or (n378,n379,n386);
xor (n379,n380,n385);
xor (n380,n381,n382);
xor (n381,n170,n175);
or (n382,n383,n384);
and (n383,n283,n289);
and (n384,n284,n285);
xor (n385,n30,n93);
or (n386,n387,n388);
and (n387,n277,n282);
and (n388,n278,n281);
not (n389,n390);
nand (n390,n379,n386);
nor (n391,n392,n393);
xor (n392,n27,n152);
or (n393,n394,n395);
and (n394,n380,n385);
and (n395,n381,n382);
nand (n396,n392,n393);
or (n397,n229,n23);
nand (n399,n3,n398);
xor (n400,n398,n401);
wire s0n401,s1n401,notn401;
or (n401,s0n401,s1n401);
not(notn401,n6);
and (s0n401,notn401,n402);
and (s1n401,n6,n8);
xor (n402,n403,n608);
xor (n403,n404,n606);
xor (n404,n405,n605);
xor (n405,n406,n596);
xor (n406,n407,n595);
xor (n407,n408,n580);
xor (n408,n409,n579);
xor (n409,n410,n559);
xor (n410,n411,n558);
xor (n411,n412,n532);
xor (n412,n413,n531);
xor (n413,n414,n502);
xor (n414,n415,n501);
xor (n415,n416,n463);
xor (n416,n417,n462);
xor (n417,n418,n421);
xor (n418,n419,n420);
and (n419,n204,n11);
and (n420,n142,n16);
or (n421,n422,n425);
and (n422,n423,n424);
and (n423,n142,n11);
and (n424,n137,n16);
and (n425,n426,n427);
xor (n426,n423,n424);
or (n427,n428,n430);
and (n428,n429,n179);
and (n429,n137,n11);
and (n430,n431,n432);
xor (n431,n429,n179);
or (n432,n433,n436);
and (n433,n434,n435);
and (n434,n160,n11);
and (n435,n90,n16);
and (n436,n437,n438);
xor (n437,n434,n435);
or (n438,n439,n442);
and (n439,n440,n441);
and (n440,n90,n11);
and (n441,n71,n16);
and (n442,n443,n444);
xor (n443,n440,n441);
or (n444,n445,n447);
and (n445,n446,n312);
and (n446,n71,n11);
and (n447,n448,n449);
xor (n448,n446,n312);
or (n449,n450,n453);
and (n450,n451,n452);
and (n451,n115,n11);
and (n452,n109,n16);
and (n453,n454,n455);
xor (n454,n451,n452);
or (n455,n456,n459);
and (n456,n457,n458);
and (n457,n109,n11);
and (n458,n10,n16);
and (n459,n460,n461);
xor (n460,n457,n458);
and (n461,n9,n14);
and (n462,n137,n79);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n426,n427);
and (n466,n160,n79);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n431,n432);
and (n472,n90,n79);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n437,n438);
and (n478,n71,n79);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n443,n444);
and (n484,n115,n79);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n448,n449);
and (n490,n109,n79);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n454,n455);
and (n496,n10,n79);
and (n497,n498,n499);
xor (n498,n495,n496);
and (n499,n500,n331);
xor (n500,n460,n461);
and (n501,n160,n67);
or (n502,n503,n505);
and (n503,n504,n89);
xor (n504,n468,n469);
and (n505,n506,n507);
xor (n506,n504,n89);
or (n507,n508,n511);
and (n508,n509,n510);
xor (n509,n474,n475);
and (n510,n71,n67);
and (n511,n512,n513);
xor (n512,n509,n510);
or (n513,n514,n516);
and (n514,n515,n247);
xor (n515,n480,n481);
and (n516,n517,n518);
xor (n517,n515,n247);
or (n518,n519,n521);
and (n519,n520,n244);
xor (n520,n486,n487);
and (n521,n522,n523);
xor (n522,n520,n244);
or (n523,n524,n526);
and (n524,n525,n304);
xor (n525,n492,n493);
and (n526,n527,n528);
xor (n527,n525,n304);
and (n528,n529,n530);
xor (n529,n498,n499);
and (n530,n15,n67);
and (n531,n90,n100);
or (n532,n533,n536);
and (n533,n534,n535);
xor (n534,n506,n507);
and (n535,n71,n100);
and (n536,n537,n538);
xor (n537,n534,n535);
or (n538,n539,n542);
and (n539,n540,n541);
xor (n540,n512,n513);
and (n541,n115,n100);
and (n542,n543,n544);
xor (n543,n540,n541);
or (n544,n545,n548);
and (n545,n546,n547);
xor (n546,n517,n518);
and (n547,n109,n100);
and (n548,n549,n550);
xor (n549,n546,n547);
or (n550,n551,n554);
and (n551,n552,n553);
xor (n552,n522,n523);
and (n553,n10,n100);
and (n554,n555,n556);
xor (n555,n552,n553);
and (n556,n557,n264);
xor (n557,n527,n528);
and (n558,n71,n49);
or (n559,n560,n563);
and (n560,n561,n562);
xor (n561,n537,n538);
and (n562,n115,n49);
and (n563,n564,n565);
xor (n564,n561,n562);
or (n565,n566,n569);
and (n566,n567,n568);
xor (n567,n543,n544);
and (n568,n109,n49);
and (n569,n570,n571);
xor (n570,n567,n568);
or (n571,n572,n574);
and (n572,n573,n253);
xor (n573,n549,n550);
and (n574,n575,n576);
xor (n575,n573,n253);
and (n576,n577,n578);
xor (n577,n555,n556);
and (n578,n15,n49);
and (n579,n115,n46);
or (n580,n581,n584);
and (n581,n582,n583);
xor (n582,n564,n565);
and (n583,n109,n46);
and (n584,n585,n586);
xor (n585,n582,n583);
or (n586,n587,n590);
and (n587,n588,n589);
xor (n588,n570,n571);
and (n589,n10,n46);
and (n590,n591,n592);
xor (n591,n588,n589);
and (n592,n593,n594);
xor (n593,n575,n576);
not (n594,n173);
and (n595,n109,n37);
or (n596,n597,n600);
and (n597,n598,n599);
xor (n598,n585,n586);
and (n599,n10,n37);
and (n600,n601,n602);
xor (n601,n598,n599);
and (n602,n603,n604);
xor (n603,n591,n592);
and (n604,n15,n37);
and (n605,n10,n125);
and (n606,n607,n608);
xor (n607,n601,n602);
and (n608,n15,n125);
endmodule
