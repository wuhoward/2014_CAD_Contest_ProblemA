module top (out,n14,n17,n18,n21,n23,n30,n33,n34,n38
        ,n46,n49,n50,n54,n64,n67,n68,n72,n79,n82
        ,n83,n87,n95,n98,n99,n103,n113,n116,n117,n122
        ,n125,n129,n389);
output out;
input n14;
input n17;
input n18;
input n21;
input n23;
input n30;
input n33;
input n34;
input n38;
input n46;
input n49;
input n50;
input n54;
input n64;
input n67;
input n68;
input n72;
input n79;
input n82;
input n83;
input n87;
input n95;
input n98;
input n99;
input n103;
input n113;
input n116;
input n117;
input n122;
input n125;
input n129;
input n389;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n16;
wire n19;
wire n20;
wire n22;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
xor (out,n0,n1044);
xor (n0,n1,n417);
xor (n1,n2,n340);
xor (n2,n3,n242);
or (n3,n4,n226,n241);
and (n4,n5,n185);
or (n5,n6,n173,n184);
and (n6,n7,n134);
or (n7,n8,n108,n133);
and (n8,n9,n59);
or (n9,n10,n42,n58);
and (n10,n11,n27);
xnor (n11,n12,n24);
nor (n12,n13,n22);
and (n13,n14,n15);
and (n15,n16,n19);
xor (n16,n17,n18);
not (n19,n20);
xor (n20,n18,n21);
and (n22,n23,n20);
and (n24,n17,n25);
not (n25,n26);
and (n26,n18,n21);
xnor (n27,n28,n39);
nor (n28,n29,n37);
and (n29,n30,n31);
and (n31,n32,n35);
xor (n32,n33,n34);
not (n35,n36);
xor (n36,n34,n17);
and (n37,n38,n36);
and (n39,n33,n40);
not (n40,n41);
and (n41,n34,n17);
and (n42,n27,n43);
xnor (n43,n44,n55);
nor (n44,n45,n53);
and (n45,n46,n47);
and (n47,n48,n51);
xor (n48,n49,n50);
not (n51,n52);
xor (n52,n50,n33);
and (n53,n54,n52);
and (n55,n49,n56);
not (n56,n57);
and (n57,n50,n33);
and (n58,n11,n43);
or (n59,n60,n91,n107);
and (n60,n61,n76);
xnor (n61,n62,n73);
nor (n62,n63,n71);
and (n63,n64,n65);
and (n65,n66,n69);
xor (n66,n67,n68);
not (n69,n70);
xor (n70,n68,n49);
and (n71,n72,n70);
and (n73,n67,n74);
not (n74,n75);
and (n75,n68,n49);
xnor (n76,n77,n88);
nor (n77,n78,n86);
and (n78,n79,n80);
and (n80,n81,n84);
xor (n81,n82,n83);
not (n84,n85);
xor (n85,n83,n67);
and (n86,n87,n85);
and (n88,n82,n89);
not (n89,n90);
and (n90,n83,n67);
and (n91,n76,n92);
xnor (n92,n93,n104);
nor (n93,n94,n102);
and (n94,n95,n96);
and (n96,n97,n100);
xor (n97,n98,n99);
not (n100,n101);
xor (n101,n99,n82);
and (n102,n103,n101);
and (n104,n98,n105);
not (n105,n106);
and (n106,n99,n82);
and (n107,n61,n92);
and (n108,n59,n109);
and (n109,n110,n119);
xnor (n110,n111,n116);
not (n111,n112);
and (n112,n113,n114);
and (n114,n115,n118);
xor (n115,n116,n117);
not (n118,n117);
xnor (n119,n120,n130);
nor (n120,n121,n128);
and (n121,n122,n123);
and (n123,n124,n126);
xor (n124,n21,n125);
not (n126,n127);
xor (n127,n125,n116);
and (n128,n129,n127);
and (n130,n21,n131);
not (n131,n132);
and (n132,n125,n116);
and (n133,n9,n109);
or (n134,n135,n160,n172);
and (n135,n136,n150);
xor (n136,n137,n146);
xor (n137,n138,n142);
xnor (n138,n139,n39);
nor (n139,n140,n141);
and (n140,n38,n31);
and (n141,n14,n36);
xnor (n142,n143,n55);
nor (n143,n144,n145);
and (n144,n54,n47);
and (n145,n30,n52);
xnor (n146,n147,n73);
nor (n147,n148,n149);
and (n148,n72,n65);
and (n149,n46,n70);
xor (n150,n151,n156);
xor (n151,n116,n152);
xnor (n152,n153,n130);
nor (n153,n154,n155);
and (n154,n129,n123);
and (n155,n113,n127);
xnor (n156,n157,n24);
nor (n157,n158,n159);
and (n158,n23,n15);
and (n159,n122,n20);
and (n160,n150,n161);
xor (n161,n162,n171);
xor (n162,n163,n167);
xnor (n163,n164,n88);
nor (n164,n165,n166);
and (n165,n87,n80);
and (n166,n64,n85);
xnor (n167,n168,n104);
nor (n168,n169,n170);
and (n169,n103,n96);
and (n170,n79,n101);
and (n171,n95,n98);
and (n172,n136,n161);
and (n173,n134,n174);
xor (n174,n175,n180);
xor (n175,n176,n177);
not (n176,n116);
xnor (n177,n178,n130);
not (n178,n179);
and (n179,n113,n123);
xnor (n180,n181,n24);
nor (n181,n182,n183);
and (n182,n122,n15);
and (n183,n129,n20);
and (n184,n7,n174);
and (n185,n186,n200);
xor (n186,n187,n196);
xor (n187,n188,n192);
or (n188,n189,n190,n191);
and (n189,n138,n142);
and (n190,n142,n146);
and (n191,n138,n146);
or (n192,n193,n194,n195);
and (n193,n116,n152);
and (n194,n152,n156);
and (n195,n116,n156);
or (n196,n197,n198,n199);
and (n197,n163,n167);
and (n198,n167,n171);
and (n199,n163,n171);
xnor (n200,n201,n212);
xor (n201,n202,n211);
xor (n202,n203,n207);
xnor (n203,n204,n88);
nor (n204,n205,n206);
and (n205,n64,n80);
and (n206,n72,n85);
xnor (n207,n208,n104);
nor (n208,n209,n210);
and (n209,n79,n96);
and (n210,n87,n101);
and (n211,n103,n98);
xor (n212,n213,n222);
xor (n213,n214,n218);
xnor (n214,n215,n39);
nor (n215,n216,n217);
and (n216,n14,n31);
and (n217,n23,n36);
xnor (n218,n219,n55);
nor (n219,n220,n221);
and (n220,n30,n47);
and (n221,n38,n52);
xnor (n222,n223,n73);
nor (n223,n224,n225);
and (n224,n46,n65);
and (n225,n54,n70);
and (n226,n185,n227);
xor (n227,n228,n237);
xor (n228,n229,n233);
or (n229,n230,n231,n232);
and (n230,n176,n177);
and (n231,n177,n180);
and (n232,n176,n180);
or (n233,n234,n235,n236);
and (n234,n203,n207);
and (n235,n207,n211);
and (n236,n203,n211);
or (n237,n238,n239,n240);
and (n238,n214,n218);
and (n239,n218,n222);
and (n240,n214,n222);
and (n241,n5,n227);
xor (n242,n243,n298);
xor (n243,n244,n287);
or (n244,n245,n251,n286);
and (n245,n246,n250);
or (n246,n247,n248,n249);
and (n247,n188,n192);
and (n248,n192,n196);
and (n249,n188,n196);
or (n250,n201,n212);
and (n251,n250,n252);
xor (n252,n253,n279);
xor (n253,n254,n265);
not (n254,n255);
xor (n255,n256,n261);
xor (n256,n130,n257);
xnor (n257,n258,n24);
nor (n258,n259,n260);
and (n259,n129,n15);
and (n260,n113,n20);
xnor (n261,n262,n39);
nor (n262,n263,n264);
and (n263,n23,n31);
and (n264,n122,n36);
xor (n265,n266,n275);
xor (n266,n267,n271);
xnor (n267,n268,n55);
nor (n268,n269,n270);
and (n269,n38,n47);
and (n270,n14,n52);
xnor (n271,n272,n73);
nor (n272,n273,n274);
and (n273,n54,n65);
and (n274,n30,n70);
xnor (n275,n276,n88);
nor (n276,n277,n278);
and (n277,n72,n80);
and (n278,n46,n85);
not (n279,n280);
xnor (n280,n281,n285);
xnor (n281,n282,n104);
nor (n282,n283,n284);
and (n283,n87,n96);
and (n284,n64,n101);
and (n285,n79,n98);
and (n286,n246,n252);
xor (n287,n288,n297);
xor (n288,n289,n293);
or (n289,n290,n291,n292);
and (n290,n130,n257);
and (n291,n257,n261);
and (n292,n130,n261);
or (n293,n294,n295,n296);
and (n294,n267,n271);
and (n295,n271,n275);
and (n296,n267,n275);
or (n297,n281,n285);
xor (n298,n299,n308);
xor (n299,n300,n304);
or (n300,n301,n302,n303);
and (n301,n229,n233);
and (n302,n233,n237);
and (n303,n229,n237);
or (n304,n305,n306,n307);
and (n305,n255,n265);
and (n306,n265,n280);
and (n307,n255,n280);
xor (n308,n309,n334);
xor (n309,n310,n320);
xor (n310,n311,n316);
xor (n311,n312,n313);
not (n312,n130);
xnor (n313,n314,n24);
not (n314,n315);
and (n315,n113,n15);
xnor (n316,n317,n39);
nor (n317,n318,n319);
and (n318,n122,n31);
and (n319,n129,n36);
xor (n320,n321,n330);
xor (n321,n322,n326);
xnor (n322,n323,n55);
nor (n323,n324,n325);
and (n324,n14,n47);
and (n325,n23,n52);
xnor (n326,n327,n73);
nor (n327,n328,n329);
and (n328,n30,n65);
and (n329,n38,n70);
xnor (n330,n331,n88);
nor (n331,n332,n333);
and (n332,n46,n80);
and (n333,n54,n85);
xor (n334,n335,n339);
xnor (n335,n336,n104);
nor (n336,n337,n338);
and (n337,n64,n96);
and (n338,n72,n101);
and (n339,n87,n98);
or (n340,n341,n413,n416);
and (n341,n342,n411);
or (n342,n343,n408,n410);
and (n343,n344,n406);
or (n344,n345,n402,n405);
and (n345,n346,n392);
or (n346,n347,n380,n391);
and (n347,n348,n364);
or (n348,n349,n358,n363);
and (n349,n350,n354);
xnor (n350,n351,n116);
nor (n351,n352,n353);
and (n352,n129,n114);
and (n353,n113,n117);
xnor (n354,n355,n130);
nor (n355,n356,n357);
and (n356,n23,n123);
and (n357,n122,n127);
and (n358,n354,n359);
xnor (n359,n360,n24);
nor (n360,n361,n362);
and (n361,n38,n15);
and (n362,n14,n20);
and (n363,n350,n359);
or (n364,n365,n374,n379);
and (n365,n366,n370);
xnor (n366,n367,n39);
nor (n367,n368,n369);
and (n368,n54,n31);
and (n369,n30,n36);
xnor (n370,n371,n55);
nor (n371,n372,n373);
and (n372,n72,n47);
and (n373,n46,n52);
and (n374,n370,n375);
xnor (n375,n376,n73);
nor (n376,n377,n378);
and (n377,n87,n65);
and (n378,n64,n70);
and (n379,n366,n375);
and (n380,n364,n381);
and (n381,n382,n386);
xnor (n382,n383,n88);
nor (n383,n384,n385);
and (n384,n103,n80);
and (n385,n79,n85);
xnor (n386,n387,n104);
nor (n387,n388,n390);
and (n388,n389,n96);
and (n390,n95,n101);
and (n391,n348,n381);
or (n392,n393,n398,n401);
and (n393,n394,n396);
not (n394,n395);
nand (n395,n389,n98);
xor (n396,n397,n43);
xor (n397,n11,n27);
and (n398,n396,n399);
xor (n399,n400,n92);
xor (n400,n61,n76);
and (n401,n394,n399);
and (n402,n392,n403);
xor (n403,n404,n161);
xor (n404,n136,n150);
and (n405,n346,n403);
xor (n406,n407,n174);
xor (n407,n7,n134);
and (n408,n406,n409);
xor (n409,n186,n200);
and (n410,n344,n409);
xor (n411,n412,n227);
xor (n412,n5,n185);
and (n413,n411,n414);
xor (n414,n415,n252);
xor (n415,n246,n250);
and (n416,n342,n414);
or (n417,n418,n495);
and (n418,n419,n421);
xor (n419,n420,n414);
xor (n420,n342,n411);
and (n421,n422,n493);
or (n422,n423,n489,n492);
and (n423,n424,n484);
or (n424,n425,n481,n483);
and (n425,n426,n472);
or (n426,n427,n454,n471);
and (n427,n428,n442);
or (n428,n429,n438,n441);
and (n429,n430,n434);
xnor (n430,n431,n73);
nor (n431,n432,n433);
and (n432,n79,n65);
and (n433,n87,n70);
xnor (n434,n435,n88);
nor (n435,n436,n437);
and (n436,n95,n80);
and (n437,n103,n85);
and (n438,n434,n439);
xnor (n439,n440,n104);
nand (n440,n389,n101);
and (n441,n430,n439);
or (n442,n443,n452,n453);
and (n443,n444,n448);
xnor (n444,n445,n116);
nor (n445,n446,n447);
and (n446,n122,n114);
and (n447,n129,n117);
xnor (n448,n449,n130);
nor (n449,n450,n451);
and (n450,n14,n123);
and (n451,n23,n127);
and (n452,n448,n104);
and (n453,n444,n104);
and (n454,n442,n455);
or (n455,n456,n465,n470);
and (n456,n457,n461);
xnor (n457,n458,n24);
nor (n458,n459,n460);
and (n459,n30,n15);
and (n460,n38,n20);
xnor (n461,n462,n39);
nor (n462,n463,n464);
and (n463,n46,n31);
and (n464,n54,n36);
and (n465,n461,n466);
xnor (n466,n467,n55);
nor (n467,n468,n469);
and (n468,n64,n47);
and (n469,n72,n52);
and (n470,n457,n466);
and (n471,n428,n455);
or (n472,n473,n478,n480);
and (n473,n474,n476);
xor (n474,n475,n359);
xor (n475,n350,n354);
xor (n476,n477,n375);
xor (n477,n366,n370);
and (n478,n476,n479);
xor (n479,n382,n386);
and (n480,n474,n479);
and (n481,n472,n482);
xor (n482,n110,n119);
and (n483,n426,n482);
and (n484,n485,n487);
xor (n485,n486,n381);
xor (n486,n348,n364);
xor (n487,n488,n399);
xor (n488,n394,n396);
and (n489,n484,n490);
xor (n490,n491,n109);
xor (n491,n9,n59);
and (n492,n424,n490);
xor (n493,n494,n409);
xor (n494,n344,n406);
and (n495,n496,n497);
xor (n496,n419,n421);
or (n497,n498,n505);
and (n498,n499,n500);
xor (n499,n422,n493);
and (n500,n501,n503);
xor (n501,n502,n490);
xor (n502,n424,n484);
xor (n503,n504,n403);
xor (n504,n346,n392);
and (n505,n506,n507);
xor (n506,n499,n500);
or (n507,n508,n571);
and (n508,n509,n515);
xor (n509,n510,n513);
xor (n510,n490,n511);
xor (n511,n504,n512);
not (n512,n150);
xor (n513,n502,n514);
xnor (n514,n136,n161);
or (n515,n516,n568,n570);
and (n516,n517,n566);
or (n517,n518,n562,n565);
and (n518,n519,n557);
or (n519,n520,n553,n556);
and (n520,n521,n537);
or (n521,n522,n531,n536);
and (n522,n523,n527);
xnor (n523,n524,n116);
nor (n524,n525,n526);
and (n525,n23,n114);
and (n526,n122,n117);
xnor (n527,n528,n130);
nor (n528,n529,n530);
and (n529,n38,n123);
and (n530,n14,n127);
and (n531,n527,n532);
xnor (n532,n533,n24);
nor (n533,n534,n535);
and (n534,n54,n15);
and (n535,n30,n20);
and (n536,n523,n532);
or (n537,n538,n547,n552);
and (n538,n539,n543);
xnor (n539,n540,n39);
nor (n540,n541,n542);
and (n541,n72,n31);
and (n542,n46,n36);
xnor (n543,n544,n55);
nor (n544,n545,n546);
and (n545,n87,n47);
and (n546,n64,n52);
and (n547,n543,n548);
xnor (n548,n549,n73);
nor (n549,n550,n551);
and (n550,n103,n65);
and (n551,n79,n70);
and (n552,n539,n548);
and (n553,n537,n554);
xor (n554,n555,n439);
xor (n555,n430,n434);
and (n556,n521,n554);
and (n557,n558,n560);
xor (n558,n559,n104);
xor (n559,n444,n448);
xor (n560,n561,n466);
xor (n561,n457,n461);
and (n562,n557,n563);
xor (n563,n564,n479);
xor (n564,n474,n476);
and (n565,n519,n563);
xor (n566,n567,n482);
xor (n567,n426,n472);
and (n568,n566,n569);
xor (n569,n485,n487);
and (n570,n517,n569);
and (n571,n572,n573);
xor (n572,n509,n515);
or (n573,n574,n628);
and (n574,n575,n577);
xor (n575,n576,n569);
xor (n576,n517,n566);
or (n577,n578,n624,n627);
and (n578,n579,n622);
or (n579,n580,n619,n621);
and (n580,n581,n617);
or (n581,n582,n611,n616);
and (n582,n583,n595);
or (n583,n584,n593,n594);
and (n584,n585,n589);
xnor (n585,n586,n116);
nor (n586,n587,n588);
and (n587,n14,n114);
and (n588,n23,n117);
xnor (n589,n590,n130);
nor (n590,n591,n592);
and (n591,n30,n123);
and (n592,n38,n127);
and (n593,n589,n88);
and (n594,n585,n88);
or (n595,n596,n605,n610);
and (n596,n597,n601);
xnor (n597,n598,n24);
nor (n598,n599,n600);
and (n599,n46,n15);
and (n600,n54,n20);
xnor (n601,n602,n39);
nor (n602,n603,n604);
and (n603,n64,n31);
and (n604,n72,n36);
and (n605,n601,n606);
xnor (n606,n607,n55);
nor (n607,n608,n609);
and (n608,n79,n47);
and (n609,n87,n52);
and (n610,n597,n606);
and (n611,n595,n612);
xnor (n612,n613,n88);
nor (n613,n614,n615);
and (n614,n389,n80);
and (n615,n95,n85);
and (n616,n583,n612);
xor (n617,n618,n554);
xor (n618,n521,n537);
and (n619,n617,n620);
xor (n620,n558,n560);
and (n621,n581,n620);
xor (n622,n623,n455);
xor (n623,n428,n442);
and (n624,n622,n625);
xor (n625,n626,n563);
xor (n626,n519,n557);
and (n627,n579,n625);
and (n628,n629,n630);
xor (n629,n575,n577);
or (n630,n631,n701);
and (n631,n632,n634);
xor (n632,n633,n625);
xor (n633,n579,n622);
or (n634,n635,n697,n700);
and (n635,n636,n692);
or (n636,n637,n688,n691);
and (n637,n638,n678);
or (n638,n639,n672,n677);
and (n639,n640,n656);
or (n640,n641,n650,n655);
and (n641,n642,n646);
xnor (n642,n643,n39);
nor (n643,n644,n645);
and (n644,n87,n31);
and (n645,n64,n36);
xnor (n646,n647,n55);
nor (n647,n648,n649);
and (n648,n103,n47);
and (n649,n79,n52);
and (n650,n646,n651);
xnor (n651,n652,n73);
nor (n652,n653,n654);
and (n653,n389,n65);
and (n654,n95,n70);
and (n655,n642,n651);
or (n656,n657,n666,n671);
and (n657,n658,n662);
xnor (n658,n659,n116);
nor (n659,n660,n661);
and (n660,n38,n114);
and (n661,n14,n117);
xnor (n662,n663,n130);
nor (n663,n664,n665);
and (n664,n54,n123);
and (n665,n30,n127);
and (n666,n662,n667);
xnor (n667,n668,n24);
nor (n668,n669,n670);
and (n669,n72,n15);
and (n670,n46,n20);
and (n671,n658,n667);
and (n672,n656,n673);
xnor (n673,n674,n73);
nor (n674,n675,n676);
and (n675,n95,n65);
and (n676,n103,n70);
and (n677,n640,n673);
or (n678,n679,n684,n687);
and (n679,n680,n682);
xnor (n680,n681,n88);
nand (n681,n389,n85);
xor (n682,n683,n88);
xor (n683,n585,n589);
and (n684,n682,n685);
xor (n685,n686,n606);
xor (n686,n597,n601);
and (n687,n680,n685);
and (n688,n678,n689);
xor (n689,n690,n548);
xor (n690,n539,n543);
and (n691,n638,n689);
and (n692,n693,n695);
xor (n693,n694,n532);
xor (n694,n523,n527);
xor (n695,n696,n612);
xor (n696,n583,n595);
and (n697,n692,n698);
xor (n698,n699,n620);
xor (n699,n581,n617);
and (n700,n636,n698);
and (n701,n702,n703);
xor (n702,n632,n634);
or (n703,n704,n756);
and (n704,n705,n707);
xor (n705,n706,n698);
xor (n706,n636,n692);
or (n707,n708,n753,n755);
and (n708,n709,n751);
or (n709,n710,n747,n750);
and (n710,n711,n745);
or (n711,n712,n741,n744);
and (n712,n713,n729);
or (n713,n714,n723,n728);
and (n714,n715,n719);
xnor (n715,n716,n24);
nor (n716,n717,n718);
and (n717,n64,n15);
and (n718,n72,n20);
xnor (n719,n720,n39);
nor (n720,n721,n722);
and (n721,n79,n31);
and (n722,n87,n36);
and (n723,n719,n724);
xnor (n724,n725,n55);
nor (n725,n726,n727);
and (n726,n95,n47);
and (n727,n103,n52);
and (n728,n715,n724);
or (n729,n730,n739,n740);
and (n730,n731,n735);
xnor (n731,n732,n116);
nor (n732,n733,n734);
and (n733,n30,n114);
and (n734,n38,n117);
xnor (n735,n736,n130);
nor (n736,n737,n738);
and (n737,n46,n123);
and (n738,n54,n127);
and (n739,n735,n73);
and (n740,n731,n73);
and (n741,n729,n742);
xor (n742,n743,n651);
xor (n743,n642,n646);
and (n744,n713,n742);
xor (n745,n746,n673);
xor (n746,n640,n656);
and (n747,n745,n748);
xor (n748,n749,n685);
xor (n749,n680,n682);
and (n750,n711,n748);
xor (n751,n752,n689);
xor (n752,n638,n678);
and (n753,n751,n754);
xor (n754,n693,n695);
and (n755,n709,n754);
and (n756,n757,n758);
xor (n757,n705,n707);
or (n758,n759,n797);
and (n759,n760,n762);
xor (n760,n761,n754);
xor (n761,n709,n751);
and (n762,n763,n795);
or (n763,n764,n791,n794);
and (n764,n765,n789);
or (n765,n766,n785,n788);
and (n766,n767,n783);
or (n767,n768,n777,n782);
and (n768,n769,n773);
xnor (n769,n770,n116);
nor (n770,n771,n772);
and (n771,n54,n114);
and (n772,n30,n117);
xnor (n773,n774,n130);
nor (n774,n775,n776);
and (n775,n72,n123);
and (n776,n46,n127);
and (n777,n773,n778);
xnor (n778,n779,n24);
nor (n779,n780,n781);
and (n780,n87,n15);
and (n781,n64,n20);
and (n782,n769,n778);
xnor (n783,n784,n73);
nand (n784,n389,n70);
and (n785,n783,n786);
xor (n786,n787,n724);
xor (n787,n715,n719);
and (n788,n767,n786);
xor (n789,n790,n667);
xor (n790,n658,n662);
and (n791,n789,n792);
xor (n792,n793,n742);
xor (n793,n713,n729);
and (n794,n765,n792);
xor (n795,n796,n748);
xor (n796,n711,n745);
and (n797,n798,n799);
xor (n798,n760,n762);
or (n799,n800,n852);
and (n800,n801,n802);
xor (n801,n763,n795);
and (n802,n803,n850);
or (n803,n804,n846,n849);
and (n804,n805,n839);
or (n805,n806,n833,n838);
and (n806,n807,n821);
or (n807,n808,n817,n820);
and (n808,n809,n813);
xnor (n809,n810,n24);
nor (n810,n811,n812);
and (n811,n79,n15);
and (n812,n87,n20);
xnor (n813,n814,n39);
nor (n814,n815,n816);
and (n815,n95,n31);
and (n816,n103,n36);
and (n817,n813,n818);
xnor (n818,n819,n55);
nand (n819,n389,n52);
and (n820,n809,n818);
or (n821,n822,n831,n832);
and (n822,n823,n827);
xnor (n823,n824,n116);
nor (n824,n825,n826);
and (n825,n46,n114);
and (n826,n54,n117);
xnor (n827,n828,n130);
nor (n828,n829,n830);
and (n829,n64,n123);
and (n830,n72,n127);
and (n831,n827,n55);
and (n832,n823,n55);
and (n833,n821,n834);
xnor (n834,n835,n39);
nor (n835,n836,n837);
and (n836,n103,n31);
and (n837,n79,n36);
and (n838,n807,n834);
and (n839,n840,n844);
xnor (n840,n841,n55);
nor (n841,n842,n843);
and (n842,n389,n47);
and (n843,n95,n52);
xor (n844,n845,n778);
xor (n845,n769,n773);
and (n846,n839,n847);
xor (n847,n848,n73);
xor (n848,n731,n735);
and (n849,n805,n847);
xor (n850,n851,n792);
xor (n851,n765,n789);
and (n852,n853,n854);
xor (n853,n801,n802);
or (n854,n855,n862);
and (n855,n856,n857);
xor (n856,n803,n850);
and (n857,n858,n860);
xor (n858,n859,n786);
xor (n859,n767,n783);
xor (n860,n861,n847);
xor (n861,n805,n839);
and (n862,n863,n864);
xor (n863,n856,n857);
or (n864,n865,n898);
and (n865,n866,n867);
xor (n866,n858,n860);
or (n867,n868,n895,n897);
and (n868,n869,n893);
or (n869,n870,n889,n892);
and (n870,n871,n887);
or (n871,n872,n881,n886);
and (n872,n873,n877);
xnor (n873,n874,n116);
nor (n874,n875,n876);
and (n875,n72,n114);
and (n876,n46,n117);
xnor (n877,n878,n130);
nor (n878,n879,n880);
and (n879,n87,n123);
and (n880,n64,n127);
and (n881,n877,n882);
xnor (n882,n883,n24);
nor (n883,n884,n885);
and (n884,n103,n15);
and (n885,n79,n20);
and (n886,n873,n882);
xor (n887,n888,n818);
xor (n888,n809,n813);
and (n889,n887,n890);
xor (n890,n891,n55);
xor (n891,n823,n827);
and (n892,n871,n890);
xor (n893,n894,n834);
xor (n894,n807,n821);
and (n895,n893,n896);
xor (n896,n840,n844);
and (n897,n869,n896);
and (n898,n899,n900);
xor (n899,n866,n867);
or (n900,n901,n934);
and (n901,n902,n904);
xor (n902,n903,n896);
xor (n903,n869,n893);
and (n904,n905,n932);
or (n905,n906,n926,n931);
and (n906,n907,n919);
or (n907,n908,n917,n918);
and (n908,n909,n913);
xnor (n909,n910,n116);
nor (n910,n911,n912);
and (n911,n64,n114);
and (n912,n72,n117);
xnor (n913,n914,n130);
nor (n914,n915,n916);
and (n915,n79,n123);
and (n916,n87,n127);
and (n917,n913,n39);
and (n918,n909,n39);
and (n919,n920,n924);
xnor (n920,n921,n24);
nor (n921,n922,n923);
and (n922,n95,n15);
and (n923,n103,n20);
xnor (n924,n925,n39);
nand (n925,n389,n36);
and (n926,n919,n927);
xnor (n927,n928,n39);
nor (n928,n929,n930);
and (n929,n389,n31);
and (n930,n95,n36);
and (n931,n907,n927);
xor (n932,n933,n890);
xor (n933,n871,n887);
and (n934,n935,n936);
xor (n935,n902,n904);
or (n936,n937,n944);
and (n937,n938,n939);
xor (n938,n905,n932);
and (n939,n940,n942);
xor (n940,n941,n882);
xor (n941,n873,n877);
xor (n942,n943,n927);
xor (n943,n907,n919);
and (n944,n945,n946);
xor (n945,n938,n939);
or (n946,n947,n972);
and (n947,n948,n949);
xor (n948,n940,n942);
or (n949,n950,n969,n971);
and (n950,n951,n967);
or (n951,n952,n961,n966);
and (n952,n953,n957);
xnor (n953,n954,n116);
nor (n954,n955,n956);
and (n955,n87,n114);
and (n956,n64,n117);
xnor (n957,n958,n130);
nor (n958,n959,n960);
and (n959,n103,n123);
and (n960,n79,n127);
and (n961,n957,n962);
xnor (n962,n963,n24);
nor (n963,n964,n965);
and (n964,n389,n15);
and (n965,n95,n20);
and (n966,n953,n962);
xor (n967,n968,n39);
xor (n968,n909,n913);
and (n969,n967,n970);
xor (n970,n920,n924);
and (n971,n951,n970);
and (n972,n973,n974);
xor (n973,n948,n949);
or (n974,n975,n993);
and (n975,n976,n978);
xor (n976,n977,n970);
xor (n977,n951,n967);
and (n978,n979,n991);
or (n979,n980,n989,n990);
and (n980,n981,n985);
xnor (n981,n982,n116);
nor (n982,n983,n984);
and (n983,n79,n114);
and (n984,n87,n117);
xnor (n985,n986,n130);
nor (n986,n987,n988);
and (n987,n95,n123);
and (n988,n103,n127);
and (n989,n985,n24);
and (n990,n981,n24);
xor (n991,n992,n962);
xor (n992,n953,n957);
and (n993,n994,n995);
xor (n994,n976,n978);
or (n995,n996,n1003);
and (n996,n997,n998);
xor (n997,n979,n991);
and (n998,n999,n1001);
xnor (n999,n1000,n24);
nand (n1000,n389,n20);
xor (n1001,n1002,n24);
xor (n1002,n981,n985);
and (n1003,n1004,n1005);
xor (n1004,n997,n998);
or (n1005,n1006,n1017);
and (n1006,n1007,n1008);
xor (n1007,n999,n1001);
and (n1008,n1009,n1013);
xnor (n1009,n1010,n116);
nor (n1010,n1011,n1012);
and (n1011,n103,n114);
and (n1012,n79,n117);
xnor (n1013,n1014,n130);
nor (n1014,n1015,n1016);
and (n1015,n389,n123);
and (n1016,n95,n127);
and (n1017,n1018,n1019);
xor (n1018,n1007,n1008);
or (n1019,n1020,n1027);
and (n1020,n1021,n1022);
xor (n1021,n1009,n1013);
and (n1022,n1023,n130);
xnor (n1023,n1024,n116);
nor (n1024,n1025,n1026);
and (n1025,n95,n114);
and (n1026,n103,n117);
and (n1027,n1028,n1029);
xor (n1028,n1021,n1022);
or (n1029,n1030,n1034);
and (n1030,n1031,n1033);
xnor (n1031,n1032,n130);
nand (n1032,n389,n127);
xor (n1033,n1023,n130);
and (n1034,n1035,n1036);
xor (n1035,n1031,n1033);
and (n1036,n1037,n1041);
xnor (n1037,n1038,n116);
nor (n1038,n1039,n1040);
and (n1039,n389,n114);
and (n1040,n95,n117);
and (n1041,n1042,n116);
xnor (n1042,n1043,n116);
nand (n1043,n389,n117);
xor (n1044,n1045,n1127);
xor (n1045,n1046,n1113);
xor (n1046,n1047,n1084);
or (n1047,n1048,n1070,n1083);
and (n1048,n1049,n1061);
or (n1049,n1050,n1052,n1060);
and (n1050,n7,n1051);
or (n1051,n136,n161);
and (n1052,n1051,n1053);
xor (n1053,n1054,n1059);
xor (n1054,n1055,n1057);
xor (n1055,n1056,n214);
xor (n1056,n177,n180);
xor (n1057,n1058,n203);
xor (n1058,n218,n222);
xnor (n1059,n207,n211);
and (n1060,n7,n1053);
xor (n1061,n1062,n1069);
xor (n1062,n1063,n1066);
or (n1063,n231,n1064,n1065);
and (n1064,n180,n214);
and (n1065,n177,n214);
or (n1066,n239,n1067,n1068);
and (n1067,n222,n203);
and (n1068,n218,n203);
or (n1069,n207,n211);
and (n1070,n1061,n1071);
xor (n1071,n1072,n252);
xor (n1072,n1073,n1079);
or (n1073,n1074,n1078,n249);
and (n1074,n188,n1075);
or (n1075,n1076,n194,n1077);
and (n1076,n176,n152);
and (n1077,n176,n156);
and (n1078,n1075,n196);
or (n1079,n1080,n1081,n1082);
and (n1080,n1055,n1057);
and (n1081,n1057,n1059);
and (n1082,n1055,n1059);
and (n1083,n1049,n1071);
xor (n1084,n1085,n1096);
xor (n1085,n1086,n1090);
or (n1086,n1087,n1088,n1089);
and (n1087,n1073,n1079);
and (n1088,n1079,n252);
and (n1089,n1073,n252);
xor (n1090,n1091,n1095);
xor (n1091,n1092,n293);
or (n1092,n1093,n291,n1094);
and (n1093,n312,n257);
and (n1094,n312,n261);
and (n1095,n281,n285);
xor (n1096,n1097,n1106);
xor (n1097,n1098,n1102);
or (n1098,n1099,n1100,n1101);
and (n1099,n1063,n1066);
and (n1100,n1066,n1069);
and (n1101,n1063,n1069);
or (n1102,n1103,n1104,n1105);
and (n1103,n254,n265);
and (n1104,n265,n279);
and (n1105,n254,n279);
xor (n1106,n1107,n1112);
xor (n1107,n1108,n1110);
xor (n1108,n1109,n322);
xor (n1109,n313,n316);
xor (n1110,n1111,n335);
xor (n1111,n326,n330);
not (n1112,n339);
and (n1113,n1114,n1125);
or (n1114,n1115,n1121,n1124);
and (n1115,n1116,n1119);
or (n1116,n345,n1117,n1118);
and (n1117,n392,n512);
and (n1118,n346,n512);
xor (n1119,n1120,n196);
xor (n1120,n188,n1075);
and (n1121,n1119,n1122);
xor (n1122,n1123,n1053);
xor (n1123,n7,n1051);
and (n1124,n1116,n1122);
xor (n1125,n1126,n1071);
xor (n1126,n1049,n1061);
or (n1127,n1128,n1136);
and (n1128,n1129,n1130);
xor (n1129,n1114,n1125);
and (n1130,n1131,n1134);
or (n1131,n423,n1132,n1133);
and (n1132,n484,n514);
and (n1133,n424,n514);
xor (n1134,n1135,n1122);
xor (n1135,n1116,n1119);
and (n1136,n1137,n1138);
xor (n1137,n1129,n1130);
or (n1138,n1139,n505);
and (n1139,n1140,n1141);
xor (n1140,n1131,n1134);
or (n1141,n1142,n1143,n1144);
and (n1142,n490,n511);
and (n1143,n511,n513);
and (n1144,n490,n513);
endmodule
