module top (out,n10,n13,n15,n16,n21,n22,n32,n33,n35
        ,n38,n39,n44,n51,n99,n150,n257,n260,n265,n274
        ,n276,n279,n336,n386);
output out;
input n10;
input n13;
input n15;
input n16;
input n21;
input n22;
input n32;
input n33;
input n35;
input n38;
input n39;
input n44;
input n51;
input n99;
input n150;
input n257;
input n260;
input n265;
input n274;
input n276;
input n279;
input n336;
input n386;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n11;
wire n12;
wire n14;
wire n17;
wire n18;
wire n19;
wire n20;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n258;
wire n259;
wire n261;
wire n262;
wire n263;
wire n264;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n275;
wire n277;
wire n278;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
xor (out,n0,n540);
xor (n0,n1,n485);
xor (n1,n2,n249);
xor (n2,n3,n135);
xor (n3,n4,n92);
xor (n4,n5,n69);
xor (n5,n6,n25);
or (n6,n7,n17,n24);
and (n7,n8,n14);
nor (n8,n9,n11);
not (n9,n10);
and (n11,n12,n10);
not (n12,n13);
and (n14,n15,n16);
and (n17,n14,n18);
nor (n18,n19,n23);
and (n19,n20,n22);
not (n20,n21);
not (n23,n22);
and (n24,n8,n18);
or (n25,n26,n55,n68);
and (n26,n27,n53);
or (n27,n28,n47,n52);
and (n28,n29,n41);
or (n29,n30,n36,n40);
and (n30,n31,n34);
and (n31,n32,n33);
and (n34,n35,n22);
and (n36,n34,n37);
and (n37,n38,n39);
and (n40,n31,n37);
xor (n41,n42,n46);
xor (n42,n43,n45);
and (n43,n32,n44);
and (n45,n35,n33);
and (n46,n38,n22);
and (n47,n41,n48);
xor (n48,n49,n50);
and (n49,n10,n16);
and (n50,n15,n51);
and (n52,n29,n48);
xor (n53,n54,n18);
xor (n54,n8,n14);
and (n55,n53,n56);
xor (n56,n57,n63);
xor (n57,n58,n62);
or (n58,n59,n60,n61);
and (n59,n43,n45);
and (n60,n45,n46);
and (n61,n43,n46);
and (n62,n49,n50);
xor (n63,n64,n67);
xor (n64,n65,n66);
and (n65,n32,n51);
and (n66,n35,n44);
and (n67,n38,n33);
and (n68,n27,n56);
xor (n69,n70,n84);
xor (n70,n71,n75);
or (n71,n72,n73,n74);
and (n72,n58,n62);
and (n73,n62,n63);
and (n74,n58,n63);
xor (n75,n76,n81);
xor (n76,n77,n80);
nor (n77,n78,n79);
not (n78,n15);
and (n79,n12,n15);
and (n80,n32,n16);
nor (n81,n82,n83);
and (n82,n20,n33);
not (n83,n33);
xor (n84,n85,n91);
xor (n85,n86,n90);
or (n86,n87,n88,n89);
and (n87,n65,n66);
and (n88,n66,n67);
and (n89,n65,n67);
and (n90,n35,n51);
and (n91,n38,n44);
or (n92,n93,n131,n134);
and (n93,n94,n112);
or (n94,n95,n107,n111);
and (n95,n96,n104);
or (n96,n97,n101,n103);
and (n97,n98,n100);
and (n98,n99,n16);
and (n100,n10,n51);
and (n101,n100,n102);
and (n102,n15,n44);
and (n103,n98,n102);
nor (n104,n105,n106);
not (n105,n99);
and (n106,n12,n99);
and (n107,n104,n108);
nor (n108,n109,n110);
and (n109,n20,n39);
not (n110,n39);
and (n111,n96,n108);
or (n112,n113,n127,n130);
and (n113,n114,n125);
or (n114,n115,n121,n124);
and (n115,n116,n119);
and (n116,n117,n118);
and (n117,n32,n22);
and (n118,n35,n39);
xor (n119,n120,n102);
xor (n120,n98,n100);
and (n121,n119,n122);
xor (n122,n123,n37);
xor (n123,n31,n34);
and (n124,n116,n122);
xor (n125,n126,n108);
xor (n126,n96,n104);
and (n127,n125,n128);
xor (n128,n129,n48);
xor (n129,n29,n41);
and (n130,n114,n128);
and (n131,n112,n132);
xor (n132,n133,n56);
xor (n133,n27,n53);
and (n134,n94,n132);
or (n135,n136,n155);
and (n136,n137,n139);
xor (n137,n138,n132);
xor (n138,n94,n112);
and (n139,n140,n153);
or (n140,n141,n147,n152);
and (n141,n142,n145);
and (n142,n143,n144);
and (n143,n15,n33);
xor (n144,n117,n118);
xor (n145,n146,n122);
xor (n146,n116,n119);
and (n147,n145,n148);
nor (n148,n149,n151);
not (n149,n150);
and (n151,n12,n150);
and (n152,n142,n148);
xor (n153,n154,n128);
xor (n154,n114,n125);
and (n155,n156,n157);
xor (n156,n137,n139);
or (n157,n158,n188);
and (n158,n159,n160);
xor (n159,n140,n153);
or (n160,n161,n184,n187);
and (n161,n162,n169);
or (n162,n163,n166,n168);
and (n163,n164,n165);
and (n164,n150,n16);
and (n165,n99,n51);
and (n166,n165,n167);
and (n167,n10,n44);
and (n168,n164,n167);
or (n169,n170,n181,n183);
and (n170,n171,n179);
or (n171,n172,n175,n178);
and (n172,n173,n174);
and (n173,n10,n22);
and (n174,n15,n39);
and (n175,n176,n177);
and (n176,n15,n22);
and (n177,n32,n39);
and (n178,n172,n177);
xor (n179,n180,n167);
xor (n180,n164,n165);
and (n181,n179,n182);
xor (n182,n143,n144);
and (n183,n171,n182);
and (n184,n169,n185);
xor (n185,n186,n148);
xor (n186,n142,n145);
and (n187,n162,n185);
and (n188,n189,n190);
xor (n189,n159,n160);
or (n190,n191,n219);
and (n191,n192,n194);
xor (n192,n193,n185);
xor (n193,n162,n169);
or (n194,n195,n215,n218);
and (n195,n196,n199);
and (n196,n197,n198);
and (n197,n99,n44);
and (n198,n10,n33);
or (n199,n200,n211,n214);
and (n200,n201,n210);
or (n201,n202,n207,n209);
and (n202,n203,n206);
and (n203,n204,n205);
and (n204,n99,n22);
and (n205,n10,n39);
and (n206,n99,n33);
and (n207,n206,n208);
xor (n208,n173,n174);
and (n209,n203,n208);
xor (n210,n197,n198);
and (n211,n210,n212);
xor (n212,n213,n177);
xor (n213,n172,n176);
and (n214,n201,n212);
and (n215,n199,n216);
xor (n216,n217,n182);
xor (n217,n171,n179);
and (n218,n196,n216);
and (n219,n220,n221);
xor (n220,n192,n194);
or (n221,n222,n244);
and (n222,n223,n225);
xor (n223,n224,n216);
xor (n224,n196,n199);
and (n225,n226,n242);
or (n226,n227,n238,n241);
and (n227,n228,n237);
or (n228,n229,n234,n236);
and (n229,n230,n233);
and (n230,n231,n232);
and (n231,n150,n22);
and (n232,n99,n39);
and (n233,n150,n33);
and (n234,n233,n235);
xor (n235,n204,n205);
and (n236,n230,n235);
and (n237,n150,n44);
and (n238,n237,n239);
xor (n239,n240,n208);
xor (n240,n203,n206);
and (n241,n228,n239);
xor (n242,n243,n212);
xor (n243,n201,n210);
and (n244,n245,n246);
xor (n245,n223,n225);
and (n246,n247,n248);
and (n247,n150,n51);
xor (n248,n226,n242);
xor (n249,n250,n371);
xor (n250,n251,n329);
xor (n251,n252,n307);
xor (n252,n253,n267);
or (n253,n254,n261,n266);
and (n254,n255,n259);
nor (n255,n256,n258);
not (n256,n257);
and (n258,n12,n257);
and (n259,n260,n16);
and (n261,n259,n262);
nor (n262,n263,n23);
and (n263,n264,n22);
not (n264,n265);
and (n266,n255,n262);
or (n267,n268,n293,n306);
and (n268,n269,n291);
or (n269,n270,n286,n290);
and (n270,n271,n281);
or (n271,n272,n277,n280);
and (n272,n273,n275);
and (n273,n274,n33);
and (n275,n276,n22);
and (n277,n275,n278);
and (n278,n279,n39);
and (n280,n273,n278);
xor (n281,n282,n285);
xor (n282,n283,n284);
and (n283,n274,n44);
and (n284,n276,n33);
and (n285,n279,n22);
and (n286,n281,n287);
xor (n287,n288,n289);
and (n288,n257,n16);
and (n289,n260,n51);
and (n290,n271,n287);
xor (n291,n292,n262);
xor (n292,n255,n259);
and (n293,n291,n294);
xor (n294,n295,n301);
xor (n295,n296,n300);
or (n296,n297,n298,n299);
and (n297,n283,n284);
and (n298,n284,n285);
and (n299,n283,n285);
and (n300,n288,n289);
xor (n301,n302,n305);
xor (n302,n303,n304);
and (n303,n274,n51);
and (n304,n276,n44);
and (n305,n279,n33);
and (n306,n269,n294);
xor (n307,n308,n321);
xor (n308,n309,n313);
or (n309,n310,n311,n312);
and (n310,n296,n300);
and (n311,n300,n301);
and (n312,n296,n301);
xor (n313,n314,n319);
xor (n314,n315,n318);
nor (n315,n316,n317);
not (n316,n260);
and (n317,n12,n260);
and (n318,n274,n16);
nor (n319,n320,n83);
and (n320,n264,n33);
xor (n321,n322,n328);
xor (n322,n323,n327);
or (n323,n324,n325,n326);
and (n324,n303,n304);
and (n325,n304,n305);
and (n326,n303,n305);
and (n327,n276,n51);
and (n328,n279,n44);
or (n329,n330,n367,n370);
and (n330,n331,n348);
or (n331,n332,n344,n347);
and (n332,n333,n341);
or (n333,n334,n338,n340);
and (n334,n335,n337);
and (n335,n336,n16);
and (n337,n257,n51);
and (n338,n337,n339);
and (n339,n260,n44);
and (n340,n335,n339);
nor (n341,n342,n343);
not (n342,n336);
and (n343,n12,n336);
and (n344,n341,n345);
nor (n345,n346,n110);
and (n346,n264,n39);
and (n347,n333,n345);
or (n348,n349,n363,n366);
and (n349,n350,n361);
or (n350,n351,n357,n360);
and (n351,n352,n355);
and (n352,n353,n354);
and (n353,n274,n22);
and (n354,n276,n39);
xor (n355,n356,n339);
xor (n356,n335,n337);
and (n357,n355,n358);
xor (n358,n359,n278);
xor (n359,n273,n275);
and (n360,n352,n358);
xor (n361,n362,n345);
xor (n362,n333,n341);
and (n363,n361,n364);
xor (n364,n365,n287);
xor (n365,n271,n281);
and (n366,n350,n364);
and (n367,n348,n368);
xor (n368,n369,n294);
xor (n369,n269,n291);
and (n370,n331,n368);
or (n371,n372,n391);
and (n372,n373,n375);
xor (n373,n374,n368);
xor (n374,n331,n348);
and (n375,n376,n389);
or (n376,n377,n383,n388);
and (n377,n378,n381);
and (n378,n379,n380);
and (n379,n260,n33);
xor (n380,n353,n354);
xor (n381,n382,n358);
xor (n382,n352,n355);
and (n383,n381,n384);
nor (n384,n385,n387);
not (n385,n386);
and (n387,n12,n386);
and (n388,n378,n384);
xor (n389,n390,n364);
xor (n390,n350,n361);
and (n391,n392,n393);
xor (n392,n373,n375);
or (n393,n394,n424);
and (n394,n395,n396);
xor (n395,n376,n389);
or (n396,n397,n420,n423);
and (n397,n398,n405);
or (n398,n399,n402,n404);
and (n399,n400,n401);
and (n400,n386,n16);
and (n401,n336,n51);
and (n402,n401,n403);
and (n403,n257,n44);
and (n404,n400,n403);
or (n405,n406,n417,n419);
and (n406,n407,n415);
or (n407,n408,n411,n414);
and (n408,n409,n410);
and (n409,n257,n22);
and (n410,n260,n39);
and (n411,n412,n413);
and (n412,n260,n22);
and (n413,n274,n39);
and (n414,n408,n413);
xor (n415,n416,n403);
xor (n416,n400,n401);
and (n417,n415,n418);
xor (n418,n379,n380);
and (n419,n407,n418);
and (n420,n405,n421);
xor (n421,n422,n384);
xor (n422,n378,n381);
and (n423,n398,n421);
and (n424,n425,n426);
xor (n425,n395,n396);
or (n426,n427,n455);
and (n427,n428,n430);
xor (n428,n429,n421);
xor (n429,n398,n405);
or (n430,n431,n451,n454);
and (n431,n432,n435);
and (n432,n433,n434);
and (n433,n336,n44);
and (n434,n257,n33);
or (n435,n436,n447,n450);
and (n436,n437,n446);
or (n437,n438,n443,n445);
and (n438,n439,n442);
and (n439,n440,n441);
and (n440,n336,n22);
and (n441,n257,n39);
and (n442,n336,n33);
and (n443,n442,n444);
xor (n444,n409,n410);
and (n445,n439,n444);
xor (n446,n433,n434);
and (n447,n446,n448);
xor (n448,n449,n413);
xor (n449,n408,n412);
and (n450,n437,n448);
and (n451,n435,n452);
xor (n452,n453,n418);
xor (n453,n407,n415);
and (n454,n432,n452);
and (n455,n456,n457);
xor (n456,n428,n430);
or (n457,n458,n480);
and (n458,n459,n461);
xor (n459,n460,n452);
xor (n460,n432,n435);
and (n461,n462,n478);
or (n462,n463,n474,n477);
and (n463,n464,n473);
or (n464,n465,n470,n472);
and (n465,n466,n469);
and (n466,n467,n468);
and (n467,n386,n22);
and (n468,n336,n39);
and (n469,n386,n33);
and (n470,n469,n471);
xor (n471,n440,n441);
and (n472,n466,n471);
and (n473,n386,n44);
and (n474,n473,n475);
xor (n475,n476,n444);
xor (n476,n439,n442);
and (n477,n464,n475);
xor (n478,n479,n448);
xor (n479,n437,n446);
and (n480,n481,n482);
xor (n481,n459,n461);
and (n482,n483,n484);
and (n483,n386,n51);
xor (n484,n462,n478);
or (n485,n486,n489,n539);
and (n486,n487,n488);
xor (n487,n156,n157);
xor (n488,n392,n393);
and (n489,n488,n490);
or (n490,n491,n494,n538);
and (n491,n492,n493);
xor (n492,n189,n190);
xor (n493,n425,n426);
and (n494,n493,n495);
or (n495,n496,n499,n537);
and (n496,n497,n498);
xor (n497,n220,n221);
xor (n498,n456,n457);
and (n499,n498,n500);
or (n500,n501,n504,n536);
and (n501,n502,n503);
xor (n502,n245,n246);
xor (n503,n481,n482);
and (n504,n503,n505);
or (n505,n506,n509,n535);
and (n506,n507,n508);
xor (n507,n247,n248);
xor (n508,n483,n484);
and (n509,n508,n510);
or (n510,n511,n516,n534);
and (n511,n512,n514);
xor (n512,n513,n239);
xor (n513,n228,n237);
xor (n514,n515,n475);
xor (n515,n464,n473);
and (n516,n514,n517);
or (n517,n518,n523,n533);
and (n518,n519,n521);
xor (n519,n520,n235);
xor (n520,n230,n233);
xor (n521,n522,n471);
xor (n522,n466,n469);
and (n523,n521,n524);
or (n524,n525,n528,n532);
and (n525,n526,n527);
xor (n526,n231,n232);
xor (n527,n467,n468);
and (n528,n527,n529);
and (n529,n530,n531);
and (n530,n150,n39);
and (n531,n386,n39);
and (n532,n526,n529);
and (n533,n519,n524);
and (n534,n512,n517);
and (n535,n507,n510);
and (n536,n502,n505);
and (n537,n497,n500);
and (n538,n492,n495);
and (n539,n487,n490);
xor (n540,n541,n698);
xor (n541,n542,n664);
xor (n542,n543,n635);
xor (n543,n544,n590);
and (n544,n545,n571);
or (n545,n546,n562,n570);
and (n546,n547,n555);
and (n547,n548,n16);
xor (n548,n549,n550);
xor (n549,n10,n257);
or (n550,n551,n552,n554);
and (n551,n99,n336);
and (n552,n336,n553);
and (n553,n150,n386);
and (n554,n99,n553);
and (n555,n556,n51);
xor (n556,n557,n558);
xor (n557,n15,n260);
or (n558,n559,n560,n561);
and (n559,n10,n257);
and (n560,n257,n550);
and (n561,n10,n550);
and (n562,n555,n563);
and (n563,n564,n44);
xor (n564,n565,n566);
xor (n565,n32,n274);
or (n566,n567,n568,n569);
and (n567,n15,n260);
and (n568,n260,n558);
and (n569,n15,n558);
and (n570,n547,n563);
nor (n571,n572,n110);
and (n572,n573,n39);
not (n573,n574);
or (n574,n575,n576,n589);
and (n575,n21,n265);
and (n576,n265,n577);
or (n577,n578,n579,n588);
and (n578,n38,n279);
and (n579,n279,n580);
or (n580,n581,n582,n587);
and (n581,n35,n276);
and (n582,n276,n583);
or (n583,n584,n585,n586);
and (n584,n32,n274);
and (n585,n274,n566);
and (n586,n32,n566);
and (n587,n35,n583);
and (n588,n38,n580);
and (n589,n21,n577);
or (n590,n591,n632,n634);
and (n591,n592,n614);
or (n592,n593,n610,n613);
and (n593,n594,n599);
nor (n594,n595,n598);
not (n595,n596);
xor (n596,n597,n553);
xor (n597,n99,n336);
and (n598,n12,n596);
xor (n599,n600,n607);
xor (n600,n601,n604);
and (n601,n602,n33);
xor (n602,n603,n583);
xor (n603,n35,n276);
and (n604,n605,n22);
xor (n605,n606,n580);
xor (n606,n38,n279);
and (n607,n608,n39);
xor (n608,n609,n577);
xor (n609,n21,n265);
and (n610,n599,n611);
xor (n611,n612,n563);
xor (n612,n547,n555);
and (n613,n594,n611);
xor (n614,n615,n625);
xor (n615,n616,n620);
or (n616,n617,n618,n619);
and (n617,n601,n604);
and (n618,n604,n607);
and (n619,n601,n607);
xor (n620,n621,n624);
xor (n621,n622,n623);
and (n622,n602,n44);
and (n623,n605,n33);
and (n624,n608,n22);
xor (n625,n626,n631);
xor (n626,n627,n630);
nor (n627,n628,n629);
not (n628,n548);
and (n629,n12,n548);
and (n630,n556,n16);
and (n631,n564,n51);
and (n632,n614,n633);
xor (n633,n545,n571);
and (n634,n592,n633);
xor (n635,n636,n649);
xor (n636,n637,n641);
or (n637,n638,n639,n640);
and (n638,n616,n620);
and (n639,n620,n625);
and (n640,n616,n625);
xor (n641,n642,n647);
xor (n642,n643,n646);
nor (n643,n644,n645);
not (n644,n556);
and (n645,n12,n556);
and (n646,n564,n16);
nor (n647,n648,n23);
and (n648,n573,n22);
xor (n649,n650,n659);
xor (n650,n651,n655);
or (n651,n652,n653,n654);
and (n652,n622,n623);
and (n653,n623,n624);
and (n654,n622,n624);
or (n655,n656,n657,n658);
and (n656,n627,n630);
and (n657,n630,n631);
and (n658,n627,n631);
xor (n659,n660,n663);
xor (n660,n661,n662);
and (n661,n602,n51);
and (n662,n605,n44);
and (n663,n608,n33);
or (n664,n665,n694,n697);
and (n665,n666,n677);
and (n666,n667,n674);
or (n667,n668,n671,n673);
and (n668,n669,n670);
and (n669,n548,n51);
and (n670,n556,n44);
and (n671,n670,n672);
and (n672,n564,n33);
and (n673,n669,n672);
and (n674,n675,n676);
and (n675,n602,n22);
and (n676,n605,n39);
or (n677,n678,n690,n693);
and (n678,n679,n689);
or (n679,n680,n686,n688);
and (n680,n681,n684);
and (n681,n682,n683);
and (n682,n564,n22);
and (n683,n602,n39);
xor (n684,n685,n672);
xor (n685,n669,n670);
and (n686,n684,n687);
xor (n687,n675,n676);
and (n688,n681,n687);
xor (n689,n667,n674);
and (n690,n689,n691);
xor (n691,n692,n611);
xor (n692,n594,n599);
and (n693,n679,n691);
and (n694,n677,n695);
xor (n695,n696,n633);
xor (n696,n592,n614);
and (n697,n666,n695);
or (n698,n699,n724);
and (n699,n700,n702);
xor (n700,n701,n695);
xor (n701,n666,n677);
or (n702,n703,n720,n723);
and (n703,n704,n710);
and (n704,n705,n709);
nor (n705,n706,n708);
not (n706,n707);
xor (n707,n150,n386);
and (n708,n12,n707);
and (n709,n596,n16);
or (n710,n711,n717,n719);
and (n711,n712,n715);
and (n712,n713,n714);
and (n713,n556,n33);
xor (n714,n682,n683);
xor (n715,n716,n687);
xor (n716,n681,n684);
and (n717,n715,n718);
xor (n718,n705,n709);
and (n719,n712,n718);
and (n720,n710,n721);
xor (n721,n722,n691);
xor (n722,n679,n689);
and (n723,n704,n721);
and (n724,n725,n726);
xor (n725,n700,n702);
or (n726,n727,n758);
and (n727,n728,n730);
xor (n728,n729,n721);
xor (n729,n704,n710);
or (n730,n731,n754,n757);
and (n731,n732,n739);
or (n732,n733,n736,n738);
and (n733,n734,n735);
and (n734,n707,n16);
and (n735,n596,n51);
and (n736,n735,n737);
and (n737,n548,n44);
and (n738,n734,n737);
or (n739,n740,n751,n753);
and (n740,n741,n749);
or (n741,n742,n745,n748);
and (n742,n743,n744);
and (n743,n548,n22);
and (n744,n556,n39);
and (n745,n746,n747);
and (n746,n556,n22);
and (n747,n564,n39);
and (n748,n742,n747);
xor (n749,n750,n737);
xor (n750,n734,n735);
and (n751,n749,n752);
xor (n752,n713,n714);
and (n753,n741,n752);
and (n754,n739,n755);
xor (n755,n756,n718);
xor (n756,n712,n715);
and (n757,n732,n755);
and (n758,n759,n760);
xor (n759,n728,n730);
or (n760,n761,n789);
and (n761,n762,n764);
xor (n762,n763,n755);
xor (n763,n732,n739);
or (n764,n765,n785,n788);
and (n765,n766,n769);
and (n766,n767,n768);
and (n767,n596,n44);
and (n768,n548,n33);
or (n769,n770,n781,n784);
and (n770,n771,n780);
or (n771,n772,n777,n779);
and (n772,n773,n776);
and (n773,n774,n775);
and (n774,n596,n22);
and (n775,n548,n39);
and (n776,n596,n33);
and (n777,n776,n778);
xor (n778,n743,n744);
and (n779,n773,n778);
xor (n780,n767,n768);
and (n781,n780,n782);
xor (n782,n783,n747);
xor (n783,n742,n746);
and (n784,n771,n782);
and (n785,n769,n786);
xor (n786,n787,n752);
xor (n787,n741,n749);
and (n788,n766,n786);
and (n789,n790,n791);
xor (n790,n762,n764);
or (n791,n792,n814);
and (n792,n793,n795);
xor (n793,n794,n786);
xor (n794,n766,n769);
and (n795,n796,n812);
or (n796,n797,n808,n811);
and (n797,n798,n807);
or (n798,n799,n804,n806);
and (n799,n800,n803);
and (n800,n801,n802);
and (n801,n707,n22);
and (n802,n596,n39);
and (n803,n707,n33);
and (n804,n803,n805);
xor (n805,n774,n775);
and (n806,n800,n805);
and (n807,n707,n44);
and (n808,n807,n809);
xor (n809,n810,n778);
xor (n810,n773,n776);
and (n811,n798,n809);
xor (n812,n813,n782);
xor (n813,n771,n780);
and (n814,n815,n816);
xor (n815,n793,n795);
and (n816,n817,n818);
and (n817,n707,n51);
xor (n818,n796,n812);
endmodule
