module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n160,n213,n260,n301
        ,n336,n365,n388,n405,n416,n442,n443,n447,n449,n456
        ,n463,n470,n477,n484,n491,n498,n505,n512,n518,n520
        ,n579,n632,n679,n720,n755,n784,n807,n824,n835,n839);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n160;
input n213;
input n260;
input n301;
input n336;
input n365;
input n388;
input n405;
input n416;
input n442;
input n443;
input n447;
input n449;
input n456;
input n463;
input n470;
input n477;
input n484;
input n491;
input n498;
input n505;
input n512;
input n518;
input n520;
input n579;
input n632;
input n679;
input n720;
input n755;
input n784;
input n807;
input n824;
input n835;
input n839;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n444;
wire n445;
wire n446;
wire n448;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n519;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n836;
wire n837;
wire n838;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
xor (out,n0,n840);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n839);
and (s0n0,notn0,n1);
and (s1n0,n839,n420);
xor (n1,n2,n417);
xor (n2,n3,n415);
xor (n3,n4,n406);
xor (n4,n5,n404);
xor (n5,n6,n389);
xor (n6,n7,n387);
xor (n7,n8,n366);
xor (n8,n9,n364);
xor (n9,n10,n337);
xor (n10,n11,n335);
xor (n11,n12,n302);
xor (n12,n13,n300);
xor (n13,n14,n261);
xor (n14,n15,n259);
xor (n15,n16,n214);
xor (n16,n17,n212);
xor (n17,n18,n161);
xor (n18,n19,n159);
xor (n19,n20,n102);
xor (n20,n21,n100);
xor (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n30,n101);
or (n102,n103,n106);
and (n103,n104,n105);
xor (n104,n32,n33);
and (n105,n37,n101);
and (n106,n107,n108);
xor (n107,n104,n105);
or (n108,n109,n112);
and (n109,n110,n111);
xor (n110,n39,n40);
and (n111,n44,n101);
and (n112,n113,n114);
xor (n113,n110,n111);
or (n114,n115,n118);
and (n115,n116,n117);
xor (n116,n46,n47);
and (n117,n51,n101);
and (n118,n119,n120);
xor (n119,n116,n117);
or (n120,n121,n124);
and (n121,n122,n123);
xor (n122,n53,n54);
and (n123,n58,n101);
and (n124,n125,n126);
xor (n125,n122,n123);
or (n126,n127,n130);
and (n127,n128,n129);
xor (n128,n60,n61);
and (n129,n65,n101);
and (n130,n131,n132);
xor (n131,n128,n129);
or (n132,n133,n136);
and (n133,n134,n135);
xor (n134,n67,n68);
and (n135,n72,n101);
and (n136,n137,n138);
xor (n137,n134,n135);
or (n138,n139,n142);
and (n139,n140,n141);
xor (n140,n74,n75);
and (n141,n79,n101);
and (n142,n143,n144);
xor (n143,n140,n141);
or (n144,n145,n148);
and (n145,n146,n147);
xor (n146,n81,n82);
and (n147,n86,n101);
and (n148,n149,n150);
xor (n149,n146,n147);
or (n150,n151,n154);
and (n151,n152,n153);
xor (n152,n88,n89);
and (n153,n93,n101);
and (n154,n155,n156);
xor (n155,n152,n153);
and (n156,n157,n158);
xor (n157,n95,n96);
and (n158,n99,n101);
and (n159,n37,n160);
or (n161,n162,n165);
and (n162,n163,n164);
xor (n163,n107,n108);
and (n164,n44,n160);
and (n165,n166,n167);
xor (n166,n163,n164);
or (n167,n168,n171);
and (n168,n169,n170);
xor (n169,n113,n114);
and (n170,n51,n160);
and (n171,n172,n173);
xor (n172,n169,n170);
or (n173,n174,n177);
and (n174,n175,n176);
xor (n175,n119,n120);
and (n176,n58,n160);
and (n177,n178,n179);
xor (n178,n175,n176);
or (n179,n180,n183);
and (n180,n181,n182);
xor (n181,n125,n126);
and (n182,n65,n160);
and (n183,n184,n185);
xor (n184,n181,n182);
or (n185,n186,n189);
and (n186,n187,n188);
xor (n187,n131,n132);
and (n188,n72,n160);
and (n189,n190,n191);
xor (n190,n187,n188);
or (n191,n192,n195);
and (n192,n193,n194);
xor (n193,n137,n138);
and (n194,n79,n160);
and (n195,n196,n197);
xor (n196,n193,n194);
or (n197,n198,n201);
and (n198,n199,n200);
xor (n199,n143,n144);
and (n200,n86,n160);
and (n201,n202,n203);
xor (n202,n199,n200);
or (n203,n204,n207);
and (n204,n205,n206);
xor (n205,n149,n150);
and (n206,n93,n160);
and (n207,n208,n209);
xor (n208,n205,n206);
and (n209,n210,n211);
xor (n210,n155,n156);
and (n211,n99,n160);
and (n212,n44,n213);
or (n214,n215,n218);
and (n215,n216,n217);
xor (n216,n166,n167);
and (n217,n51,n213);
and (n218,n219,n220);
xor (n219,n216,n217);
or (n220,n221,n224);
and (n221,n222,n223);
xor (n222,n172,n173);
and (n223,n58,n213);
and (n224,n225,n226);
xor (n225,n222,n223);
or (n226,n227,n230);
and (n227,n228,n229);
xor (n228,n178,n179);
and (n229,n65,n213);
and (n230,n231,n232);
xor (n231,n228,n229);
or (n232,n233,n236);
and (n233,n234,n235);
xor (n234,n184,n185);
and (n235,n72,n213);
and (n236,n237,n238);
xor (n237,n234,n235);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n190,n191);
and (n241,n79,n213);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n196,n197);
and (n247,n86,n213);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n202,n203);
and (n253,n93,n213);
and (n254,n255,n256);
xor (n255,n252,n253);
and (n256,n257,n258);
xor (n257,n208,n209);
and (n258,n99,n213);
and (n259,n51,n260);
or (n261,n262,n265);
and (n262,n263,n264);
xor (n263,n219,n220);
and (n264,n58,n260);
and (n265,n266,n267);
xor (n266,n263,n264);
or (n267,n268,n271);
and (n268,n269,n270);
xor (n269,n225,n226);
and (n270,n65,n260);
and (n271,n272,n273);
xor (n272,n269,n270);
or (n273,n274,n277);
and (n274,n275,n276);
xor (n275,n231,n232);
and (n276,n72,n260);
and (n277,n278,n279);
xor (n278,n275,n276);
or (n279,n280,n283);
and (n280,n281,n282);
xor (n281,n237,n238);
and (n282,n79,n260);
and (n283,n284,n285);
xor (n284,n281,n282);
or (n285,n286,n289);
and (n286,n287,n288);
xor (n287,n243,n244);
and (n288,n86,n260);
and (n289,n290,n291);
xor (n290,n287,n288);
or (n291,n292,n295);
and (n292,n293,n294);
xor (n293,n249,n250);
and (n294,n93,n260);
and (n295,n296,n297);
xor (n296,n293,n294);
and (n297,n298,n299);
xor (n298,n255,n256);
and (n299,n99,n260);
and (n300,n58,n301);
or (n302,n303,n306);
and (n303,n304,n305);
xor (n304,n266,n267);
and (n305,n65,n301);
and (n306,n307,n308);
xor (n307,n304,n305);
or (n308,n309,n312);
and (n309,n310,n311);
xor (n310,n272,n273);
and (n311,n72,n301);
and (n312,n313,n314);
xor (n313,n310,n311);
or (n314,n315,n318);
and (n315,n316,n317);
xor (n316,n278,n279);
and (n317,n79,n301);
and (n318,n319,n320);
xor (n319,n316,n317);
or (n320,n321,n324);
and (n321,n322,n323);
xor (n322,n284,n285);
and (n323,n86,n301);
and (n324,n325,n326);
xor (n325,n322,n323);
or (n326,n327,n330);
and (n327,n328,n329);
xor (n328,n290,n291);
and (n329,n93,n301);
and (n330,n331,n332);
xor (n331,n328,n329);
and (n332,n333,n334);
xor (n333,n296,n297);
and (n334,n99,n301);
and (n335,n65,n336);
or (n337,n338,n341);
and (n338,n339,n340);
xor (n339,n307,n308);
and (n340,n72,n336);
and (n341,n342,n343);
xor (n342,n339,n340);
or (n343,n344,n347);
and (n344,n345,n346);
xor (n345,n313,n314);
and (n346,n79,n336);
and (n347,n348,n349);
xor (n348,n345,n346);
or (n349,n350,n353);
and (n350,n351,n352);
xor (n351,n319,n320);
and (n352,n86,n336);
and (n353,n354,n355);
xor (n354,n351,n352);
or (n355,n356,n359);
and (n356,n357,n358);
xor (n357,n325,n326);
and (n358,n93,n336);
and (n359,n360,n361);
xor (n360,n357,n358);
and (n361,n362,n363);
xor (n362,n331,n332);
and (n363,n99,n336);
and (n364,n72,n365);
or (n366,n367,n370);
and (n367,n368,n369);
xor (n368,n342,n343);
and (n369,n79,n365);
and (n370,n371,n372);
xor (n371,n368,n369);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n348,n349);
and (n375,n86,n365);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n354,n355);
and (n381,n93,n365);
and (n382,n383,n384);
xor (n383,n380,n381);
and (n384,n385,n386);
xor (n385,n360,n361);
and (n386,n99,n365);
and (n387,n79,n388);
or (n389,n390,n393);
and (n390,n391,n392);
xor (n391,n371,n372);
and (n392,n86,n388);
and (n393,n394,n395);
xor (n394,n391,n392);
or (n395,n396,n399);
and (n396,n397,n398);
xor (n397,n377,n378);
and (n398,n93,n388);
and (n399,n400,n401);
xor (n400,n397,n398);
and (n401,n402,n403);
xor (n402,n383,n384);
and (n403,n99,n388);
and (n404,n86,n405);
or (n406,n407,n410);
and (n407,n408,n409);
xor (n408,n394,n395);
and (n409,n93,n405);
and (n410,n411,n412);
xor (n411,n408,n409);
and (n412,n413,n414);
xor (n413,n400,n401);
and (n414,n99,n405);
and (n415,n93,n416);
and (n417,n418,n419);
xor (n418,n411,n412);
and (n419,n99,n416);
xor (n420,n421,n836);
xor (n421,n422,n834);
xor (n422,n423,n825);
xor (n423,n424,n823);
xor (n424,n425,n808);
xor (n425,n426,n806);
xor (n426,n427,n785);
xor (n427,n428,n783);
xor (n428,n429,n756);
xor (n429,n430,n754);
xor (n430,n431,n721);
xor (n431,n432,n719);
xor (n432,n433,n680);
xor (n433,n434,n678);
xor (n434,n435,n633);
xor (n435,n436,n631);
xor (n436,n437,n580);
xor (n437,n438,n578);
xor (n438,n439,n521);
xor (n439,n440,n519);
xor (n440,n441,n444);
and (n441,n442,n443);
or (n444,n445,n450);
and (n445,n446,n448);
and (n446,n442,n447);
and (n448,n449,n443);
and (n450,n451,n452);
xor (n451,n446,n448);
or (n452,n453,n457);
and (n453,n454,n455);
and (n454,n449,n447);
and (n455,n456,n443);
and (n457,n458,n459);
xor (n458,n454,n455);
or (n459,n460,n464);
and (n460,n461,n462);
and (n461,n456,n447);
and (n462,n463,n443);
and (n464,n465,n466);
xor (n465,n461,n462);
or (n466,n467,n471);
and (n467,n468,n469);
and (n468,n463,n447);
and (n469,n470,n443);
and (n471,n472,n473);
xor (n472,n468,n469);
or (n473,n474,n478);
and (n474,n475,n476);
and (n475,n470,n447);
and (n476,n477,n443);
and (n478,n479,n480);
xor (n479,n475,n476);
or (n480,n481,n485);
and (n481,n482,n483);
and (n482,n477,n447);
and (n483,n484,n443);
and (n485,n486,n487);
xor (n486,n482,n483);
or (n487,n488,n492);
and (n488,n489,n490);
and (n489,n484,n447);
and (n490,n491,n443);
and (n492,n493,n494);
xor (n493,n489,n490);
or (n494,n495,n499);
and (n495,n496,n497);
and (n496,n491,n447);
and (n497,n498,n443);
and (n499,n500,n501);
xor (n500,n496,n497);
or (n501,n502,n506);
and (n502,n503,n504);
and (n503,n498,n447);
and (n504,n505,n443);
and (n506,n507,n508);
xor (n507,n503,n504);
or (n508,n509,n513);
and (n509,n510,n511);
and (n510,n505,n447);
and (n511,n512,n443);
and (n513,n514,n515);
xor (n514,n510,n511);
and (n515,n516,n517);
and (n516,n512,n447);
and (n517,n518,n443);
and (n519,n449,n520);
or (n521,n522,n525);
and (n522,n523,n524);
xor (n523,n451,n452);
and (n524,n456,n520);
and (n525,n526,n527);
xor (n526,n523,n524);
or (n527,n528,n531);
and (n528,n529,n530);
xor (n529,n458,n459);
and (n530,n463,n520);
and (n531,n532,n533);
xor (n532,n529,n530);
or (n533,n534,n537);
and (n534,n535,n536);
xor (n535,n465,n466);
and (n536,n470,n520);
and (n537,n538,n539);
xor (n538,n535,n536);
or (n539,n540,n543);
and (n540,n541,n542);
xor (n541,n472,n473);
and (n542,n477,n520);
and (n543,n544,n545);
xor (n544,n541,n542);
or (n545,n546,n549);
and (n546,n547,n548);
xor (n547,n479,n480);
and (n548,n484,n520);
and (n549,n550,n551);
xor (n550,n547,n548);
or (n551,n552,n555);
and (n552,n553,n554);
xor (n553,n486,n487);
and (n554,n491,n520);
and (n555,n556,n557);
xor (n556,n553,n554);
or (n557,n558,n561);
and (n558,n559,n560);
xor (n559,n493,n494);
and (n560,n498,n520);
and (n561,n562,n563);
xor (n562,n559,n560);
or (n563,n564,n567);
and (n564,n565,n566);
xor (n565,n500,n501);
and (n566,n505,n520);
and (n567,n568,n569);
xor (n568,n565,n566);
or (n569,n570,n573);
and (n570,n571,n572);
xor (n571,n507,n508);
and (n572,n512,n520);
and (n573,n574,n575);
xor (n574,n571,n572);
and (n575,n576,n577);
xor (n576,n514,n515);
and (n577,n518,n520);
and (n578,n456,n579);
or (n580,n581,n584);
and (n581,n582,n583);
xor (n582,n526,n527);
and (n583,n463,n579);
and (n584,n585,n586);
xor (n585,n582,n583);
or (n586,n587,n590);
and (n587,n588,n589);
xor (n588,n532,n533);
and (n589,n470,n579);
and (n590,n591,n592);
xor (n591,n588,n589);
or (n592,n593,n596);
and (n593,n594,n595);
xor (n594,n538,n539);
and (n595,n477,n579);
and (n596,n597,n598);
xor (n597,n594,n595);
or (n598,n599,n602);
and (n599,n600,n601);
xor (n600,n544,n545);
and (n601,n484,n579);
and (n602,n603,n604);
xor (n603,n600,n601);
or (n604,n605,n608);
and (n605,n606,n607);
xor (n606,n550,n551);
and (n607,n491,n579);
and (n608,n609,n610);
xor (n609,n606,n607);
or (n610,n611,n614);
and (n611,n612,n613);
xor (n612,n556,n557);
and (n613,n498,n579);
and (n614,n615,n616);
xor (n615,n612,n613);
or (n616,n617,n620);
and (n617,n618,n619);
xor (n618,n562,n563);
and (n619,n505,n579);
and (n620,n621,n622);
xor (n621,n618,n619);
or (n622,n623,n626);
and (n623,n624,n625);
xor (n624,n568,n569);
and (n625,n512,n579);
and (n626,n627,n628);
xor (n627,n624,n625);
and (n628,n629,n630);
xor (n629,n574,n575);
and (n630,n518,n579);
and (n631,n463,n632);
or (n633,n634,n637);
and (n634,n635,n636);
xor (n635,n585,n586);
and (n636,n470,n632);
and (n637,n638,n639);
xor (n638,n635,n636);
or (n639,n640,n643);
and (n640,n641,n642);
xor (n641,n591,n592);
and (n642,n477,n632);
and (n643,n644,n645);
xor (n644,n641,n642);
or (n645,n646,n649);
and (n646,n647,n648);
xor (n647,n597,n598);
and (n648,n484,n632);
and (n649,n650,n651);
xor (n650,n647,n648);
or (n651,n652,n655);
and (n652,n653,n654);
xor (n653,n603,n604);
and (n654,n491,n632);
and (n655,n656,n657);
xor (n656,n653,n654);
or (n657,n658,n661);
and (n658,n659,n660);
xor (n659,n609,n610);
and (n660,n498,n632);
and (n661,n662,n663);
xor (n662,n659,n660);
or (n663,n664,n667);
and (n664,n665,n666);
xor (n665,n615,n616);
and (n666,n505,n632);
and (n667,n668,n669);
xor (n668,n665,n666);
or (n669,n670,n673);
and (n670,n671,n672);
xor (n671,n621,n622);
and (n672,n512,n632);
and (n673,n674,n675);
xor (n674,n671,n672);
and (n675,n676,n677);
xor (n676,n627,n628);
and (n677,n518,n632);
and (n678,n470,n679);
or (n680,n681,n684);
and (n681,n682,n683);
xor (n682,n638,n639);
and (n683,n477,n679);
and (n684,n685,n686);
xor (n685,n682,n683);
or (n686,n687,n690);
and (n687,n688,n689);
xor (n688,n644,n645);
and (n689,n484,n679);
and (n690,n691,n692);
xor (n691,n688,n689);
or (n692,n693,n696);
and (n693,n694,n695);
xor (n694,n650,n651);
and (n695,n491,n679);
and (n696,n697,n698);
xor (n697,n694,n695);
or (n698,n699,n702);
and (n699,n700,n701);
xor (n700,n656,n657);
and (n701,n498,n679);
and (n702,n703,n704);
xor (n703,n700,n701);
or (n704,n705,n708);
and (n705,n706,n707);
xor (n706,n662,n663);
and (n707,n505,n679);
and (n708,n709,n710);
xor (n709,n706,n707);
or (n710,n711,n714);
and (n711,n712,n713);
xor (n712,n668,n669);
and (n713,n512,n679);
and (n714,n715,n716);
xor (n715,n712,n713);
and (n716,n717,n718);
xor (n717,n674,n675);
and (n718,n518,n679);
and (n719,n477,n720);
or (n721,n722,n725);
and (n722,n723,n724);
xor (n723,n685,n686);
and (n724,n484,n720);
and (n725,n726,n727);
xor (n726,n723,n724);
or (n727,n728,n731);
and (n728,n729,n730);
xor (n729,n691,n692);
and (n730,n491,n720);
and (n731,n732,n733);
xor (n732,n729,n730);
or (n733,n734,n737);
and (n734,n735,n736);
xor (n735,n697,n698);
and (n736,n498,n720);
and (n737,n738,n739);
xor (n738,n735,n736);
or (n739,n740,n743);
and (n740,n741,n742);
xor (n741,n703,n704);
and (n742,n505,n720);
and (n743,n744,n745);
xor (n744,n741,n742);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n709,n710);
and (n748,n512,n720);
and (n749,n750,n751);
xor (n750,n747,n748);
and (n751,n752,n753);
xor (n752,n715,n716);
and (n753,n518,n720);
and (n754,n484,n755);
or (n756,n757,n760);
and (n757,n758,n759);
xor (n758,n726,n727);
and (n759,n491,n755);
and (n760,n761,n762);
xor (n761,n758,n759);
or (n762,n763,n766);
and (n763,n764,n765);
xor (n764,n732,n733);
and (n765,n498,n755);
and (n766,n767,n768);
xor (n767,n764,n765);
or (n768,n769,n772);
and (n769,n770,n771);
xor (n770,n738,n739);
and (n771,n505,n755);
and (n772,n773,n774);
xor (n773,n770,n771);
or (n774,n775,n778);
and (n775,n776,n777);
xor (n776,n744,n745);
and (n777,n512,n755);
and (n778,n779,n780);
xor (n779,n776,n777);
and (n780,n781,n782);
xor (n781,n750,n751);
and (n782,n518,n755);
and (n783,n491,n784);
or (n785,n786,n789);
and (n786,n787,n788);
xor (n787,n761,n762);
and (n788,n498,n784);
and (n789,n790,n791);
xor (n790,n787,n788);
or (n791,n792,n795);
and (n792,n793,n794);
xor (n793,n767,n768);
and (n794,n505,n784);
and (n795,n796,n797);
xor (n796,n793,n794);
or (n797,n798,n801);
and (n798,n799,n800);
xor (n799,n773,n774);
and (n800,n512,n784);
and (n801,n802,n803);
xor (n802,n799,n800);
and (n803,n804,n805);
xor (n804,n779,n780);
and (n805,n518,n784);
and (n806,n498,n807);
or (n808,n809,n812);
and (n809,n810,n811);
xor (n810,n790,n791);
and (n811,n505,n807);
and (n812,n813,n814);
xor (n813,n810,n811);
or (n814,n815,n818);
and (n815,n816,n817);
xor (n816,n796,n797);
and (n817,n512,n807);
and (n818,n819,n820);
xor (n819,n816,n817);
and (n820,n821,n822);
xor (n821,n802,n803);
and (n822,n518,n807);
and (n823,n505,n824);
or (n825,n826,n829);
and (n826,n827,n828);
xor (n827,n813,n814);
and (n828,n512,n824);
and (n829,n830,n831);
xor (n830,n827,n828);
and (n831,n832,n833);
xor (n832,n819,n820);
and (n833,n518,n824);
and (n834,n512,n835);
and (n836,n837,n838);
xor (n837,n830,n831);
and (n838,n518,n835);
xor (n840,n841,n1256);
xor (n841,n842,n1254);
xor (n842,n843,n1245);
xor (n843,n844,n1243);
xor (n844,n845,n1228);
xor (n845,n846,n1226);
xor (n846,n847,n1205);
xor (n847,n848,n1203);
xor (n848,n849,n1176);
xor (n849,n850,n1174);
xor (n850,n851,n1141);
xor (n851,n852,n1139);
xor (n852,n853,n1100);
xor (n853,n854,n1098);
xor (n854,n855,n1053);
xor (n855,n856,n1051);
xor (n856,n857,n1000);
xor (n857,n858,n998);
xor (n858,n859,n941);
xor (n859,n860,n939);
xor (n860,n861,n864);
and (n861,n862,n863);
wire s0n862,s1n862,notn862;
or (n862,s0n862,s1n862);
not(notn862,n839);
and (s0n862,notn862,n23);
and (s1n862,n839,n442);
wire s0n863,s1n863,notn863;
or (n863,s0n863,s1n863);
not(notn863,n839);
and (s0n863,notn863,n24);
and (s1n863,n839,n443);
or (n864,n865,n870);
and (n865,n866,n868);
and (n866,n862,n867);
wire s0n867,s1n867,notn867;
or (n867,s0n867,s1n867);
not(notn867,n839);
and (s0n867,notn867,n28);
and (s1n867,n839,n447);
and (n868,n869,n863);
wire s0n869,s1n869,notn869;
or (n869,s0n869,s1n869);
not(notn869,n839);
and (s0n869,notn869,n30);
and (s1n869,n839,n449);
and (n870,n871,n872);
xor (n871,n866,n868);
or (n872,n873,n877);
and (n873,n874,n875);
and (n874,n869,n867);
and (n875,n876,n863);
wire s0n876,s1n876,notn876;
or (n876,s0n876,s1n876);
not(notn876,n839);
and (s0n876,notn876,n37);
and (s1n876,n839,n456);
and (n877,n878,n879);
xor (n878,n874,n875);
or (n879,n880,n884);
and (n880,n881,n882);
and (n881,n876,n867);
and (n882,n883,n863);
wire s0n883,s1n883,notn883;
or (n883,s0n883,s1n883);
not(notn883,n839);
and (s0n883,notn883,n44);
and (s1n883,n839,n463);
and (n884,n885,n886);
xor (n885,n881,n882);
or (n886,n887,n891);
and (n887,n888,n889);
and (n888,n883,n867);
and (n889,n890,n863);
wire s0n890,s1n890,notn890;
or (n890,s0n890,s1n890);
not(notn890,n839);
and (s0n890,notn890,n51);
and (s1n890,n839,n470);
and (n891,n892,n893);
xor (n892,n888,n889);
or (n893,n894,n898);
and (n894,n895,n896);
and (n895,n890,n867);
and (n896,n897,n863);
wire s0n897,s1n897,notn897;
or (n897,s0n897,s1n897);
not(notn897,n839);
and (s0n897,notn897,n58);
and (s1n897,n839,n477);
and (n898,n899,n900);
xor (n899,n895,n896);
or (n900,n901,n905);
and (n901,n902,n903);
and (n902,n897,n867);
and (n903,n904,n863);
wire s0n904,s1n904,notn904;
or (n904,s0n904,s1n904);
not(notn904,n839);
and (s0n904,notn904,n65);
and (s1n904,n839,n484);
and (n905,n906,n907);
xor (n906,n902,n903);
or (n907,n908,n912);
and (n908,n909,n910);
and (n909,n904,n867);
and (n910,n911,n863);
wire s0n911,s1n911,notn911;
or (n911,s0n911,s1n911);
not(notn911,n839);
and (s0n911,notn911,n72);
and (s1n911,n839,n491);
and (n912,n913,n914);
xor (n913,n909,n910);
or (n914,n915,n919);
and (n915,n916,n917);
and (n916,n911,n867);
and (n917,n918,n863);
wire s0n918,s1n918,notn918;
or (n918,s0n918,s1n918);
not(notn918,n839);
and (s0n918,notn918,n79);
and (s1n918,n839,n498);
and (n919,n920,n921);
xor (n920,n916,n917);
or (n921,n922,n926);
and (n922,n923,n924);
and (n923,n918,n867);
and (n924,n925,n863);
wire s0n925,s1n925,notn925;
or (n925,s0n925,s1n925);
not(notn925,n839);
and (s0n925,notn925,n86);
and (s1n925,n839,n505);
and (n926,n927,n928);
xor (n927,n923,n924);
or (n928,n929,n933);
and (n929,n930,n931);
and (n930,n925,n867);
and (n931,n932,n863);
wire s0n932,s1n932,notn932;
or (n932,s0n932,s1n932);
not(notn932,n839);
and (s0n932,notn932,n93);
and (s1n932,n839,n512);
and (n933,n934,n935);
xor (n934,n930,n931);
and (n935,n936,n937);
and (n936,n932,n867);
and (n937,n938,n863);
wire s0n938,s1n938,notn938;
or (n938,s0n938,s1n938);
not(notn938,n839);
and (s0n938,notn938,n99);
and (s1n938,n839,n518);
and (n939,n869,n940);
wire s0n940,s1n940,notn940;
or (n940,s0n940,s1n940);
not(notn940,n839);
and (s0n940,notn940,n101);
and (s1n940,n839,n520);
or (n941,n942,n945);
and (n942,n943,n944);
xor (n943,n871,n872);
and (n944,n876,n940);
and (n945,n946,n947);
xor (n946,n943,n944);
or (n947,n948,n951);
and (n948,n949,n950);
xor (n949,n878,n879);
and (n950,n883,n940);
and (n951,n952,n953);
xor (n952,n949,n950);
or (n953,n954,n957);
and (n954,n955,n956);
xor (n955,n885,n886);
and (n956,n890,n940);
and (n957,n958,n959);
xor (n958,n955,n956);
or (n959,n960,n963);
and (n960,n961,n962);
xor (n961,n892,n893);
and (n962,n897,n940);
and (n963,n964,n965);
xor (n964,n961,n962);
or (n965,n966,n969);
and (n966,n967,n968);
xor (n967,n899,n900);
and (n968,n904,n940);
and (n969,n970,n971);
xor (n970,n967,n968);
or (n971,n972,n975);
and (n972,n973,n974);
xor (n973,n906,n907);
and (n974,n911,n940);
and (n975,n976,n977);
xor (n976,n973,n974);
or (n977,n978,n981);
and (n978,n979,n980);
xor (n979,n913,n914);
and (n980,n918,n940);
and (n981,n982,n983);
xor (n982,n979,n980);
or (n983,n984,n987);
and (n984,n985,n986);
xor (n985,n920,n921);
and (n986,n925,n940);
and (n987,n988,n989);
xor (n988,n985,n986);
or (n989,n990,n993);
and (n990,n991,n992);
xor (n991,n927,n928);
and (n992,n932,n940);
and (n993,n994,n995);
xor (n994,n991,n992);
and (n995,n996,n997);
xor (n996,n934,n935);
and (n997,n938,n940);
and (n998,n876,n999);
wire s0n999,s1n999,notn999;
or (n999,s0n999,s1n999);
not(notn999,n839);
and (s0n999,notn999,n160);
and (s1n999,n839,n579);
or (n1000,n1001,n1004);
and (n1001,n1002,n1003);
xor (n1002,n946,n947);
and (n1003,n883,n999);
and (n1004,n1005,n1006);
xor (n1005,n1002,n1003);
or (n1006,n1007,n1010);
and (n1007,n1008,n1009);
xor (n1008,n952,n953);
and (n1009,n890,n999);
and (n1010,n1011,n1012);
xor (n1011,n1008,n1009);
or (n1012,n1013,n1016);
and (n1013,n1014,n1015);
xor (n1014,n958,n959);
and (n1015,n897,n999);
and (n1016,n1017,n1018);
xor (n1017,n1014,n1015);
or (n1018,n1019,n1022);
and (n1019,n1020,n1021);
xor (n1020,n964,n965);
and (n1021,n904,n999);
and (n1022,n1023,n1024);
xor (n1023,n1020,n1021);
or (n1024,n1025,n1028);
and (n1025,n1026,n1027);
xor (n1026,n970,n971);
and (n1027,n911,n999);
and (n1028,n1029,n1030);
xor (n1029,n1026,n1027);
or (n1030,n1031,n1034);
and (n1031,n1032,n1033);
xor (n1032,n976,n977);
and (n1033,n918,n999);
and (n1034,n1035,n1036);
xor (n1035,n1032,n1033);
or (n1036,n1037,n1040);
and (n1037,n1038,n1039);
xor (n1038,n982,n983);
and (n1039,n925,n999);
and (n1040,n1041,n1042);
xor (n1041,n1038,n1039);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n988,n989);
and (n1045,n932,n999);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
and (n1048,n1049,n1050);
xor (n1049,n994,n995);
and (n1050,n938,n999);
and (n1051,n883,n1052);
wire s0n1052,s1n1052,notn1052;
or (n1052,s0n1052,s1n1052);
not(notn1052,n839);
and (s0n1052,notn1052,n213);
and (s1n1052,n839,n632);
or (n1053,n1054,n1057);
and (n1054,n1055,n1056);
xor (n1055,n1005,n1006);
and (n1056,n890,n1052);
and (n1057,n1058,n1059);
xor (n1058,n1055,n1056);
or (n1059,n1060,n1063);
and (n1060,n1061,n1062);
xor (n1061,n1011,n1012);
and (n1062,n897,n1052);
and (n1063,n1064,n1065);
xor (n1064,n1061,n1062);
or (n1065,n1066,n1069);
and (n1066,n1067,n1068);
xor (n1067,n1017,n1018);
and (n1068,n904,n1052);
and (n1069,n1070,n1071);
xor (n1070,n1067,n1068);
or (n1071,n1072,n1075);
and (n1072,n1073,n1074);
xor (n1073,n1023,n1024);
and (n1074,n911,n1052);
and (n1075,n1076,n1077);
xor (n1076,n1073,n1074);
or (n1077,n1078,n1081);
and (n1078,n1079,n1080);
xor (n1079,n1029,n1030);
and (n1080,n918,n1052);
and (n1081,n1082,n1083);
xor (n1082,n1079,n1080);
or (n1083,n1084,n1087);
and (n1084,n1085,n1086);
xor (n1085,n1035,n1036);
and (n1086,n925,n1052);
and (n1087,n1088,n1089);
xor (n1088,n1085,n1086);
or (n1089,n1090,n1093);
and (n1090,n1091,n1092);
xor (n1091,n1041,n1042);
and (n1092,n932,n1052);
and (n1093,n1094,n1095);
xor (n1094,n1091,n1092);
and (n1095,n1096,n1097);
xor (n1096,n1047,n1048);
and (n1097,n938,n1052);
and (n1098,n890,n1099);
wire s0n1099,s1n1099,notn1099;
or (n1099,s0n1099,s1n1099);
not(notn1099,n839);
and (s0n1099,notn1099,n260);
and (s1n1099,n839,n679);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
xor (n1102,n1058,n1059);
and (n1103,n897,n1099);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1064,n1065);
and (n1109,n904,n1099);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1070,n1071);
and (n1115,n911,n1099);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1076,n1077);
and (n1121,n918,n1099);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1082,n1083);
and (n1127,n925,n1099);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1088,n1089);
and (n1133,n932,n1099);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
and (n1136,n1137,n1138);
xor (n1137,n1094,n1095);
and (n1138,n938,n1099);
and (n1139,n897,n1140);
wire s0n1140,s1n1140,notn1140;
or (n1140,s0n1140,s1n1140);
not(notn1140,n839);
and (s0n1140,notn1140,n301);
and (s1n1140,n839,n720);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
xor (n1143,n1105,n1106);
and (n1144,n904,n1140);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
xor (n1149,n1111,n1112);
and (n1150,n911,n1140);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
xor (n1155,n1117,n1118);
and (n1156,n918,n1140);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1163);
and (n1160,n1161,n1162);
xor (n1161,n1123,n1124);
and (n1162,n925,n1140);
and (n1163,n1164,n1165);
xor (n1164,n1161,n1162);
or (n1165,n1166,n1169);
and (n1166,n1167,n1168);
xor (n1167,n1129,n1130);
and (n1168,n932,n1140);
and (n1169,n1170,n1171);
xor (n1170,n1167,n1168);
and (n1171,n1172,n1173);
xor (n1172,n1135,n1136);
and (n1173,n938,n1140);
and (n1174,n904,n1175);
wire s0n1175,s1n1175,notn1175;
or (n1175,s0n1175,s1n1175);
not(notn1175,n839);
and (s0n1175,notn1175,n336);
and (s1n1175,n839,n755);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1146,n1147);
and (n1179,n911,n1175);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1152,n1153);
and (n1185,n918,n1175);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1158,n1159);
and (n1191,n925,n1175);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1164,n1165);
and (n1197,n932,n1175);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
and (n1200,n1201,n1202);
xor (n1201,n1170,n1171);
and (n1202,n938,n1175);
and (n1203,n911,n1204);
wire s0n1204,s1n1204,notn1204;
or (n1204,s0n1204,s1n1204);
not(notn1204,n839);
and (s0n1204,notn1204,n365);
and (s1n1204,n839,n784);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1181,n1182);
and (n1208,n918,n1204);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1187,n1188);
and (n1214,n925,n1204);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1193,n1194);
and (n1220,n932,n1204);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
and (n1223,n1224,n1225);
xor (n1224,n1199,n1200);
and (n1225,n938,n1204);
and (n1226,n918,n1227);
wire s0n1227,s1n1227,notn1227;
or (n1227,s0n1227,s1n1227);
not(notn1227,n839);
and (s0n1227,notn1227,n388);
and (s1n1227,n839,n807);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1210,n1211);
and (n1231,n925,n1227);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1216,n1217);
and (n1237,n932,n1227);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
and (n1240,n1241,n1242);
xor (n1241,n1222,n1223);
and (n1242,n938,n1227);
and (n1243,n925,n1244);
wire s0n1244,s1n1244,notn1244;
or (n1244,s0n1244,s1n1244);
not(notn1244,n839);
and (s0n1244,notn1244,n405);
and (s1n1244,n839,n824);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1233,n1234);
and (n1248,n932,n1244);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
and (n1251,n1252,n1253);
xor (n1252,n1239,n1240);
and (n1253,n938,n1244);
and (n1254,n932,n1255);
wire s0n1255,s1n1255,notn1255;
or (n1255,s0n1255,s1n1255);
not(notn1255,n839);
and (s0n1255,notn1255,n416);
and (s1n1255,n839,n835);
and (n1256,n1257,n1258);
xor (n1257,n1250,n1251);
and (n1258,n938,n1255);
endmodule
