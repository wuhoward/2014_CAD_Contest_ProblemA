module top (out,n3,n11,n13,n14,n16,n18,n19,n24,n30
        ,n33,n34,n40,n41,n56,n58,n59,n68,n69,n71
        ,n72,n82,n91,n104,n105,n112,n118,n131,n137,n156
        ,n162);
output out;
input n3;
input n11;
input n13;
input n14;
input n16;
input n18;
input n19;
input n24;
input n30;
input n33;
input n34;
input n40;
input n41;
input n56;
input n58;
input n59;
input n68;
input n69;
input n71;
input n72;
input n82;
input n91;
input n104;
input n105;
input n112;
input n118;
input n131;
input n137;
input n156;
input n162;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n12;
wire n15;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n70;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
xor (out,n0,n516);
nand (n0,n1,n42);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
xor (n5,n6,n38);
xor (n6,n7,n35);
xor (n7,n8,n31);
xor (n8,n9,n20);
xor (n9,n10,n15);
and (n10,n11,n12);
wire s0n12,s1n12,notn12;
or (n12,s0n12,s1n12);
not(notn12,n3);
and (s0n12,notn12,n13);
and (s1n12,n3,n14);
and (n15,n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n3);
and (s0n17,notn17,n18);
and (s1n17,n3,n19);
or (n20,n21,n25);
and (n21,n22,n23);
and (n22,n16,n12);
and (n23,n24,n17);
and (n25,n26,n27);
xor (n26,n22,n23);
and (n27,n28,n29);
and (n28,n24,n12);
and (n29,n30,n17);
and (n31,n24,n32);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n3);
and (s0n32,notn32,n33);
and (s1n32,n3,n34);
and (n35,n36,n37);
xor (n36,n26,n27);
and (n37,n30,n32);
and (n38,n30,n39);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n3);
and (s0n39,notn39,n40);
and (s1n39,n3,n41);
nand (n42,n43,n2);
xnor (n43,n44,n265);
nand (n44,n45,n264);
nand (n45,n46,n223);
not (n46,n47);
xor (n47,n48,n200);
xor (n48,n49,n121);
xor (n49,n50,n96);
xor (n50,n51,n85);
nand (n51,n52,n78);
or (n52,n53,n63);
not (n53,n54);
nor (n54,n55,n60);
and (n55,n56,n57);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n3);
and (s0n57,notn57,n58);
and (s1n57,n3,n59);
and (n60,n61,n62);
not (n61,n56);
not (n62,n57);
nand (n63,n64,n75);
nor (n64,n65,n73);
and (n65,n66,n70);
not (n66,n67);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n3);
and (s0n67,notn67,n68);
and (s1n67,n3,n69);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n3);
and (s0n70,notn70,n71);
and (s1n70,n3,n72);
and (n73,n67,n74);
not (n74,n70);
nand (n75,n76,n77);
or (n76,n66,n57);
nand (n77,n57,n66);
nand (n78,n79,n80);
not (n79,n64);
nor (n80,n81,n83);
and (n81,n82,n57);
and (n83,n84,n62);
not (n84,n82);
nor (n85,n86,n92);
nand (n86,n57,n87);
not (n87,n88);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n3);
and (s0n88,notn88,1'b0);
and (s1n88,n3,n90);
and (n90,n91,n59);
nor (n92,n93,n95);
and (n93,n88,n94);
not (n94,n11);
and (n95,n87,n11);
nand (n96,n97,n115);
or (n97,n98,n110);
nand (n98,n99,n107);
not (n99,n100);
nand (n100,n101,n106);
or (n101,n102,n39);
not (n102,n103);
wire s0n103,s1n103,notn103;
or (n103,s0n103,s1n103);
not(notn103,n3);
and (s0n103,notn103,n104);
and (s1n103,n3,n105);
nand (n106,n39,n102);
nand (n107,n108,n109);
or (n108,n102,n70);
nand (n109,n70,n102);
nor (n110,n111,n113);
and (n111,n74,n112);
and (n113,n70,n114);
not (n114,n112);
or (n115,n99,n116);
nor (n116,n117,n119);
and (n117,n74,n118);
and (n119,n70,n120);
not (n120,n118);
xor (n121,n122,n178);
xor (n122,n123,n165);
xor (n123,n124,n141);
nand (n124,n125,n134);
or (n125,n126,n129);
not (n126,n127);
nor (n127,n128,n12);
not (n128,n17);
nor (n129,n130,n132);
and (n130,n128,n131);
and (n132,n17,n133);
not (n133,n131);
or (n134,n135,n140);
nor (n135,n136,n138);
and (n136,n128,n137);
and (n138,n17,n139);
not (n139,n137);
not (n140,n12);
nand (n141,n142,n159);
or (n142,n143,n153);
not (n143,n144);
and (n144,n145,n149);
nand (n145,n146,n148);
or (n146,n147,n39);
not (n147,n32);
nand (n148,n39,n147);
not (n149,n150);
nand (n150,n151,n152);
or (n151,n147,n17);
nand (n152,n17,n147);
nor (n153,n154,n157);
and (n154,n155,n156);
not (n155,n39);
and (n157,n39,n158);
not (n158,n156);
or (n159,n149,n160);
nor (n160,n161,n163);
and (n161,n155,n162);
and (n163,n39,n164);
not (n164,n162);
and (n165,n166,n172);
nand (n166,n167,n171);
or (n167,n126,n168);
nor (n168,n169,n170);
and (n169,n128,n162);
and (n170,n17,n164);
or (n171,n129,n140);
nand (n172,n173,n177);
or (n173,n143,n174);
nor (n174,n175,n176);
and (n175,n155,n118);
and (n176,n39,n120);
or (n177,n153,n149);
or (n178,n179,n199);
and (n179,n180,n193);
xor (n180,n181,n188);
nand (n181,n182,n187);
or (n182,n183,n63);
not (n183,n184);
nor (n184,n185,n186);
and (n185,n11,n57);
and (n186,n94,n62);
nand (n187,n79,n54);
nor (n188,n86,n189);
nor (n189,n190,n192);
and (n190,n88,n191);
not (n191,n16);
and (n192,n87,n16);
nand (n193,n194,n198);
or (n194,n98,n195);
nor (n195,n196,n197);
and (n196,n74,n82);
and (n197,n70,n84);
or (n198,n99,n110);
and (n199,n181,n188);
and (n200,n201,n202);
xor (n201,n166,n172);
or (n202,n203,n222);
and (n203,n204,n216);
xor (n204,n205,n211);
nand (n205,n206,n210);
or (n206,n207,n63);
nor (n207,n208,n209);
and (n208,n16,n62);
and (n209,n191,n57);
nand (n210,n184,n79);
nor (n211,n86,n212);
nor (n212,n213,n215);
and (n213,n88,n214);
not (n214,n24);
and (n215,n87,n24);
nand (n216,n217,n221);
or (n217,n126,n218);
nor (n218,n219,n220);
and (n219,n128,n156);
and (n220,n17,n158);
or (n221,n168,n140);
and (n222,n205,n211);
not (n223,n224);
or (n224,n225,n263);
and (n225,n226,n229);
xor (n226,n227,n228);
xor (n227,n180,n193);
xor (n228,n201,n202);
or (n229,n230,n262);
and (n230,n231,n244);
xor (n231,n232,n238);
nand (n232,n233,n237);
or (n233,n98,n234);
nor (n234,n235,n236);
and (n235,n74,n56);
and (n236,n70,n61);
or (n237,n99,n195);
nand (n238,n239,n243);
or (n239,n143,n240);
nor (n240,n241,n242);
and (n241,n155,n112);
and (n242,n39,n114);
or (n243,n174,n149);
or (n244,n245,n261);
and (n245,n246,n255);
xor (n246,n247,n249);
and (n247,n248,n30);
not (n248,n86);
nand (n249,n250,n254);
or (n250,n126,n251);
nor (n251,n252,n253);
and (n252,n120,n17);
and (n253,n118,n128);
or (n254,n218,n140);
nand (n255,n256,n260);
or (n256,n63,n257);
nor (n257,n258,n259);
and (n258,n24,n62);
and (n259,n214,n57);
or (n260,n64,n207);
and (n261,n247,n249);
and (n262,n232,n238);
and (n263,n227,n228);
nand (n264,n47,n224);
nand (n265,n266,n515);
or (n266,n267,n307);
nor (n267,n268,n269);
xor (n268,n226,n229);
or (n269,n270,n306);
and (n270,n271,n305);
xor (n271,n272,n273);
xor (n272,n204,n216);
or (n273,n274,n304);
and (n274,n275,n289);
xor (n275,n276,n283);
nand (n276,n277,n282);
or (n277,n143,n278);
not (n278,n279);
nor (n279,n280,n281);
and (n280,n82,n39);
and (n281,n84,n155);
or (n282,n149,n240);
nand (n283,n284,n288);
or (n284,n98,n285);
nor (n285,n286,n287);
and (n286,n74,n11);
and (n287,n70,n94);
or (n288,n99,n234);
and (n289,n290,n296);
nor (n290,n291,n62);
nor (n291,n292,n294);
and (n292,n74,n293);
nand (n293,n67,n30);
and (n294,n66,n295);
not (n295,n30);
nand (n296,n297,n302);
or (n297,n298,n126);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n112,n17);
and (n301,n114,n128);
nand (n302,n303,n12);
not (n303,n251);
and (n304,n276,n283);
xor (n305,n231,n244);
and (n306,n272,n273);
not (n307,n308);
nand (n308,n309,n510);
not (n309,n310);
nor (n310,n311,n491);
nor (n311,n312,n489);
and (n312,n313,n463);
or (n313,n314,n462);
and (n314,n315,n379);
xor (n315,n316,n356);
or (n316,n317,n355);
and (n317,n318,n340);
xor (n318,n319,n329);
nand (n319,n320,n325);
or (n320,n321,n143);
not (n321,n322);
nor (n322,n323,n324);
and (n323,n191,n155);
and (n324,n16,n39);
nand (n325,n150,n326);
nor (n326,n327,n328);
and (n327,n11,n39);
and (n328,n155,n94);
nand (n329,n330,n335);
or (n330,n331,n99);
not (n331,n332);
nor (n332,n333,n334);
and (n333,n24,n70);
and (n334,n214,n74);
nand (n335,n336,n337);
not (n336,n98);
nand (n337,n338,n339);
or (n338,n74,n30);
or (n339,n70,n295);
xor (n340,n341,n346);
and (n341,n342,n70);
nand (n342,n343,n345);
or (n343,n39,n344);
and (n344,n30,n103);
or (n345,n103,n30);
nand (n346,n347,n351);
or (n347,n126,n348);
nor (n348,n349,n350);
and (n349,n128,n56);
and (n350,n17,n61);
or (n351,n352,n140);
nor (n352,n353,n354);
and (n353,n82,n128);
and (n354,n84,n17);
and (n355,n319,n329);
xor (n356,n357,n365);
xor (n357,n358,n364);
nand (n358,n359,n360);
or (n359,n331,n98);
or (n360,n99,n361);
nor (n361,n362,n363);
and (n362,n74,n16);
and (n363,n70,n191);
and (n364,n341,n346);
xor (n365,n366,n372);
xor (n366,n367,n368);
and (n367,n79,n30);
nand (n368,n369,n370);
or (n369,n140,n298);
nand (n370,n371,n127);
not (n371,n352);
nand (n372,n373,n375);
or (n373,n374,n143);
not (n374,n326);
nand (n375,n150,n376);
nand (n376,n377,n378);
or (n377,n39,n61);
or (n378,n155,n56);
or (n379,n380,n461);
and (n380,n381,n402);
xor (n381,n382,n401);
or (n382,n383,n400);
and (n383,n384,n393);
xor (n384,n385,n386);
and (n385,n100,n30);
nand (n386,n387,n392);
or (n387,n388,n143);
not (n388,n389);
nor (n389,n390,n391);
and (n390,n24,n39);
and (n391,n214,n155);
nand (n392,n322,n150);
nand (n393,n394,n399);
or (n394,n126,n395);
not (n395,n396);
nor (n396,n397,n398);
and (n397,n94,n128);
and (n398,n11,n17);
or (n399,n348,n140);
and (n400,n385,n386);
xor (n401,n318,n340);
or (n402,n403,n460);
and (n403,n404,n459);
xor (n404,n405,n418);
nor (n405,n406,n414);
not (n406,n407);
nand (n407,n408,n413);
or (n408,n409,n126);
not (n409,n410);
nand (n410,n411,n412);
or (n411,n191,n17);
nand (n412,n17,n191);
nand (n413,n396,n12);
nand (n414,n415,n39);
nand (n415,n416,n417);
or (n416,n17,n37);
or (n417,n32,n30);
nand (n418,n419,n457);
or (n419,n420,n443);
not (n420,n421);
nand (n421,n422,n442);
or (n422,n423,n432);
nor (n423,n424,n431);
nand (n424,n425,n430);
or (n425,n426,n126);
not (n426,n427);
nand (n427,n428,n429);
or (n428,n214,n17);
nand (n429,n17,n214);
nand (n430,n410,n12);
nor (n431,n149,n295);
nand (n432,n433,n440);
nand (n433,n434,n439);
or (n434,n435,n126);
not (n435,n436);
nand (n436,n437,n438);
or (n437,n128,n30);
or (n438,n17,n295);
nand (n439,n427,n12);
nor (n440,n441,n128);
and (n441,n30,n12);
nand (n442,n424,n431);
not (n443,n444);
nand (n444,n445,n453);
not (n445,n446);
nand (n446,n447,n452);
or (n447,n448,n143);
not (n448,n449);
nand (n449,n450,n451);
or (n450,n155,n30);
or (n451,n39,n295);
nand (n452,n150,n389);
nor (n453,n454,n456);
and (n454,n406,n455);
not (n455,n414);
and (n456,n407,n414);
nand (n457,n458,n446);
not (n458,n453);
xor (n459,n384,n393);
and (n460,n405,n418);
and (n461,n382,n401);
and (n462,n316,n356);
or (n463,n464,n486);
xor (n464,n465,n470);
xor (n465,n466,n467);
xor (n466,n290,n296);
or (n467,n468,n469);
and (n468,n366,n372);
and (n469,n367,n368);
xor (n470,n471,n483);
xor (n471,n472,n479);
nand (n472,n473,n478);
or (n473,n474,n63);
not (n474,n475);
nand (n475,n476,n477);
or (n476,n62,n30);
or (n477,n57,n295);
or (n478,n64,n257);
nand (n479,n480,n482);
or (n480,n481,n143);
not (n481,n376);
nand (n482,n150,n279);
nand (n483,n484,n485);
or (n484,n98,n361);
or (n485,n99,n285);
or (n486,n487,n488);
and (n487,n357,n365);
and (n488,n358,n364);
not (n489,n490);
nand (n490,n464,n486);
nand (n491,n492,n504);
not (n492,n493);
nor (n493,n494,n501);
xor (n494,n495,n500);
xor (n495,n496,n499);
or (n496,n497,n498);
and (n497,n471,n483);
and (n498,n472,n479);
xor (n499,n246,n255);
xor (n500,n275,n289);
or (n501,n502,n503);
and (n502,n465,n470);
and (n503,n466,n467);
not (n504,n505);
nor (n505,n506,n509);
or (n506,n507,n508);
and (n507,n495,n500);
and (n508,n496,n499);
xor (n509,n271,n305);
nor (n510,n511,n514);
and (n511,n504,n512);
not (n512,n513);
nand (n513,n494,n501);
and (n514,n506,n509);
nand (n515,n268,n269);
wire s0n516,s1n516,notn516;
or (n516,s0n516,s1n516);
not(notn516,n3);
and (s0n516,notn516,n517);
and (s1n516,n3,n5);
xor (n517,n518,n804);
xor (n518,n519,n812);
xor (n519,n520,n799);
xor (n520,n521,n805);
xor (n521,n522,n793);
xor (n522,n523,n790);
xor (n523,n524,n789);
xor (n524,n525,n769);
xor (n525,n526,n55);
xor (n526,n527,n742);
xor (n527,n528,n741);
xor (n528,n529,n709);
xor (n529,n530,n708);
xor (n530,n531,n670);
xor (n531,n532,n669);
xor (n532,n533,n630);
xor (n533,n534,n629);
xor (n534,n535,n584);
xor (n535,n536,n583);
xor (n536,n537,n540);
xor (n537,n538,n539);
and (n538,n137,n12);
and (n539,n131,n17);
or (n540,n541,n544);
and (n541,n542,n543);
and (n542,n131,n12);
and (n543,n162,n17);
and (n544,n545,n546);
xor (n545,n542,n543);
or (n546,n547,n550);
and (n547,n548,n549);
and (n548,n162,n12);
and (n549,n156,n17);
and (n550,n551,n552);
xor (n551,n548,n549);
or (n552,n553,n556);
and (n553,n554,n555);
and (n554,n156,n12);
and (n555,n118,n17);
and (n556,n557,n558);
xor (n557,n554,n555);
or (n558,n559,n561);
and (n559,n560,n300);
and (n560,n118,n12);
and (n561,n562,n563);
xor (n562,n560,n300);
or (n563,n564,n567);
and (n564,n565,n566);
and (n565,n112,n12);
and (n566,n82,n17);
and (n567,n568,n569);
xor (n568,n565,n566);
or (n569,n570,n573);
and (n570,n571,n572);
and (n571,n82,n12);
and (n572,n56,n17);
and (n573,n574,n575);
xor (n574,n571,n572);
or (n575,n576,n578);
and (n576,n577,n398);
and (n577,n56,n12);
and (n578,n579,n580);
xor (n579,n577,n398);
or (n580,n581,n582);
and (n581,n10,n15);
and (n582,n9,n20);
and (n583,n162,n32);
or (n584,n585,n588);
and (n585,n586,n587);
xor (n586,n545,n546);
and (n587,n156,n32);
and (n588,n589,n590);
xor (n589,n586,n587);
or (n590,n591,n594);
and (n591,n592,n593);
xor (n592,n551,n552);
and (n593,n118,n32);
and (n594,n595,n596);
xor (n595,n592,n593);
or (n596,n597,n600);
and (n597,n598,n599);
xor (n598,n557,n558);
and (n599,n112,n32);
and (n600,n601,n602);
xor (n601,n598,n599);
or (n602,n603,n606);
and (n603,n604,n605);
xor (n604,n562,n563);
and (n605,n82,n32);
and (n606,n607,n608);
xor (n607,n604,n605);
or (n608,n609,n612);
and (n609,n610,n611);
xor (n610,n568,n569);
and (n611,n56,n32);
and (n612,n613,n614);
xor (n613,n610,n611);
or (n614,n615,n618);
and (n615,n616,n617);
xor (n616,n574,n575);
and (n617,n11,n32);
and (n618,n619,n620);
xor (n619,n616,n617);
or (n620,n621,n624);
and (n621,n622,n623);
xor (n622,n579,n580);
and (n623,n16,n32);
and (n624,n625,n626);
xor (n625,n622,n623);
or (n626,n627,n628);
and (n627,n8,n31);
and (n628,n7,n35);
and (n629,n156,n39);
or (n630,n631,n634);
and (n631,n632,n633);
xor (n632,n589,n590);
and (n633,n118,n39);
and (n634,n635,n636);
xor (n635,n632,n633);
or (n636,n637,n640);
and (n637,n638,n639);
xor (n638,n595,n596);
and (n639,n112,n39);
and (n640,n641,n642);
xor (n641,n638,n639);
or (n642,n643,n645);
and (n643,n644,n280);
xor (n644,n601,n602);
and (n645,n646,n647);
xor (n646,n644,n280);
or (n647,n648,n651);
and (n648,n649,n650);
xor (n649,n607,n608);
and (n650,n56,n39);
and (n651,n652,n653);
xor (n652,n649,n650);
or (n653,n654,n656);
and (n654,n655,n327);
xor (n655,n613,n614);
and (n656,n657,n658);
xor (n657,n655,n327);
or (n658,n659,n661);
and (n659,n660,n324);
xor (n660,n619,n620);
and (n661,n662,n663);
xor (n662,n660,n324);
or (n663,n664,n666);
and (n664,n665,n390);
xor (n665,n625,n626);
and (n666,n667,n668);
xor (n667,n665,n390);
and (n668,n6,n38);
and (n669,n118,n103);
or (n670,n671,n674);
and (n671,n672,n673);
xor (n672,n635,n636);
and (n673,n112,n103);
and (n674,n675,n676);
xor (n675,n672,n673);
or (n676,n677,n680);
and (n677,n678,n679);
xor (n678,n641,n642);
and (n679,n82,n103);
and (n680,n681,n682);
xor (n681,n678,n679);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n646,n647);
and (n685,n56,n103);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n652,n653);
and (n691,n11,n103);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n698);
and (n695,n696,n697);
xor (n696,n657,n658);
and (n697,n16,n103);
and (n698,n699,n700);
xor (n699,n696,n697);
or (n700,n701,n704);
and (n701,n702,n703);
xor (n702,n662,n663);
and (n703,n24,n103);
and (n704,n705,n706);
xor (n705,n702,n703);
and (n706,n707,n344);
xor (n707,n667,n668);
and (n708,n112,n70);
or (n709,n710,n713);
and (n710,n711,n712);
xor (n711,n675,n676);
and (n712,n82,n70);
and (n713,n714,n715);
xor (n714,n711,n712);
or (n715,n716,n719);
and (n716,n717,n718);
xor (n717,n681,n682);
and (n718,n56,n70);
and (n719,n720,n721);
xor (n720,n717,n718);
or (n721,n722,n725);
and (n722,n723,n724);
xor (n723,n687,n688);
and (n724,n11,n70);
and (n725,n726,n727);
xor (n726,n723,n724);
or (n727,n728,n731);
and (n728,n729,n730);
xor (n729,n693,n694);
and (n730,n16,n70);
and (n731,n732,n733);
xor (n732,n729,n730);
or (n733,n734,n736);
and (n734,n735,n333);
xor (n735,n699,n700);
and (n736,n737,n738);
xor (n737,n735,n333);
and (n738,n739,n740);
xor (n739,n705,n706);
and (n740,n30,n70);
and (n741,n82,n67);
or (n742,n743,n746);
and (n743,n744,n745);
xor (n744,n714,n715);
and (n745,n56,n67);
and (n746,n747,n748);
xor (n747,n744,n745);
or (n748,n749,n752);
and (n749,n750,n751);
xor (n750,n720,n721);
and (n751,n11,n67);
and (n752,n753,n754);
xor (n753,n750,n751);
or (n754,n755,n758);
and (n755,n756,n757);
xor (n756,n726,n727);
and (n757,n16,n67);
and (n758,n759,n760);
xor (n759,n756,n757);
or (n760,n761,n764);
and (n761,n762,n763);
xor (n762,n732,n733);
and (n763,n24,n67);
and (n764,n765,n766);
xor (n765,n762,n763);
and (n766,n767,n768);
xor (n767,n737,n738);
not (n768,n293);
or (n769,n770,n772);
and (n770,n771,n185);
xor (n771,n747,n748);
and (n772,n773,n774);
xor (n773,n771,n185);
or (n774,n775,n778);
and (n775,n776,n777);
xor (n776,n753,n754);
and (n777,n16,n57);
and (n778,n779,n780);
xor (n779,n776,n777);
or (n780,n781,n784);
and (n781,n782,n783);
xor (n782,n759,n760);
and (n783,n24,n57);
and (n784,n785,n786);
xor (n785,n782,n783);
and (n786,n787,n788);
xor (n787,n765,n766);
and (n788,n30,n57);
and (n789,n11,n88);
or (n790,n791,n794);
and (n791,n792,n793);
xor (n792,n773,n774);
and (n793,n16,n88);
and (n794,n795,n796);
xor (n795,n792,n793);
or (n796,n797,n800);
and (n797,n798,n799);
xor (n798,n779,n780);
and (n799,n24,n88);
and (n800,n801,n802);
xor (n801,n798,n799);
and (n802,n803,n804);
xor (n803,n785,n786);
and (n804,n30,n88);
or (n805,n806,n808);
and (n806,n807,n799);
xor (n807,n795,n796);
and (n808,n809,n810);
xor (n809,n807,n799);
and (n810,n811,n804);
xor (n811,n801,n802);
and (n812,n813,n804);
xor (n813,n809,n810);
endmodule
