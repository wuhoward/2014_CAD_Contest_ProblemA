module top (out,n4,n5,n22,n23,n29,n31,n38,n52,n53
        ,n59,n63,n69,n78,n79,n87,n93,n104,n105,n110
        ,n121,n128,n134,n145,n151,n155,n161,n169,n175,n179
        ,n185,n193,n203,n208,n243,n987);
output out;
input n4;
input n5;
input n22;
input n23;
input n29;
input n31;
input n38;
input n52;
input n53;
input n59;
input n63;
input n69;
input n78;
input n79;
input n87;
input n93;
input n104;
input n105;
input n110;
input n121;
input n128;
input n134;
input n145;
input n151;
input n155;
input n161;
input n169;
input n175;
input n179;
input n185;
input n193;
input n203;
input n208;
input n243;
input n987;
wire n0;
wire n1;
wire n2;
wire n3;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
xor (out,n0,n989);
or (n0,n1,n986);
and (n1,n2,n6);
nor (n2,n3,n5);
not (n3,n4);
nor (n6,n7,n983);
and (n7,n8,n479);
nor (n8,n9,n478);
not (n9,n10);
nand (n10,n11,n416);
xor (n11,n12,n351);
xor (n12,n13,n211);
xor (n13,n14,n138);
xor (n14,n15,n96);
xor (n15,n16,n72);
xor (n16,n17,n46);
nand (n17,n18,n34);
or (n18,n19,n26);
nor (n19,n20,n24);
and (n20,n21,n23);
not (n21,n22);
and (n24,n22,n25);
not (n25,n23);
not (n26,n27);
nand (n27,n28,n32);
or (n28,n29,n30);
not (n30,n31);
or (n32,n33,n31);
not (n33,n29);
nand (n34,n35,n41);
not (n35,n36);
nor (n36,n37,n39);
and (n37,n38,n33);
and (n39,n40,n29);
not (n40,n38);
not (n41,n42);
nand (n42,n19,n43);
nand (n43,n44,n45);
or (n44,n22,n33);
nand (n45,n33,n22);
nand (n46,n47,n66);
or (n47,n48,n61);
nand (n48,n49,n56);
nor (n49,n50,n54);
and (n50,n51,n53);
not (n51,n52);
and (n54,n52,n55);
not (n55,n53);
nand (n56,n57,n60);
nand (n57,n58,n53);
not (n58,n59);
nand (n60,n59,n55);
nor (n61,n62,n64);
and (n62,n63,n58);
and (n64,n59,n65);
not (n65,n63);
or (n66,n67,n49);
nor (n67,n68,n70);
and (n68,n69,n58);
and (n70,n59,n71);
not (n71,n69);
nand (n72,n73,n90);
or (n73,n74,n85);
nand (n74,n75,n82);
or (n75,n76,n80);
and (n76,n77,n79);
not (n77,n78);
and (n80,n78,n81);
not (n81,n79);
nor (n82,n83,n84);
and (n83,n59,n77);
and (n84,n58,n78);
nor (n85,n86,n88);
and (n86,n87,n81);
and (n88,n79,n89);
not (n89,n87);
or (n90,n91,n82);
nor (n91,n92,n94);
and (n92,n93,n81);
and (n94,n79,n95);
not (n95,n93);
nand (n96,n97,n137);
or (n97,n98,n113);
not (n98,n99);
nand (n99,n100,n106);
or (n100,n101,n104);
not (n101,n102);
nand (n102,n103,n105);
not (n103,n104);
not (n106,n107);
nor (n107,n108,n111);
and (n108,n109,n110);
not (n109,n105);
and (n111,n105,n112);
not (n112,n110);
not (n113,n114);
nand (n114,n115,n131);
or (n115,n116,n126);
nand (n116,n117,n123);
not (n117,n118);
nand (n118,n119,n122);
or (n119,n120,n105);
not (n120,n121);
nand (n122,n120,n105);
nand (n123,n124,n125);
or (n124,n120,n23);
nand (n125,n23,n120);
nor (n126,n127,n129);
and (n127,n25,n128);
and (n129,n23,n130);
not (n130,n128);
or (n131,n117,n132);
nor (n132,n133,n135);
and (n133,n25,n134);
and (n135,n23,n136);
not (n136,n134);
nand (n137,n98,n113);
xor (n138,n139,n188);
xor (n139,n140,n164);
nand (n140,n141,n158);
or (n141,n142,n153);
nand (n142,n143,n148);
nor (n143,n144,n146);
and (n144,n81,n145);
and (n146,n79,n147);
not (n147,n145);
nand (n148,n149,n152);
or (n149,n150,n145);
not (n150,n151);
nand (n152,n150,n145);
nor (n153,n154,n156);
and (n154,n155,n150);
and (n156,n157,n151);
not (n157,n155);
or (n158,n159,n143);
nor (n159,n160,n162);
and (n160,n161,n150);
and (n162,n151,n163);
not (n163,n161);
nand (n164,n165,n182);
or (n165,n166,n177);
nand (n166,n167,n172);
nor (n167,n168,n170);
and (n168,n33,n169);
and (n170,n29,n171);
not (n171,n169);
nand (n172,n173,n176);
or (n173,n169,n174);
not (n174,n175);
nand (n176,n174,n169);
nor (n177,n178,n180);
and (n178,n174,n179);
and (n180,n175,n181);
not (n181,n179);
or (n182,n167,n183);
nor (n183,n184,n186);
and (n184,n174,n185);
and (n186,n175,n187);
not (n187,n185);
nand (n188,n189,n205);
or (n189,n190,n199);
nand (n190,n191,n196);
nor (n191,n192,n194);
and (n192,n174,n193);
and (n194,n175,n195);
not (n195,n193);
nand (n196,n197,n198);
or (n197,n51,n193);
nand (n198,n51,n193);
not (n199,n200);
nor (n200,n201,n204);
and (n201,n202,n51);
not (n202,n203);
and (n204,n203,n52);
or (n205,n206,n191);
nor (n206,n207,n209);
and (n207,n51,n208);
and (n209,n52,n210);
not (n210,n208);
or (n211,n212,n350);
and (n212,n213,n290);
xor (n213,n214,n256);
or (n214,n215,n255);
and (n215,n216,n238);
xor (n216,n217,n226);
nand (n217,n218,n222);
or (n218,n48,n219);
nor (n219,n220,n221);
and (n220,n87,n58);
and (n221,n59,n89);
or (n222,n49,n223);
nor (n223,n224,n225);
and (n224,n58,n93);
and (n225,n59,n95);
nand (n226,n227,n232);
or (n227,n82,n228);
not (n228,n229);
nand (n229,n230,n231);
or (n230,n163,n79);
or (n231,n81,n161);
nand (n232,n233,n237);
not (n233,n234);
nor (n234,n235,n236);
and (n235,n81,n155);
and (n236,n157,n79);
not (n237,n74);
and (n238,n239,n246);
nor (n239,n240,n81);
nor (n240,n241,n244);
and (n241,n242,n58);
nand (n242,n78,n243);
and (n244,n245,n77);
not (n245,n243);
nand (n246,n247,n251);
or (n247,n248,n102);
nor (n248,n249,n250);
and (n249,n109,n31);
and (n250,n105,n30);
or (n251,n252,n103);
nor (n252,n253,n254);
and (n253,n105,n130);
nor (n254,n105,n130);
and (n255,n217,n226);
xor (n256,n257,n273);
xor (n257,n258,n261);
nand (n258,n259,n260);
or (n259,n74,n228);
or (n260,n85,n82);
xor (n261,n262,n267);
nor (n262,n263,n150);
nor (n263,n264,n266);
and (n264,n265,n81);
nand (n265,n243,n145);
and (n266,n245,n147);
nand (n267,n268,n272);
or (n268,n269,n102);
nor (n269,n270,n271);
and (n270,n134,n109);
and (n271,n136,n105);
or (n272,n107,n103);
or (n273,n274,n289);
and (n274,n275,n280);
xor (n275,n276,n277);
nor (n276,n143,n245);
nand (n277,n278,n279);
or (n278,n252,n102);
or (n279,n269,n103);
nand (n280,n281,n285);
or (n281,n116,n282);
nor (n282,n283,n284);
and (n283,n25,n38);
and (n284,n23,n40);
or (n285,n117,n286);
nor (n286,n287,n288);
and (n287,n25,n31);
and (n288,n23,n30);
and (n289,n276,n277);
or (n290,n291,n349);
and (n291,n292,n348);
xor (n292,n293,n323);
or (n293,n294,n322);
and (n294,n295,n312);
xor (n295,n296,n302);
nand (n296,n297,n301);
or (n297,n116,n298);
nor (n298,n299,n300);
and (n299,n185,n25);
and (n300,n187,n23);
or (n301,n117,n282);
nand (n302,n303,n308);
or (n303,n304,n166);
not (n304,n305);
nand (n305,n306,n307);
or (n306,n175,n71);
or (n307,n174,n69);
or (n308,n309,n167);
nor (n309,n310,n311);
and (n310,n203,n174);
and (n311,n175,n202);
nand (n312,n313,n318);
or (n313,n190,n314);
not (n314,n315);
nor (n315,n316,n317);
and (n316,n95,n51);
and (n317,n93,n52);
or (n318,n319,n191);
nor (n319,n320,n321);
and (n320,n51,n63);
and (n321,n52,n65);
and (n322,n296,n302);
or (n323,n324,n347);
and (n324,n325,n341);
xor (n325,n326,n335);
nand (n326,n327,n331);
or (n327,n42,n328);
nor (n328,n329,n330);
and (n329,n33,n208);
and (n330,n29,n210);
or (n331,n19,n332);
nor (n332,n333,n334);
and (n333,n33,n179);
and (n334,n29,n181);
nand (n335,n336,n340);
or (n336,n48,n337);
nor (n337,n338,n339);
and (n338,n161,n58);
and (n339,n59,n163);
or (n340,n219,n49);
nand (n341,n342,n346);
or (n342,n74,n343);
nor (n343,n344,n345);
and (n344,n245,n79);
and (n345,n243,n81);
or (n346,n234,n82);
and (n347,n326,n335);
xor (n348,n275,n280);
and (n349,n293,n323);
and (n350,n214,n256);
xor (n351,n352,n397);
xor (n352,n353,n356);
or (n353,n354,n355);
and (n354,n257,n273);
and (n355,n258,n261);
xor (n356,n357,n378);
xor (n357,n358,n359);
and (n358,n262,n267);
or (n359,n360,n377);
and (n360,n361,n371);
xor (n361,n362,n365);
nand (n362,n363,n364);
or (n363,n116,n286);
or (n364,n117,n126);
nand (n365,n366,n370);
or (n366,n142,n367);
nor (n367,n368,n369);
and (n368,n245,n151);
and (n369,n243,n150);
or (n370,n153,n143);
nand (n371,n372,n376);
or (n372,n166,n373);
nor (n373,n374,n375);
and (n374,n174,n208);
and (n375,n175,n210);
or (n376,n167,n177);
and (n377,n362,n365);
or (n378,n379,n396);
and (n379,n380,n393);
xor (n380,n381,n387);
nand (n381,n382,n383);
or (n382,n191,n199);
or (n383,n190,n384);
nor (n384,n385,n386);
and (n385,n51,n69);
and (n386,n52,n71);
nand (n387,n388,n392);
or (n388,n42,n389);
nor (n389,n390,n391);
and (n390,n33,n185);
and (n391,n29,n187);
or (n392,n19,n36);
nand (n393,n394,n395);
or (n394,n48,n223);
or (n395,n49,n61);
and (n396,n381,n387);
or (n397,n398,n415);
and (n398,n399,n414);
xor (n399,n400,n413);
or (n400,n401,n412);
and (n401,n402,n409);
xor (n402,n403,n406);
nand (n403,n404,n405);
or (n404,n166,n309);
or (n405,n373,n167);
nand (n406,n407,n408);
or (n407,n190,n319);
or (n408,n384,n191);
nand (n409,n410,n411);
or (n410,n42,n332);
or (n411,n19,n389);
and (n412,n403,n406);
xor (n413,n380,n393);
xor (n414,n361,n371);
and (n415,n400,n413);
or (n416,n417,n477);
and (n417,n418,n476);
xor (n418,n419,n420);
xor (n419,n399,n414);
or (n420,n421,n475);
and (n421,n422,n425);
xor (n422,n423,n424);
xor (n423,n402,n409);
xor (n424,n216,n238);
or (n425,n426,n474);
and (n426,n427,n450);
xor (n427,n428,n429);
xor (n428,n239,n246);
or (n429,n430,n449);
and (n430,n431,n442);
xor (n431,n432,n434);
and (n432,n433,n243);
not (n433,n82);
nand (n434,n435,n440);
or (n435,n436,n116);
not (n436,n437);
nand (n437,n438,n439);
or (n438,n23,n181);
or (n439,n25,n179);
nand (n440,n441,n118);
not (n441,n298);
nand (n442,n443,n448);
or (n443,n166,n444);
not (n444,n445);
nand (n445,n446,n447);
or (n446,n175,n65);
or (n447,n174,n63);
or (n448,n167,n304);
and (n449,n432,n434);
or (n450,n451,n473);
and (n451,n452,n467);
xor (n452,n453,n461);
nand (n453,n454,n459);
or (n454,n455,n190);
not (n455,n456);
nand (n456,n457,n458);
or (n457,n52,n89);
or (n458,n51,n87);
nand (n459,n315,n460);
not (n460,n191);
nand (n461,n462,n463);
or (n462,n103,n248);
or (n463,n464,n102);
nor (n464,n465,n466);
and (n465,n109,n38);
and (n466,n105,n40);
nand (n467,n468,n472);
or (n468,n469,n48);
nor (n469,n470,n471);
and (n470,n155,n58);
and (n471,n59,n157);
or (n472,n337,n49);
and (n473,n453,n461);
and (n474,n428,n429);
and (n475,n423,n424);
xor (n476,n213,n290);
and (n477,n419,n420);
nor (n478,n416,n11);
or (n479,n480,n982);
and (n480,n481,n545);
xor (n481,n482,n544);
or (n482,n483,n543);
and (n483,n484,n487);
xor (n484,n485,n486);
xor (n485,n292,n348);
xor (n486,n422,n425);
or (n487,n488,n542);
and (n488,n489,n492);
xor (n489,n490,n491);
xor (n490,n325,n341);
xor (n491,n295,n312);
or (n492,n493,n541);
and (n493,n494,n515);
xor (n494,n495,n501);
nand (n495,n496,n500);
or (n496,n42,n497);
nor (n497,n498,n499);
and (n498,n33,n203);
and (n499,n29,n202);
or (n500,n19,n328);
nor (n501,n502,n509);
not (n502,n503);
nand (n503,n504,n508);
or (n504,n505,n116);
nor (n505,n506,n507);
and (n506,n208,n25);
and (n507,n210,n23);
nand (n508,n118,n437);
nand (n509,n510,n59);
nand (n510,n511,n512);
or (n511,n243,n53);
nand (n512,n513,n51);
not (n513,n514);
and (n514,n243,n53);
or (n515,n516,n540);
and (n516,n517,n533);
xor (n517,n518,n526);
nand (n518,n519,n520);
or (n519,n167,n444);
nand (n520,n521,n525);
not (n521,n522);
nor (n522,n523,n524);
and (n523,n95,n175);
and (n524,n93,n174);
not (n525,n166);
nand (n526,n527,n532);
or (n527,n528,n190);
not (n528,n529);
nor (n529,n530,n531);
and (n530,n51,n163);
and (n531,n161,n52);
nand (n532,n460,n456);
nand (n533,n534,n539);
or (n534,n535,n102);
not (n535,n536);
or (n536,n537,n538);
and (n537,n187,n105);
and (n538,n185,n109);
or (n539,n464,n103);
and (n540,n518,n526);
and (n541,n495,n501);
and (n542,n490,n491);
and (n543,n485,n486);
xor (n544,n418,n476);
or (n545,n546,n981);
and (n546,n547,n581);
xor (n547,n548,n580);
or (n548,n549,n579);
and (n549,n550,n578);
xor (n550,n551,n552);
xor (n551,n427,n450);
or (n552,n553,n577);
and (n553,n554,n557);
xor (n554,n555,n556);
xor (n555,n452,n467);
xor (n556,n431,n442);
or (n557,n558,n576);
and (n558,n559,n572);
xor (n559,n560,n566);
nand (n560,n561,n565);
or (n561,n48,n562);
nor (n562,n563,n564);
and (n563,n245,n59);
and (n564,n243,n58);
or (n565,n469,n49);
nand (n566,n567,n571);
or (n567,n42,n568);
nor (n568,n569,n570);
and (n569,n33,n69);
and (n570,n29,n71);
or (n571,n19,n497);
nand (n572,n573,n575);
or (n573,n574,n502);
not (n574,n509);
or (n575,n503,n509);
and (n576,n560,n566);
and (n577,n555,n556);
xor (n578,n489,n492);
and (n579,n551,n552);
xor (n580,n484,n487);
nand (n581,n582,n977);
or (n582,n583,n955);
nor (n583,n584,n954);
and (n584,n585,n935);
or (n585,n586,n934);
and (n586,n587,n730);
xor (n587,n588,n699);
or (n588,n589,n698);
and (n589,n590,n660);
xor (n590,n591,n621);
xor (n591,n592,n611);
xor (n592,n593,n602);
nand (n593,n594,n598);
or (n594,n166,n595);
nor (n595,n596,n597);
and (n596,n161,n174);
and (n597,n163,n175);
or (n598,n599,n167);
nor (n599,n600,n601);
and (n600,n174,n87);
and (n601,n175,n89);
nand (n602,n603,n607);
or (n603,n190,n604);
nor (n604,n605,n606);
and (n605,n245,n52);
and (n606,n243,n51);
or (n607,n608,n191);
nor (n608,n609,n610);
and (n609,n155,n51);
and (n610,n157,n52);
nand (n611,n612,n617);
or (n612,n102,n613);
not (n613,n614);
nor (n614,n615,n616);
and (n615,n208,n105);
and (n616,n210,n109);
or (n617,n618,n103);
nor (n618,n619,n620);
and (n619,n179,n109);
and (n620,n181,n105);
or (n621,n622,n659);
and (n622,n623,n642);
xor (n623,n624,n633);
nand (n624,n625,n629);
or (n625,n116,n626);
nor (n626,n627,n628);
and (n627,n25,n63);
and (n628,n23,n65);
or (n629,n117,n630);
nor (n630,n631,n632);
and (n631,n71,n23);
and (n632,n69,n25);
nand (n633,n634,n638);
or (n634,n42,n635);
nor (n635,n636,n637);
and (n636,n87,n33);
and (n637,n29,n89);
or (n638,n19,n639);
nor (n639,n640,n641);
and (n640,n33,n93);
and (n641,n29,n95);
and (n642,n643,n649);
nor (n643,n644,n174);
nor (n644,n645,n648);
and (n645,n646,n33);
not (n646,n647);
and (n647,n243,n169);
and (n648,n245,n171);
nand (n649,n650,n655);
or (n650,n651,n102);
not (n651,n652);
nor (n652,n653,n654);
and (n653,n71,n109);
and (n654,n69,n105);
or (n655,n656,n103);
nor (n656,n657,n658);
and (n657,n203,n109);
and (n658,n202,n105);
and (n659,n624,n633);
xor (n660,n661,n683);
xor (n661,n662,n668);
nand (n662,n663,n664);
or (n663,n42,n639);
or (n664,n19,n665);
nor (n665,n666,n667);
and (n666,n33,n63);
and (n667,n29,n65);
xor (n668,n669,n674);
nor (n669,n670,n51);
nor (n670,n671,n673);
and (n671,n672,n174);
nand (n672,n243,n193);
and (n673,n245,n195);
nand (n674,n675,n680);
or (n675,n117,n676);
not (n676,n677);
nand (n677,n678,n679);
or (n678,n23,n202);
or (n679,n25,n203);
nand (n680,n681,n682);
not (n681,n630);
not (n682,n116);
or (n683,n684,n697);
and (n684,n685,n690);
xor (n685,n686,n687);
nor (n686,n191,n245);
nand (n687,n688,n689);
or (n688,n103,n613);
or (n689,n656,n102);
nand (n690,n691,n692);
or (n691,n167,n595);
nand (n692,n693,n525);
not (n693,n694);
or (n694,n695,n696);
and (n695,n157,n174);
and (n696,n155,n175);
and (n697,n686,n687);
and (n698,n591,n621);
xor (n699,n700,n715);
xor (n700,n701,n712);
xor (n701,n702,n709);
xor (n702,n703,n706);
nand (n703,n704,n705);
or (n704,n191,n528);
or (n705,n190,n608);
nand (n706,n707,n708);
or (n707,n618,n102);
nand (n708,n536,n104);
nand (n709,n710,n711);
or (n710,n42,n665);
or (n711,n19,n568);
or (n712,n713,n714);
and (n713,n661,n683);
and (n714,n662,n668);
xor (n715,n716,n721);
xor (n716,n717,n718);
and (n717,n669,n674);
or (n718,n719,n720);
and (n719,n592,n611);
and (n720,n593,n602);
xor (n721,n722,n727);
xor (n722,n723,n724);
nor (n723,n49,n245);
nand (n724,n725,n726);
or (n725,n676,n116);
or (n726,n117,n505);
nand (n727,n728,n729);
or (n728,n166,n599);
or (n729,n167,n522);
nand (n730,n731,n930,n933);
nand (n731,n732,n787,n923);
not (n732,n733);
nor (n733,n734,n761);
xor (n734,n735,n760);
xor (n735,n736,n759);
or (n736,n737,n758);
and (n737,n738,n752);
xor (n738,n739,n745);
nand (n739,n740,n744);
or (n740,n166,n741);
nor (n741,n742,n743);
and (n742,n245,n175);
and (n743,n243,n174);
or (n744,n694,n167);
nand (n745,n746,n751);
or (n746,n747,n116);
not (n747,n748);
nor (n748,n749,n750);
and (n749,n93,n23);
and (n750,n95,n25);
or (n751,n117,n626);
nand (n752,n753,n757);
or (n753,n42,n754);
nor (n754,n755,n756);
and (n755,n161,n33);
and (n756,n29,n163);
or (n757,n19,n635);
and (n758,n739,n745);
xor (n759,n685,n690);
xor (n760,n623,n642);
or (n761,n762,n786);
and (n762,n763,n785);
xor (n763,n764,n765);
xor (n764,n643,n649);
or (n765,n766,n784);
and (n766,n767,n777);
xor (n767,n768,n770);
and (n768,n769,n243);
not (n769,n167);
nand (n770,n771,n776);
or (n771,n102,n772);
not (n772,n773);
nor (n773,n774,n775);
and (n774,n65,n109);
and (n775,n63,n105);
nand (n776,n652,n104);
nand (n777,n778,n783);
or (n778,n779,n116);
not (n779,n780);
nor (n780,n781,n782);
and (n781,n89,n25);
and (n782,n87,n23);
nand (n783,n748,n118);
and (n784,n768,n770);
xor (n785,n738,n752);
and (n786,n764,n765);
or (n787,n788,n922);
and (n788,n789,n815);
xor (n789,n790,n814);
or (n790,n791,n813);
and (n791,n792,n812);
xor (n792,n793,n799);
nand (n793,n794,n798);
or (n794,n42,n795);
nor (n795,n796,n797);
and (n796,n33,n155);
and (n797,n29,n157);
or (n798,n754,n19);
and (n799,n800,n806);
and (n800,n801,n29);
nand (n801,n802,n803);
or (n802,n243,n22);
nand (n803,n804,n25);
not (n804,n805);
and (n805,n243,n22);
nand (n806,n807,n808);
or (n807,n103,n772);
or (n808,n809,n102);
nor (n809,n810,n811);
and (n810,n109,n93);
and (n811,n105,n95);
xor (n812,n767,n777);
and (n813,n793,n799);
xor (n814,n763,n785);
nand (n815,n816,n921);
or (n816,n817,n916);
nor (n817,n818,n915);
and (n818,n819,n894);
nand (n819,n820,n892);
or (n820,n821,n875);
not (n821,n822);
or (n822,n823,n874);
and (n823,n824,n853);
xor (n824,n825,n834);
nand (n825,n826,n830);
or (n826,n116,n827);
nor (n827,n828,n829);
and (n828,n23,n245);
and (n829,n243,n25);
or (n830,n117,n831);
nor (n831,n832,n833);
and (n832,n157,n23);
and (n833,n155,n25);
nand (n834,n835,n852);
or (n835,n836,n842);
not (n836,n837);
nand (n837,n838,n23);
nand (n838,n839,n841);
or (n839,n840,n105);
and (n840,n243,n121);
nand (n841,n245,n120);
not (n842,n843);
nand (n843,n844,n848);
or (n844,n845,n102);
or (n845,n846,n847);
and (n846,n161,n105);
and (n847,n163,n109);
or (n848,n849,n103);
nor (n849,n850,n851);
and (n850,n89,n105);
and (n851,n87,n109);
or (n852,n843,n837);
or (n853,n854,n873);
and (n854,n855,n863);
xor (n855,n856,n857);
nor (n856,n117,n245);
nand (n857,n858,n862);
or (n858,n859,n102);
nor (n859,n860,n861);
and (n860,n157,n105);
and (n861,n155,n109);
or (n862,n845,n103);
nor (n863,n864,n871);
nor (n864,n865,n867);
and (n865,n866,n104);
not (n866,n859);
and (n867,n868,n101);
nand (n868,n869,n870);
or (n869,n245,n105);
nand (n870,n105,n245);
or (n871,n872,n109);
and (n872,n243,n104);
and (n873,n856,n857);
and (n874,n825,n834);
not (n875,n876);
nand (n876,n877,n891);
not (n877,n878);
xor (n878,n879,n888);
xor (n879,n880,n882);
and (n880,n881,n243);
not (n881,n19);
nand (n882,n883,n884);
or (n883,n831,n116);
nand (n884,n885,n118);
nor (n885,n886,n887);
and (n886,n163,n25);
and (n887,n161,n23);
nand (n888,n889,n890);
or (n889,n849,n102);
or (n890,n809,n103);
nand (n891,n836,n843);
nand (n892,n893,n878);
not (n893,n891);
nand (n894,n895,n911);
not (n895,n896);
xor (n896,n897,n910);
xor (n897,n898,n902);
nand (n898,n899,n901);
or (n899,n900,n116);
not (n900,n885);
nand (n901,n780,n118);
nand (n902,n903,n908);
or (n903,n904,n42);
not (n904,n905);
nand (n905,n906,n907);
or (n906,n243,n33);
or (n907,n245,n29);
nand (n908,n909,n881);
not (n909,n795);
xor (n910,n800,n806);
not (n911,n912);
or (n912,n913,n914);
and (n913,n879,n888);
and (n914,n880,n882);
nor (n915,n895,n911);
nor (n916,n917,n918);
xor (n917,n792,n812);
or (n918,n919,n920);
and (n919,n897,n910);
and (n920,n898,n902);
nand (n921,n917,n918);
and (n922,n790,n814);
nand (n923,n924,n928);
not (n924,n925);
or (n925,n926,n927);
and (n926,n735,n760);
and (n927,n736,n759);
not (n928,n929);
xor (n929,n590,n660);
nand (n930,n931,n923);
not (n931,n932);
nand (n932,n734,n761);
nand (n933,n929,n925);
and (n934,n588,n699);
or (n935,n936,n951);
xor (n936,n937,n948);
xor (n937,n938,n939);
xor (n938,n559,n572);
xor (n939,n940,n947);
xor (n940,n941,n944);
or (n941,n942,n943);
and (n942,n722,n727);
and (n943,n723,n724);
or (n944,n945,n946);
and (n945,n702,n709);
and (n946,n703,n706);
xor (n947,n517,n533);
or (n948,n949,n950);
and (n949,n716,n721);
and (n950,n717,n718);
or (n951,n952,n953);
and (n952,n700,n715);
and (n953,n701,n712);
and (n954,n936,n951);
nand (n955,n956,n970);
not (n956,n957);
and (n957,n958,n966);
not (n958,n959);
xor (n959,n960,n965);
xor (n960,n961,n962);
xor (n961,n494,n515);
or (n962,n963,n964);
and (n963,n940,n947);
and (n964,n941,n944);
xor (n965,n554,n557);
not (n966,n967);
or (n967,n968,n969);
and (n968,n937,n948);
and (n969,n938,n939);
nand (n970,n971,n973);
not (n971,n972);
xor (n972,n550,n578);
not (n973,n974);
or (n974,n975,n976);
and (n975,n960,n965);
and (n976,n961,n962);
nor (n977,n978,n980);
and (n978,n970,n979);
nor (n979,n958,n966);
nor (n980,n971,n973);
and (n981,n548,n580);
and (n982,n482,n544);
and (n983,n984,n985);
not (n984,n8);
not (n985,n479);
and (n986,n987,n988);
not (n988,n2);
or (n989,n990,n986);
and (n990,n991,n2);
xor (n991,n992,n1696);
xor (n992,n993,n1694);
xor (n993,n994,n1693);
xor (n994,n995,n1684);
xor (n995,n996,n1683);
xor (n996,n997,n1668);
xor (n997,n998,n1667);
xor (n998,n999,n1646);
xor (n999,n1000,n1645);
xor (n1000,n1001,n1618);
xor (n1001,n1002,n1617);
xor (n1002,n1003,n1585);
xor (n1003,n1004,n1584);
xor (n1004,n1005,n1547);
xor (n1005,n1006,n204);
xor (n1006,n1007,n1502);
xor (n1007,n1008,n1501);
xor (n1008,n1009,n1451);
xor (n1009,n1010,n1450);
xor (n1010,n1011,n1394);
xor (n1011,n1012,n1393);
xor (n1012,n1013,n1330);
xor (n1013,n1014,n1329);
xor (n1014,n1015,n1261);
xor (n1015,n1016,n1260);
xor (n1016,n1017,n1188);
xor (n1017,n1018,n1187);
xor (n1018,n1019,n1107);
xor (n1019,n1020,n1106);
xor (n1020,n1021,n1024);
xor (n1021,n1022,n1023);
and (n1022,n110,n104);
and (n1023,n110,n105);
or (n1024,n1025,n1027);
and (n1025,n1022,n1026);
and (n1026,n134,n105);
and (n1027,n1028,n1029);
xor (n1028,n1022,n1026);
or (n1029,n1030,n1033);
and (n1030,n1031,n1032);
and (n1031,n134,n104);
and (n1032,n128,n105);
and (n1033,n1034,n1035);
xor (n1034,n1031,n1032);
or (n1035,n1036,n1039);
and (n1036,n1037,n1038);
and (n1037,n128,n104);
and (n1038,n31,n105);
and (n1039,n1040,n1041);
xor (n1040,n1037,n1038);
or (n1041,n1042,n1045);
and (n1042,n1043,n1044);
and (n1043,n31,n104);
and (n1044,n38,n105);
and (n1045,n1046,n1047);
xor (n1046,n1043,n1044);
or (n1047,n1048,n1051);
and (n1048,n1049,n1050);
and (n1049,n38,n104);
and (n1050,n185,n105);
and (n1051,n1052,n1053);
xor (n1052,n1049,n1050);
or (n1053,n1054,n1057);
and (n1054,n1055,n1056);
and (n1055,n185,n104);
and (n1056,n179,n105);
and (n1057,n1058,n1059);
xor (n1058,n1055,n1056);
or (n1059,n1060,n1062);
and (n1060,n1061,n615);
and (n1061,n179,n104);
and (n1062,n1063,n1064);
xor (n1063,n1061,n615);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
and (n1066,n208,n104);
and (n1067,n203,n105);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1073);
and (n1071,n1072,n654);
and (n1072,n203,n104);
and (n1073,n1074,n1075);
xor (n1074,n1072,n654);
or (n1075,n1076,n1078);
and (n1076,n1077,n775);
and (n1077,n69,n104);
and (n1078,n1079,n1080);
xor (n1079,n1077,n775);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
and (n1082,n63,n104);
and (n1083,n93,n105);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
and (n1088,n93,n104);
and (n1089,n87,n105);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1095);
and (n1093,n1094,n846);
and (n1094,n87,n104);
and (n1095,n1096,n1097);
xor (n1096,n1094,n846);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
and (n1099,n161,n104);
and (n1100,n155,n105);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
and (n1103,n1104,n1105);
and (n1104,n155,n104);
and (n1105,n243,n105);
and (n1106,n134,n121);
or (n1107,n1108,n1111);
and (n1108,n1109,n1110);
xor (n1109,n1028,n1029);
and (n1110,n128,n121);
and (n1111,n1112,n1113);
xor (n1112,n1109,n1110);
or (n1113,n1114,n1117);
and (n1114,n1115,n1116);
xor (n1115,n1034,n1035);
and (n1116,n31,n121);
and (n1117,n1118,n1119);
xor (n1118,n1115,n1116);
or (n1119,n1120,n1123);
and (n1120,n1121,n1122);
xor (n1121,n1040,n1041);
and (n1122,n38,n121);
and (n1123,n1124,n1125);
xor (n1124,n1121,n1122);
or (n1125,n1126,n1129);
and (n1126,n1127,n1128);
xor (n1127,n1046,n1047);
and (n1128,n185,n121);
and (n1129,n1130,n1131);
xor (n1130,n1127,n1128);
or (n1131,n1132,n1135);
and (n1132,n1133,n1134);
xor (n1133,n1052,n1053);
and (n1134,n179,n121);
and (n1135,n1136,n1137);
xor (n1136,n1133,n1134);
or (n1137,n1138,n1141);
and (n1138,n1139,n1140);
xor (n1139,n1058,n1059);
and (n1140,n208,n121);
and (n1141,n1142,n1143);
xor (n1142,n1139,n1140);
or (n1143,n1144,n1147);
and (n1144,n1145,n1146);
xor (n1145,n1063,n1064);
and (n1146,n203,n121);
and (n1147,n1148,n1149);
xor (n1148,n1145,n1146);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
xor (n1151,n1069,n1070);
and (n1152,n69,n121);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
xor (n1157,n1074,n1075);
and (n1158,n63,n121);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n1079,n1080);
and (n1164,n93,n121);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1085,n1086);
and (n1170,n87,n121);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1091,n1092);
and (n1176,n161,n121);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1096,n1097);
and (n1182,n155,n121);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
and (n1185,n1186,n840);
xor (n1186,n1102,n1103);
and (n1187,n128,n23);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1112,n1113);
and (n1191,n31,n23);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1118,n1119);
and (n1197,n38,n23);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1124,n1125);
and (n1203,n185,n23);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1130,n1131);
and (n1209,n179,n23);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1136,n1137);
and (n1215,n208,n23);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1142,n1143);
and (n1221,n203,n23);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1148,n1149);
and (n1227,n69,n23);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1154,n1155);
and (n1233,n63,n23);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
or (n1236,n1237,n1239);
and (n1237,n1238,n749);
xor (n1238,n1160,n1161);
and (n1239,n1240,n1241);
xor (n1240,n1238,n749);
or (n1241,n1242,n1244);
and (n1242,n1243,n782);
xor (n1243,n1166,n1167);
and (n1244,n1245,n1246);
xor (n1245,n1243,n782);
or (n1246,n1247,n1249);
and (n1247,n1248,n887);
xor (n1248,n1172,n1173);
and (n1249,n1250,n1251);
xor (n1250,n1248,n887);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1178,n1179);
and (n1254,n155,n23);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
and (n1257,n1258,n1259);
xor (n1258,n1184,n1185);
and (n1259,n243,n23);
and (n1260,n31,n22);
or (n1261,n1262,n1265);
and (n1262,n1263,n1264);
xor (n1263,n1193,n1194);
and (n1264,n38,n22);
and (n1265,n1266,n1267);
xor (n1266,n1263,n1264);
or (n1267,n1268,n1271);
and (n1268,n1269,n1270);
xor (n1269,n1199,n1200);
and (n1270,n185,n22);
and (n1271,n1272,n1273);
xor (n1272,n1269,n1270);
or (n1273,n1274,n1277);
and (n1274,n1275,n1276);
xor (n1275,n1205,n1206);
and (n1276,n179,n22);
and (n1277,n1278,n1279);
xor (n1278,n1275,n1276);
or (n1279,n1280,n1283);
and (n1280,n1281,n1282);
xor (n1281,n1211,n1212);
and (n1282,n208,n22);
and (n1283,n1284,n1285);
xor (n1284,n1281,n1282);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1217,n1218);
and (n1288,n203,n22);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1223,n1224);
and (n1294,n69,n22);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
or (n1297,n1298,n1301);
and (n1298,n1299,n1300);
xor (n1299,n1229,n1230);
and (n1300,n63,n22);
and (n1301,n1302,n1303);
xor (n1302,n1299,n1300);
or (n1303,n1304,n1307);
and (n1304,n1305,n1306);
xor (n1305,n1235,n1236);
and (n1306,n93,n22);
and (n1307,n1308,n1309);
xor (n1308,n1305,n1306);
or (n1309,n1310,n1313);
and (n1310,n1311,n1312);
xor (n1311,n1240,n1241);
and (n1312,n87,n22);
and (n1313,n1314,n1315);
xor (n1314,n1311,n1312);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1245,n1246);
and (n1318,n161,n22);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1250,n1251);
and (n1324,n155,n22);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
and (n1327,n1328,n805);
xor (n1328,n1256,n1257);
and (n1329,n38,n29);
or (n1330,n1331,n1334);
and (n1331,n1332,n1333);
xor (n1332,n1266,n1267);
and (n1333,n185,n29);
and (n1334,n1335,n1336);
xor (n1335,n1332,n1333);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1272,n1273);
and (n1339,n179,n29);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1278,n1279);
and (n1345,n208,n29);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
or (n1348,n1349,n1352);
and (n1349,n1350,n1351);
xor (n1350,n1284,n1285);
and (n1351,n203,n29);
and (n1352,n1353,n1354);
xor (n1353,n1350,n1351);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1290,n1291);
and (n1357,n69,n29);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1296,n1297);
and (n1363,n63,n29);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1302,n1303);
and (n1369,n93,n29);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1308,n1309);
and (n1375,n87,n29);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1314,n1315);
and (n1381,n161,n29);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1320,n1321);
and (n1387,n155,n29);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
and (n1390,n1391,n1392);
xor (n1391,n1326,n1327);
and (n1392,n243,n29);
and (n1393,n185,n169);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1335,n1336);
and (n1397,n179,n169);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
or (n1400,n1401,n1404);
and (n1401,n1402,n1403);
xor (n1402,n1341,n1342);
and (n1403,n208,n169);
and (n1404,n1405,n1406);
xor (n1405,n1402,n1403);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1347,n1348);
and (n1409,n203,n169);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1353,n1354);
and (n1415,n69,n169);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1359,n1360);
and (n1421,n63,n169);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1365,n1366);
and (n1427,n93,n169);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1371,n1372);
and (n1433,n87,n169);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1377,n1378);
and (n1439,n161,n169);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1383,n1384);
and (n1445,n155,n169);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
and (n1448,n1449,n647);
xor (n1449,n1389,n1390);
and (n1450,n179,n175);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1399,n1400);
and (n1454,n208,n175);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
or (n1457,n1458,n1461);
and (n1458,n1459,n1460);
xor (n1459,n1405,n1406);
and (n1460,n203,n175);
and (n1461,n1462,n1463);
xor (n1462,n1459,n1460);
or (n1463,n1464,n1467);
and (n1464,n1465,n1466);
xor (n1465,n1411,n1412);
and (n1466,n69,n175);
and (n1467,n1468,n1469);
xor (n1468,n1465,n1466);
or (n1469,n1470,n1473);
and (n1470,n1471,n1472);
xor (n1471,n1417,n1418);
and (n1472,n63,n175);
and (n1473,n1474,n1475);
xor (n1474,n1471,n1472);
or (n1475,n1476,n1479);
and (n1476,n1477,n1478);
xor (n1477,n1423,n1424);
and (n1478,n93,n175);
and (n1479,n1480,n1481);
xor (n1480,n1477,n1478);
or (n1481,n1482,n1485);
and (n1482,n1483,n1484);
xor (n1483,n1429,n1430);
and (n1484,n87,n175);
and (n1485,n1486,n1487);
xor (n1486,n1483,n1484);
or (n1487,n1488,n1491);
and (n1488,n1489,n1490);
xor (n1489,n1435,n1436);
and (n1490,n161,n175);
and (n1491,n1492,n1493);
xor (n1492,n1489,n1490);
or (n1493,n1494,n1496);
and (n1494,n1495,n696);
xor (n1495,n1441,n1442);
and (n1496,n1497,n1498);
xor (n1497,n1495,n696);
and (n1498,n1499,n1500);
xor (n1499,n1447,n1448);
and (n1500,n243,n175);
and (n1501,n208,n193);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1456,n1457);
and (n1505,n203,n193);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1462,n1463);
and (n1511,n69,n193);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1468,n1469);
and (n1517,n63,n193);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
or (n1520,n1521,n1524);
and (n1521,n1522,n1523);
xor (n1522,n1474,n1475);
and (n1523,n93,n193);
and (n1524,n1525,n1526);
xor (n1525,n1522,n1523);
or (n1526,n1527,n1530);
and (n1527,n1528,n1529);
xor (n1528,n1480,n1481);
and (n1529,n87,n193);
and (n1530,n1531,n1532);
xor (n1531,n1528,n1529);
or (n1532,n1533,n1536);
and (n1533,n1534,n1535);
xor (n1534,n1486,n1487);
and (n1535,n161,n193);
and (n1536,n1537,n1538);
xor (n1537,n1534,n1535);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1492,n1493);
and (n1541,n155,n193);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
and (n1544,n1545,n1546);
xor (n1545,n1497,n1498);
not (n1546,n672);
or (n1547,n1548,n1551);
and (n1548,n1549,n1550);
xor (n1549,n1507,n1508);
and (n1550,n69,n52);
and (n1551,n1552,n1553);
xor (n1552,n1549,n1550);
or (n1553,n1554,n1557);
and (n1554,n1555,n1556);
xor (n1555,n1513,n1514);
and (n1556,n63,n52);
and (n1557,n1558,n1559);
xor (n1558,n1555,n1556);
or (n1559,n1560,n1562);
and (n1560,n1561,n317);
xor (n1561,n1519,n1520);
and (n1562,n1563,n1564);
xor (n1563,n1561,n317);
or (n1564,n1565,n1568);
and (n1565,n1566,n1567);
xor (n1566,n1525,n1526);
and (n1567,n87,n52);
and (n1568,n1569,n1570);
xor (n1569,n1566,n1567);
or (n1570,n1571,n1573);
and (n1571,n1572,n531);
xor (n1572,n1531,n1532);
and (n1573,n1574,n1575);
xor (n1574,n1572,n531);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1537,n1538);
and (n1578,n155,n52);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
and (n1581,n1582,n1583);
xor (n1582,n1543,n1544);
and (n1583,n243,n52);
and (n1584,n69,n53);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1552,n1553);
and (n1588,n63,n53);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1558,n1559);
and (n1594,n93,n53);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
or (n1597,n1598,n1601);
and (n1598,n1599,n1600);
xor (n1599,n1563,n1564);
and (n1600,n87,n53);
and (n1601,n1602,n1603);
xor (n1602,n1599,n1600);
or (n1603,n1604,n1607);
and (n1604,n1605,n1606);
xor (n1605,n1569,n1570);
and (n1606,n161,n53);
and (n1607,n1608,n1609);
xor (n1608,n1605,n1606);
or (n1609,n1610,n1613);
and (n1610,n1611,n1612);
xor (n1611,n1574,n1575);
and (n1612,n155,n53);
and (n1613,n1614,n1615);
xor (n1614,n1611,n1612);
and (n1615,n1616,n514);
xor (n1616,n1580,n1581);
and (n1617,n63,n59);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1590,n1591);
and (n1621,n93,n59);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1596,n1597);
and (n1627,n87,n59);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1602,n1603);
and (n1633,n161,n59);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1608,n1609);
and (n1639,n155,n59);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
and (n1642,n1643,n1644);
xor (n1643,n1614,n1615);
and (n1644,n243,n59);
and (n1645,n93,n78);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1623,n1624);
and (n1649,n87,n78);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1629,n1630);
and (n1655,n161,n78);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1635,n1636);
and (n1661,n155,n78);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
and (n1664,n1665,n1666);
xor (n1665,n1641,n1642);
not (n1666,n242);
and (n1667,n87,n79);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1651,n1652);
and (n1671,n161,n79);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1657,n1658);
and (n1677,n155,n79);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
and (n1680,n1681,n1682);
xor (n1681,n1663,n1664);
and (n1682,n243,n79);
and (n1683,n161,n145);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1673,n1674);
and (n1687,n155,n145);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
and (n1690,n1691,n1692);
xor (n1691,n1679,n1680);
not (n1692,n265);
and (n1693,n155,n151);
and (n1694,n1695,n1696);
xor (n1695,n1689,n1690);
and (n1696,n243,n151);
endmodule
