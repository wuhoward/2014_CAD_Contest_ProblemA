module top (out,n17,n18,n24,n28,n34,n44,n45,n53,n59
        ,n71,n72,n80,n86,n100,n106,n110,n116,n131,n146
        ,n147,n155,n161,n212,n213,n323,n329,n354,n402,n410
        ,n414,n436,n470);
output out;
input n17;
input n18;
input n24;
input n28;
input n34;
input n44;
input n45;
input n53;
input n59;
input n71;
input n72;
input n80;
input n86;
input n100;
input n106;
input n110;
input n116;
input n131;
input n146;
input n147;
input n155;
input n161;
input n212;
input n213;
input n323;
input n329;
input n354;
input n402;
input n410;
input n414;
input n436;
input n470;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n411;
wire n412;
wire n413;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
xor (out,n0,n1424);
nand (n0,n1,n1423);
or (n1,n2,n282);
not (n2,n3);
nand (n3,n4,n281);
or (n4,n5,n241);
or (n5,n6,n240);
and (n6,n7,n199);
xor (n7,n8,n121);
or (n8,n9,n120);
and (n9,n10,n62);
xor (n10,n11,n37);
nand (n11,n12,n31);
or (n12,n13,n26);
nand (n13,n14,n21);
nor (n14,n15,n19);
and (n15,n16,n18);
not (n16,n17);
and (n19,n17,n20);
not (n20,n18);
nand (n21,n22,n25);
nand (n22,n23,n18);
not (n23,n24);
nand (n25,n24,n20);
nor (n26,n27,n29);
and (n27,n23,n28);
and (n29,n24,n30);
not (n30,n28);
or (n31,n14,n32);
nor (n32,n33,n35);
and (n33,n23,n34);
and (n35,n24,n36);
not (n36,n34);
not (n37,n38);
nand (n38,n39,n56);
or (n39,n40,n51);
nand (n40,n41,n48);
nor (n41,n42,n46);
and (n42,n43,n45);
not (n43,n44);
and (n46,n44,n47);
not (n47,n45);
nand (n48,n49,n50);
or (n49,n16,n45);
nand (n50,n16,n45);
nor (n51,n52,n54);
and (n52,n16,n53);
and (n54,n17,n55);
not (n55,n53);
or (n56,n41,n57);
nor (n57,n58,n60);
and (n58,n16,n59);
and (n60,n17,n61);
not (n61,n59);
or (n62,n63,n119);
and (n63,n64,n95);
xor (n64,n65,n89);
nand (n65,n66,n83);
or (n66,n67,n78);
nand (n67,n68,n75);
or (n68,n69,n73);
and (n69,n70,n72);
not (n70,n71);
and (n73,n71,n74);
not (n74,n72);
nor (n75,n76,n77);
and (n76,n24,n70);
and (n77,n23,n71);
nor (n78,n79,n81);
and (n79,n74,n80);
and (n81,n72,n82);
not (n82,n80);
or (n83,n84,n75);
nor (n84,n85,n87);
and (n85,n86,n74);
and (n87,n72,n88);
not (n88,n86);
nand (n89,n90,n94);
or (n90,n40,n91);
nor (n91,n92,n93);
and (n92,n16,n34);
and (n93,n17,n36);
or (n94,n41,n51);
nand (n95,n96,n113);
or (n96,n97,n108);
nand (n97,n98,n103);
nor (n98,n99,n101);
and (n99,n74,n100);
and (n101,n72,n102);
not (n102,n100);
nand (n103,n104,n107);
or (n104,n105,n100);
not (n105,n106);
nand (n107,n105,n100);
nor (n108,n109,n111);
and (n109,n110,n105);
and (n111,n106,n112);
not (n112,n110);
or (n113,n114,n98);
nor (n114,n115,n117);
and (n115,n116,n105);
and (n117,n106,n118);
not (n118,n116);
and (n119,n65,n89);
and (n120,n11,n37);
xor (n121,n122,n185);
xor (n122,n123,n165);
or (n123,n124,n164);
and (n124,n125,n140);
xor (n125,n126,n134);
nand (n126,n127,n128);
or (n127,n67,n84);
or (n128,n129,n75);
nor (n129,n130,n132);
and (n130,n74,n131);
and (n132,n72,n133);
not (n133,n131);
nand (n134,n135,n136);
or (n135,n97,n114);
or (n136,n98,n137);
nor (n137,n138,n139);
and (n138,n105,n80);
and (n139,n106,n82);
nand (n140,n141,n158);
or (n141,n142,n153);
nand (n142,n143,n150);
nor (n143,n144,n148);
and (n144,n145,n147);
not (n145,n146);
and (n148,n146,n149);
not (n149,n147);
nand (n150,n151,n152);
or (n151,n147,n43);
nand (n152,n43,n147);
nor (n153,n154,n156);
and (n154,n43,n155);
and (n156,n44,n157);
not (n157,n155);
or (n158,n143,n159);
nor (n159,n160,n162);
and (n160,n43,n161);
and (n162,n44,n163);
not (n163,n161);
and (n164,n126,n134);
xor (n165,n166,n178);
xor (n166,n167,n172);
nand (n167,n168,n171);
or (n168,n169,n170);
not (n169,n143);
not (n170,n142);
not (n171,n159);
nand (n172,n173,n174);
or (n173,n40,n57);
or (n174,n41,n175);
nor (n175,n176,n177);
and (n176,n16,n155);
and (n177,n17,n157);
nand (n178,n179,n184);
or (n179,n75,n180);
not (n180,n181);
nand (n181,n182,n183);
or (n182,n72,n30);
or (n183,n74,n28);
or (n184,n67,n129);
xor (n185,n186,n38);
xor (n186,n187,n193);
nand (n187,n188,n189);
or (n188,n97,n137);
or (n189,n190,n98);
nor (n190,n191,n192);
and (n191,n105,n86);
and (n192,n106,n88);
nand (n193,n194,n195);
or (n194,n13,n32);
or (n195,n14,n196);
nor (n196,n197,n198);
and (n197,n23,n53);
and (n198,n24,n55);
or (n199,n200,n239);
and (n200,n201,n238);
xor (n201,n202,n237);
or (n202,n203,n236);
and (n203,n204,n230);
xor (n204,n205,n224);
nand (n205,n206,n220);
or (n206,n207,n219);
not (n207,n208);
nand (n208,n209,n216);
nor (n209,n210,n214);
and (n210,n211,n213);
not (n211,n212);
and (n214,n212,n215);
not (n215,n213);
nand (n216,n217,n218);
or (n217,n212,n145);
nand (n218,n145,n212);
not (n219,n209);
not (n220,n221);
nor (n221,n222,n223);
and (n222,n145,n161);
and (n223,n146,n163);
nand (n224,n225,n229);
or (n225,n142,n226);
nor (n226,n227,n228);
and (n227,n43,n59);
and (n228,n44,n61);
or (n229,n143,n153);
nand (n230,n231,n235);
or (n231,n13,n232);
nor (n232,n233,n234);
and (n233,n23,n131);
and (n234,n24,n133);
or (n235,n14,n26);
and (n236,n205,n224);
xor (n237,n125,n140);
xor (n238,n10,n62);
and (n239,n202,n237);
and (n240,n8,n121);
xor (n241,n242,n278);
xor (n242,n243,n246);
or (n243,n244,n245);
and (n244,n186,n38);
and (n245,n187,n193);
xor (n246,n247,n258);
xor (n247,n248,n255);
not (n248,n249);
nand (n249,n250,n251);
or (n250,n40,n175);
or (n251,n41,n252);
nor (n252,n253,n254);
and (n253,n16,n161);
and (n254,n17,n163);
or (n255,n256,n257);
and (n256,n166,n178);
and (n257,n167,n172);
xor (n258,n259,n272);
xor (n259,n260,n266);
nand (n260,n261,n262);
or (n261,n97,n190);
or (n262,n98,n263);
nor (n263,n264,n265);
and (n264,n105,n131);
and (n265,n106,n133);
nand (n266,n267,n268);
or (n267,n13,n196);
or (n268,n14,n269);
nor (n269,n270,n271);
and (n270,n23,n59);
and (n271,n24,n61);
nand (n272,n273,n274);
or (n273,n180,n67);
or (n274,n275,n75);
nor (n275,n276,n277);
and (n276,n74,n34);
and (n277,n72,n36);
or (n278,n279,n280);
and (n279,n122,n185);
and (n280,n123,n165);
nand (n281,n5,n241);
not (n282,n283);
nand (n283,n284,n1422);
or (n284,n285,n1417);
nor (n285,n286,n1413);
and (n286,n287,n1375);
nand (n287,n288,n1364);
or (n288,n289,n863);
nand (n289,n290,n742,n858);
nor (n290,n291,n678);
nor (n291,n292,n586);
xor (n292,n293,n538);
xor (n293,n294,n384);
xor (n294,n295,n361);
xor (n295,n296,n333);
or (n296,n297,n332);
and (n297,n298,n319);
xor (n298,n299,n310);
nand (n299,n300,n305);
or (n300,n209,n301);
not (n301,n302);
nand (n302,n303,n304);
or (n303,n146,n55);
or (n304,n145,n53);
nand (n305,n306,n207);
not (n306,n307);
nor (n307,n308,n309);
and (n308,n34,n145);
and (n309,n36,n146);
nand (n310,n311,n315);
or (n311,n13,n312);
nor (n312,n313,n314);
and (n313,n110,n23);
and (n314,n24,n112);
or (n315,n316,n14);
nor (n316,n317,n318);
and (n317,n116,n23);
and (n318,n24,n118);
nand (n319,n320,n326);
or (n320,n67,n321);
nor (n321,n322,n324);
and (n322,n323,n74);
and (n324,n72,n325);
not (n325,n323);
or (n326,n327,n75);
nor (n327,n328,n330);
and (n328,n329,n74);
and (n330,n72,n331);
not (n331,n329);
and (n332,n299,n310);
xor (n333,n334,n350);
xor (n334,n335,n344);
nand (n335,n336,n340);
or (n336,n142,n337);
nor (n337,n338,n339);
and (n338,n43,n28);
and (n339,n44,n30);
or (n340,n143,n341);
nor (n341,n342,n343);
and (n342,n43,n34);
and (n343,n44,n36);
nand (n344,n345,n346);
or (n345,n67,n327);
or (n346,n347,n75);
nor (n347,n348,n349);
and (n348,n110,n74);
and (n349,n72,n112);
nand (n350,n351,n357);
or (n351,n97,n352);
nor (n352,n353,n355);
and (n353,n354,n105);
and (n355,n106,n356);
not (n356,n354);
or (n357,n358,n98);
nor (n358,n359,n360);
and (n359,n323,n105);
and (n360,n106,n325);
xor (n361,n362,n378);
xor (n362,n363,n369);
nand (n363,n364,n365);
or (n364,n301,n208);
or (n365,n209,n366);
nor (n366,n367,n368);
and (n367,n145,n59);
and (n368,n146,n61);
nand (n369,n370,n374);
or (n370,n40,n371);
nor (n371,n372,n373);
and (n372,n16,n86);
and (n373,n17,n88);
or (n374,n41,n375);
nor (n375,n376,n377);
and (n376,n16,n131);
and (n377,n17,n133);
nand (n378,n379,n380);
or (n379,n13,n316);
or (n380,n14,n381);
nor (n381,n382,n383);
and (n382,n80,n23);
and (n383,n24,n82);
or (n384,n385,n537);
and (n385,n386,n509);
xor (n386,n387,n450);
or (n387,n388,n449);
and (n388,n389,n419);
xor (n389,n390,n397);
nand (n390,n391,n396);
or (n391,n67,n392);
not (n392,n393);
nand (n393,n394,n395);
or (n394,n356,n72);
or (n395,n74,n354);
or (n396,n321,n75);
xor (n397,n398,n405);
nor (n398,n399,n105);
nor (n399,n400,n403);
and (n400,n401,n74);
nand (n401,n402,n100);
and (n403,n404,n102);
not (n404,n402);
nand (n405,n406,n415);
or (n406,n407,n412);
nor (n407,n408,n411);
and (n408,n155,n409);
not (n409,n410);
and (n411,n157,n410);
nand (n412,n413,n410);
not (n413,n414);
or (n415,n416,n413);
nor (n416,n417,n418);
and (n417,n409,n161);
and (n418,n410,n163);
or (n419,n420,n448);
and (n420,n421,n429);
xor (n421,n422,n423);
nor (n422,n98,n404);
nand (n423,n424,n428);
or (n424,n425,n412);
nor (n425,n426,n427);
and (n426,n410,n61);
nor (n427,n410,n61);
or (n428,n407,n413);
nand (n429,n430,n444);
or (n430,n431,n441);
nand (n431,n432,n438);
not (n432,n433);
nand (n433,n434,n437);
or (n434,n435,n410);
not (n435,n436);
nand (n437,n435,n410);
nand (n438,n439,n440);
or (n439,n435,n213);
nand (n440,n213,n435);
nor (n441,n442,n443);
and (n442,n215,n34);
and (n443,n213,n36);
or (n444,n432,n445);
nor (n445,n446,n447);
and (n446,n215,n53);
and (n447,n213,n55);
and (n448,n422,n423);
and (n449,n390,n397);
xor (n450,n451,n483);
xor (n451,n452,n453);
and (n452,n398,n405);
or (n453,n454,n482);
and (n454,n455,n473);
xor (n455,n456,n462);
nand (n456,n457,n458);
or (n457,n431,n445);
or (n458,n432,n459);
nor (n459,n460,n461);
and (n460,n215,n59);
and (n461,n213,n61);
nand (n462,n463,n467);
or (n463,n97,n464);
nor (n464,n465,n466);
and (n465,n404,n106);
and (n466,n402,n105);
or (n467,n468,n98);
nor (n468,n469,n471);
and (n469,n470,n105);
and (n471,n472,n106);
not (n472,n470);
nand (n473,n474,n478);
or (n474,n142,n475);
nor (n475,n476,n477);
and (n476,n43,n86);
and (n477,n44,n88);
or (n478,n143,n479);
nor (n479,n480,n481);
and (n480,n43,n131);
and (n481,n44,n133);
and (n482,n456,n462);
or (n483,n484,n508);
and (n484,n485,n502);
xor (n485,n486,n496);
nand (n486,n487,n492);
or (n487,n41,n488);
not (n488,n489);
nor (n489,n490,n491);
and (n490,n82,n16);
and (n491,n80,n17);
or (n492,n40,n493);
nor (n493,n494,n495);
and (n494,n16,n116);
and (n495,n17,n118);
nand (n496,n497,n501);
or (n497,n208,n498);
nor (n498,n499,n500);
and (n499,n145,n28);
and (n500,n146,n30);
or (n501,n209,n307);
nand (n502,n503,n507);
or (n503,n13,n504);
nor (n504,n505,n506);
and (n505,n23,n329);
and (n506,n24,n331);
or (n507,n14,n312);
and (n508,n486,n496);
or (n509,n510,n536);
and (n510,n511,n535);
xor (n511,n512,n534);
or (n512,n513,n533);
and (n513,n514,n527);
xor (n514,n515,n521);
nand (n515,n516,n520);
or (n516,n142,n517);
nor (n517,n518,n519);
and (n518,n80,n43);
and (n519,n44,n82);
or (n520,n475,n143);
nand (n521,n522,n526);
or (n522,n40,n523);
nor (n523,n524,n525);
and (n524,n16,n110);
and (n525,n17,n112);
or (n526,n493,n41);
nand (n527,n528,n532);
or (n528,n208,n529);
nor (n529,n530,n531);
and (n530,n145,n131);
and (n531,n146,n133);
or (n532,n209,n498);
and (n533,n515,n521);
xor (n534,n485,n502);
xor (n535,n455,n473);
and (n536,n512,n534);
and (n537,n387,n450);
xor (n538,n539,n578);
xor (n539,n540,n543);
or (n540,n541,n542);
and (n541,n451,n483);
and (n542,n452,n453);
xor (n543,n544,n565);
xor (n544,n545,n555);
not (n545,n546);
nand (n546,n547,n551);
or (n547,n431,n548);
nor (n548,n549,n550);
and (n549,n215,n155);
and (n550,n213,n157);
or (n551,n432,n552);
nor (n552,n553,n554);
and (n553,n215,n161);
and (n554,n213,n163);
nand (n555,n556,n561);
not (n556,n557);
nand (n557,n558,n560);
or (n558,n559,n414);
not (n559,n412);
not (n560,n416);
not (n561,n562);
nand (n562,n563,n564);
or (n563,n431,n459);
or (n564,n432,n548);
or (n565,n566,n577);
and (n566,n567,n574);
xor (n567,n568,n571);
nand (n568,n569,n570);
or (n569,n97,n468);
or (n570,n352,n98);
nand (n571,n572,n573);
or (n572,n142,n479);
or (n573,n143,n337);
nand (n574,n575,n576);
or (n575,n40,n488);
or (n576,n371,n41);
and (n577,n568,n571);
or (n578,n579,n585);
and (n579,n580,n584);
xor (n580,n581,n582);
xor (n581,n298,n319);
nand (n582,n583,n555);
or (n583,n556,n561);
xor (n584,n567,n574);
and (n585,n581,n582);
or (n586,n587,n677);
and (n587,n588,n676);
xor (n588,n589,n590);
xor (n589,n580,n584);
or (n590,n591,n675);
and (n591,n592,n624);
xor (n592,n593,n623);
or (n593,n594,n622);
and (n594,n595,n610);
xor (n595,n596,n602);
nand (n596,n597,n601);
or (n597,n13,n598);
nor (n598,n599,n600);
and (n599,n323,n23);
and (n600,n24,n325);
or (n601,n14,n504);
nand (n602,n603,n604);
or (n603,n75,n392);
nand (n604,n605,n609);
not (n605,n606);
nor (n606,n607,n608);
and (n607,n74,n470);
and (n608,n472,n72);
not (n609,n67);
and (n610,n611,n616);
nor (n611,n612,n74);
nor (n612,n613,n615);
and (n613,n614,n23);
nand (n614,n71,n402);
and (n615,n404,n70);
nand (n616,n617,n621);
or (n617,n618,n412);
nor (n618,n619,n620);
and (n619,n409,n53);
and (n620,n410,n55);
or (n621,n425,n413);
and (n622,n596,n602);
xor (n623,n389,n419);
or (n624,n625,n674);
and (n625,n626,n673);
xor (n626,n627,n651);
or (n627,n628,n650);
and (n628,n629,n643);
xor (n629,n630,n636);
nand (n630,n631,n635);
or (n631,n431,n632);
nor (n632,n633,n634);
and (n633,n28,n215);
and (n634,n30,n213);
or (n635,n432,n441);
nand (n636,n637,n642);
or (n637,n638,n142);
not (n638,n639);
nand (n639,n640,n641);
or (n640,n44,n118);
or (n641,n43,n116);
or (n642,n517,n143);
nand (n643,n644,n649);
or (n644,n40,n645);
not (n645,n646);
nor (n646,n647,n648);
and (n647,n331,n16);
and (n648,n329,n17);
or (n649,n523,n41);
and (n650,n630,n636);
or (n651,n652,n672);
and (n652,n653,n666);
xor (n653,n654,n660);
nand (n654,n655,n659);
or (n655,n208,n656);
nor (n656,n657,n658);
and (n657,n145,n86);
and (n658,n146,n88);
or (n659,n209,n529);
nand (n660,n661,n665);
or (n661,n13,n662);
nor (n662,n663,n664);
and (n663,n354,n23);
and (n664,n24,n356);
or (n665,n598,n14);
nand (n666,n667,n671);
or (n667,n67,n668);
nor (n668,n669,n670);
and (n669,n404,n72);
and (n670,n402,n74);
or (n671,n606,n75);
and (n672,n654,n660);
xor (n673,n421,n429);
and (n674,n627,n651);
and (n675,n593,n623);
xor (n676,n386,n509);
and (n677,n589,n590);
nor (n678,n679,n741);
or (n679,n680,n740);
and (n680,n681,n739);
xor (n681,n682,n683);
xor (n682,n511,n535);
or (n683,n684,n738);
and (n684,n685,n688);
xor (n685,n686,n687);
xor (n686,n514,n527);
xor (n687,n595,n610);
or (n688,n689,n737);
and (n689,n690,n713);
xor (n690,n691,n692);
xor (n691,n611,n616);
or (n692,n693,n712);
and (n693,n694,n705);
xor (n694,n695,n697);
and (n695,n696,n402);
not (n696,n75);
nand (n697,n698,n703);
or (n698,n699,n431);
not (n699,n700);
nand (n700,n701,n702);
or (n701,n213,n133);
or (n702,n215,n131);
nand (n703,n704,n433);
not (n704,n632);
nand (n705,n706,n711);
or (n706,n142,n707);
not (n707,n708);
nand (n708,n709,n710);
or (n709,n44,n112);
or (n710,n43,n110);
or (n711,n143,n638);
and (n712,n695,n697);
or (n713,n714,n736);
and (n714,n715,n730);
xor (n715,n716,n724);
nand (n716,n717,n722);
or (n717,n718,n40);
not (n718,n719);
nand (n719,n720,n721);
or (n720,n17,n325);
or (n721,n16,n323);
nand (n722,n646,n723);
not (n723,n41);
nand (n724,n725,n726);
or (n725,n413,n618);
or (n726,n727,n412);
nor (n727,n728,n729);
and (n728,n409,n34);
and (n729,n410,n36);
nand (n730,n731,n735);
or (n731,n732,n13);
nor (n732,n733,n734);
and (n733,n470,n23);
and (n734,n24,n472);
or (n735,n662,n14);
and (n736,n716,n724);
and (n737,n691,n692);
and (n738,n686,n687);
xor (n739,n592,n624);
and (n740,n682,n683);
xor (n741,n588,n676);
or (n742,n743,n813);
or (n743,n744,n812);
and (n744,n745,n809);
xor (n745,n746,n790);
xor (n746,n747,n771);
xor (n747,n748,n751);
or (n748,n749,n750);
and (n749,n334,n350);
and (n750,n335,n344);
xor (n751,n752,n765);
xor (n752,n753,n759);
nand (n753,n754,n755);
or (n754,n13,n381);
or (n755,n756,n14);
nor (n756,n757,n758);
and (n757,n86,n23);
and (n758,n24,n88);
nand (n759,n760,n761);
or (n760,n142,n341);
or (n761,n143,n762);
nor (n762,n763,n764);
and (n763,n43,n53);
and (n764,n44,n55);
nand (n765,n766,n767);
or (n766,n67,n347);
or (n767,n768,n75);
nor (n768,n769,n770);
and (n769,n116,n74);
and (n770,n72,n118);
xor (n771,n772,n783);
xor (n772,n773,n777);
nand (n773,n774,n776);
or (n774,n433,n775);
not (n775,n431);
not (n776,n552);
nand (n777,n778,n779);
or (n778,n208,n366);
or (n779,n209,n780);
nor (n780,n781,n782);
and (n781,n145,n155);
and (n782,n146,n157);
nand (n783,n784,n789);
or (n784,n785,n41);
not (n785,n786);
nand (n786,n787,n788);
or (n787,n17,n30);
or (n788,n16,n28);
or (n789,n40,n375);
xor (n790,n791,n806);
xor (n791,n792,n803);
xor (n792,n793,n800);
xor (n793,n794,n546);
nand (n794,n795,n796);
or (n795,n97,n358);
or (n796,n797,n98);
nor (n797,n798,n799);
and (n798,n105,n329);
and (n799,n106,n331);
or (n800,n801,n802);
and (n801,n362,n378);
and (n802,n363,n369);
or (n803,n804,n805);
and (n804,n544,n565);
and (n805,n545,n555);
or (n806,n807,n808);
and (n807,n295,n361);
and (n808,n296,n333);
or (n809,n810,n811);
and (n810,n539,n578);
and (n811,n540,n543);
and (n812,n746,n790);
xor (n813,n814,n855);
xor (n814,n815,n834);
xor (n815,n816,n823);
xor (n816,n817,n820);
or (n817,n818,n819);
and (n818,n752,n765);
and (n819,n753,n759);
or (n820,n821,n822);
and (n821,n772,n783);
and (n822,n773,n777);
xor (n823,n824,n831);
xor (n824,n825,n828);
nand (n825,n826,n827);
or (n826,n13,n756);
or (n827,n14,n232);
nand (n828,n829,n830);
or (n829,n67,n768);
or (n830,n78,n75);
nand (n831,n832,n833);
or (n832,n208,n780);
or (n833,n209,n221);
xor (n834,n835,n852);
xor (n835,n836,n849);
xor (n836,n837,n845);
xor (n837,n838,n841);
nand (n838,n839,n840);
or (n839,n97,n797);
or (n840,n108,n98);
nand (n841,n842,n843);
or (n842,n785,n40);
nand (n843,n844,n723);
not (n844,n91);
not (n845,n846);
nand (n846,n847,n848);
or (n847,n142,n762);
or (n848,n143,n226);
or (n849,n850,n851);
and (n850,n793,n800);
and (n851,n794,n546);
or (n852,n853,n854);
and (n853,n747,n771);
and (n854,n748,n751);
or (n855,n856,n857);
and (n856,n791,n806);
and (n857,n792,n803);
or (n858,n859,n860);
xor (n859,n745,n809);
or (n860,n861,n862);
and (n861,n293,n538);
and (n862,n294,n384);
not (n863,n864);
or (n864,n865,n1363);
and (n865,n866,n929);
xor (n866,n867,n928);
or (n867,n868,n927);
and (n868,n869,n872);
xor (n869,n870,n871);
xor (n870,n626,n673);
xor (n871,n685,n688);
or (n872,n873,n926);
and (n873,n874,n877);
xor (n874,n875,n876);
xor (n875,n653,n666);
xor (n876,n629,n643);
or (n877,n878,n925);
and (n878,n879,n900);
xor (n879,n880,n886);
nand (n880,n881,n885);
or (n881,n208,n882);
nor (n882,n883,n884);
and (n883,n145,n80);
and (n884,n146,n82);
or (n885,n209,n656);
nor (n886,n887,n894);
not (n887,n888);
nand (n888,n889,n893);
or (n889,n890,n431);
nor (n890,n891,n892);
and (n891,n86,n215);
and (n892,n88,n213);
nand (n893,n433,n700);
nand (n894,n895,n24);
nand (n895,n896,n897);
or (n896,n402,n18);
nand (n897,n898,n16);
not (n898,n899);
and (n899,n402,n18);
or (n900,n901,n924);
and (n901,n902,n917);
xor (n902,n903,n910);
nand (n903,n904,n905);
or (n904,n143,n707);
nand (n905,n906,n170);
not (n906,n907);
nor (n907,n908,n909);
and (n908,n331,n44);
and (n909,n329,n43);
nand (n910,n911,n916);
or (n911,n912,n40);
not (n912,n913);
nor (n913,n914,n915);
and (n914,n16,n356);
and (n915,n354,n17);
nand (n916,n723,n719);
nand (n917,n918,n923);
or (n918,n919,n412);
not (n919,n920);
or (n920,n921,n922);
and (n921,n30,n410);
and (n922,n28,n409);
or (n923,n727,n413);
and (n924,n903,n910);
and (n925,n880,n886);
and (n926,n875,n876);
and (n927,n870,n871);
xor (n928,n681,n739);
or (n929,n930,n1362);
and (n930,n931,n965);
xor (n931,n932,n964);
or (n932,n933,n963);
and (n933,n934,n962);
xor (n934,n935,n936);
xor (n935,n690,n713);
or (n936,n937,n961);
and (n937,n938,n941);
xor (n938,n939,n940);
xor (n939,n715,n730);
xor (n940,n694,n705);
or (n941,n942,n960);
and (n942,n943,n956);
xor (n943,n944,n950);
nand (n944,n945,n949);
or (n945,n13,n946);
nor (n946,n947,n948);
and (n947,n404,n24);
and (n948,n402,n23);
or (n949,n732,n14);
nand (n950,n951,n955);
or (n951,n208,n952);
nor (n952,n953,n954);
and (n953,n145,n116);
and (n954,n146,n118);
or (n955,n209,n882);
nand (n956,n957,n959);
or (n957,n958,n887);
not (n958,n894);
or (n959,n888,n894);
and (n960,n944,n950);
and (n961,n939,n940);
xor (n962,n874,n877);
and (n963,n935,n936);
xor (n964,n869,n872);
nand (n965,n966,n1358);
or (n966,n967,n1336);
nor (n967,n968,n1335);
and (n968,n969,n1316);
or (n969,n970,n1315);
and (n970,n971,n1113);
xor (n971,n972,n1082);
or (n972,n973,n1081);
and (n973,n974,n1044);
xor (n974,n975,n1005);
xor (n975,n976,n995);
xor (n976,n977,n986);
nand (n977,n978,n982);
or (n978,n142,n979);
nor (n979,n980,n981);
and (n980,n354,n43);
and (n981,n356,n44);
or (n982,n983,n143);
nor (n983,n984,n985);
and (n984,n43,n323);
and (n985,n44,n325);
nand (n986,n987,n991);
or (n987,n40,n988);
nor (n988,n989,n990);
and (n989,n404,n17);
and (n990,n402,n16);
or (n991,n992,n41);
nor (n992,n993,n994);
and (n993,n470,n16);
and (n994,n472,n17);
nand (n995,n996,n1001);
or (n996,n412,n997);
not (n997,n998);
nor (n998,n999,n1000);
and (n999,n86,n410);
and (n1000,n88,n409);
or (n1001,n1002,n413);
nor (n1002,n1003,n1004);
and (n1003,n131,n409);
and (n1004,n133,n410);
or (n1005,n1006,n1043);
and (n1006,n1007,n1026);
xor (n1007,n1008,n1017);
nand (n1008,n1009,n1013);
or (n1009,n431,n1010);
nor (n1010,n1011,n1012);
and (n1011,n215,n110);
and (n1012,n213,n112);
or (n1013,n432,n1014);
nor (n1014,n1015,n1016);
and (n1015,n118,n213);
and (n1016,n116,n215);
nand (n1017,n1018,n1022);
or (n1018,n208,n1019);
nor (n1019,n1020,n1021);
and (n1020,n323,n145);
and (n1021,n146,n325);
or (n1022,n209,n1023);
nor (n1023,n1024,n1025);
and (n1024,n145,n329);
and (n1025,n146,n331);
and (n1026,n1027,n1033);
nor (n1027,n1028,n43);
nor (n1028,n1029,n1032);
and (n1029,n1030,n145);
not (n1030,n1031);
and (n1031,n402,n147);
and (n1032,n404,n149);
nand (n1033,n1034,n1039);
or (n1034,n1035,n412);
not (n1035,n1036);
nor (n1036,n1037,n1038);
and (n1037,n118,n409);
and (n1038,n116,n410);
or (n1039,n1040,n413);
nor (n1040,n1041,n1042);
and (n1041,n80,n409);
and (n1042,n82,n410);
and (n1043,n1008,n1017);
xor (n1044,n1045,n1066);
xor (n1045,n1046,n1052);
nand (n1046,n1047,n1048);
or (n1047,n208,n1023);
or (n1048,n209,n1049);
nor (n1049,n1050,n1051);
and (n1050,n145,n110);
and (n1051,n146,n112);
xor (n1052,n1053,n1058);
nor (n1053,n1054,n16);
nor (n1054,n1055,n1057);
and (n1055,n1056,n43);
nand (n1056,n402,n45);
and (n1057,n404,n47);
nand (n1058,n1059,n1064);
or (n1059,n432,n1060);
not (n1060,n1061);
nand (n1061,n1062,n1063);
or (n1062,n213,n82);
or (n1063,n215,n80);
nand (n1064,n1065,n775);
not (n1065,n1014);
or (n1066,n1067,n1080);
and (n1067,n1068,n1073);
xor (n1068,n1069,n1070);
nor (n1069,n41,n404);
nand (n1070,n1071,n1072);
or (n1071,n413,n997);
or (n1072,n1040,n412);
nand (n1073,n1074,n1075);
or (n1074,n143,n979);
nand (n1075,n1076,n170);
not (n1076,n1077);
or (n1077,n1078,n1079);
and (n1078,n472,n43);
and (n1079,n470,n44);
and (n1080,n1069,n1070);
and (n1081,n975,n1005);
xor (n1082,n1083,n1098);
xor (n1083,n1084,n1095);
xor (n1084,n1085,n1092);
xor (n1085,n1086,n1089);
nand (n1086,n1087,n1088);
or (n1087,n41,n912);
or (n1088,n40,n992);
nand (n1089,n1090,n1091);
or (n1090,n1002,n412);
nand (n1091,n920,n414);
nand (n1092,n1093,n1094);
or (n1093,n208,n1049);
or (n1094,n209,n952);
or (n1095,n1096,n1097);
and (n1096,n1045,n1066);
and (n1097,n1046,n1052);
xor (n1098,n1099,n1104);
xor (n1099,n1100,n1101);
and (n1100,n1053,n1058);
or (n1101,n1102,n1103);
and (n1102,n976,n995);
and (n1103,n977,n986);
xor (n1104,n1105,n1110);
xor (n1105,n1106,n1107);
nor (n1106,n14,n404);
nand (n1107,n1108,n1109);
or (n1108,n1060,n431);
or (n1109,n432,n890);
nand (n1110,n1111,n1112);
or (n1111,n142,n983);
or (n1112,n143,n907);
nand (n1113,n1114,n1311,n1314);
nand (n1114,n1115,n1169,n1304);
not (n1115,n1116);
nor (n1116,n1117,n1144);
xor (n1117,n1118,n1143);
xor (n1118,n1119,n1142);
or (n1119,n1120,n1141);
and (n1120,n1121,n1135);
xor (n1121,n1122,n1128);
nand (n1122,n1123,n1127);
or (n1123,n142,n1124);
nor (n1124,n1125,n1126);
and (n1125,n404,n44);
and (n1126,n402,n43);
or (n1127,n1077,n143);
nand (n1128,n1129,n1134);
or (n1129,n1130,n431);
not (n1130,n1131);
nor (n1131,n1132,n1133);
and (n1132,n329,n213);
and (n1133,n331,n215);
or (n1134,n432,n1010);
nand (n1135,n1136,n1140);
or (n1136,n208,n1137);
nor (n1137,n1138,n1139);
and (n1138,n354,n145);
and (n1139,n146,n356);
or (n1140,n209,n1019);
and (n1141,n1122,n1128);
xor (n1142,n1068,n1073);
xor (n1143,n1007,n1026);
or (n1144,n1145,n1168);
and (n1145,n1146,n1167);
xor (n1146,n1147,n1148);
xor (n1147,n1027,n1033);
or (n1148,n1149,n1166);
and (n1149,n1150,n1159);
xor (n1150,n1151,n1152);
and (n1151,n169,n402);
nand (n1152,n1153,n1158);
or (n1153,n412,n1154);
not (n1154,n1155);
nor (n1155,n1156,n1157);
and (n1156,n112,n409);
and (n1157,n110,n410);
nand (n1158,n1036,n414);
nand (n1159,n1160,n1165);
or (n1160,n1161,n431);
not (n1161,n1162);
nor (n1162,n1163,n1164);
and (n1163,n325,n215);
and (n1164,n323,n213);
nand (n1165,n1131,n433);
and (n1166,n1151,n1152);
xor (n1167,n1121,n1135);
and (n1168,n1147,n1148);
or (n1169,n1170,n1303);
and (n1170,n1171,n1197);
xor (n1171,n1172,n1196);
or (n1172,n1173,n1195);
and (n1173,n1174,n1194);
xor (n1174,n1175,n1181);
nand (n1175,n1176,n1180);
or (n1176,n208,n1177);
nor (n1177,n1178,n1179);
and (n1178,n145,n470);
and (n1179,n146,n472);
or (n1180,n1137,n209);
and (n1181,n1182,n1188);
and (n1182,n1183,n146);
nand (n1183,n1184,n1185);
or (n1184,n402,n212);
nand (n1185,n1186,n215);
not (n1186,n1187);
and (n1187,n402,n212);
nand (n1188,n1189,n1190);
or (n1189,n413,n1154);
or (n1190,n1191,n412);
nor (n1191,n1192,n1193);
and (n1192,n409,n329);
and (n1193,n410,n331);
xor (n1194,n1150,n1159);
and (n1195,n1175,n1181);
xor (n1196,n1146,n1167);
nand (n1197,n1198,n1302);
or (n1198,n1199,n1297);
nor (n1199,n1200,n1296);
and (n1200,n1201,n1275);
nand (n1201,n1202,n1273);
or (n1202,n1203,n1257);
not (n1203,n1204);
or (n1204,n1205,n1256);
and (n1205,n1206,n1235);
xor (n1206,n1207,n1216);
nand (n1207,n1208,n1212);
or (n1208,n431,n1209);
nor (n1209,n1210,n1211);
and (n1210,n213,n404);
and (n1211,n402,n215);
or (n1212,n432,n1213);
nor (n1213,n1214,n1215);
and (n1214,n472,n213);
and (n1215,n470,n215);
nand (n1216,n1217,n1234);
or (n1217,n1218,n1224);
not (n1218,n1219);
nand (n1219,n1220,n213);
nand (n1220,n1221,n1223);
or (n1221,n1222,n410);
and (n1222,n402,n436);
nand (n1223,n404,n435);
not (n1224,n1225);
nand (n1225,n1226,n1230);
or (n1226,n1227,n412);
or (n1227,n1228,n1229);
and (n1228,n354,n410);
and (n1229,n356,n409);
or (n1230,n1231,n413);
nor (n1231,n1232,n1233);
and (n1232,n325,n410);
and (n1233,n323,n409);
or (n1234,n1225,n1219);
or (n1235,n1236,n1255);
and (n1236,n1237,n1245);
xor (n1237,n1238,n1239);
nor (n1238,n432,n404);
nand (n1239,n1240,n1244);
or (n1240,n1241,n412);
nor (n1241,n1242,n1243);
and (n1242,n472,n410);
and (n1243,n470,n409);
or (n1244,n1227,n413);
nor (n1245,n1246,n1253);
nor (n1246,n1247,n1249);
and (n1247,n1248,n414);
not (n1248,n1241);
and (n1249,n1250,n559);
nand (n1250,n1251,n1252);
or (n1251,n404,n410);
nand (n1252,n410,n404);
or (n1253,n1254,n409);
and (n1254,n402,n414);
and (n1255,n1238,n1239);
and (n1256,n1207,n1216);
not (n1257,n1258);
nand (n1258,n1259,n1272);
not (n1259,n1260);
xor (n1260,n1261,n1269);
xor (n1261,n1262,n1263);
and (n1262,n219,n402);
nand (n1263,n1264,n1265);
or (n1264,n1213,n431);
nand (n1265,n1266,n433);
nor (n1266,n1267,n1268);
and (n1267,n356,n215);
and (n1268,n354,n213);
nand (n1269,n1270,n1271);
or (n1270,n1231,n412);
or (n1271,n1191,n413);
nand (n1272,n1218,n1225);
nand (n1273,n1274,n1260);
not (n1274,n1272);
nand (n1275,n1276,n1292);
not (n1276,n1277);
xor (n1277,n1278,n1291);
xor (n1278,n1279,n1283);
nand (n1279,n1280,n1282);
or (n1280,n1281,n431);
not (n1281,n1266);
nand (n1282,n1162,n433);
nand (n1283,n1284,n1289);
or (n1284,n1285,n208);
not (n1285,n1286);
nand (n1286,n1287,n1288);
or (n1287,n402,n145);
or (n1288,n404,n146);
nand (n1289,n1290,n219);
not (n1290,n1177);
xor (n1291,n1182,n1188);
not (n1292,n1293);
or (n1293,n1294,n1295);
and (n1294,n1261,n1269);
and (n1295,n1262,n1263);
nor (n1296,n1276,n1292);
nor (n1297,n1298,n1299);
xor (n1298,n1174,n1194);
or (n1299,n1300,n1301);
and (n1300,n1278,n1291);
and (n1301,n1279,n1283);
nand (n1302,n1298,n1299);
and (n1303,n1172,n1196);
nand (n1304,n1305,n1309);
not (n1305,n1306);
or (n1306,n1307,n1308);
and (n1307,n1118,n1143);
and (n1308,n1119,n1142);
not (n1309,n1310);
xor (n1310,n974,n1044);
nand (n1311,n1312,n1304);
not (n1312,n1313);
nand (n1313,n1117,n1144);
nand (n1314,n1310,n1306);
and (n1315,n972,n1082);
or (n1316,n1317,n1332);
xor (n1317,n1318,n1329);
xor (n1318,n1319,n1320);
xor (n1319,n943,n956);
xor (n1320,n1321,n1328);
xor (n1321,n1322,n1325);
or (n1322,n1323,n1324);
and (n1323,n1105,n1110);
and (n1324,n1106,n1107);
or (n1325,n1326,n1327);
and (n1326,n1085,n1092);
and (n1327,n1086,n1089);
xor (n1328,n902,n917);
or (n1329,n1330,n1331);
and (n1330,n1099,n1104);
and (n1331,n1100,n1101);
or (n1332,n1333,n1334);
and (n1333,n1083,n1098);
and (n1334,n1084,n1095);
and (n1335,n1317,n1332);
nand (n1336,n1337,n1351);
not (n1337,n1338);
and (n1338,n1339,n1347);
not (n1339,n1340);
xor (n1340,n1341,n1346);
xor (n1341,n1342,n1343);
xor (n1342,n879,n900);
or (n1343,n1344,n1345);
and (n1344,n1321,n1328);
and (n1345,n1322,n1325);
xor (n1346,n938,n941);
not (n1347,n1348);
or (n1348,n1349,n1350);
and (n1349,n1318,n1329);
and (n1350,n1319,n1320);
nand (n1351,n1352,n1354);
not (n1352,n1353);
xor (n1353,n934,n962);
not (n1354,n1355);
or (n1355,n1356,n1357);
and (n1356,n1341,n1346);
and (n1357,n1342,n1343);
nor (n1358,n1359,n1361);
and (n1359,n1351,n1360);
nor (n1360,n1339,n1347);
nor (n1361,n1352,n1354);
and (n1362,n932,n964);
and (n1363,n867,n928);
nor (n1364,n1365,n1374);
and (n1365,n1366,n742);
nand (n1366,n1367,n1369);
not (n1367,n1368);
and (n1368,n859,n860);
nand (n1369,n1370,n858);
nand (n1370,n1371,n1373);
or (n1371,n291,n1372);
nand (n1372,n741,n679);
nand (n1373,n292,n586);
and (n1374,n813,n743);
nor (n1375,n1376,n1400);
nor (n1376,n1377,n1380);
or (n1377,n1378,n1379);
and (n1378,n814,n855);
and (n1379,n815,n834);
xor (n1380,n1381,n1397);
xor (n1381,n1382,n1385);
or (n1382,n1383,n1384);
and (n1383,n816,n823);
and (n1384,n817,n820);
xor (n1385,n1386,n1391);
xor (n1386,n1387,n1388);
xor (n1387,n204,n230);
or (n1388,n1389,n1390);
and (n1389,n837,n845);
and (n1390,n838,n841);
xor (n1391,n1392,n1396);
xor (n1392,n846,n1393);
or (n1393,n1394,n1395);
and (n1394,n824,n831);
and (n1395,n825,n828);
xor (n1396,n64,n95);
or (n1397,n1398,n1399);
and (n1398,n835,n852);
and (n1399,n836,n849);
nor (n1400,n1401,n1404);
or (n1401,n1402,n1403);
and (n1402,n1381,n1397);
and (n1403,n1382,n1385);
xor (n1404,n1405,n1410);
xor (n1405,n1406,n1409);
or (n1406,n1407,n1408);
and (n1407,n1392,n1396);
and (n1408,n846,n1393);
xor (n1409,n201,n238);
or (n1410,n1411,n1412);
and (n1411,n1386,n1391);
and (n1412,n1387,n1388);
nand (n1413,n1414,n1416);
or (n1414,n1415,n1400);
nand (n1415,n1377,n1380);
nand (n1416,n1401,n1404);
nor (n1417,n1418,n1419);
xor (n1418,n7,n199);
or (n1419,n1420,n1421);
and (n1420,n1405,n1410);
and (n1421,n1406,n1409);
nand (n1422,n1419,n1418);
or (n1423,n283,n3);
xor (n1424,n1425,n2631);
xor (n1425,n1426,n2749);
xor (n1426,n1427,n2626);
xor (n1427,n1428,n2742);
xor (n1428,n1429,n2620);
xor (n1429,n1430,n2730);
xor (n1430,n1431,n2614);
xor (n1431,n1432,n2713);
xor (n1432,n1433,n2608);
xor (n1433,n1434,n2691);
xor (n1434,n1435,n2602);
xor (n1435,n1436,n2664);
xor (n1436,n1437,n2596);
xor (n1437,n1438,n2632);
xor (n1438,n1439,n2590);
xor (n1439,n1440,n2587);
xor (n1440,n1441,n2586);
xor (n1441,n1442,n2535);
xor (n1442,n1443,n2534);
xor (n1443,n1444,n2477);
xor (n1444,n1445,n2476);
xor (n1445,n1446,n2413);
xor (n1446,n1447,n2412);
xor (n1447,n1448,n2343);
xor (n1448,n1449,n2342);
xor (n1449,n1450,n2268);
xor (n1450,n1451,n2267);
xor (n1451,n1452,n2189);
xor (n1452,n1453,n2188);
xor (n1453,n1454,n2101);
xor (n1454,n1455,n2100);
xor (n1455,n1456,n2009);
xor (n1456,n1457,n2008);
xor (n1457,n1458,n1912);
xor (n1458,n1459,n1911);
xor (n1459,n1460,n1479);
xor (n1460,n1461,n1478);
xor (n1461,n1462,n1477);
xor (n1462,n1463,n1476);
xor (n1463,n1464,n1475);
xor (n1464,n1465,n1474);
xor (n1465,n1466,n1473);
xor (n1466,n1467,n1472);
xor (n1467,n1468,n1471);
xor (n1468,n1469,n1470);
and (n1469,n161,n414);
and (n1470,n161,n410);
and (n1471,n1469,n1470);
and (n1472,n161,n436);
and (n1473,n1467,n1472);
and (n1474,n161,n213);
and (n1475,n1465,n1474);
and (n1476,n161,n212);
and (n1477,n1463,n1476);
and (n1478,n161,n146);
or (n1479,n1480,n1481);
and (n1480,n1461,n1478);
and (n1481,n1460,n1482);
or (n1482,n1480,n1483);
and (n1483,n1460,n1484);
or (n1484,n1480,n1485);
and (n1485,n1460,n1486);
or (n1486,n1487,n1828);
and (n1487,n1488,n1827);
xor (n1488,n1462,n1489);
or (n1489,n1490,n1745);
and (n1490,n1491,n1744);
xor (n1491,n1464,n1492);
or (n1492,n1493,n1664);
and (n1493,n1494,n1663);
xor (n1494,n1466,n1495);
or (n1495,n1496,n1581);
and (n1496,n1497,n1580);
xor (n1497,n1468,n1498);
or (n1498,n1499,n1501);
and (n1499,n1469,n1500);
and (n1500,n155,n410);
and (n1501,n1502,n1503);
xor (n1502,n1469,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
and (n1505,n155,n414);
and (n1506,n59,n410);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
and (n1511,n59,n414);
and (n1512,n53,n410);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
and (n1517,n53,n414);
and (n1518,n34,n410);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
and (n1523,n34,n414);
and (n1524,n28,n410);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
and (n1529,n28,n414);
and (n1530,n131,n410);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1536);
and (n1534,n1535,n999);
and (n1535,n131,n414);
and (n1536,n1537,n1538);
xor (n1537,n1535,n999);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
and (n1540,n86,n414);
and (n1541,n80,n410);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
or (n1544,n1545,n1547);
and (n1545,n1546,n1038);
and (n1546,n80,n414);
and (n1547,n1548,n1549);
xor (n1548,n1546,n1038);
or (n1549,n1550,n1552);
and (n1550,n1551,n1157);
and (n1551,n116,n414);
and (n1552,n1553,n1554);
xor (n1553,n1551,n1157);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
and (n1556,n110,n414);
and (n1557,n329,n410);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
and (n1562,n329,n414);
and (n1563,n323,n410);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
or (n1566,n1567,n1569);
and (n1567,n1568,n1228);
and (n1568,n323,n414);
and (n1569,n1570,n1571);
xor (n1570,n1568,n1228);
or (n1571,n1572,n1575);
and (n1572,n1573,n1574);
and (n1573,n354,n414);
and (n1574,n470,n410);
and (n1575,n1576,n1577);
xor (n1576,n1573,n1574);
and (n1577,n1578,n1579);
and (n1578,n470,n414);
and (n1579,n402,n410);
and (n1580,n155,n436);
and (n1581,n1582,n1583);
xor (n1582,n1497,n1580);
or (n1583,n1584,n1587);
and (n1584,n1585,n1586);
xor (n1585,n1502,n1503);
and (n1586,n59,n436);
and (n1587,n1588,n1589);
xor (n1588,n1585,n1586);
or (n1589,n1590,n1593);
and (n1590,n1591,n1592);
xor (n1591,n1508,n1509);
and (n1592,n53,n436);
and (n1593,n1594,n1595);
xor (n1594,n1591,n1592);
or (n1595,n1596,n1599);
and (n1596,n1597,n1598);
xor (n1597,n1514,n1515);
and (n1598,n34,n436);
and (n1599,n1600,n1601);
xor (n1600,n1597,n1598);
or (n1601,n1602,n1605);
and (n1602,n1603,n1604);
xor (n1603,n1520,n1521);
and (n1604,n28,n436);
and (n1605,n1606,n1607);
xor (n1606,n1603,n1604);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1526,n1527);
and (n1610,n131,n436);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1532,n1533);
and (n1616,n86,n436);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1537,n1538);
and (n1622,n80,n436);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1543,n1544);
and (n1628,n116,n436);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1548,n1549);
and (n1634,n110,n436);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1553,n1554);
and (n1640,n329,n436);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1559,n1560);
and (n1646,n323,n436);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1565,n1566);
and (n1652,n354,n436);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1570,n1571);
and (n1658,n470,n436);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
and (n1661,n1662,n1222);
xor (n1662,n1576,n1577);
and (n1663,n155,n213);
and (n1664,n1665,n1666);
xor (n1665,n1494,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1582,n1583);
and (n1669,n59,n213);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1588,n1589);
and (n1675,n53,n213);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1594,n1595);
and (n1681,n34,n213);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1600,n1601);
and (n1687,n28,n213);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
or (n1690,n1691,n1694);
and (n1691,n1692,n1693);
xor (n1692,n1606,n1607);
and (n1693,n131,n213);
and (n1694,n1695,n1696);
xor (n1695,n1692,n1693);
or (n1696,n1697,n1700);
and (n1697,n1698,n1699);
xor (n1698,n1612,n1613);
and (n1699,n86,n213);
and (n1700,n1701,n1702);
xor (n1701,n1698,n1699);
or (n1702,n1703,n1706);
and (n1703,n1704,n1705);
xor (n1704,n1618,n1619);
and (n1705,n80,n213);
and (n1706,n1707,n1708);
xor (n1707,n1704,n1705);
or (n1708,n1709,n1712);
and (n1709,n1710,n1711);
xor (n1710,n1624,n1625);
and (n1711,n116,n213);
and (n1712,n1713,n1714);
xor (n1713,n1710,n1711);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
xor (n1716,n1630,n1631);
and (n1717,n110,n213);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1723);
and (n1721,n1722,n1132);
xor (n1722,n1636,n1637);
and (n1723,n1724,n1725);
xor (n1724,n1722,n1132);
or (n1725,n1726,n1728);
and (n1726,n1727,n1164);
xor (n1727,n1642,n1643);
and (n1728,n1729,n1730);
xor (n1729,n1727,n1164);
or (n1730,n1731,n1733);
and (n1731,n1732,n1268);
xor (n1732,n1648,n1649);
and (n1733,n1734,n1735);
xor (n1734,n1732,n1268);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1654,n1655);
and (n1738,n470,n213);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
and (n1741,n1742,n1743);
xor (n1742,n1660,n1661);
and (n1743,n402,n213);
and (n1744,n155,n212);
and (n1745,n1746,n1747);
xor (n1746,n1491,n1744);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1665,n1666);
and (n1750,n59,n212);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1671,n1672);
and (n1756,n53,n212);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1677,n1678);
and (n1762,n34,n212);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1683,n1684);
and (n1768,n28,n212);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1689,n1690);
and (n1774,n131,n212);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1695,n1696);
and (n1780,n86,n212);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1701,n1702);
and (n1786,n80,n212);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1707,n1708);
and (n1792,n116,n212);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1713,n1714);
and (n1798,n110,n212);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1719,n1720);
and (n1804,n329,n212);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1724,n1725);
and (n1810,n323,n212);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1729,n1730);
and (n1816,n354,n212);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1734,n1735);
and (n1822,n470,n212);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
and (n1825,n1826,n1187);
xor (n1826,n1740,n1741);
and (n1827,n155,n146);
and (n1828,n1829,n1830);
xor (n1829,n1488,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1746,n1747);
and (n1833,n59,n146);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1752,n1753);
and (n1839,n53,n146);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1758,n1759);
and (n1845,n34,n146);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1764,n1765);
and (n1851,n28,n146);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1770,n1771);
and (n1857,n131,n146);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1776,n1777);
and (n1863,n86,n146);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1782,n1783);
and (n1869,n80,n146);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1788,n1789);
and (n1875,n116,n146);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1794,n1795);
and (n1881,n110,n146);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1800,n1801);
and (n1887,n329,n146);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1806,n1807);
and (n1893,n323,n146);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1812,n1813);
and (n1899,n354,n146);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1818,n1819);
and (n1905,n470,n146);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
and (n1908,n1909,n1910);
xor (n1909,n1824,n1825);
and (n1910,n402,n146);
and (n1911,n161,n147);
or (n1912,n1913,n1915);
and (n1913,n1914,n1911);
xor (n1914,n1460,n1482);
and (n1915,n1916,n1917);
xor (n1916,n1914,n1911);
or (n1917,n1918,n1920);
and (n1918,n1919,n1911);
xor (n1919,n1460,n1484);
and (n1920,n1921,n1922);
xor (n1921,n1919,n1911);
or (n1922,n1923,n1926);
and (n1923,n1924,n1925);
xor (n1924,n1460,n1486);
and (n1925,n155,n147);
and (n1926,n1927,n1928);
xor (n1927,n1924,n1925);
or (n1928,n1929,n1932);
and (n1929,n1930,n1931);
xor (n1930,n1829,n1830);
and (n1931,n59,n147);
and (n1932,n1933,n1934);
xor (n1933,n1930,n1931);
or (n1934,n1935,n1938);
and (n1935,n1936,n1937);
xor (n1936,n1835,n1836);
and (n1937,n53,n147);
and (n1938,n1939,n1940);
xor (n1939,n1936,n1937);
or (n1940,n1941,n1944);
and (n1941,n1942,n1943);
xor (n1942,n1841,n1842);
and (n1943,n34,n147);
and (n1944,n1945,n1946);
xor (n1945,n1942,n1943);
or (n1946,n1947,n1950);
and (n1947,n1948,n1949);
xor (n1948,n1847,n1848);
and (n1949,n28,n147);
and (n1950,n1951,n1952);
xor (n1951,n1948,n1949);
or (n1952,n1953,n1956);
and (n1953,n1954,n1955);
xor (n1954,n1853,n1854);
and (n1955,n131,n147);
and (n1956,n1957,n1958);
xor (n1957,n1954,n1955);
or (n1958,n1959,n1962);
and (n1959,n1960,n1961);
xor (n1960,n1859,n1860);
and (n1961,n86,n147);
and (n1962,n1963,n1964);
xor (n1963,n1960,n1961);
or (n1964,n1965,n1968);
and (n1965,n1966,n1967);
xor (n1966,n1865,n1866);
and (n1967,n80,n147);
and (n1968,n1969,n1970);
xor (n1969,n1966,n1967);
or (n1970,n1971,n1974);
and (n1971,n1972,n1973);
xor (n1972,n1871,n1872);
and (n1973,n116,n147);
and (n1974,n1975,n1976);
xor (n1975,n1972,n1973);
or (n1976,n1977,n1980);
and (n1977,n1978,n1979);
xor (n1978,n1877,n1878);
and (n1979,n110,n147);
and (n1980,n1981,n1982);
xor (n1981,n1978,n1979);
or (n1982,n1983,n1986);
and (n1983,n1984,n1985);
xor (n1984,n1883,n1884);
and (n1985,n329,n147);
and (n1986,n1987,n1988);
xor (n1987,n1984,n1985);
or (n1988,n1989,n1992);
and (n1989,n1990,n1991);
xor (n1990,n1889,n1890);
and (n1991,n323,n147);
and (n1992,n1993,n1994);
xor (n1993,n1990,n1991);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1895,n1896);
and (n1997,n354,n147);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
or (n2000,n2001,n2004);
and (n2001,n2002,n2003);
xor (n2002,n1901,n1902);
and (n2003,n470,n147);
and (n2004,n2005,n2006);
xor (n2005,n2002,n2003);
and (n2006,n2007,n1031);
xor (n2007,n1907,n1908);
and (n2008,n161,n44);
or (n2009,n2010,n2012);
and (n2010,n2011,n2008);
xor (n2011,n1916,n1917);
and (n2012,n2013,n2014);
xor (n2013,n2011,n2008);
or (n2014,n2015,n2018);
and (n2015,n2016,n2017);
xor (n2016,n1921,n1922);
and (n2017,n155,n44);
and (n2018,n2019,n2020);
xor (n2019,n2016,n2017);
or (n2020,n2021,n2024);
and (n2021,n2022,n2023);
xor (n2022,n1927,n1928);
and (n2023,n59,n44);
and (n2024,n2025,n2026);
xor (n2025,n2022,n2023);
or (n2026,n2027,n2030);
and (n2027,n2028,n2029);
xor (n2028,n1933,n1934);
and (n2029,n53,n44);
and (n2030,n2031,n2032);
xor (n2031,n2028,n2029);
or (n2032,n2033,n2036);
and (n2033,n2034,n2035);
xor (n2034,n1939,n1940);
and (n2035,n34,n44);
and (n2036,n2037,n2038);
xor (n2037,n2034,n2035);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
xor (n2040,n1945,n1946);
and (n2041,n28,n44);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
or (n2044,n2045,n2048);
and (n2045,n2046,n2047);
xor (n2046,n1951,n1952);
and (n2047,n131,n44);
and (n2048,n2049,n2050);
xor (n2049,n2046,n2047);
or (n2050,n2051,n2054);
and (n2051,n2052,n2053);
xor (n2052,n1957,n1958);
and (n2053,n86,n44);
and (n2054,n2055,n2056);
xor (n2055,n2052,n2053);
or (n2056,n2057,n2060);
and (n2057,n2058,n2059);
xor (n2058,n1963,n1964);
and (n2059,n80,n44);
and (n2060,n2061,n2062);
xor (n2061,n2058,n2059);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
xor (n2064,n1969,n1970);
and (n2065,n116,n44);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n1975,n1976);
and (n2071,n110,n44);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2078);
and (n2075,n2076,n2077);
xor (n2076,n1981,n1982);
and (n2077,n329,n44);
and (n2078,n2079,n2080);
xor (n2079,n2076,n2077);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n1987,n1988);
and (n2083,n323,n44);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n1993,n1994);
and (n2089,n354,n44);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2095);
and (n2093,n2094,n1079);
xor (n2094,n1999,n2000);
and (n2095,n2096,n2097);
xor (n2096,n2094,n1079);
and (n2097,n2098,n2099);
xor (n2098,n2005,n2006);
and (n2099,n402,n44);
and (n2100,n161,n45);
or (n2101,n2102,n2105);
and (n2102,n2103,n2104);
xor (n2103,n2013,n2014);
and (n2104,n155,n45);
and (n2105,n2106,n2107);
xor (n2106,n2103,n2104);
or (n2107,n2108,n2111);
and (n2108,n2109,n2110);
xor (n2109,n2019,n2020);
and (n2110,n59,n45);
and (n2111,n2112,n2113);
xor (n2112,n2109,n2110);
or (n2113,n2114,n2117);
and (n2114,n2115,n2116);
xor (n2115,n2025,n2026);
and (n2116,n53,n45);
and (n2117,n2118,n2119);
xor (n2118,n2115,n2116);
or (n2119,n2120,n2123);
and (n2120,n2121,n2122);
xor (n2121,n2031,n2032);
and (n2122,n34,n45);
and (n2123,n2124,n2125);
xor (n2124,n2121,n2122);
or (n2125,n2126,n2129);
and (n2126,n2127,n2128);
xor (n2127,n2037,n2038);
and (n2128,n28,n45);
and (n2129,n2130,n2131);
xor (n2130,n2127,n2128);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2043,n2044);
and (n2134,n131,n45);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2049,n2050);
and (n2140,n86,n45);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2055,n2056);
and (n2146,n80,n45);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2061,n2062);
and (n2152,n116,n45);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2067,n2068);
and (n2158,n110,n45);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2073,n2074);
and (n2164,n329,n45);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
or (n2167,n2168,n2171);
and (n2168,n2169,n2170);
xor (n2169,n2079,n2080);
and (n2170,n323,n45);
and (n2171,n2172,n2173);
xor (n2172,n2169,n2170);
or (n2173,n2174,n2177);
and (n2174,n2175,n2176);
xor (n2175,n2085,n2086);
and (n2176,n354,n45);
and (n2177,n2178,n2179);
xor (n2178,n2175,n2176);
or (n2179,n2180,n2183);
and (n2180,n2181,n2182);
xor (n2181,n2091,n2092);
and (n2182,n470,n45);
and (n2183,n2184,n2185);
xor (n2184,n2181,n2182);
and (n2185,n2186,n2187);
xor (n2186,n2096,n2097);
not (n2187,n1056);
and (n2188,n155,n17);
or (n2189,n2190,n2193);
and (n2190,n2191,n2192);
xor (n2191,n2106,n2107);
and (n2192,n59,n17);
and (n2193,n2194,n2195);
xor (n2194,n2191,n2192);
or (n2195,n2196,n2199);
and (n2196,n2197,n2198);
xor (n2197,n2112,n2113);
and (n2198,n53,n17);
and (n2199,n2200,n2201);
xor (n2200,n2197,n2198);
or (n2201,n2202,n2205);
and (n2202,n2203,n2204);
xor (n2203,n2118,n2119);
and (n2204,n34,n17);
and (n2205,n2206,n2207);
xor (n2206,n2203,n2204);
or (n2207,n2208,n2211);
and (n2208,n2209,n2210);
xor (n2209,n2124,n2125);
and (n2210,n28,n17);
and (n2211,n2212,n2213);
xor (n2212,n2209,n2210);
or (n2213,n2214,n2217);
and (n2214,n2215,n2216);
xor (n2215,n2130,n2131);
and (n2216,n131,n17);
and (n2217,n2218,n2219);
xor (n2218,n2215,n2216);
or (n2219,n2220,n2223);
and (n2220,n2221,n2222);
xor (n2221,n2136,n2137);
and (n2222,n86,n17);
and (n2223,n2224,n2225);
xor (n2224,n2221,n2222);
or (n2225,n2226,n2228);
and (n2226,n2227,n491);
xor (n2227,n2142,n2143);
and (n2228,n2229,n2230);
xor (n2229,n2227,n491);
or (n2230,n2231,n2234);
and (n2231,n2232,n2233);
xor (n2232,n2148,n2149);
and (n2233,n116,n17);
and (n2234,n2235,n2236);
xor (n2235,n2232,n2233);
or (n2236,n2237,n2240);
and (n2237,n2238,n2239);
xor (n2238,n2154,n2155);
and (n2239,n110,n17);
and (n2240,n2241,n2242);
xor (n2241,n2238,n2239);
or (n2242,n2243,n2245);
and (n2243,n2244,n648);
xor (n2244,n2160,n2161);
and (n2245,n2246,n2247);
xor (n2246,n2244,n648);
or (n2247,n2248,n2251);
and (n2248,n2249,n2250);
xor (n2249,n2166,n2167);
and (n2250,n323,n17);
and (n2251,n2252,n2253);
xor (n2252,n2249,n2250);
or (n2253,n2254,n2256);
and (n2254,n2255,n915);
xor (n2255,n2172,n2173);
and (n2256,n2257,n2258);
xor (n2257,n2255,n915);
or (n2258,n2259,n2262);
and (n2259,n2260,n2261);
xor (n2260,n2178,n2179);
and (n2261,n470,n17);
and (n2262,n2263,n2264);
xor (n2263,n2260,n2261);
and (n2264,n2265,n2266);
xor (n2265,n2184,n2185);
and (n2266,n402,n17);
and (n2267,n59,n18);
or (n2268,n2269,n2272);
and (n2269,n2270,n2271);
xor (n2270,n2194,n2195);
and (n2271,n53,n18);
and (n2272,n2273,n2274);
xor (n2273,n2270,n2271);
or (n2274,n2275,n2278);
and (n2275,n2276,n2277);
xor (n2276,n2200,n2201);
and (n2277,n34,n18);
and (n2278,n2279,n2280);
xor (n2279,n2276,n2277);
or (n2280,n2281,n2284);
and (n2281,n2282,n2283);
xor (n2282,n2206,n2207);
and (n2283,n28,n18);
and (n2284,n2285,n2286);
xor (n2285,n2282,n2283);
or (n2286,n2287,n2290);
and (n2287,n2288,n2289);
xor (n2288,n2212,n2213);
and (n2289,n131,n18);
and (n2290,n2291,n2292);
xor (n2291,n2288,n2289);
or (n2292,n2293,n2296);
and (n2293,n2294,n2295);
xor (n2294,n2218,n2219);
and (n2295,n86,n18);
and (n2296,n2297,n2298);
xor (n2297,n2294,n2295);
or (n2298,n2299,n2302);
and (n2299,n2300,n2301);
xor (n2300,n2224,n2225);
and (n2301,n80,n18);
and (n2302,n2303,n2304);
xor (n2303,n2300,n2301);
or (n2304,n2305,n2308);
and (n2305,n2306,n2307);
xor (n2306,n2229,n2230);
and (n2307,n116,n18);
and (n2308,n2309,n2310);
xor (n2309,n2306,n2307);
or (n2310,n2311,n2314);
and (n2311,n2312,n2313);
xor (n2312,n2235,n2236);
and (n2313,n110,n18);
and (n2314,n2315,n2316);
xor (n2315,n2312,n2313);
or (n2316,n2317,n2320);
and (n2317,n2318,n2319);
xor (n2318,n2241,n2242);
and (n2319,n329,n18);
and (n2320,n2321,n2322);
xor (n2321,n2318,n2319);
or (n2322,n2323,n2326);
and (n2323,n2324,n2325);
xor (n2324,n2246,n2247);
and (n2325,n323,n18);
and (n2326,n2327,n2328);
xor (n2327,n2324,n2325);
or (n2328,n2329,n2332);
and (n2329,n2330,n2331);
xor (n2330,n2252,n2253);
and (n2331,n354,n18);
and (n2332,n2333,n2334);
xor (n2333,n2330,n2331);
or (n2334,n2335,n2338);
and (n2335,n2336,n2337);
xor (n2336,n2257,n2258);
and (n2337,n470,n18);
and (n2338,n2339,n2340);
xor (n2339,n2336,n2337);
and (n2340,n2341,n899);
xor (n2341,n2263,n2264);
and (n2342,n53,n24);
or (n2343,n2344,n2347);
and (n2344,n2345,n2346);
xor (n2345,n2273,n2274);
and (n2346,n34,n24);
and (n2347,n2348,n2349);
xor (n2348,n2345,n2346);
or (n2349,n2350,n2353);
and (n2350,n2351,n2352);
xor (n2351,n2279,n2280);
and (n2352,n28,n24);
and (n2353,n2354,n2355);
xor (n2354,n2351,n2352);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2285,n2286);
and (n2358,n131,n24);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2291,n2292);
and (n2364,n86,n24);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2297,n2298);
and (n2370,n80,n24);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2303,n2304);
and (n2376,n116,n24);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2309,n2310);
and (n2382,n110,n24);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2315,n2316);
and (n2388,n329,n24);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2321,n2322);
and (n2394,n323,n24);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2327,n2328);
and (n2400,n354,n24);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
or (n2403,n2404,n2407);
and (n2404,n2405,n2406);
xor (n2405,n2333,n2334);
and (n2406,n470,n24);
and (n2407,n2408,n2409);
xor (n2408,n2405,n2406);
and (n2409,n2410,n2411);
xor (n2410,n2339,n2340);
and (n2411,n402,n24);
and (n2412,n34,n71);
or (n2413,n2414,n2417);
and (n2414,n2415,n2416);
xor (n2415,n2348,n2349);
and (n2416,n28,n71);
and (n2417,n2418,n2419);
xor (n2418,n2415,n2416);
or (n2419,n2420,n2423);
and (n2420,n2421,n2422);
xor (n2421,n2354,n2355);
and (n2422,n131,n71);
and (n2423,n2424,n2425);
xor (n2424,n2421,n2422);
or (n2425,n2426,n2429);
and (n2426,n2427,n2428);
xor (n2427,n2360,n2361);
and (n2428,n86,n71);
and (n2429,n2430,n2431);
xor (n2430,n2427,n2428);
or (n2431,n2432,n2435);
and (n2432,n2433,n2434);
xor (n2433,n2366,n2367);
and (n2434,n80,n71);
and (n2435,n2436,n2437);
xor (n2436,n2433,n2434);
or (n2437,n2438,n2441);
and (n2438,n2439,n2440);
xor (n2439,n2372,n2373);
and (n2440,n116,n71);
and (n2441,n2442,n2443);
xor (n2442,n2439,n2440);
or (n2443,n2444,n2447);
and (n2444,n2445,n2446);
xor (n2445,n2378,n2379);
and (n2446,n110,n71);
and (n2447,n2448,n2449);
xor (n2448,n2445,n2446);
or (n2449,n2450,n2453);
and (n2450,n2451,n2452);
xor (n2451,n2384,n2385);
and (n2452,n329,n71);
and (n2453,n2454,n2455);
xor (n2454,n2451,n2452);
or (n2455,n2456,n2459);
and (n2456,n2457,n2458);
xor (n2457,n2390,n2391);
and (n2458,n323,n71);
and (n2459,n2460,n2461);
xor (n2460,n2457,n2458);
or (n2461,n2462,n2465);
and (n2462,n2463,n2464);
xor (n2463,n2396,n2397);
and (n2464,n354,n71);
and (n2465,n2466,n2467);
xor (n2466,n2463,n2464);
or (n2467,n2468,n2471);
and (n2468,n2469,n2470);
xor (n2469,n2402,n2403);
and (n2470,n470,n71);
and (n2471,n2472,n2473);
xor (n2472,n2469,n2470);
and (n2473,n2474,n2475);
xor (n2474,n2408,n2409);
not (n2475,n614);
and (n2476,n28,n72);
or (n2477,n2478,n2481);
and (n2478,n2479,n2480);
xor (n2479,n2418,n2419);
and (n2480,n131,n72);
and (n2481,n2482,n2483);
xor (n2482,n2479,n2480);
or (n2483,n2484,n2487);
and (n2484,n2485,n2486);
xor (n2485,n2424,n2425);
and (n2486,n86,n72);
and (n2487,n2488,n2489);
xor (n2488,n2485,n2486);
or (n2489,n2490,n2493);
and (n2490,n2491,n2492);
xor (n2491,n2430,n2431);
and (n2492,n80,n72);
and (n2493,n2494,n2495);
xor (n2494,n2491,n2492);
or (n2495,n2496,n2499);
and (n2496,n2497,n2498);
xor (n2497,n2436,n2437);
and (n2498,n116,n72);
and (n2499,n2500,n2501);
xor (n2500,n2497,n2498);
or (n2501,n2502,n2505);
and (n2502,n2503,n2504);
xor (n2503,n2442,n2443);
and (n2504,n110,n72);
and (n2505,n2506,n2507);
xor (n2506,n2503,n2504);
or (n2507,n2508,n2511);
and (n2508,n2509,n2510);
xor (n2509,n2448,n2449);
and (n2510,n329,n72);
and (n2511,n2512,n2513);
xor (n2512,n2509,n2510);
or (n2513,n2514,n2517);
and (n2514,n2515,n2516);
xor (n2515,n2454,n2455);
and (n2516,n323,n72);
and (n2517,n2518,n2519);
xor (n2518,n2515,n2516);
or (n2519,n2520,n2523);
and (n2520,n2521,n2522);
xor (n2521,n2460,n2461);
and (n2522,n354,n72);
and (n2523,n2524,n2525);
xor (n2524,n2521,n2522);
or (n2525,n2526,n2529);
and (n2526,n2527,n2528);
xor (n2527,n2466,n2467);
and (n2528,n470,n72);
and (n2529,n2530,n2531);
xor (n2530,n2527,n2528);
and (n2531,n2532,n2533);
xor (n2532,n2472,n2473);
and (n2533,n402,n72);
and (n2534,n131,n100);
or (n2535,n2536,n2539);
and (n2536,n2537,n2538);
xor (n2537,n2482,n2483);
and (n2538,n86,n100);
and (n2539,n2540,n2541);
xor (n2540,n2537,n2538);
or (n2541,n2542,n2545);
and (n2542,n2543,n2544);
xor (n2543,n2488,n2489);
and (n2544,n80,n100);
and (n2545,n2546,n2547);
xor (n2546,n2543,n2544);
or (n2547,n2548,n2551);
and (n2548,n2549,n2550);
xor (n2549,n2494,n2495);
and (n2550,n116,n100);
and (n2551,n2552,n2553);
xor (n2552,n2549,n2550);
or (n2553,n2554,n2557);
and (n2554,n2555,n2556);
xor (n2555,n2500,n2501);
and (n2556,n110,n100);
and (n2557,n2558,n2559);
xor (n2558,n2555,n2556);
or (n2559,n2560,n2563);
and (n2560,n2561,n2562);
xor (n2561,n2506,n2507);
and (n2562,n329,n100);
and (n2563,n2564,n2565);
xor (n2564,n2561,n2562);
or (n2565,n2566,n2569);
and (n2566,n2567,n2568);
xor (n2567,n2512,n2513);
and (n2568,n323,n100);
and (n2569,n2570,n2571);
xor (n2570,n2567,n2568);
or (n2571,n2572,n2575);
and (n2572,n2573,n2574);
xor (n2573,n2518,n2519);
and (n2574,n354,n100);
and (n2575,n2576,n2577);
xor (n2576,n2573,n2574);
or (n2577,n2578,n2581);
and (n2578,n2579,n2580);
xor (n2579,n2524,n2525);
and (n2580,n470,n100);
and (n2581,n2582,n2583);
xor (n2582,n2579,n2580);
and (n2583,n2584,n2585);
xor (n2584,n2530,n2531);
not (n2585,n401);
and (n2586,n86,n106);
or (n2587,n2588,n2591);
and (n2588,n2589,n2590);
xor (n2589,n2540,n2541);
and (n2590,n80,n106);
and (n2591,n2592,n2593);
xor (n2592,n2589,n2590);
or (n2593,n2594,n2597);
and (n2594,n2595,n2596);
xor (n2595,n2546,n2547);
and (n2596,n116,n106);
and (n2597,n2598,n2599);
xor (n2598,n2595,n2596);
or (n2599,n2600,n2603);
and (n2600,n2601,n2602);
xor (n2601,n2552,n2553);
and (n2602,n110,n106);
and (n2603,n2604,n2605);
xor (n2604,n2601,n2602);
or (n2605,n2606,n2609);
and (n2606,n2607,n2608);
xor (n2607,n2558,n2559);
and (n2608,n329,n106);
and (n2609,n2610,n2611);
xor (n2610,n2607,n2608);
or (n2611,n2612,n2615);
and (n2612,n2613,n2614);
xor (n2613,n2564,n2565);
and (n2614,n323,n106);
and (n2615,n2616,n2617);
xor (n2616,n2613,n2614);
or (n2617,n2618,n2621);
and (n2618,n2619,n2620);
xor (n2619,n2570,n2571);
and (n2620,n354,n106);
and (n2621,n2622,n2623);
xor (n2622,n2619,n2620);
or (n2623,n2624,n2627);
and (n2624,n2625,n2626);
xor (n2625,n2576,n2577);
and (n2626,n470,n106);
and (n2627,n2628,n2629);
xor (n2628,n2625,n2626);
and (n2629,n2630,n2631);
xor (n2630,n2582,n2583);
and (n2631,n402,n106);
or (n2632,n2633,n2635);
and (n2633,n2634,n2596);
xor (n2634,n2592,n2593);
and (n2635,n2636,n2637);
xor (n2636,n2634,n2596);
or (n2637,n2638,n2640);
and (n2638,n2639,n2602);
xor (n2639,n2598,n2599);
and (n2640,n2641,n2642);
xor (n2641,n2639,n2602);
or (n2642,n2643,n2645);
and (n2643,n2644,n2608);
xor (n2644,n2604,n2605);
and (n2645,n2646,n2647);
xor (n2646,n2644,n2608);
or (n2647,n2648,n2650);
and (n2648,n2649,n2614);
xor (n2649,n2610,n2611);
and (n2650,n2651,n2652);
xor (n2651,n2649,n2614);
or (n2652,n2653,n2655);
and (n2653,n2654,n2620);
xor (n2654,n2616,n2617);
and (n2655,n2656,n2657);
xor (n2656,n2654,n2620);
or (n2657,n2658,n2660);
and (n2658,n2659,n2626);
xor (n2659,n2622,n2623);
and (n2660,n2661,n2662);
xor (n2661,n2659,n2626);
and (n2662,n2663,n2631);
xor (n2663,n2628,n2629);
or (n2664,n2665,n2667);
and (n2665,n2666,n2602);
xor (n2666,n2636,n2637);
and (n2667,n2668,n2669);
xor (n2668,n2666,n2602);
or (n2669,n2670,n2672);
and (n2670,n2671,n2608);
xor (n2671,n2641,n2642);
and (n2672,n2673,n2674);
xor (n2673,n2671,n2608);
or (n2674,n2675,n2677);
and (n2675,n2676,n2614);
xor (n2676,n2646,n2647);
and (n2677,n2678,n2679);
xor (n2678,n2676,n2614);
or (n2679,n2680,n2682);
and (n2680,n2681,n2620);
xor (n2681,n2651,n2652);
and (n2682,n2683,n2684);
xor (n2683,n2681,n2620);
or (n2684,n2685,n2687);
and (n2685,n2686,n2626);
xor (n2686,n2656,n2657);
and (n2687,n2688,n2689);
xor (n2688,n2686,n2626);
and (n2689,n2690,n2631);
xor (n2690,n2661,n2662);
or (n2691,n2692,n2694);
and (n2692,n2693,n2608);
xor (n2693,n2668,n2669);
and (n2694,n2695,n2696);
xor (n2695,n2693,n2608);
or (n2696,n2697,n2699);
and (n2697,n2698,n2614);
xor (n2698,n2673,n2674);
and (n2699,n2700,n2701);
xor (n2700,n2698,n2614);
or (n2701,n2702,n2704);
and (n2702,n2703,n2620);
xor (n2703,n2678,n2679);
and (n2704,n2705,n2706);
xor (n2705,n2703,n2620);
or (n2706,n2707,n2709);
and (n2707,n2708,n2626);
xor (n2708,n2683,n2684);
and (n2709,n2710,n2711);
xor (n2710,n2708,n2626);
and (n2711,n2712,n2631);
xor (n2712,n2688,n2689);
or (n2713,n2714,n2716);
and (n2714,n2715,n2614);
xor (n2715,n2695,n2696);
and (n2716,n2717,n2718);
xor (n2717,n2715,n2614);
or (n2718,n2719,n2721);
and (n2719,n2720,n2620);
xor (n2720,n2700,n2701);
and (n2721,n2722,n2723);
xor (n2722,n2720,n2620);
or (n2723,n2724,n2726);
and (n2724,n2725,n2626);
xor (n2725,n2705,n2706);
and (n2726,n2727,n2728);
xor (n2727,n2725,n2626);
and (n2728,n2729,n2631);
xor (n2729,n2710,n2711);
or (n2730,n2731,n2733);
and (n2731,n2732,n2620);
xor (n2732,n2717,n2718);
and (n2733,n2734,n2735);
xor (n2734,n2732,n2620);
or (n2735,n2736,n2738);
and (n2736,n2737,n2626);
xor (n2737,n2722,n2723);
and (n2738,n2739,n2740);
xor (n2739,n2737,n2626);
and (n2740,n2741,n2631);
xor (n2741,n2727,n2728);
or (n2742,n2743,n2745);
and (n2743,n2744,n2626);
xor (n2744,n2734,n2735);
and (n2745,n2746,n2747);
xor (n2746,n2744,n2626);
and (n2747,n2748,n2631);
xor (n2748,n2739,n2740);
and (n2749,n2750,n2631);
xor (n2750,n2746,n2747);
endmodule
