module top (out,n17,n19,n22,n24,n28,n30,n35,n37,n40
        ,n42,n57,n63,n119,n148,n206,n323,n326,n330,n335
        ,n338,n356,n436,n492);
output out;
input n17;
input n19;
input n22;
input n24;
input n28;
input n30;
input n35;
input n37;
input n40;
input n42;
input n57;
input n63;
input n119;
input n148;
input n206;
input n323;
input n326;
input n330;
input n335;
input n338;
input n356;
input n436;
input n492;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n20;
wire n21;
wire n23;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n38;
wire n39;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n327;
wire n328;
wire n329;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
xor (out,n0,n697);
buf (n0,n1);
xor (n1,n2,n595);
xor (n2,n3,n309);
buf (n3,n4);
buf (n4,n5);
xor (n5,n6,n136);
xor (n6,n7,n95);
xor (n7,n8,n78);
xor (n8,n9,n75);
or (n9,n10,n65,n74);
and (n10,n11,n50);
or (n11,n12,n43,n49);
and (n12,n13,n32);
or (n13,n14,n25,n31);
and (n14,n15,n20);
and (n15,n16,n18);
buf (n16,n17);
buf (n18,n19);
and (n20,n21,n23);
buf (n21,n22);
buf (n23,n24);
and (n25,n20,n26);
and (n26,n27,n29);
buf (n27,n28);
buf (n29,n30);
and (n31,n15,n26);
and (n32,n33,n38);
and (n33,n34,n36);
buf (n34,n35);
buf (n36,n37);
and (n38,n39,n41);
buf (n39,n40);
buf (n41,n42);
and (n43,n32,n44);
xor (n44,n45,n48);
xor (n45,n46,n47);
and (n46,n16,n41);
and (n47,n21,n18);
and (n48,n27,n23);
and (n49,n13,n44);
xor (n50,n51,n59);
xor (n51,n52,n58);
nor (n52,n53,n54);
not (n53,n39);
and (n54,n55,n39);
not (n55,n56);
buf (n56,n57);
and (n58,n16,n36);
nor (n59,n60,n64);
and (n60,n61,n23);
not (n61,n62);
buf (n62,n63);
not (n64,n23);
and (n65,n50,n66);
xor (n66,n67,n73);
xor (n67,n68,n72);
or (n68,n69,n70,n71);
and (n69,n46,n47);
and (n70,n47,n48);
and (n71,n46,n48);
and (n72,n21,n41);
and (n73,n27,n18);
and (n74,n11,n66);
nor (n75,n76,n77);
and (n76,n61,n18);
not (n77,n18);
xor (n78,n79,n88);
xor (n79,n80,n84);
or (n80,n81,n82,n83);
and (n81,n52,n58);
and (n82,n58,n59);
and (n83,n52,n59);
or (n84,n85,n86,n87);
and (n85,n68,n72);
and (n86,n72,n73);
and (n87,n68,n73);
xor (n88,n89,n94);
xor (n89,n90,n93);
nor (n90,n91,n92);
not (n91,n16);
and (n92,n55,n16);
and (n93,n21,n36);
and (n94,n27,n41);
or (n95,n96,n132,n135);
and (n96,n97,n108);
or (n97,n98,n103,n107);
and (n98,n99,n102);
nor (n99,n100,n101);
not (n100,n34);
and (n101,n55,n34);
and (n102,n39,n36);
and (n103,n102,n104);
nor (n104,n105,n106);
and (n105,n61,n29);
not (n106,n29);
and (n107,n99,n104);
or (n108,n109,n128,n131);
and (n109,n110,n126);
or (n110,n111,n123,n125);
and (n111,n112,n121);
or (n112,n113,n116,n120);
and (n113,n114,n115);
and (n114,n16,n23);
and (n115,n21,n29);
and (n116,n115,n117);
and (n117,n27,n118);
buf (n118,n119);
and (n120,n114,n117);
xor (n121,n122,n26);
xor (n122,n15,n20);
and (n123,n121,n124);
xor (n124,n33,n38);
and (n125,n112,n124);
xor (n126,n127,n104);
xor (n127,n99,n102);
and (n128,n126,n129);
xor (n129,n130,n44);
xor (n130,n13,n32);
and (n131,n110,n129);
and (n132,n108,n133);
xor (n133,n134,n66);
xor (n134,n11,n50);
and (n135,n97,n133);
or (n136,n137,n186);
and (n137,n138,n140);
xor (n138,n139,n133);
xor (n139,n97,n108);
or (n140,n141,n182,n185);
and (n141,n142,n161);
or (n142,n143,n156,n160);
and (n143,n144,n153);
or (n144,n145,n150,n152);
and (n145,n146,n149);
and (n146,n147,n36);
buf (n147,n148);
and (n149,n34,n41);
and (n150,n149,n151);
and (n151,n39,n18);
and (n152,n146,n151);
nor (n153,n154,n155);
not (n154,n147);
and (n155,n55,n147);
and (n156,n153,n157);
nor (n157,n158,n159);
and (n158,n61,n118);
not (n159,n118);
and (n160,n144,n157);
or (n161,n162,n178,n181);
and (n162,n163,n176);
or (n163,n164,n172,n175);
and (n164,n165,n170);
or (n165,n166,1'b0,1'b0);
and (n166,n167,n168);
and (n167,n16,n29);
and (n168,n21,n118);
xor (n170,n171,n151);
xor (n171,n146,n149);
and (n172,n170,n173);
xor (n173,n174,n117);
xor (n174,n114,n115);
and (n175,n165,n173);
xor (n176,n177,n157);
xor (n177,n144,n153);
and (n178,n176,n179);
xor (n179,n180,n124);
xor (n180,n112,n121);
and (n181,n163,n179);
and (n182,n161,n183);
xor (n183,n184,n129);
xor (n184,n110,n126);
and (n185,n142,n183);
and (n186,n187,n188);
xor (n187,n138,n140);
or (n188,n189,n211);
and (n189,n190,n192);
xor (n190,n191,n183);
xor (n191,n142,n161);
or (n192,1'b0,n193,1'b0);
and (n193,n194,n209);
or (n194,n195,n202,n208);
and (n195,n196,n200);
or (n196,1'b0,n197,1'b0);
and (n197,n198,n199);
and (n198,n39,n23);
xor (n199,n167,n168);
xor (n200,n201,n173);
xor (n201,n165,n170);
and (n202,n200,n203);
nor (n203,n204,n207);
not (n204,n205);
buf (n205,n206);
and (n207,n55,n205);
and (n208,n196,n203);
xor (n209,n210,n179);
xor (n210,n163,n176);
and (n211,n212,n213);
xor (n212,n190,n192);
or (n213,n214,n246);
and (n214,n215,n216);
xor (n215,n194,n209);
or (n216,n217,n242,n245);
and (n217,n218,n225);
or (n218,n219,n222,n224);
and (n219,n220,n221);
and (n220,n205,n36);
and (n221,n147,n41);
and (n222,n221,n223);
and (n223,n34,n18);
and (n224,n220,n223);
or (n225,n226,n239,n241);
and (n226,n227,n237);
or (n227,n228,n234,n236);
and (n228,n229,n233);
or (n229,n230,1'b0,1'b0);
and (n230,n231,n232);
and (n231,n34,n29);
and (n232,n39,n118);
and (n233,n39,n29);
and (n234,n233,n235);
and (n235,n16,n118);
and (n236,n229,n235);
xor (n237,n238,n223);
xor (n238,n220,n221);
and (n239,n237,n240);
xor (n240,n198,n199);
and (n241,n227,n240);
and (n242,n225,n243);
xor (n243,n244,n203);
xor (n244,n196,n200);
and (n245,n218,n243);
and (n246,n247,n248);
xor (n247,n215,n216);
or (n248,n249,n278);
and (n249,n250,n252);
xor (n250,n251,n243);
xor (n251,n218,n225);
or (n252,n253,n274,n277);
and (n253,n254,n257);
and (n254,n255,n256);
and (n255,n147,n18);
and (n256,n34,n23);
or (n257,n258,n270,n273);
and (n258,n259,n269);
or (n259,n260,n266,n268);
and (n260,n261,n265);
or (n261,n262,1'b0,1'b0);
and (n262,n263,n264);
and (n263,n147,n29);
and (n264,n34,n118);
and (n265,n147,n23);
and (n266,n265,n267);
xor (n267,n231,n232);
and (n268,n261,n267);
xor (n269,n255,n256);
and (n270,n269,n271);
xor (n271,n272,n235);
xor (n272,n229,n233);
and (n273,n259,n271);
and (n274,n257,n275);
xor (n275,n276,n240);
xor (n276,n227,n237);
and (n277,n254,n275);
and (n278,n279,n280);
xor (n279,n250,n252);
or (n280,n281,n304);
and (n281,n282,n284);
xor (n282,n283,n275);
xor (n283,n254,n257);
and (n284,n285,n302);
or (n285,n286,n298,n301);
and (n286,n287,n297);
or (n287,n288,n294,n296);
and (n288,n289,n293);
or (n289,n290,1'b0,1'b0);
and (n290,n291,n292);
and (n291,n205,n29);
and (n292,n147,n118);
and (n293,n205,n23);
and (n294,n293,n295);
xor (n295,n263,n264);
and (n296,n289,n295);
and (n297,n205,n18);
and (n298,n297,n299);
xor (n299,n300,n267);
xor (n300,n261,n265);
and (n301,n287,n299);
xor (n302,n303,n271);
xor (n303,n259,n269);
and (n304,n305,n306);
xor (n305,n282,n284);
and (n306,n307,n308);
and (n307,n205,n41);
xor (n308,n285,n302);
buf (n309,n310);
buf (n310,n311);
xor (n311,n312,n424);
xor (n312,n313,n386);
xor (n313,n314,n369);
xor (n314,n315,n367);
or (n315,n316,n357,n366);
and (n316,n317,n346);
or (n317,n318,n339,n345);
and (n318,n319,n332);
or (n319,n320,n327,n331);
and (n320,n321,n324);
and (n321,n322,n18);
buf (n322,n323);
and (n324,n325,n23);
buf (n325,n326);
and (n327,n324,n328);
and (n328,n329,n29);
buf (n329,n330);
and (n331,n321,n328);
and (n332,n333,n336);
and (n333,n334,n36);
buf (n334,n335);
and (n336,n337,n41);
buf (n337,n338);
and (n339,n332,n340);
xor (n340,n341,n344);
xor (n341,n342,n343);
and (n342,n322,n41);
and (n343,n325,n18);
and (n344,n329,n23);
and (n345,n319,n340);
xor (n346,n347,n352);
xor (n347,n348,n351);
nor (n348,n349,n350);
not (n349,n337);
and (n350,n55,n337);
and (n351,n322,n36);
nor (n352,n353,n64);
and (n353,n354,n23);
not (n354,n355);
buf (n355,n356);
and (n357,n346,n358);
xor (n358,n359,n365);
xor (n359,n360,n364);
or (n360,n361,n362,n363);
and (n361,n342,n343);
and (n362,n343,n344);
and (n363,n342,n344);
and (n364,n325,n41);
and (n365,n329,n18);
and (n366,n317,n358);
nor (n367,n368,n77);
and (n368,n354,n18);
xor (n369,n370,n379);
xor (n370,n371,n375);
or (n371,n372,n373,n374);
and (n372,n348,n351);
and (n373,n351,n352);
and (n374,n348,n352);
or (n375,n376,n377,n378);
and (n376,n360,n364);
and (n377,n364,n365);
and (n378,n360,n365);
xor (n379,n380,n385);
xor (n380,n381,n384);
nor (n381,n382,n383);
not (n382,n322);
and (n383,n55,n322);
and (n384,n325,n36);
and (n385,n329,n41);
or (n386,n387,n420,n423);
and (n387,n388,n398);
or (n388,n389,n394,n397);
and (n389,n390,n393);
nor (n390,n391,n392);
not (n391,n334);
and (n392,n55,n334);
and (n393,n337,n36);
and (n394,n393,n395);
nor (n395,n396,n106);
and (n396,n354,n29);
and (n397,n390,n395);
or (n398,n399,n416,n419);
and (n399,n400,n414);
or (n400,n401,n411,n413);
and (n401,n402,n409);
or (n402,n403,n406,n408);
and (n403,n404,n405);
and (n404,n322,n23);
and (n405,n325,n29);
and (n406,n405,n407);
and (n407,n329,n118);
and (n408,n404,n407);
xor (n409,n410,n328);
xor (n410,n321,n324);
and (n411,n409,n412);
xor (n412,n333,n336);
and (n413,n402,n412);
xor (n414,n415,n395);
xor (n415,n390,n393);
and (n416,n414,n417);
xor (n417,n418,n340);
xor (n418,n319,n332);
and (n419,n400,n417);
and (n420,n398,n421);
xor (n421,n422,n358);
xor (n422,n317,n346);
and (n423,n388,n421);
or (n424,n425,n472);
and (n425,n426,n428);
xor (n426,n427,n421);
xor (n427,n388,n398);
or (n428,n429,n468,n471);
and (n429,n430,n448);
or (n430,n431,n444,n447);
and (n431,n432,n441);
or (n432,n433,n438,n440);
and (n433,n434,n437);
and (n434,n435,n36);
buf (n435,n436);
and (n437,n334,n41);
and (n438,n437,n439);
and (n439,n337,n18);
and (n440,n434,n439);
nor (n441,n442,n443);
not (n442,n435);
and (n443,n55,n435);
and (n444,n441,n445);
nor (n445,n446,n159);
and (n446,n354,n118);
and (n447,n432,n445);
or (n448,n449,n464,n467);
and (n449,n450,n462);
or (n450,n451,n458,n461);
and (n451,n452,n456);
or (n452,n453,1'b0,1'b0);
and (n453,n454,n455);
and (n454,n322,n29);
and (n455,n325,n118);
xor (n456,n457,n439);
xor (n457,n434,n437);
and (n458,n456,n459);
xor (n459,n460,n407);
xor (n460,n404,n405);
and (n461,n452,n459);
xor (n462,n463,n445);
xor (n463,n432,n441);
and (n464,n462,n465);
xor (n465,n466,n412);
xor (n466,n402,n409);
and (n467,n450,n465);
and (n468,n448,n469);
xor (n469,n470,n417);
xor (n470,n400,n414);
and (n471,n430,n469);
and (n472,n473,n474);
xor (n473,n426,n428);
or (n474,n475,n497);
and (n475,n476,n478);
xor (n476,n477,n469);
xor (n477,n430,n448);
or (n478,1'b0,n479,1'b0);
and (n479,n480,n495);
or (n480,n481,n488,n494);
and (n481,n482,n486);
or (n482,1'b0,n483,1'b0);
and (n483,n484,n485);
and (n484,n337,n23);
xor (n485,n454,n455);
xor (n486,n487,n459);
xor (n487,n452,n456);
and (n488,n486,n489);
nor (n489,n490,n493);
not (n490,n491);
buf (n491,n492);
and (n493,n55,n491);
and (n494,n482,n489);
xor (n495,n496,n465);
xor (n496,n450,n462);
and (n497,n498,n499);
xor (n498,n476,n478);
or (n499,n500,n532);
and (n500,n501,n502);
xor (n501,n480,n495);
or (n502,n503,n528,n531);
and (n503,n504,n511);
or (n504,n505,n508,n510);
and (n505,n506,n507);
and (n506,n491,n36);
and (n507,n435,n41);
and (n508,n507,n509);
and (n509,n334,n18);
and (n510,n506,n509);
or (n511,n512,n525,n527);
and (n512,n513,n523);
or (n513,n514,n520,n522);
and (n514,n515,n519);
or (n515,n516,1'b0,1'b0);
and (n516,n517,n518);
and (n517,n334,n29);
and (n518,n337,n118);
and (n519,n337,n29);
and (n520,n519,n521);
and (n521,n322,n118);
and (n522,n515,n521);
xor (n523,n524,n509);
xor (n524,n506,n507);
and (n525,n523,n526);
xor (n526,n484,n485);
and (n527,n513,n526);
and (n528,n511,n529);
xor (n529,n530,n489);
xor (n530,n482,n486);
and (n531,n504,n529);
and (n532,n533,n534);
xor (n533,n501,n502);
or (n534,n535,n564);
and (n535,n536,n538);
xor (n536,n537,n529);
xor (n537,n504,n511);
or (n538,n539,n560,n563);
and (n539,n540,n543);
and (n540,n541,n542);
and (n541,n435,n18);
and (n542,n334,n23);
or (n543,n544,n556,n559);
and (n544,n545,n555);
or (n545,n546,n552,n554);
and (n546,n547,n551);
or (n547,n548,1'b0,1'b0);
and (n548,n549,n550);
and (n549,n435,n29);
and (n550,n334,n118);
and (n551,n435,n23);
and (n552,n551,n553);
xor (n553,n517,n518);
and (n554,n547,n553);
xor (n555,n541,n542);
and (n556,n555,n557);
xor (n557,n558,n521);
xor (n558,n515,n519);
and (n559,n545,n557);
and (n560,n543,n561);
xor (n561,n562,n526);
xor (n562,n513,n523);
and (n563,n540,n561);
and (n564,n565,n566);
xor (n565,n536,n538);
or (n566,n567,n590);
and (n567,n568,n570);
xor (n568,n569,n561);
xor (n569,n540,n543);
and (n570,n571,n588);
or (n571,n572,n584,n587);
and (n572,n573,n583);
or (n573,n574,n580,n582);
and (n574,n575,n579);
or (n575,n576,1'b0,1'b0);
and (n576,n577,n578);
and (n577,n491,n29);
and (n578,n435,n118);
and (n579,n491,n23);
and (n580,n579,n581);
xor (n581,n549,n550);
and (n582,n575,n581);
and (n583,n491,n18);
and (n584,n583,n585);
xor (n585,n586,n553);
xor (n586,n547,n551);
and (n587,n573,n585);
xor (n588,n589,n557);
xor (n589,n545,n555);
and (n590,n591,n592);
xor (n591,n568,n570);
and (n592,n593,n594);
and (n593,n491,n41);
xor (n594,n571,n588);
or (n595,n596,n603,n696);
and (n596,n597,n600);
buf (n597,n598);
buf (n598,n599);
xor (n599,n187,n188);
buf (n600,n601);
buf (n601,n602);
xor (n602,n473,n474);
and (n603,n600,n604);
or (n604,n605,n612,n695);
and (n605,n606,n609);
buf (n606,n607);
buf (n607,n608);
xor (n608,n212,n213);
buf (n609,n610);
buf (n610,n611);
xor (n611,n498,n499);
and (n612,n609,n613);
or (n613,n614,n621,n694);
and (n614,n615,n618);
buf (n615,n616);
buf (n616,n617);
xor (n617,n247,n248);
buf (n618,n619);
buf (n619,n620);
xor (n620,n533,n534);
and (n621,n618,n622);
or (n622,n623,n630,n693);
and (n623,n624,n627);
buf (n624,n625);
buf (n625,n626);
xor (n626,n279,n280);
buf (n627,n628);
buf (n628,n629);
xor (n629,n565,n566);
and (n630,n627,n631);
or (n631,n632,n639,n692);
and (n632,n633,n636);
buf (n633,n634);
buf (n634,n635);
xor (n635,n305,n306);
buf (n636,n637);
buf (n637,n638);
xor (n638,n591,n592);
and (n639,n636,n640);
or (n640,n641,n648,n691);
and (n641,n642,n645);
buf (n642,n643);
buf (n643,n644);
xor (n644,n307,n308);
buf (n645,n646);
buf (n646,n647);
xor (n647,n593,n594);
and (n648,n645,n649);
or (n649,n650,n659,n690);
and (n650,n651,n655);
buf (n651,n652);
buf (n652,n653);
xor (n653,n654,n299);
xor (n654,n287,n297);
buf (n655,n656);
buf (n656,n657);
xor (n657,n658,n585);
xor (n658,n573,n583);
and (n659,n655,n660);
or (n660,n661,n670,n689);
and (n661,n662,n666);
buf (n662,n663);
buf (n663,n664);
xor (n664,n665,n295);
xor (n665,n289,n293);
buf (n666,n667);
buf (n667,n668);
xor (n668,n669,n581);
xor (n669,n575,n579);
and (n670,n666,n671);
or (n671,n672,n679,n688);
and (n672,n673,n676);
buf (n673,n674);
buf (n674,n675);
xor (n675,n291,n292);
buf (n676,n677);
buf (n677,n678);
xor (n678,n577,n578);
and (n679,n676,n680);
or (n680,n681,1'b0,1'b0);
and (n681,n682,n685);
buf (n682,n683);
buf (n683,n684);
and (n684,n205,n118);
buf (n685,n686);
buf (n686,n687);
and (n687,n491,n118);
and (n688,n673,n680);
and (n689,n662,n671);
and (n690,n651,n660);
and (n691,n642,n649);
and (n692,n633,n640);
and (n693,n624,n631);
and (n694,n615,n622);
and (n695,n606,n613);
and (n696,n597,n604);
buf (n697,n698);
xor (n698,n699,n856);
xor (n699,n700,n820);
xor (n700,n701,n798);
xor (n701,n702,n746);
or (n702,n703,n725,n745);
and (n703,n704,n718);
nor (n704,n705,n717);
not (n705,n706);
xor (n706,n707,n708);
xor (n707,n39,n337);
or (n708,n709,n710,n716);
and (n709,n34,n334);
and (n710,n334,n711);
or (n711,n712,n713,n715);
and (n712,n147,n435);
and (n713,n435,n714);
and (n714,n205,n491);
and (n715,n147,n714);
and (n716,n34,n711);
and (n717,n55,n706);
and (n718,n719,n36);
xor (n719,n720,n721);
xor (n720,n16,n322);
or (n721,n722,n723,n724);
and (n722,n39,n337);
and (n723,n337,n708);
and (n724,n39,n708);
and (n725,n718,n726);
nor (n726,n727,n106);
and (n727,n728,n29);
not (n728,n729);
or (n729,n730,n731,n744);
and (n730,n62,n355);
and (n731,n355,n732);
or (n732,n733,n734,n743);
and (n733,n27,n329);
and (n734,n329,n735);
or (n735,n736,n737,n742);
and (n736,n21,n325);
and (n737,n325,n738);
or (n738,n739,n740,n741);
and (n739,n16,n322);
and (n740,n322,n721);
and (n741,n16,n721);
and (n742,n21,n738);
and (n743,n27,n735);
and (n744,n62,n732);
and (n745,n704,n726);
or (n746,n747,n781,n797);
and (n747,n748,n779);
or (n748,n749,n768,n778);
and (n749,n750,n763);
or (n750,n751,n758,n762);
and (n751,n752,n755);
and (n752,n753,n23);
xor (n753,n754,n738);
xor (n754,n21,n325);
and (n755,n756,n29);
xor (n756,n757,n735);
xor (n757,n27,n329);
and (n758,n755,n759);
and (n759,n760,n118);
xor (n760,n761,n732);
xor (n761,n62,n355);
and (n762,n752,n759);
xor (n763,n764,n767);
xor (n764,n765,n766);
and (n765,n753,n18);
and (n766,n756,n23);
and (n767,n760,n29);
and (n768,n763,n769);
xor (n769,n770,n777);
xor (n770,n771,n776);
nor (n771,n772,n775);
not (n772,n773);
xor (n773,n774,n711);
xor (n774,n34,n334);
and (n775,n55,n773);
and (n776,n706,n36);
and (n777,n719,n41);
and (n778,n750,n769);
xor (n779,n780,n726);
xor (n780,n704,n718);
and (n781,n779,n782);
xor (n782,n783,n792);
xor (n783,n784,n788);
or (n784,n785,n786,n787);
and (n785,n765,n766);
and (n786,n766,n767);
and (n787,n765,n767);
or (n788,n789,n790,n791);
and (n789,n771,n776);
and (n790,n776,n777);
and (n791,n771,n777);
xor (n792,n793,n796);
xor (n793,n794,n795);
and (n794,n753,n41);
and (n795,n756,n18);
and (n796,n760,n23);
and (n797,n748,n782);
xor (n798,n799,n812);
xor (n799,n800,n804);
or (n800,n801,n802,n803);
and (n801,n784,n788);
and (n802,n788,n792);
and (n803,n784,n792);
xor (n804,n805,n810);
xor (n805,n806,n809);
nor (n806,n807,n808);
not (n807,n719);
and (n808,n55,n719);
and (n809,n753,n36);
nor (n810,n811,n64);
and (n811,n728,n23);
xor (n812,n813,n819);
xor (n813,n814,n818);
or (n814,n815,n816,n817);
and (n815,n794,n795);
and (n816,n795,n796);
and (n817,n794,n796);
and (n818,n756,n41);
and (n819,n760,n18);
or (n820,n821,n852,n855);
and (n821,n822,n832);
and (n822,n823,n830);
or (n823,n824,n827,n829);
and (n824,n825,n826);
and (n825,n773,n36);
and (n826,n706,n41);
and (n827,n826,n828);
and (n828,n719,n18);
and (n829,n825,n828);
nor (n830,n831,n159);
and (n831,n728,n118);
or (n832,n833,n849,n851);
and (n833,n834,n847);
or (n834,n835,n843,n846);
and (n835,n836,n841);
nor (n836,n837,n840);
not (n837,n838);
xor (n838,n839,n714);
xor (n839,n147,n435);
and (n840,n55,n838);
xor (n841,n842,n759);
xor (n842,n752,n755);
and (n843,n841,n844);
xor (n844,n845,n828);
xor (n845,n825,n826);
and (n846,n836,n844);
xor (n847,n848,n769);
xor (n848,n750,n763);
and (n849,n847,n850);
xor (n850,n823,n830);
and (n851,n834,n850);
and (n852,n832,n853);
xor (n853,n854,n782);
xor (n854,n748,n779);
and (n855,n822,n853);
or (n856,n857,n894);
and (n857,n858,n860);
xor (n858,n859,n853);
xor (n859,n822,n832);
or (n860,n861,n890,n893);
and (n861,n862,n873);
and (n862,n863,n870);
or (n863,n864,n867,n869);
and (n864,n865,n866);
and (n865,n773,n41);
and (n866,n706,n18);
and (n867,n866,n868);
and (n868,n719,n23);
and (n869,n865,n868);
and (n870,n871,n872);
and (n871,n753,n29);
and (n872,n756,n118);
or (n873,n874,n886,n889);
and (n874,n875,n885);
or (n875,n876,n882,n884);
and (n876,n877,n880);
and (n877,n878,n879);
and (n878,n719,n29);
and (n879,n753,n118);
xor (n880,n881,n868);
xor (n881,n865,n866);
and (n882,n880,n883);
xor (n883,n871,n872);
and (n884,n877,n883);
xor (n885,n863,n870);
and (n886,n885,n887);
xor (n887,n888,n844);
xor (n888,n836,n841);
and (n889,n875,n887);
and (n890,n873,n891);
xor (n891,n892,n850);
xor (n892,n834,n847);
and (n893,n862,n891);
and (n894,n895,n896);
xor (n895,n858,n860);
or (n896,n897,n922);
and (n897,n898,n900);
xor (n898,n899,n891);
xor (n899,n862,n873);
or (n900,n901,n918,n921);
and (n901,n902,n908);
and (n902,n903,n907);
nor (n903,n904,n906);
not (n904,n905);
xor (n905,n205,n491);
and (n906,n55,n905);
and (n907,n838,n36);
or (n908,n909,n915,n917);
and (n909,n910,n913);
and (n910,n911,n912);
and (n911,n706,n23);
xor (n912,n878,n879);
xor (n913,n914,n883);
xor (n914,n877,n880);
and (n915,n913,n916);
xor (n916,n903,n907);
and (n917,n910,n916);
and (n918,n908,n919);
xor (n919,n920,n887);
xor (n920,n875,n885);
and (n921,n902,n919);
and (n922,n923,n924);
xor (n923,n898,n900);
or (n924,n925,n957);
and (n925,n926,n928);
xor (n926,n927,n919);
xor (n927,n902,n908);
or (n928,n929,n953,n956);
and (n929,n930,n937);
or (n930,n931,n934,n936);
and (n931,n932,n933);
and (n932,n905,n36);
and (n933,n838,n41);
and (n934,n933,n935);
and (n935,n773,n18);
and (n936,n932,n935);
or (n937,n938,n950,n952);
and (n938,n939,n948);
or (n939,n940,n945,n947);
and (n940,n941,n944);
and (n941,n942,n943);
and (n942,n773,n29);
and (n943,n706,n118);
and (n944,n706,n29);
and (n945,n944,n946);
and (n946,n719,n118);
and (n947,n941,n946);
xor (n948,n949,n935);
xor (n949,n932,n933);
and (n950,n948,n951);
xor (n951,n911,n912);
and (n952,n939,n951);
and (n953,n937,n954);
xor (n954,n955,n916);
xor (n955,n910,n913);
and (n956,n930,n954);
and (n957,n958,n959);
xor (n958,n926,n928);
or (n959,n960,n988);
and (n960,n961,n963);
xor (n961,n962,n954);
xor (n962,n930,n937);
or (n963,n964,n984,n987);
and (n964,n965,n968);
and (n965,n966,n967);
and (n966,n838,n18);
and (n967,n773,n23);
or (n968,n969,n980,n983);
and (n969,n970,n979);
or (n970,n971,n976,n978);
and (n971,n972,n975);
and (n972,n973,n974);
and (n973,n838,n29);
and (n974,n773,n118);
and (n975,n838,n23);
and (n976,n975,n977);
xor (n977,n942,n943);
and (n978,n972,n977);
xor (n979,n966,n967);
and (n980,n979,n981);
xor (n981,n982,n946);
xor (n982,n941,n944);
and (n983,n970,n981);
and (n984,n968,n985);
xor (n985,n986,n951);
xor (n986,n939,n948);
and (n987,n965,n985);
and (n988,n989,n990);
xor (n989,n961,n963);
or (n990,n991,n1013);
and (n991,n992,n994);
xor (n992,n993,n985);
xor (n993,n965,n968);
and (n994,n995,n1011);
or (n995,n996,n1007,n1010);
and (n996,n997,n1006);
or (n997,n998,n1003,n1005);
and (n998,n999,n1002);
and (n999,n1000,n1001);
and (n1000,n905,n29);
and (n1001,n838,n118);
and (n1002,n905,n23);
and (n1003,n1002,n1004);
xor (n1004,n973,n974);
and (n1005,n999,n1004);
and (n1006,n905,n18);
and (n1007,n1006,n1008);
xor (n1008,n1009,n977);
xor (n1009,n972,n975);
and (n1010,n997,n1008);
xor (n1011,n1012,n981);
xor (n1012,n970,n979);
and (n1013,n1014,n1015);
xor (n1014,n992,n994);
and (n1015,n1016,n1017);
and (n1016,n905,n41);
xor (n1017,n995,n1011);
endmodule
