module top (out,n13,n15,n16,n17,n26,n27,n29,n30,n40
        ,n49,n53,n63,n64,n66,n67,n74,n80,n92,n93
        ,n95,n96,n99,n105,n117,n118,n127,n133,n163,n187
        ,n222);
output out;
input n13;
input n15;
input n16;
input n17;
input n26;
input n27;
input n29;
input n30;
input n40;
input n49;
input n53;
input n63;
input n64;
input n66;
input n67;
input n74;
input n80;
input n92;
input n93;
input n95;
input n96;
input n99;
input n105;
input n117;
input n118;
input n127;
input n133;
input n163;
input n187;
input n222;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n28;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n65;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n94;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
xor (out,n0,n491);
xnor (n0,n1,n239);
nand (n1,n2,n238);
nand (n2,n3,n196);
not (n3,n4);
xor (n4,n5,n172);
xor (n5,n6,n83);
xor (n6,n7,n55);
xor (n7,n8,n43);
nand (n8,n9,n36);
or (n9,n10,n21);
not (n10,n11);
nor (n11,n12,n18);
and (n12,n13,n14);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n17);
and (s0n14,notn14,n15);
and (s1n14,n17,n16);
and (n18,n19,n20);
not (n19,n13);
not (n20,n14);
nand (n21,n22,n33);
nor (n22,n23,n31);
and (n23,n24,n28);
not (n24,n25);
wire s0n25,s1n25,notn25;
or (n25,s0n25,s1n25);
not(notn25,n17);
and (s0n25,notn25,n26);
and (s1n25,n17,n27);
wire s0n28,s1n28,notn28;
or (n28,s0n28,s1n28);
not(notn28,n17);
and (s0n28,notn28,n29);
and (s1n28,n17,n30);
and (n31,n25,n32);
not (n32,n28);
nand (n33,n34,n35);
or (n34,n24,n14);
nand (n35,n14,n24);
nand (n36,n37,n38);
not (n37,n22);
nor (n38,n39,n41);
and (n39,n40,n14);
and (n41,n42,n20);
not (n42,n40);
nor (n43,n44,n50);
nand (n44,n14,n45);
not (n45,n46);
wire s0n46,s1n46,notn46;
or (n46,s0n46,s1n46);
not(notn46,n17);
and (s0n46,notn46,1'b0);
and (s1n46,n17,n48);
and (n48,n49,n16);
nor (n50,n51,n54);
and (n51,n46,n52);
not (n52,n53);
and (n54,n45,n53);
nand (n55,n56,n77);
or (n56,n57,n72);
nand (n57,n58,n69);
not (n58,n59);
nand (n59,n60,n68);
or (n60,n61,n65);
not (n61,n62);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n17);
and (s0n62,notn62,n63);
and (s1n62,n17,n64);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n17);
and (s0n65,notn65,n66);
and (s1n65,n17,n67);
nand (n68,n65,n61);
nand (n69,n70,n71);
or (n70,n61,n28);
nand (n71,n28,n61);
nor (n72,n73,n75);
and (n73,n32,n74);
and (n75,n28,n76);
not (n76,n74);
or (n77,n58,n78);
nor (n78,n79,n81);
and (n79,n32,n80);
and (n81,n28,n82);
not (n82,n80);
xor (n83,n84,n149);
xor (n84,n85,n136);
xor (n85,n86,n109);
nand (n86,n87,n102);
or (n87,n88,n97);
not (n88,n89);
nor (n89,n90,n94);
not (n90,n91);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n17);
and (s0n91,notn91,n92);
and (s1n91,n17,n93);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n17);
and (s0n94,notn94,n95);
and (s1n94,n17,n96);
nor (n97,n98,n100);
and (n98,n90,n99);
and (n100,n91,n101);
not (n101,n99);
or (n102,n103,n108);
nor (n103,n104,n106);
and (n104,n90,n105);
and (n106,n91,n107);
not (n107,n105);
not (n108,n94);
nand (n109,n110,n130);
or (n110,n111,n124);
not (n111,n112);
and (n112,n113,n120);
nand (n113,n114,n119);
or (n114,n115,n65);
not (n115,n116);
wire s0n116,s1n116,notn116;
or (n116,s0n116,s1n116);
not(notn116,n17);
and (s0n116,notn116,n117);
and (s1n116,n17,n118);
nand (n119,n65,n115);
not (n120,n121);
nand (n121,n122,n123);
or (n122,n115,n91);
nand (n123,n91,n115);
nor (n124,n125,n128);
and (n125,n126,n127);
not (n126,n65);
and (n128,n65,n129);
not (n129,n127);
or (n130,n120,n131);
nor (n131,n132,n134);
and (n132,n126,n133);
and (n134,n65,n135);
not (n135,n133);
and (n136,n137,n143);
nand (n137,n138,n142);
or (n138,n88,n139);
nor (n139,n140,n141);
and (n140,n90,n133);
and (n141,n91,n135);
or (n142,n97,n108);
nand (n143,n144,n148);
or (n144,n111,n145);
nor (n145,n146,n147);
and (n146,n126,n80);
and (n147,n65,n82);
or (n148,n124,n120);
or (n149,n150,n171);
and (n150,n151,n165);
xor (n151,n152,n159);
nand (n152,n153,n158);
or (n153,n154,n21);
not (n154,n155);
nor (n155,n156,n157);
and (n156,n53,n14);
and (n157,n52,n20);
nand (n158,n37,n11);
nor (n159,n44,n160);
nor (n160,n161,n164);
and (n161,n46,n162);
not (n162,n163);
and (n164,n45,n163);
nand (n165,n166,n170);
or (n166,n57,n167);
nor (n167,n168,n169);
and (n168,n32,n40);
and (n169,n28,n42);
or (n170,n58,n72);
and (n171,n152,n159);
and (n172,n173,n174);
xor (n173,n137,n143);
or (n174,n175,n195);
and (n175,n176,n189);
xor (n176,n177,n183);
nand (n177,n178,n182);
or (n178,n179,n21);
nor (n179,n180,n181);
and (n180,n163,n20);
and (n181,n162,n14);
nand (n182,n155,n37);
nor (n183,n44,n184);
nor (n184,n185,n188);
and (n185,n46,n186);
not (n186,n187);
and (n188,n45,n187);
nand (n189,n190,n194);
or (n190,n88,n191);
nor (n191,n192,n193);
and (n192,n90,n127);
and (n193,n91,n129);
or (n194,n139,n108);
and (n195,n177,n183);
not (n196,n197);
or (n197,n198,n237);
and (n198,n199,n202);
xor (n199,n200,n201);
xor (n200,n151,n165);
xor (n201,n173,n174);
or (n202,n203,n236);
and (n203,n204,n217);
xor (n204,n205,n211);
nand (n205,n206,n210);
or (n206,n57,n207);
nor (n207,n208,n209);
and (n208,n32,n13);
and (n209,n28,n19);
or (n210,n58,n167);
nand (n211,n212,n216);
or (n212,n111,n213);
nor (n213,n214,n215);
and (n214,n126,n74);
and (n215,n65,n76);
or (n216,n145,n120);
or (n217,n218,n235);
and (n218,n219,n229);
xor (n219,n220,n223);
and (n220,n221,n222);
not (n221,n44);
nand (n223,n224,n228);
or (n224,n88,n225);
nor (n225,n226,n227);
and (n226,n82,n91);
and (n227,n80,n90);
or (n228,n191,n108);
nand (n229,n230,n234);
or (n230,n21,n231);
nor (n231,n232,n233);
and (n232,n187,n20);
and (n233,n186,n14);
or (n234,n22,n179);
and (n235,n220,n223);
and (n236,n205,n211);
and (n237,n200,n201);
nand (n238,n4,n197);
nand (n239,n240,n490);
or (n240,n241,n281);
nor (n241,n242,n243);
xor (n242,n199,n202);
or (n243,n244,n280);
and (n244,n245,n279);
xor (n245,n246,n247);
xor (n246,n176,n189);
or (n247,n248,n278);
and (n248,n249,n263);
xor (n249,n250,n257);
nand (n250,n251,n256);
or (n251,n111,n252);
not (n252,n253);
nor (n253,n254,n255);
and (n254,n40,n65);
and (n255,n42,n126);
or (n256,n120,n213);
nand (n257,n258,n262);
or (n258,n57,n259);
nor (n259,n260,n261);
and (n260,n32,n53);
and (n261,n28,n52);
or (n262,n58,n207);
and (n263,n264,n270);
nor (n264,n265,n20);
nor (n265,n266,n268);
and (n266,n32,n267);
nand (n267,n25,n222);
and (n268,n24,n269);
not (n269,n222);
nand (n270,n271,n276);
or (n271,n272,n88);
not (n272,n273);
nor (n273,n274,n275);
and (n274,n74,n91);
and (n275,n76,n90);
nand (n276,n277,n94);
not (n277,n225);
and (n278,n250,n257);
xor (n279,n204,n217);
and (n280,n246,n247);
not (n281,n282);
nand (n282,n283,n485);
not (n283,n284);
nor (n284,n285,n466);
nor (n285,n286,n464);
and (n286,n287,n438);
or (n287,n288,n437);
and (n288,n289,n353);
xor (n289,n290,n330);
or (n290,n291,n329);
and (n291,n292,n314);
xor (n292,n293,n303);
nand (n293,n294,n299);
or (n294,n295,n111);
not (n295,n296);
nor (n296,n297,n298);
and (n297,n162,n126);
and (n298,n163,n65);
nand (n299,n121,n300);
nor (n300,n301,n302);
and (n301,n53,n65);
and (n302,n126,n52);
nand (n303,n304,n309);
or (n304,n305,n58);
not (n305,n306);
nor (n306,n307,n308);
and (n307,n187,n28);
and (n308,n186,n32);
nand (n309,n310,n311);
not (n310,n57);
nand (n311,n312,n313);
or (n312,n32,n222);
or (n313,n28,n269);
xor (n314,n315,n320);
and (n315,n316,n28);
nand (n316,n317,n319);
or (n317,n65,n318);
and (n318,n222,n62);
or (n319,n62,n222);
nand (n320,n321,n325);
or (n321,n88,n322);
nor (n322,n323,n324);
and (n323,n90,n13);
and (n324,n91,n19);
or (n325,n326,n108);
nor (n326,n327,n328);
and (n327,n40,n90);
and (n328,n42,n91);
and (n329,n293,n303);
xor (n330,n331,n339);
xor (n331,n332,n338);
nand (n332,n333,n334);
or (n333,n305,n57);
or (n334,n58,n335);
nor (n335,n336,n337);
and (n336,n32,n163);
and (n337,n28,n162);
and (n338,n315,n320);
xor (n339,n340,n346);
xor (n340,n341,n342);
and (n341,n37,n222);
nand (n342,n343,n344);
or (n343,n108,n272);
nand (n344,n345,n89);
not (n345,n326);
nand (n346,n347,n349);
or (n347,n348,n111);
not (n348,n300);
nand (n349,n121,n350);
nand (n350,n351,n352);
or (n351,n65,n19);
or (n352,n126,n13);
or (n353,n354,n436);
and (n354,n355,n376);
xor (n355,n356,n375);
or (n356,n357,n374);
and (n357,n358,n367);
xor (n358,n359,n360);
and (n359,n59,n222);
nand (n360,n361,n366);
or (n361,n362,n111);
not (n362,n363);
nor (n363,n364,n365);
and (n364,n187,n65);
and (n365,n186,n126);
nand (n366,n296,n121);
nand (n367,n368,n373);
or (n368,n88,n369);
not (n369,n370);
nor (n370,n371,n372);
and (n371,n52,n90);
and (n372,n53,n91);
or (n373,n322,n108);
and (n374,n359,n360);
xor (n375,n292,n314);
or (n376,n377,n435);
and (n377,n378,n434);
xor (n378,n379,n393);
nor (n379,n380,n388);
not (n380,n381);
nand (n381,n382,n387);
or (n382,n383,n88);
not (n383,n384);
nand (n384,n385,n386);
or (n385,n162,n91);
nand (n386,n91,n162);
nand (n387,n370,n94);
nand (n388,n389,n65);
nand (n389,n390,n392);
or (n390,n91,n391);
and (n391,n222,n116);
or (n392,n116,n222);
nand (n393,n394,n432);
or (n394,n395,n418);
not (n395,n396);
nand (n396,n397,n417);
or (n397,n398,n407);
nor (n398,n399,n406);
nand (n399,n400,n405);
or (n400,n401,n88);
not (n401,n402);
nand (n402,n403,n404);
or (n403,n186,n91);
nand (n404,n91,n186);
nand (n405,n384,n94);
nor (n406,n120,n269);
nand (n407,n408,n415);
nand (n408,n409,n414);
or (n409,n410,n88);
not (n410,n411);
nand (n411,n412,n413);
or (n412,n90,n222);
or (n413,n91,n269);
nand (n414,n402,n94);
nor (n415,n416,n90);
and (n416,n222,n94);
nand (n417,n399,n406);
not (n418,n419);
nand (n419,n420,n428);
not (n420,n421);
nand (n421,n422,n427);
or (n422,n423,n111);
not (n423,n424);
nand (n424,n425,n426);
or (n425,n126,n222);
or (n426,n65,n269);
nand (n427,n121,n363);
nor (n428,n429,n431);
and (n429,n380,n430);
not (n430,n388);
and (n431,n381,n388);
nand (n432,n433,n421);
not (n433,n428);
xor (n434,n358,n367);
and (n435,n379,n393);
and (n436,n356,n375);
and (n437,n290,n330);
or (n438,n439,n461);
xor (n439,n440,n445);
xor (n440,n441,n442);
xor (n441,n264,n270);
or (n442,n443,n444);
and (n443,n340,n346);
and (n444,n341,n342);
xor (n445,n446,n458);
xor (n446,n447,n454);
nand (n447,n448,n453);
or (n448,n449,n21);
not (n449,n450);
nand (n450,n451,n452);
or (n451,n20,n222);
or (n452,n14,n269);
or (n453,n22,n231);
nand (n454,n455,n457);
or (n455,n456,n111);
not (n456,n350);
nand (n457,n121,n253);
nand (n458,n459,n460);
or (n459,n57,n335);
or (n460,n58,n259);
or (n461,n462,n463);
and (n462,n331,n339);
and (n463,n332,n338);
not (n464,n465);
nand (n465,n439,n461);
nand (n466,n467,n479);
not (n467,n468);
nor (n468,n469,n476);
xor (n469,n470,n475);
xor (n470,n471,n474);
or (n471,n472,n473);
and (n472,n446,n458);
and (n473,n447,n454);
xor (n474,n219,n229);
xor (n475,n249,n263);
or (n476,n477,n478);
and (n477,n440,n445);
and (n478,n441,n442);
not (n479,n480);
nor (n480,n481,n484);
or (n481,n482,n483);
and (n482,n470,n475);
and (n483,n471,n474);
xor (n484,n245,n279);
nor (n485,n486,n489);
and (n486,n479,n487);
not (n487,n488);
nand (n488,n469,n476);
and (n489,n481,n484);
nand (n490,n242,n243);
xor (n491,n492,n797);
xor (n492,n493,n805);
xor (n493,n494,n792);
xor (n494,n495,n798);
xor (n495,n496,n786);
xor (n496,n497,n783);
xor (n497,n498,n782);
xor (n498,n499,n762);
xor (n499,n500,n12);
xor (n500,n501,n735);
xor (n501,n502,n734);
xor (n502,n503,n702);
xor (n503,n504,n701);
xor (n504,n505,n663);
xor (n505,n506,n662);
xor (n506,n507,n621);
xor (n507,n508,n620);
xor (n508,n509,n570);
xor (n509,n510,n569);
xor (n510,n511,n514);
xor (n511,n512,n513);
and (n512,n105,n94);
and (n513,n99,n91);
or (n514,n515,n518);
and (n515,n516,n517);
and (n516,n99,n94);
and (n517,n133,n91);
and (n518,n519,n520);
xor (n519,n516,n517);
or (n520,n521,n524);
and (n521,n522,n523);
and (n522,n133,n94);
and (n523,n127,n91);
and (n524,n525,n526);
xor (n525,n522,n523);
or (n526,n527,n530);
and (n527,n528,n529);
and (n528,n127,n94);
and (n529,n80,n91);
and (n530,n531,n532);
xor (n531,n528,n529);
or (n532,n533,n535);
and (n533,n534,n274);
and (n534,n80,n94);
and (n535,n536,n537);
xor (n536,n534,n274);
or (n537,n538,n541);
and (n538,n539,n540);
and (n539,n74,n94);
and (n540,n40,n91);
and (n541,n542,n543);
xor (n542,n539,n540);
or (n543,n544,n547);
and (n544,n545,n546);
and (n545,n40,n94);
and (n546,n13,n91);
and (n547,n548,n549);
xor (n548,n545,n546);
or (n549,n550,n552);
and (n550,n551,n372);
and (n551,n13,n94);
and (n552,n553,n554);
xor (n553,n551,n372);
or (n554,n555,n558);
and (n555,n556,n557);
and (n556,n53,n94);
and (n557,n163,n91);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
and (n562,n163,n94);
and (n563,n187,n91);
and (n564,n565,n566);
xor (n565,n562,n563);
and (n566,n567,n568);
and (n567,n187,n94);
and (n568,n222,n91);
and (n569,n133,n116);
or (n570,n571,n574);
and (n571,n572,n573);
xor (n572,n519,n520);
and (n573,n127,n116);
and (n574,n575,n576);
xor (n575,n572,n573);
or (n576,n577,n580);
and (n577,n578,n579);
xor (n578,n525,n526);
and (n579,n80,n116);
and (n580,n581,n582);
xor (n581,n578,n579);
or (n582,n583,n586);
and (n583,n584,n585);
xor (n584,n531,n532);
and (n585,n74,n116);
and (n586,n587,n588);
xor (n587,n584,n585);
or (n588,n589,n592);
and (n589,n590,n591);
xor (n590,n536,n537);
and (n591,n40,n116);
and (n592,n593,n594);
xor (n593,n590,n591);
or (n594,n595,n598);
and (n595,n596,n597);
xor (n596,n542,n543);
and (n597,n13,n116);
and (n598,n599,n600);
xor (n599,n596,n597);
or (n600,n601,n604);
and (n601,n602,n603);
xor (n602,n548,n549);
and (n603,n53,n116);
and (n604,n605,n606);
xor (n605,n602,n603);
or (n606,n607,n610);
and (n607,n608,n609);
xor (n608,n553,n554);
and (n609,n163,n116);
and (n610,n611,n612);
xor (n611,n608,n609);
or (n612,n613,n616);
and (n613,n614,n615);
xor (n614,n559,n560);
and (n615,n187,n116);
and (n616,n617,n618);
xor (n617,n614,n615);
and (n618,n619,n391);
xor (n619,n565,n566);
and (n620,n127,n65);
or (n621,n622,n625);
and (n622,n623,n624);
xor (n623,n575,n576);
and (n624,n80,n65);
and (n625,n626,n627);
xor (n626,n623,n624);
or (n627,n628,n631);
and (n628,n629,n630);
xor (n629,n581,n582);
and (n630,n74,n65);
and (n631,n632,n633);
xor (n632,n629,n630);
or (n633,n634,n636);
and (n634,n635,n254);
xor (n635,n587,n588);
and (n636,n637,n638);
xor (n637,n635,n254);
or (n638,n639,n642);
and (n639,n640,n641);
xor (n640,n593,n594);
and (n641,n13,n65);
and (n642,n643,n644);
xor (n643,n640,n641);
or (n644,n645,n647);
and (n645,n646,n301);
xor (n646,n599,n600);
and (n647,n648,n649);
xor (n648,n646,n301);
or (n649,n650,n652);
and (n650,n651,n298);
xor (n651,n605,n606);
and (n652,n653,n654);
xor (n653,n651,n298);
or (n654,n655,n657);
and (n655,n656,n364);
xor (n656,n611,n612);
and (n657,n658,n659);
xor (n658,n656,n364);
and (n659,n660,n661);
xor (n660,n617,n618);
and (n661,n222,n65);
and (n662,n80,n62);
or (n663,n664,n667);
and (n664,n665,n666);
xor (n665,n626,n627);
and (n666,n74,n62);
and (n667,n668,n669);
xor (n668,n665,n666);
or (n669,n670,n673);
and (n670,n671,n672);
xor (n671,n632,n633);
and (n672,n40,n62);
and (n673,n674,n675);
xor (n674,n671,n672);
or (n675,n676,n679);
and (n676,n677,n678);
xor (n677,n637,n638);
and (n678,n13,n62);
and (n679,n680,n681);
xor (n680,n677,n678);
or (n681,n682,n685);
and (n682,n683,n684);
xor (n683,n643,n644);
and (n684,n53,n62);
and (n685,n686,n687);
xor (n686,n683,n684);
or (n687,n688,n691);
and (n688,n689,n690);
xor (n689,n648,n649);
and (n690,n163,n62);
and (n691,n692,n693);
xor (n692,n689,n690);
or (n693,n694,n697);
and (n694,n695,n696);
xor (n695,n653,n654);
and (n696,n187,n62);
and (n697,n698,n699);
xor (n698,n695,n696);
and (n699,n700,n318);
xor (n700,n658,n659);
and (n701,n74,n28);
or (n702,n703,n706);
and (n703,n704,n705);
xor (n704,n668,n669);
and (n705,n40,n28);
and (n706,n707,n708);
xor (n707,n704,n705);
or (n708,n709,n712);
and (n709,n710,n711);
xor (n710,n674,n675);
and (n711,n13,n28);
and (n712,n713,n714);
xor (n713,n710,n711);
or (n714,n715,n718);
and (n715,n716,n717);
xor (n716,n680,n681);
and (n717,n53,n28);
and (n718,n719,n720);
xor (n719,n716,n717);
or (n720,n721,n724);
and (n721,n722,n723);
xor (n722,n686,n687);
and (n723,n163,n28);
and (n724,n725,n726);
xor (n725,n722,n723);
or (n726,n727,n729);
and (n727,n728,n307);
xor (n728,n692,n693);
and (n729,n730,n731);
xor (n730,n728,n307);
and (n731,n732,n733);
xor (n732,n698,n699);
and (n733,n222,n28);
and (n734,n40,n25);
or (n735,n736,n739);
and (n736,n737,n738);
xor (n737,n707,n708);
and (n738,n13,n25);
and (n739,n740,n741);
xor (n740,n737,n738);
or (n741,n742,n745);
and (n742,n743,n744);
xor (n743,n713,n714);
and (n744,n53,n25);
and (n745,n746,n747);
xor (n746,n743,n744);
or (n747,n748,n751);
and (n748,n749,n750);
xor (n749,n719,n720);
and (n750,n163,n25);
and (n751,n752,n753);
xor (n752,n749,n750);
or (n753,n754,n757);
and (n754,n755,n756);
xor (n755,n725,n726);
and (n756,n187,n25);
and (n757,n758,n759);
xor (n758,n755,n756);
and (n759,n760,n761);
xor (n760,n730,n731);
not (n761,n267);
or (n762,n763,n765);
and (n763,n764,n156);
xor (n764,n740,n741);
and (n765,n766,n767);
xor (n766,n764,n156);
or (n767,n768,n771);
and (n768,n769,n770);
xor (n769,n746,n747);
and (n770,n163,n14);
and (n771,n772,n773);
xor (n772,n769,n770);
or (n773,n774,n777);
and (n774,n775,n776);
xor (n775,n752,n753);
and (n776,n187,n14);
and (n777,n778,n779);
xor (n778,n775,n776);
and (n779,n780,n781);
xor (n780,n758,n759);
and (n781,n222,n14);
and (n782,n53,n46);
or (n783,n784,n787);
and (n784,n785,n786);
xor (n785,n766,n767);
and (n786,n163,n46);
and (n787,n788,n789);
xor (n788,n785,n786);
or (n789,n790,n793);
and (n790,n791,n792);
xor (n791,n772,n773);
and (n792,n187,n46);
and (n793,n794,n795);
xor (n794,n791,n792);
and (n795,n796,n797);
xor (n796,n778,n779);
and (n797,n222,n46);
or (n798,n799,n801);
and (n799,n800,n792);
xor (n800,n788,n789);
and (n801,n802,n803);
xor (n802,n800,n792);
and (n803,n804,n797);
xor (n804,n794,n795);
and (n805,n806,n797);
xor (n806,n802,n803);
endmodule
