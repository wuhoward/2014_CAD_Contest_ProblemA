module top (out,n16,n18,n24,n33,n38,n42,n48,n52,n53
        ,n61,n70,n76,n89,n118,n119,n184,n186,n206,n225
        ,n231,n239,n245,n287,n292,n315,n380,n442,n489,n519);
output out;
input n16;
input n18;
input n24;
input n33;
input n38;
input n42;
input n48;
input n52;
input n53;
input n61;
input n70;
input n76;
input n89;
input n118;
input n119;
input n184;
input n186;
input n206;
input n225;
input n231;
input n239;
input n245;
input n287;
input n292;
input n315;
input n380;
input n442;
input n489;
input n519;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n17;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n288;
wire n289;
wire n290;
wire n291;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
xor (out,n0,n1381);
nand (n0,n1,n1380);
or (n1,n2,n165);
not (n2,n3);
nor (n3,n4,n164);
and (n4,n5,n143);
or (n5,n6,n142);
and (n6,n7,n104);
xor (n7,n8,n54);
xor (n8,n9,n51);
xor (n9,n10,n26);
nand (n10,n11,n18);
or (n11,n12,n21);
not (n12,n13);
nand (n13,n14,n20);
nand (n14,n15,n19);
or (n15,n16,n17);
not (n17,n18);
nand (n19,n17,n16);
not (n20,n21);
nand (n21,n22,n25);
or (n22,n23,n16);
not (n23,n24);
nand (n25,n23,n16);
nand (n26,n27,n45);
or (n27,n28,n40);
not (n28,n29);
and (n29,n30,n35);
not (n30,n31);
nand (n31,n32,n34);
or (n32,n33,n17);
nand (n34,n33,n17);
nand (n35,n36,n39);
or (n36,n33,n37);
not (n37,n38);
nand (n39,n37,n33);
nor (n40,n41,n43);
and (n41,n37,n42);
and (n43,n38,n44);
not (n44,n42);
or (n45,n30,n46);
nor (n46,n47,n49);
and (n47,n37,n48);
and (n49,n38,n50);
not (n50,n48);
and (n51,n52,n53);
xor (n54,n55,n85);
xor (n55,n56,n79);
nand (n56,n57,n73);
or (n57,n58,n67);
nand (n58,n59,n64);
nor (n59,n60,n62);
and (n60,n37,n61);
and (n62,n38,n63);
not (n63,n61);
nand (n64,n65,n66);
or (n65,n63,n52);
nand (n66,n63,n52);
nor (n67,n68,n71);
and (n68,n69,n70);
not (n69,n52);
and (n71,n52,n72);
not (n72,n70);
or (n73,n59,n74);
nor (n74,n75,n77);
and (n75,n69,n76);
and (n77,n52,n78);
not (n78,n76);
nand (n79,n80,n84);
or (n80,n13,n81);
nor (n81,n82,n83);
and (n82,n17,n48);
and (n83,n18,n50);
or (n84,n20,n17);
or (n85,n86,n103);
and (n86,n87,n96);
xor (n87,n88,n90);
and (n88,n52,n89);
nand (n90,n91,n95);
or (n91,n28,n92);
nor (n92,n93,n94);
and (n93,n37,n76);
and (n94,n38,n78);
or (n95,n30,n40);
nand (n96,n97,n102);
or (n97,n58,n98);
nor (n98,n99,n100);
and (n99,n69,n53);
and (n100,n52,n101);
not (n101,n53);
or (n102,n59,n67);
and (n103,n88,n90);
or (n104,n105,n141);
and (n105,n106,n140);
xor (n106,n107,n108);
not (n107,n79);
or (n108,n109,n139);
and (n109,n110,n132);
xor (n110,n111,n126);
nand (n111,n112,n24);
or (n112,n113,n125);
not (n113,n114);
nand (n114,n115,n122);
nor (n115,n116,n120);
and (n116,n117,n119);
not (n117,n118);
and (n120,n118,n121);
not (n121,n119);
nand (n122,n123,n124);
or (n123,n119,n23);
nand (n124,n23,n119);
not (n125,n115);
nand (n126,n127,n131);
or (n127,n13,n128);
nor (n128,n129,n130);
and (n129,n17,n42);
and (n130,n18,n44);
or (n131,n20,n81);
nand (n132,n133,n138);
or (n133,n58,n134);
nor (n134,n135,n136);
and (n135,n69,n89);
and (n136,n52,n137);
not (n137,n89);
or (n138,n59,n98);
and (n139,n111,n126);
xor (n140,n87,n96);
and (n141,n107,n108);
and (n142,n8,n54);
xor (n143,n144,n161);
xor (n144,n145,n148);
or (n145,n146,n147);
and (n146,n9,n51);
and (n147,n10,n26);
xor (n148,n149,n157);
xor (n149,n150,n156);
nand (n150,n151,n152);
or (n151,n58,n74);
or (n152,n59,n153);
nor (n153,n154,n155);
and (n154,n69,n42);
and (n155,n52,n44);
and (n156,n52,n70);
nor (n157,n158,n160);
and (n158,n29,n159);
not (n159,n46);
and (n160,n31,n38);
or (n161,n162,n163);
and (n162,n55,n85);
and (n163,n56,n79);
nor (n164,n143,n5);
nand (n165,n166,n855,n1379);
nand (n166,n167,n849);
nand (n167,n168,n835);
or (n168,n169,n694);
not (n169,n170);
nand (n170,n171,n689);
or (n171,n172,n563);
not (n172,n173);
nand (n173,n174,n562);
or (n174,n175,n494);
nor (n175,n176,n425);
xor (n176,n177,n365);
xor (n177,n178,n279);
xor (n178,n179,n257);
xor (n179,n180,n216);
and (n180,n181,n196);
nand (n181,n182,n192);
or (n182,n183,n187);
nand (n183,n184,n185);
not (n185,n186);
not (n187,n188);
nor (n188,n189,n190);
and (n189,n42,n184);
and (n190,n44,n191);
not (n191,n184);
or (n192,n193,n185);
nor (n193,n194,n195);
and (n194,n191,n48);
and (n195,n184,n50);
nand (n196,n197,n212);
or (n197,n198,n202);
not (n198,n199);
nand (n199,n200,n201);
or (n200,n118,n72);
or (n201,n117,n70);
not (n202,n203);
nor (n203,n204,n208);
nand (n204,n205,n207);
or (n205,n191,n206);
nand (n207,n191,n206);
nor (n208,n209,n210);
and (n209,n117,n206);
and (n210,n118,n211);
not (n211,n206);
nand (n212,n204,n213);
nor (n213,n214,n215);
and (n214,n118,n76);
and (n215,n78,n117);
or (n216,n217,n256);
and (n217,n218,n247);
xor (n218,n219,n233);
nand (n219,n220,n227);
or (n220,n221,n13);
not (n221,n222);
nor (n222,n223,n226);
and (n223,n224,n17);
not (n224,n225);
and (n226,n225,n18);
nand (n227,n21,n228);
nor (n228,n229,n232);
and (n229,n230,n17);
not (n230,n231);
and (n232,n18,n231);
nand (n233,n234,n241);
or (n234,n235,n28);
not (n235,n236);
nor (n236,n237,n240);
and (n237,n238,n37);
not (n238,n239);
and (n240,n239,n38);
nand (n241,n31,n242);
nand (n242,n243,n246);
or (n243,n38,n244);
not (n244,n245);
or (n246,n37,n245);
nand (n247,n248,n252);
or (n248,n114,n249);
nor (n249,n250,n251);
and (n250,n23,n89);
and (n251,n24,n137);
or (n252,n115,n253);
nor (n253,n254,n255);
and (n254,n23,n53);
and (n255,n24,n101);
and (n256,n219,n233);
xor (n257,n258,n273);
xor (n258,n259,n266);
nand (n259,n260,n262);
or (n260,n261,n13);
not (n261,n228);
nand (n262,n21,n263);
nor (n263,n264,n265);
and (n264,n137,n17);
and (n265,n18,n89);
nand (n266,n267,n269);
or (n267,n268,n28);
not (n268,n242);
nand (n269,n31,n270);
nor (n270,n271,n272);
and (n271,n224,n37);
and (n272,n38,n225);
nand (n273,n274,n275);
or (n274,n114,n253);
or (n275,n276,n115);
nor (n276,n277,n278);
and (n277,n23,n70);
and (n278,n24,n72);
xor (n279,n280,n318);
xor (n280,n281,n304);
xor (n281,n282,n293);
xor (n282,n283,n291);
nand (n283,n284,n288);
or (n284,n285,n58);
not (n285,n286);
xor (n286,n287,n52);
nand (n288,n289,n290);
not (n289,n59);
xor (n290,n239,n52);
and (n291,n52,n292);
xor (n293,n294,n297);
nand (n294,n295,n296);
or (n295,n193,n183);
or (n296,n191,n185);
nand (n297,n298,n300);
or (n298,n299,n202);
not (n299,n213);
nand (n300,n204,n301);
nor (n301,n302,n303);
and (n302,n44,n117);
and (n303,n118,n42);
or (n304,n305,n317);
and (n305,n306,n316);
xor (n306,n307,n314);
nand (n307,n308,n313);
or (n308,n309,n58);
nor (n309,n310,n311);
and (n310,n292,n69);
and (n311,n52,n312);
not (n312,n292);
nand (n313,n289,n286);
and (n314,n52,n315);
xor (n316,n181,n196);
and (n317,n307,n314);
or (n318,n319,n364);
and (n319,n320,n363);
xor (n320,n321,n338);
and (n321,n322,n330);
nand (n322,n323,n324);
or (n323,n185,n187);
nand (n324,n325,n329);
not (n325,n326);
nor (n326,n327,n328);
and (n327,n191,n76);
and (n328,n184,n78);
not (n329,n183);
nand (n330,n331,n333);
or (n331,n332,n198);
not (n332,n204);
nand (n333,n334,n203);
not (n334,n335);
nor (n335,n336,n337);
and (n336,n117,n53);
and (n337,n118,n101);
or (n338,n339,n362);
and (n339,n340,n356);
xor (n340,n341,n348);
nand (n341,n342,n347);
or (n342,n343,n13);
not (n343,n344);
nor (n344,n345,n346);
and (n345,n244,n17);
and (n346,n18,n245);
nand (n347,n222,n21);
nand (n348,n349,n355);
or (n349,n350,n28);
not (n350,n351);
nand (n351,n352,n354);
or (n352,n38,n353);
not (n353,n287);
or (n354,n37,n287);
nand (n355,n31,n236);
nand (n356,n357,n361);
or (n357,n114,n358);
nor (n358,n359,n360);
and (n359,n231,n23);
and (n360,n24,n230);
or (n361,n249,n115);
and (n362,n341,n348);
xor (n363,n218,n247);
and (n364,n321,n338);
or (n365,n366,n424);
and (n366,n367,n383);
xor (n367,n368,n369);
xor (n368,n306,n316);
or (n369,n370,n382);
and (n370,n371,n381);
xor (n371,n372,n379);
nand (n372,n373,n378);
or (n373,n58,n374);
nor (n374,n375,n376);
and (n375,n315,n69);
and (n376,n52,n377);
not (n377,n315);
or (n378,n309,n59);
and (n379,n52,n380);
xor (n381,n322,n330);
and (n382,n372,n379);
or (n383,n384,n423);
and (n384,n385,n422);
xor (n385,n386,n399);
and (n386,n387,n393);
nand (n387,n388,n392);
or (n388,n183,n389);
nor (n389,n390,n391);
and (n390,n191,n70);
and (n391,n184,n72);
or (n392,n326,n185);
nand (n393,n394,n398);
or (n394,n202,n395);
nor (n395,n396,n397);
and (n396,n117,n89);
and (n397,n118,n137);
or (n398,n332,n335);
or (n399,n400,n421);
and (n400,n401,n415);
xor (n401,n402,n409);
nand (n402,n403,n408);
or (n403,n404,n13);
not (n404,n405);
nor (n405,n406,n407);
and (n406,n238,n17);
and (n407,n18,n239);
nand (n408,n21,n344);
nand (n409,n410,n414);
or (n410,n28,n411);
nor (n411,n412,n413);
and (n412,n37,n292);
and (n413,n38,n312);
nand (n414,n31,n351);
nand (n415,n416,n420);
or (n416,n114,n417);
nor (n417,n418,n419);
and (n418,n225,n23);
and (n419,n24,n224);
or (n420,n115,n358);
and (n421,n402,n409);
xor (n422,n340,n356);
and (n423,n386,n399);
and (n424,n368,n369);
or (n425,n426,n493);
and (n426,n427,n492);
xor (n427,n428,n429);
xor (n428,n320,n363);
or (n429,n430,n491);
and (n430,n431,n445);
xor (n431,n432,n433);
xor (n432,n371,n381);
or (n433,n434,n444);
and (n434,n435,n443);
xor (n435,n436,n441);
nand (n436,n437,n440);
or (n437,n438,n58);
not (n438,n439);
xor (n439,n380,n52);
or (n440,n59,n374);
and (n441,n52,n442);
xor (n443,n387,n393);
and (n444,n436,n441);
and (n445,n446,n470);
or (n446,n447,n469);
and (n447,n448,n463);
xor (n448,n449,n457);
nand (n449,n450,n455);
or (n450,n451,n202);
not (n451,n452);
nand (n452,n453,n454);
or (n453,n118,n230);
or (n454,n117,n231);
nand (n455,n456,n204);
not (n456,n395);
nand (n457,n458,n462);
or (n458,n13,n459);
nor (n459,n460,n461);
and (n460,n17,n287);
and (n461,n18,n353);
or (n462,n20,n404);
nand (n463,n464,n468);
or (n464,n28,n465);
nor (n465,n466,n467);
and (n466,n37,n315);
and (n467,n38,n377);
or (n468,n30,n411);
and (n469,n449,n457);
or (n470,n471,n490);
and (n471,n472,n488);
xor (n472,n473,n479);
nand (n473,n474,n478);
or (n474,n114,n475);
nor (n475,n476,n477);
and (n476,n23,n245);
and (n477,n24,n244);
or (n478,n417,n115);
nand (n479,n480,n481);
or (n480,n438,n59);
nand (n481,n482,n487);
not (n482,n483);
nor (n483,n484,n485);
and (n484,n442,n69);
and (n485,n486,n52);
not (n486,n442);
not (n487,n58);
and (n488,n52,n489);
and (n490,n473,n479);
and (n491,n432,n433);
xor (n492,n367,n383);
and (n493,n428,n429);
nand (n494,n495,n496);
xor (n495,n427,n492);
or (n496,n497,n561);
and (n497,n498,n501);
xor (n498,n499,n500);
xor (n499,n385,n422);
xor (n500,n431,n445);
or (n501,n502,n560);
and (n502,n503,n506);
xor (n503,n504,n505);
xor (n504,n401,n415);
xor (n505,n435,n443);
or (n506,n507,n559);
and (n507,n508,n533);
xor (n508,n509,n515);
nand (n509,n510,n514);
or (n510,n183,n511);
nor (n511,n512,n513);
and (n512,n191,n53);
and (n513,n184,n101);
or (n514,n389,n185);
or (n515,n516,n532);
and (n516,n517,n526);
xor (n517,n518,n520);
and (n518,n52,n519);
nand (n520,n521,n522);
or (n521,n332,n451);
nand (n522,n203,n523);
nand (n523,n524,n525);
or (n524,n118,n224);
or (n525,n117,n225);
nand (n526,n527,n531);
or (n527,n13,n528);
nor (n528,n529,n530);
and (n529,n17,n292);
and (n530,n18,n312);
or (n531,n459,n20);
and (n532,n518,n520);
or (n533,n534,n558);
and (n534,n535,n551);
xor (n535,n536,n545);
nand (n536,n537,n543);
or (n537,n538,n28);
not (n538,n539);
nor (n539,n540,n542);
and (n540,n541,n37);
not (n541,n380);
and (n542,n38,n380);
nand (n543,n544,n31);
not (n544,n465);
nand (n545,n546,n550);
or (n546,n547,n183);
nor (n547,n548,n549);
and (n548,n191,n89);
and (n549,n184,n137);
or (n550,n511,n185);
nand (n551,n552,n557);
or (n552,n58,n553);
nor (n553,n554,n555);
and (n554,n69,n489);
and (n555,n52,n556);
not (n556,n489);
or (n557,n59,n483);
and (n558,n536,n545);
and (n559,n509,n515);
and (n560,n504,n505);
and (n561,n499,n500);
nand (n562,n176,n425);
not (n563,n564);
nor (n564,n565,n684);
nor (n565,n566,n675);
xor (n566,n567,n664);
xor (n567,n568,n624);
xor (n568,n569,n603);
xor (n569,n570,n595);
or (n570,n571,n594);
and (n571,n572,n588);
xor (n572,n573,n581);
nand (n573,n574,n576);
or (n574,n575,n13);
not (n575,n263);
nand (n576,n577,n21);
not (n577,n578);
nor (n578,n579,n580);
and (n579,n17,n53);
and (n580,n18,n101);
nand (n581,n582,n584);
or (n582,n583,n28);
not (n583,n270);
nand (n584,n31,n585);
nand (n585,n586,n587);
or (n586,n38,n230);
or (n587,n37,n231);
nand (n588,n589,n590);
or (n589,n114,n276);
or (n590,n115,n591);
nor (n591,n592,n593);
and (n592,n23,n76);
and (n593,n24,n78);
and (n594,n573,n581);
nand (n595,n596,n597);
not (n596,n191);
nor (n597,n598,n599);
and (n598,n203,n301);
nor (n599,n332,n600);
nor (n600,n601,n602);
and (n601,n50,n118);
and (n602,n48,n117);
xor (n603,n604,n621);
xor (n604,n605,n612);
nand (n605,n606,n608);
or (n606,n607,n28);
not (n607,n585);
nand (n608,n31,n609);
nor (n609,n610,n611);
and (n610,n137,n37);
and (n611,n38,n89);
nand (n612,n613,n616);
or (n613,n59,n614);
not (n614,n615);
xor (n615,n225,n52);
nand (n616,n617,n487);
not (n617,n618);
nor (n618,n619,n620);
and (n619,n69,n245);
and (n620,n52,n244);
nand (n621,n622,n623);
or (n622,n202,n600);
or (n623,n332,n117);
xor (n624,n625,n654);
xor (n625,n626,n644);
xor (n626,n627,n636);
xor (n627,n628,n629);
and (n628,n52,n239);
nand (n629,n630,n631);
or (n630,n13,n578);
or (n631,n20,n632);
not (n632,n633);
nor (n633,n634,n635);
and (n634,n18,n70);
and (n635,n72,n17);
not (n636,n637);
nand (n637,n638,n639);
or (n638,n591,n114);
nand (n639,n640,n125);
not (n640,n641);
nor (n641,n642,n643);
and (n642,n44,n24);
and (n643,n42,n23);
or (n644,n645,n653);
and (n645,n646,n652);
xor (n646,n647,n651);
nand (n647,n648,n650);
or (n648,n58,n649);
not (n649,n290);
or (n650,n59,n618);
and (n651,n52,n287);
and (n652,n294,n297);
and (n653,n647,n651);
or (n654,n655,n663);
and (n655,n656,n662);
xor (n656,n657,n660);
or (n657,n658,n659);
and (n658,n258,n273);
and (n659,n259,n266);
nand (n660,n661,n595);
or (n661,n596,n597);
xor (n662,n572,n588);
and (n663,n657,n660);
or (n664,n665,n674);
and (n665,n666,n671);
xor (n666,n667,n668);
xor (n667,n646,n652);
or (n668,n669,n670);
and (n669,n282,n293);
and (n670,n283,n291);
or (n671,n672,n673);
and (n672,n179,n257);
and (n673,n180,n216);
and (n674,n667,n668);
or (n675,n676,n683);
and (n676,n677,n680);
xor (n677,n678,n679);
xor (n678,n656,n662);
xor (n679,n666,n671);
or (n680,n681,n682);
and (n681,n280,n318);
and (n682,n281,n304);
and (n683,n678,n679);
nor (n684,n685,n686);
xor (n685,n677,n680);
or (n686,n687,n688);
and (n687,n177,n365);
and (n688,n178,n279);
nor (n689,n690,n693);
and (n690,n691,n692);
not (n691,n565);
and (n692,n685,n686);
and (n693,n566,n675);
not (n694,n695);
and (n695,n696,n798,n813,n820);
not (n696,n697);
nor (n697,n698,n777);
or (n698,n699,n776);
and (n699,n700,n767);
xor (n700,n701,n721);
or (n701,n702,n720);
and (n702,n703,n707);
xor (n703,n637,n704);
or (n704,n705,n706);
and (n705,n604,n621);
and (n706,n605,n612);
xor (n707,n708,n719);
xor (n708,n709,n713);
nand (n709,n710,n711);
or (n710,n614,n58);
nand (n711,n289,n712);
xor (n712,n231,n52);
nand (n713,n714,n715);
or (n714,n632,n13);
nand (n715,n21,n716);
nor (n716,n717,n718);
and (n717,n78,n17);
and (n718,n18,n76);
and (n719,n52,n245);
and (n720,n637,n704);
xor (n721,n722,n752);
xor (n722,n723,n742);
or (n723,n724,n741);
and (n724,n725,n734);
xor (n725,n726,n728);
nand (n726,n727,n118);
or (n727,n203,n204);
nand (n728,n729,n730);
or (n729,n114,n641);
or (n730,n115,n731);
nor (n731,n732,n733);
and (n732,n23,n48);
and (n733,n24,n50);
nand (n734,n735,n737);
or (n735,n28,n736);
not (n736,n609);
or (n737,n30,n738);
nor (n738,n739,n740);
and (n739,n37,n53);
and (n740,n101,n38);
and (n741,n726,n728);
xor (n742,n743,n749);
xor (n743,n744,n748);
nand (n744,n745,n747);
or (n745,n58,n746);
not (n746,n712);
or (n747,n59,n134);
and (n748,n52,n225);
nand (n749,n750,n751);
or (n750,n114,n731);
or (n751,n115,n23);
xor (n752,n753,n764);
xor (n753,n754,n760);
nand (n754,n755,n756);
or (n755,n28,n738);
or (n756,n30,n757);
nor (n757,n758,n759);
and (n758,n37,n70);
and (n759,n38,n72);
nor (n760,n761,n763);
and (n761,n762,n21);
not (n762,n128);
and (n763,n12,n716);
or (n764,n765,n766);
and (n765,n708,n719);
and (n766,n709,n713);
or (n767,n768,n775);
and (n768,n769,n774);
xor (n769,n770,n771);
xor (n770,n725,n734);
or (n771,n772,n773);
and (n772,n627,n636);
and (n773,n628,n629);
xor (n774,n703,n707);
and (n775,n770,n771);
and (n776,n701,n721);
xor (n777,n778,n795);
xor (n778,n779,n782);
or (n779,n780,n781);
and (n780,n753,n764);
and (n781,n754,n760);
xor (n782,n783,n788);
xor (n783,n784,n787);
or (n784,n785,n786);
and (n785,n743,n749);
and (n786,n744,n748);
xor (n787,n110,n132);
xor (n788,n789,n794);
xor (n789,n790,n791);
and (n790,n52,n231);
nand (n791,n792,n793);
or (n792,n28,n757);
or (n793,n92,n30);
not (n794,n760);
or (n795,n796,n797);
and (n796,n722,n752);
and (n797,n723,n742);
nand (n798,n799,n811);
not (n799,n800);
or (n800,n801,n810);
and (n801,n802,n807);
xor (n802,n803,n806);
or (n803,n804,n805);
and (n804,n569,n603);
and (n805,n570,n595);
xor (n806,n769,n774);
or (n807,n808,n809);
and (n808,n625,n654);
and (n809,n626,n644);
and (n810,n803,n806);
not (n811,n812);
xor (n812,n700,n767);
nand (n813,n814,n818);
not (n814,n815);
or (n815,n816,n817);
and (n816,n567,n664);
and (n817,n568,n624);
not (n818,n819);
xor (n819,n802,n807);
nand (n820,n821,n831);
not (n821,n822);
xor (n822,n823,n828);
xor (n823,n824,n827);
or (n824,n825,n826);
and (n825,n789,n794);
and (n826,n790,n791);
xor (n827,n106,n140);
or (n828,n829,n830);
and (n829,n783,n788);
and (n830,n784,n787);
not (n831,n832);
or (n832,n833,n834);
and (n833,n778,n795);
and (n834,n779,n782);
and (n835,n836,n845);
nand (n836,n837,n843);
nand (n837,n838,n842);
or (n838,n839,n840);
not (n839,n798);
not (n840,n841);
nor (n841,n814,n818);
nand (n842,n812,n800);
nor (n843,n697,n844);
not (n844,n820);
nor (n845,n846,n848);
and (n846,n847,n820);
and (n847,n698,n777);
nor (n848,n831,n821);
not (n849,n850);
nor (n850,n851,n854);
or (n851,n852,n853);
and (n852,n823,n828);
and (n853,n824,n827);
xor (n854,n7,n104);
nand (n855,n856,n862);
not (n856,n857);
nand (n857,n695,n858);
and (n858,n691,n859,n860);
not (n859,n684);
nor (n860,n861,n175);
nor (n861,n495,n496);
and (n862,n863,n849);
nand (n863,n864,n1086);
not (n864,n865);
nand (n865,n866,n1079);
or (n866,n867,n1057);
not (n867,n868);
nand (n868,n869,n1056);
or (n869,n870,n1005);
nor (n870,n871,n951);
xor (n871,n872,n917);
xor (n872,n873,n874);
xor (n873,n508,n533);
or (n874,n875,n916);
and (n875,n876,n879);
xor (n876,n877,n878);
xor (n877,n535,n551);
xor (n878,n517,n526);
or (n879,n880,n915);
and (n880,n881,n898);
xor (n881,n882,n889);
nand (n882,n883,n888);
or (n883,n58,n884);
nor (n884,n885,n886);
and (n885,n519,n69);
and (n886,n887,n52);
not (n887,n519);
or (n888,n59,n553);
nand (n889,n890,n894);
or (n890,n114,n891);
nor (n891,n892,n893);
and (n892,n23,n287);
and (n893,n24,n353);
or (n894,n115,n895);
nor (n895,n896,n897);
and (n896,n23,n239);
and (n897,n24,n238);
nand (n898,n899,n914);
or (n899,n900,n906);
not (n900,n901);
nand (n901,n902,n52);
nand (n902,n903,n904);
or (n903,n38,n61);
nand (n904,n905,n887);
or (n905,n63,n37);
not (n906,n907);
nand (n907,n908,n913);
or (n908,n909,n202);
not (n909,n910);
nand (n910,n911,n912);
or (n911,n118,n244);
or (n912,n117,n245);
nand (n913,n204,n523);
or (n914,n907,n901);
and (n915,n882,n889);
and (n916,n877,n878);
xor (n917,n918,n921);
xor (n918,n919,n920);
xor (n919,n472,n488);
xor (n920,n448,n463);
or (n921,n922,n950);
and (n922,n923,n928);
xor (n923,n924,n927);
nand (n924,n925,n926);
or (n925,n114,n895);
or (n926,n115,n475);
nor (n927,n906,n901);
or (n928,n929,n949);
and (n929,n930,n943);
xor (n930,n931,n937);
nand (n931,n932,n936);
or (n932,n13,n933);
nor (n933,n934,n935);
and (n934,n17,n315);
and (n935,n18,n377);
or (n936,n20,n528);
nand (n937,n938,n942);
or (n938,n28,n939);
nor (n939,n940,n941);
and (n940,n37,n442);
and (n941,n38,n486);
or (n942,n30,n538);
nand (n943,n944,n948);
or (n944,n945,n183);
nor (n945,n946,n947);
and (n946,n191,n231);
and (n947,n184,n230);
or (n948,n547,n185);
and (n949,n931,n937);
and (n950,n924,n927);
or (n951,n952,n1004);
and (n952,n953,n1003);
xor (n953,n954,n955);
xor (n954,n923,n928);
or (n955,n956,n1002);
and (n956,n957,n1001);
xor (n957,n958,n977);
or (n958,n959,n976);
and (n959,n960,n968);
xor (n960,n961,n962);
nor (n961,n59,n887);
nand (n962,n963,n967);
or (n963,n964,n202);
nor (n964,n965,n966);
and (n965,n238,n118);
and (n966,n239,n117);
nand (n967,n910,n204);
nand (n968,n969,n974);
or (n969,n970,n13);
not (n970,n971);
nand (n971,n972,n973);
or (n972,n18,n541);
or (n973,n17,n380);
nand (n974,n975,n21);
not (n975,n933);
and (n976,n961,n962);
or (n977,n978,n1000);
and (n978,n979,n994);
xor (n979,n980,n988);
nand (n980,n981,n986);
or (n981,n982,n28);
not (n982,n983);
nand (n983,n984,n985);
or (n984,n38,n556);
or (n985,n37,n489);
nand (n986,n987,n31);
not (n987,n939);
nand (n988,n989,n993);
or (n989,n990,n183);
nor (n990,n991,n992);
and (n991,n191,n225);
and (n992,n184,n224);
or (n993,n945,n185);
nand (n994,n995,n999);
or (n995,n114,n996);
nor (n996,n997,n998);
and (n997,n23,n292);
and (n998,n24,n312);
or (n999,n115,n891);
and (n1000,n980,n988);
xor (n1001,n930,n943);
and (n1002,n958,n977);
xor (n1003,n876,n879);
and (n1004,n954,n955);
nand (n1005,n1006,n1007);
xor (n1006,n953,n1003);
or (n1007,n1008,n1055);
and (n1008,n1009,n1012);
xor (n1009,n1010,n1011);
xor (n1010,n881,n898);
xor (n1011,n957,n1001);
or (n1012,n1013,n1054);
and (n1013,n1014,n1053);
xor (n1014,n1015,n1029);
and (n1015,n1016,n1022);
and (n1016,n1017,n38);
nand (n1017,n1018,n1019);
or (n1018,n18,n33);
nand (n1019,n1020,n887);
or (n1020,n1021,n17);
not (n1021,n33);
nand (n1022,n1023,n1028);
or (n1023,n1024,n202);
not (n1024,n1025);
nand (n1025,n1026,n1027);
or (n1026,n118,n353);
or (n1027,n117,n287);
or (n1028,n332,n964);
or (n1029,n1030,n1052);
and (n1030,n1031,n1045);
xor (n1031,n1032,n1038);
nand (n1032,n1033,n1034);
or (n1033,n20,n970);
or (n1034,n1035,n13);
nor (n1035,n1036,n1037);
and (n1036,n486,n18);
and (n1037,n442,n17);
nand (n1038,n1039,n1044);
or (n1039,n1040,n28);
not (n1040,n1041);
nand (n1041,n1042,n1043);
or (n1042,n38,n887);
or (n1043,n37,n519);
nand (n1044,n983,n31);
nand (n1045,n1046,n1051);
or (n1046,n1047,n183);
not (n1047,n1048);
nor (n1048,n1049,n1050);
and (n1049,n244,n191);
and (n1050,n184,n245);
or (n1051,n990,n185);
and (n1052,n1032,n1038);
xor (n1053,n960,n968);
and (n1054,n1015,n1029);
and (n1055,n1010,n1011);
nand (n1056,n871,n951);
not (n1057,n1058);
nor (n1058,n1059,n1074);
nor (n1059,n1060,n1071);
xor (n1060,n1061,n1068);
xor (n1061,n1062,n1067);
nand (n1062,n1063,n1065);
or (n1063,n470,n1064);
not (n1064,n446);
or (n1065,n446,n1066);
not (n1066,n470);
xor (n1067,n503,n506);
or (n1068,n1069,n1070);
and (n1069,n918,n921);
and (n1070,n919,n920);
or (n1071,n1072,n1073);
and (n1072,n872,n917);
and (n1073,n873,n874);
nor (n1074,n1075,n1076);
xor (n1075,n498,n501);
or (n1076,n1077,n1078);
and (n1077,n1061,n1068);
and (n1078,n1062,n1067);
nor (n1079,n1080,n1085);
and (n1080,n1081,n1082);
not (n1081,n1074);
nor (n1082,n1083,n1084);
not (n1083,n1060);
not (n1084,n1071);
and (n1085,n1075,n1076);
nand (n1086,n1058,n1087,n1376);
nand (n1087,n1088,n1364,n1375);
nand (n1088,n1089,n1127,n1226);
nand (n1089,n1090,n1092);
not (n1090,n1091);
xor (n1091,n1009,n1012);
not (n1092,n1093);
or (n1093,n1094,n1126);
and (n1094,n1095,n1125);
xor (n1095,n1096,n1097);
xor (n1096,n979,n994);
or (n1097,n1098,n1124);
and (n1098,n1099,n1107);
xor (n1099,n1100,n1106);
nand (n1100,n1101,n1105);
or (n1101,n114,n1102);
nor (n1102,n1103,n1104);
and (n1103,n23,n315);
and (n1104,n24,n377);
or (n1105,n996,n115);
xor (n1106,n1016,n1022);
or (n1107,n1108,n1123);
and (n1108,n1109,n1117);
xor (n1109,n1110,n1111);
and (n1110,n31,n519);
nand (n1111,n1112,n1113);
or (n1112,n185,n1047);
or (n1113,n1114,n183);
nor (n1114,n1115,n1116);
and (n1115,n191,n239);
and (n1116,n184,n238);
nand (n1117,n1118,n1122);
or (n1118,n13,n1119);
nor (n1119,n1120,n1121);
and (n1120,n17,n489);
and (n1121,n18,n556);
or (n1122,n20,n1035);
and (n1123,n1110,n1111);
and (n1124,n1100,n1106);
xor (n1125,n1014,n1053);
and (n1126,n1096,n1097);
nor (n1127,n1128,n1221);
not (n1128,n1129);
nor (n1129,n1130,n1194);
nor (n1130,n1131,n1166);
xor (n1131,n1132,n1165);
xor (n1132,n1133,n1134);
xor (n1133,n1031,n1045);
or (n1134,n1135,n1164);
and (n1135,n1136,n1150);
xor (n1136,n1137,n1144);
nand (n1137,n1138,n1143);
or (n1138,n1139,n202);
not (n1139,n1140);
nand (n1140,n1141,n1142);
or (n1141,n118,n312);
or (n1142,n117,n292);
nand (n1143,n204,n1025);
nand (n1144,n1145,n1149);
or (n1145,n114,n1146);
nor (n1146,n1147,n1148);
and (n1147,n380,n23);
and (n1148,n24,n541);
or (n1149,n115,n1102);
and (n1150,n1151,n1157);
nor (n1151,n1152,n17);
nor (n1152,n1153,n1155);
and (n1153,n1154,n887);
nand (n1154,n24,n16);
and (n1155,n23,n1156);
not (n1156,n16);
nand (n1157,n1158,n1163);
or (n1158,n183,n1159);
not (n1159,n1160);
nor (n1160,n1161,n1162);
and (n1161,n184,n287);
and (n1162,n353,n191);
or (n1163,n1114,n185);
and (n1164,n1137,n1144);
xor (n1165,n1099,n1107);
or (n1166,n1167,n1193);
and (n1167,n1168,n1192);
xor (n1168,n1169,n1191);
or (n1169,n1170,n1190);
and (n1170,n1171,n1184);
xor (n1171,n1172,n1178);
nand (n1172,n1173,n1177);
or (n1173,n13,n1174);
nor (n1174,n1175,n1176);
and (n1175,n17,n519);
and (n1176,n18,n887);
or (n1177,n1119,n20);
nand (n1178,n1179,n1180);
or (n1179,n1139,n332);
nand (n1180,n203,n1181);
nand (n1181,n1182,n1183);
or (n1182,n118,n377);
or (n1183,n117,n315);
nand (n1184,n1185,n1189);
or (n1185,n114,n1186);
nor (n1186,n1187,n1188);
and (n1187,n23,n442);
and (n1188,n24,n486);
or (n1189,n115,n1146);
and (n1190,n1172,n1178);
xor (n1191,n1109,n1117);
xor (n1192,n1136,n1150);
and (n1193,n1169,n1191);
nor (n1194,n1195,n1196);
xor (n1195,n1168,n1192);
or (n1196,n1197,n1220);
and (n1197,n1198,n1219);
xor (n1198,n1199,n1200);
xor (n1199,n1151,n1157);
or (n1200,n1201,n1218);
and (n1201,n1202,n1211);
xor (n1202,n1203,n1204);
and (n1203,n21,n519);
nand (n1204,n1205,n1206);
or (n1205,n185,n1159);
or (n1206,n1207,n183);
not (n1207,n1208);
nand (n1208,n1209,n1210);
or (n1209,n292,n191);
nand (n1210,n191,n292);
nand (n1211,n1212,n1217);
or (n1212,n1213,n202);
not (n1213,n1214);
nor (n1214,n1215,n1216);
and (n1215,n118,n380);
and (n1216,n541,n117);
nand (n1217,n204,n1181);
and (n1218,n1203,n1204);
xor (n1219,n1171,n1184);
and (n1220,n1199,n1200);
nor (n1221,n1222,n1223);
xor (n1222,n1095,n1125);
or (n1223,n1224,n1225);
and (n1224,n1132,n1165);
and (n1225,n1133,n1134);
or (n1226,n1227,n1363);
and (n1227,n1228,n1255);
xor (n1228,n1229,n1254);
or (n1229,n1230,n1253);
and (n1230,n1231,n1252);
xor (n1231,n1232,n1238);
nand (n1232,n1233,n1237);
or (n1233,n114,n1234);
nor (n1234,n1235,n1236);
and (n1235,n23,n489);
and (n1236,n24,n556);
or (n1237,n115,n1186);
and (n1238,n1239,n1246);
nand (n1239,n1240,n1245);
or (n1240,n183,n1241);
not (n1241,n1242);
nor (n1242,n1243,n1244);
and (n1243,n184,n315);
and (n1244,n377,n191);
nand (n1245,n1208,n186);
not (n1246,n1247);
nand (n1247,n1248,n24);
nand (n1248,n1249,n1250);
or (n1249,n118,n119);
nand (n1250,n1251,n887);
or (n1251,n121,n117);
xor (n1252,n1202,n1211);
and (n1253,n1232,n1238);
xor (n1254,n1198,n1219);
or (n1255,n1256,n1362);
and (n1256,n1257,n1281);
xor (n1257,n1258,n1280);
or (n1258,n1259,n1279);
and (n1259,n1260,n1275);
xor (n1260,n1261,n1268);
nand (n1261,n1262,n1267);
or (n1262,n1263,n202);
not (n1263,n1264);
nand (n1264,n1265,n1266);
or (n1265,n118,n486);
or (n1266,n117,n442);
nand (n1267,n204,n1214);
nand (n1268,n1269,n1274);
or (n1269,n1270,n114);
not (n1270,n1271);
nand (n1271,n1272,n1273);
or (n1272,n887,n24);
or (n1273,n23,n519);
or (n1274,n115,n1234);
nand (n1275,n1276,n1278);
or (n1276,n1246,n1277);
not (n1277,n1239);
or (n1278,n1239,n1247);
and (n1279,n1261,n1268);
xor (n1280,n1231,n1252);
or (n1281,n1282,n1361);
and (n1282,n1283,n1304);
xor (n1283,n1284,n1303);
or (n1284,n1285,n1302);
and (n1285,n1286,n1295);
xor (n1286,n1287,n1288);
nor (n1287,n115,n887);
nand (n1288,n1289,n1294);
or (n1289,n1290,n202);
not (n1290,n1291);
nor (n1291,n1292,n1293);
and (n1292,n556,n117);
and (n1293,n118,n489);
nand (n1294,n204,n1264);
nand (n1295,n1296,n1301);
or (n1296,n183,n1297);
not (n1297,n1298);
nor (n1298,n1299,n1300);
and (n1299,n541,n191);
and (n1300,n184,n380);
or (n1301,n1241,n185);
and (n1302,n1287,n1288);
xor (n1303,n1260,n1275);
or (n1304,n1305,n1360);
and (n1305,n1306,n1359);
xor (n1306,n1307,n1320);
nor (n1307,n1308,n1315);
not (n1308,n1309);
nand (n1309,n1310,n1311);
or (n1310,n185,n1297);
nand (n1311,n1312,n329);
nor (n1312,n1313,n1314);
and (n1313,n486,n191);
and (n1314,n184,n442);
nand (n1315,n1316,n118);
nand (n1316,n1317,n1318);
or (n1317,n206,n184);
or (n1318,n1319,n519);
and (n1319,n184,n206);
nand (n1320,n1321,n1358);
or (n1321,n1322,n1346);
not (n1322,n1323);
nand (n1323,n1324,n1345);
or (n1324,n1325,n1334);
nor (n1325,n1326,n1327);
and (n1326,n204,n519);
nand (n1327,n1328,n1330);
or (n1328,n185,n1329);
not (n1329,n1312);
nand (n1330,n1331,n329);
nand (n1331,n1332,n1333);
or (n1332,n556,n184);
or (n1333,n191,n489);
nand (n1334,n1335,n1338);
not (n1335,n1336);
nand (n1336,n1337,n184);
nand (n1337,n519,n186);
nand (n1338,n1339,n1341);
or (n1339,n185,n1340);
not (n1340,n1331);
nand (n1341,n1342,n329);
nor (n1342,n1343,n1344);
and (n1343,n887,n191);
and (n1344,n184,n519);
nand (n1345,n1326,n1327);
not (n1346,n1347);
nand (n1347,n1348,n1352);
nor (n1348,n1349,n1350);
and (n1349,n1315,n1309);
and (n1350,n1351,n1308);
not (n1351,n1315);
nor (n1352,n1353,n1357);
and (n1353,n203,n1354);
nand (n1354,n1355,n1356);
or (n1355,n118,n887);
or (n1356,n117,n519);
and (n1357,n204,n1291);
or (n1358,n1348,n1352);
xor (n1359,n1286,n1295);
and (n1360,n1307,n1320);
and (n1361,n1284,n1303);
and (n1362,n1258,n1280);
and (n1363,n1229,n1254);
nand (n1364,n1365,n1089);
nand (n1365,n1366,n1374);
or (n1366,n1221,n1367);
nand (n1367,n1368,n1373);
or (n1368,n1369,n1371);
not (n1369,n1370);
nand (n1370,n1195,n1196);
not (n1371,n1372);
nand (n1372,n1131,n1166);
not (n1373,n1130);
nand (n1374,n1222,n1223);
nand (n1375,n1091,n1093);
nor (n1376,n1377,n870);
not (n1377,n1378);
or (n1378,n1007,n1006);
nand (n1379,n851,n854);
nand (n1380,n2,n165);
xor (n1381,n1382,n2355);
xor (n1382,n1383,n2354);
xor (n1383,n1384,n2299);
xor (n1384,n1385,n2298);
xor (n1385,n1386,n2237);
xor (n1386,n1387,n2236);
or (n1387,n1388,n2172);
and (n1388,n1389,n156);
or (n1389,n1390,n2107);
and (n1390,n1391,n51);
or (n1391,n1392,n2044);
and (n1392,n1393,n88);
or (n1393,n1394,n1980);
and (n1394,n1395,n790);
or (n1395,n1396,n1917);
and (n1396,n1397,n748);
or (n1397,n1398,n1854);
and (n1398,n1399,n719);
or (n1399,n1400,n1791);
and (n1400,n1401,n628);
or (n1401,n1402,n1727);
and (n1402,n1403,n651);
or (n1403,n1404,n1662);
and (n1404,n1405,n291);
or (n1405,n1406,n1598);
and (n1406,n1407,n314);
or (n1407,n1408,n1536);
and (n1408,n1409,n379);
or (n1409,n1410,n1472);
and (n1410,n1411,n441);
and (n1411,n488,n1412);
or (n1412,n1413,n1415);
and (n1413,n518,n1414);
and (n1414,n61,n489);
and (n1415,n1416,n1417);
xor (n1416,n518,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
and (n1419,n61,n519);
and (n1420,n38,n489);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
and (n1425,n38,n519);
and (n1426,n33,n489);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
and (n1431,n33,n519);
and (n1432,n18,n489);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
and (n1437,n18,n519);
and (n1438,n16,n489);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
and (n1443,n16,n519);
and (n1444,n24,n489);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
and (n1449,n24,n519);
and (n1450,n119,n489);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1456);
and (n1454,n1455,n1293);
and (n1455,n119,n519);
and (n1456,n1457,n1458);
xor (n1457,n1455,n1293);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
and (n1460,n118,n519);
and (n1461,n206,n489);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
and (n1466,n206,n519);
and (n1467,n184,n489);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
and (n1470,n1344,n1471);
and (n1471,n186,n489);
and (n1472,n1473,n1474);
xor (n1473,n1411,n441);
or (n1474,n1475,n1478);
and (n1475,n1476,n1477);
xor (n1476,n488,n1412);
and (n1477,n61,n442);
and (n1478,n1479,n1480);
xor (n1479,n1476,n1477);
or (n1480,n1481,n1484);
and (n1481,n1482,n1483);
xor (n1482,n1416,n1417);
and (n1483,n38,n442);
and (n1484,n1485,n1486);
xor (n1485,n1482,n1483);
or (n1486,n1487,n1490);
and (n1487,n1488,n1489);
xor (n1488,n1422,n1423);
and (n1489,n33,n442);
and (n1490,n1491,n1492);
xor (n1491,n1488,n1489);
or (n1492,n1493,n1496);
and (n1493,n1494,n1495);
xor (n1494,n1428,n1429);
and (n1495,n18,n442);
and (n1496,n1497,n1498);
xor (n1497,n1494,n1495);
or (n1498,n1499,n1502);
and (n1499,n1500,n1501);
xor (n1500,n1434,n1435);
and (n1501,n16,n442);
and (n1502,n1503,n1504);
xor (n1503,n1500,n1501);
or (n1504,n1505,n1508);
and (n1505,n1506,n1507);
xor (n1506,n1440,n1441);
and (n1507,n24,n442);
and (n1508,n1509,n1510);
xor (n1509,n1506,n1507);
or (n1510,n1511,n1514);
and (n1511,n1512,n1513);
xor (n1512,n1446,n1447);
and (n1513,n119,n442);
and (n1514,n1515,n1516);
xor (n1515,n1512,n1513);
or (n1516,n1517,n1520);
and (n1517,n1518,n1519);
xor (n1518,n1452,n1453);
and (n1519,n118,n442);
and (n1520,n1521,n1522);
xor (n1521,n1518,n1519);
or (n1522,n1523,n1526);
and (n1523,n1524,n1525);
xor (n1524,n1457,n1458);
and (n1525,n206,n442);
and (n1526,n1527,n1528);
xor (n1527,n1524,n1525);
or (n1528,n1529,n1531);
and (n1529,n1530,n1314);
xor (n1530,n1463,n1464);
and (n1531,n1532,n1533);
xor (n1532,n1530,n1314);
and (n1533,n1534,n1535);
xor (n1534,n1469,n1470);
and (n1535,n186,n442);
and (n1536,n1537,n1538);
xor (n1537,n1409,n379);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1473,n1474);
and (n1541,n61,n380);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
or (n1544,n1545,n1547);
and (n1545,n1546,n542);
xor (n1546,n1479,n1480);
and (n1547,n1548,n1549);
xor (n1548,n1546,n542);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1485,n1486);
and (n1552,n33,n380);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1491,n1492);
and (n1558,n18,n380);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1497,n1498);
and (n1564,n16,n380);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1503,n1504);
and (n1570,n24,n380);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1509,n1510);
and (n1576,n119,n380);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1582);
and (n1580,n1581,n1215);
xor (n1581,n1515,n1516);
and (n1582,n1583,n1584);
xor (n1583,n1581,n1215);
or (n1584,n1585,n1588);
and (n1585,n1586,n1587);
xor (n1586,n1521,n1522);
and (n1587,n206,n380);
and (n1588,n1589,n1590);
xor (n1589,n1586,n1587);
or (n1590,n1591,n1593);
and (n1591,n1592,n1300);
xor (n1592,n1527,n1528);
and (n1593,n1594,n1595);
xor (n1594,n1592,n1300);
and (n1595,n1596,n1597);
xor (n1596,n1532,n1533);
and (n1597,n186,n380);
and (n1598,n1599,n1600);
xor (n1599,n1407,n314);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1537,n1538);
and (n1603,n61,n315);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1543,n1544);
and (n1609,n38,n315);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1548,n1549);
and (n1615,n33,n315);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1554,n1555);
and (n1621,n18,n315);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1560,n1561);
and (n1627,n16,n315);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1566,n1567);
and (n1633,n24,n315);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1572,n1573);
and (n1639,n119,n315);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1578,n1579);
and (n1645,n118,n315);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1583,n1584);
and (n1651,n206,n315);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1657);
and (n1655,n1656,n1243);
xor (n1656,n1589,n1590);
and (n1657,n1658,n1659);
xor (n1658,n1656,n1243);
and (n1659,n1660,n1661);
xor (n1660,n1594,n1595);
and (n1661,n186,n315);
and (n1662,n1663,n1664);
xor (n1663,n1405,n291);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1599,n1600);
and (n1667,n61,n292);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
or (n1670,n1671,n1674);
and (n1671,n1672,n1673);
xor (n1672,n1605,n1606);
and (n1673,n38,n292);
and (n1674,n1675,n1676);
xor (n1675,n1672,n1673);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1611,n1612);
and (n1679,n33,n292);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1617,n1618);
and (n1685,n18,n292);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1623,n1624);
and (n1691,n16,n292);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1629,n1630);
and (n1697,n24,n292);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1635,n1636);
and (n1703,n119,n292);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1641,n1642);
and (n1709,n118,n292);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1716);
and (n1713,n1714,n1715);
xor (n1714,n1647,n1648);
and (n1715,n206,n292);
and (n1716,n1717,n1718);
xor (n1717,n1714,n1715);
or (n1718,n1719,n1722);
and (n1719,n1720,n1721);
xor (n1720,n1653,n1654);
and (n1721,n184,n292);
and (n1722,n1723,n1724);
xor (n1723,n1720,n1721);
and (n1724,n1725,n1726);
xor (n1725,n1658,n1659);
and (n1726,n186,n292);
and (n1727,n1728,n1729);
xor (n1728,n1403,n651);
or (n1729,n1730,n1733);
and (n1730,n1731,n1732);
xor (n1731,n1663,n1664);
and (n1732,n61,n287);
and (n1733,n1734,n1735);
xor (n1734,n1731,n1732);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1669,n1670);
and (n1738,n38,n287);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
or (n1741,n1742,n1745);
and (n1742,n1743,n1744);
xor (n1743,n1675,n1676);
and (n1744,n33,n287);
and (n1745,n1746,n1747);
xor (n1746,n1743,n1744);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1681,n1682);
and (n1750,n18,n287);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1687,n1688);
and (n1756,n16,n287);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1693,n1694);
and (n1762,n24,n287);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1699,n1700);
and (n1768,n119,n287);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1705,n1706);
and (n1774,n118,n287);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1711,n1712);
and (n1780,n206,n287);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1786);
and (n1784,n1785,n1161);
xor (n1785,n1717,n1718);
and (n1786,n1787,n1788);
xor (n1787,n1785,n1161);
and (n1788,n1789,n1790);
xor (n1789,n1723,n1724);
and (n1790,n186,n287);
and (n1791,n1792,n1793);
xor (n1792,n1401,n628);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1728,n1729);
and (n1796,n61,n239);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1802);
and (n1800,n1801,n240);
xor (n1801,n1734,n1735);
and (n1802,n1803,n1804);
xor (n1803,n1801,n240);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1740,n1741);
and (n1807,n33,n239);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1813);
and (n1811,n1812,n407);
xor (n1812,n1746,n1747);
and (n1813,n1814,n1815);
xor (n1814,n1812,n407);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1752,n1753);
and (n1818,n16,n239);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1825);
and (n1822,n1823,n1824);
xor (n1823,n1758,n1759);
and (n1824,n24,n239);
and (n1825,n1826,n1827);
xor (n1826,n1823,n1824);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1764,n1765);
and (n1830,n119,n239);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
or (n1833,n1834,n1837);
and (n1834,n1835,n1836);
xor (n1835,n1770,n1771);
and (n1836,n118,n239);
and (n1837,n1838,n1839);
xor (n1838,n1835,n1836);
or (n1839,n1840,n1843);
and (n1840,n1841,n1842);
xor (n1841,n1776,n1777);
and (n1842,n206,n239);
and (n1843,n1844,n1845);
xor (n1844,n1841,n1842);
or (n1845,n1846,n1849);
and (n1846,n1847,n1848);
xor (n1847,n1782,n1783);
and (n1848,n184,n239);
and (n1849,n1850,n1851);
xor (n1850,n1847,n1848);
and (n1851,n1852,n1853);
xor (n1852,n1787,n1788);
and (n1853,n186,n239);
and (n1854,n1855,n1856);
xor (n1855,n1399,n719);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n1792,n1793);
and (n1859,n61,n245);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1798,n1799);
and (n1865,n38,n245);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
or (n1868,n1869,n1872);
and (n1869,n1870,n1871);
xor (n1870,n1803,n1804);
and (n1871,n33,n245);
and (n1872,n1873,n1874);
xor (n1873,n1870,n1871);
or (n1874,n1875,n1877);
and (n1875,n1876,n346);
xor (n1876,n1809,n1810);
and (n1877,n1878,n1879);
xor (n1878,n1876,n346);
or (n1879,n1880,n1883);
and (n1880,n1881,n1882);
xor (n1881,n1814,n1815);
and (n1882,n16,n245);
and (n1883,n1884,n1885);
xor (n1884,n1881,n1882);
or (n1885,n1886,n1889);
and (n1886,n1887,n1888);
xor (n1887,n1820,n1821);
and (n1888,n24,n245);
and (n1889,n1890,n1891);
xor (n1890,n1887,n1888);
or (n1891,n1892,n1895);
and (n1892,n1893,n1894);
xor (n1893,n1826,n1827);
and (n1894,n119,n245);
and (n1895,n1896,n1897);
xor (n1896,n1893,n1894);
or (n1897,n1898,n1901);
and (n1898,n1899,n1900);
xor (n1899,n1832,n1833);
and (n1900,n118,n245);
and (n1901,n1902,n1903);
xor (n1902,n1899,n1900);
or (n1903,n1904,n1907);
and (n1904,n1905,n1906);
xor (n1905,n1838,n1839);
and (n1906,n206,n245);
and (n1907,n1908,n1909);
xor (n1908,n1905,n1906);
or (n1909,n1910,n1912);
and (n1910,n1911,n1050);
xor (n1911,n1844,n1845);
and (n1912,n1913,n1914);
xor (n1913,n1911,n1050);
and (n1914,n1915,n1916);
xor (n1915,n1850,n1851);
and (n1916,n186,n245);
and (n1917,n1918,n1919);
xor (n1918,n1397,n748);
or (n1919,n1920,n1923);
and (n1920,n1921,n1922);
xor (n1921,n1855,n1856);
and (n1922,n61,n225);
and (n1923,n1924,n1925);
xor (n1924,n1921,n1922);
or (n1925,n1926,n1928);
and (n1926,n1927,n272);
xor (n1927,n1861,n1862);
and (n1928,n1929,n1930);
xor (n1929,n1927,n272);
or (n1930,n1931,n1934);
and (n1931,n1932,n1933);
xor (n1932,n1867,n1868);
and (n1933,n33,n225);
and (n1934,n1935,n1936);
xor (n1935,n1932,n1933);
or (n1936,n1937,n1939);
and (n1937,n1938,n226);
xor (n1938,n1873,n1874);
and (n1939,n1940,n1941);
xor (n1940,n1938,n226);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1878,n1879);
and (n1944,n16,n225);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1884,n1885);
and (n1950,n24,n225);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1890,n1891);
and (n1956,n119,n225);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1963);
and (n1960,n1961,n1962);
xor (n1961,n1896,n1897);
and (n1962,n118,n225);
and (n1963,n1964,n1965);
xor (n1964,n1961,n1962);
or (n1965,n1966,n1969);
and (n1966,n1967,n1968);
xor (n1967,n1902,n1903);
and (n1968,n206,n225);
and (n1969,n1970,n1971);
xor (n1970,n1967,n1968);
or (n1971,n1972,n1975);
and (n1972,n1973,n1974);
xor (n1973,n1908,n1909);
and (n1974,n184,n225);
and (n1975,n1976,n1977);
xor (n1976,n1973,n1974);
and (n1977,n1978,n1979);
xor (n1978,n1913,n1914);
and (n1979,n186,n225);
and (n1980,n1981,n1982);
xor (n1981,n1395,n790);
or (n1982,n1983,n1986);
and (n1983,n1984,n1985);
xor (n1984,n1918,n1919);
and (n1985,n61,n231);
and (n1986,n1987,n1988);
xor (n1987,n1984,n1985);
or (n1988,n1989,n1992);
and (n1989,n1990,n1991);
xor (n1990,n1924,n1925);
and (n1991,n38,n231);
and (n1992,n1993,n1994);
xor (n1993,n1990,n1991);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1929,n1930);
and (n1997,n33,n231);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
or (n2000,n2001,n2003);
and (n2001,n2002,n232);
xor (n2002,n1935,n1936);
and (n2003,n2004,n2005);
xor (n2004,n2002,n232);
or (n2005,n2006,n2009);
and (n2006,n2007,n2008);
xor (n2007,n1940,n1941);
and (n2008,n16,n231);
and (n2009,n2010,n2011);
xor (n2010,n2007,n2008);
or (n2011,n2012,n2015);
and (n2012,n2013,n2014);
xor (n2013,n1946,n1947);
and (n2014,n24,n231);
and (n2015,n2016,n2017);
xor (n2016,n2013,n2014);
or (n2017,n2018,n2021);
and (n2018,n2019,n2020);
xor (n2019,n1952,n1953);
and (n2020,n119,n231);
and (n2021,n2022,n2023);
xor (n2022,n2019,n2020);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
xor (n2025,n1958,n1959);
and (n2026,n118,n231);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1964,n1965);
and (n2032,n206,n231);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1970,n1971);
and (n2038,n184,n231);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
and (n2041,n2042,n2043);
xor (n2042,n1976,n1977);
and (n2043,n186,n231);
and (n2044,n2045,n2046);
xor (n2045,n1393,n88);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1981,n1982);
and (n2049,n61,n89);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
or (n2052,n2053,n2055);
and (n2053,n2054,n611);
xor (n2054,n1987,n1988);
and (n2055,n2056,n2057);
xor (n2056,n2054,n611);
or (n2057,n2058,n2061);
and (n2058,n2059,n2060);
xor (n2059,n1993,n1994);
and (n2060,n33,n89);
and (n2061,n2062,n2063);
xor (n2062,n2059,n2060);
or (n2063,n2064,n2066);
and (n2064,n2065,n265);
xor (n2065,n1999,n2000);
and (n2066,n2067,n2068);
xor (n2067,n2065,n265);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n2004,n2005);
and (n2071,n16,n89);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2078);
and (n2075,n2076,n2077);
xor (n2076,n2010,n2011);
and (n2077,n24,n89);
and (n2078,n2079,n2080);
xor (n2079,n2076,n2077);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n2016,n2017);
and (n2083,n119,n89);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n2022,n2023);
and (n2089,n118,n89);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2028,n2029);
and (n2095,n206,n89);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2034,n2035);
and (n2101,n184,n89);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
and (n2104,n2105,n2106);
xor (n2105,n2040,n2041);
and (n2106,n186,n89);
and (n2107,n2108,n2109);
xor (n2108,n1391,n51);
or (n2109,n2110,n2113);
and (n2110,n2111,n2112);
xor (n2111,n2045,n2046);
and (n2112,n61,n53);
and (n2113,n2114,n2115);
xor (n2114,n2111,n2112);
or (n2115,n2116,n2119);
and (n2116,n2117,n2118);
xor (n2117,n2051,n2052);
and (n2118,n38,n53);
and (n2119,n2120,n2121);
xor (n2120,n2117,n2118);
or (n2121,n2122,n2125);
and (n2122,n2123,n2124);
xor (n2123,n2056,n2057);
and (n2124,n33,n53);
and (n2125,n2126,n2127);
xor (n2126,n2123,n2124);
or (n2127,n2128,n2131);
and (n2128,n2129,n2130);
xor (n2129,n2062,n2063);
and (n2130,n18,n53);
and (n2131,n2132,n2133);
xor (n2132,n2129,n2130);
or (n2133,n2134,n2137);
and (n2134,n2135,n2136);
xor (n2135,n2067,n2068);
and (n2136,n16,n53);
and (n2137,n2138,n2139);
xor (n2138,n2135,n2136);
or (n2139,n2140,n2143);
and (n2140,n2141,n2142);
xor (n2141,n2073,n2074);
and (n2142,n24,n53);
and (n2143,n2144,n2145);
xor (n2144,n2141,n2142);
or (n2145,n2146,n2149);
and (n2146,n2147,n2148);
xor (n2147,n2079,n2080);
and (n2148,n119,n53);
and (n2149,n2150,n2151);
xor (n2150,n2147,n2148);
or (n2151,n2152,n2155);
and (n2152,n2153,n2154);
xor (n2153,n2085,n2086);
and (n2154,n118,n53);
and (n2155,n2156,n2157);
xor (n2156,n2153,n2154);
or (n2157,n2158,n2161);
and (n2158,n2159,n2160);
xor (n2159,n2091,n2092);
and (n2160,n206,n53);
and (n2161,n2162,n2163);
xor (n2162,n2159,n2160);
or (n2163,n2164,n2167);
and (n2164,n2165,n2166);
xor (n2165,n2097,n2098);
and (n2166,n184,n53);
and (n2167,n2168,n2169);
xor (n2168,n2165,n2166);
and (n2169,n2170,n2171);
xor (n2170,n2103,n2104);
and (n2171,n186,n53);
and (n2172,n2173,n2174);
xor (n2173,n1389,n156);
or (n2174,n2175,n2178);
and (n2175,n2176,n2177);
xor (n2176,n2108,n2109);
and (n2177,n61,n70);
and (n2178,n2179,n2180);
xor (n2179,n2176,n2177);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2114,n2115);
and (n2183,n38,n70);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2120,n2121);
and (n2189,n33,n70);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2195);
and (n2193,n2194,n634);
xor (n2194,n2126,n2127);
and (n2195,n2196,n2197);
xor (n2196,n2194,n634);
or (n2197,n2198,n2201);
and (n2198,n2199,n2200);
xor (n2199,n2132,n2133);
and (n2200,n16,n70);
and (n2201,n2202,n2203);
xor (n2202,n2199,n2200);
or (n2203,n2204,n2207);
and (n2204,n2205,n2206);
xor (n2205,n2138,n2139);
and (n2206,n24,n70);
and (n2207,n2208,n2209);
xor (n2208,n2205,n2206);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2144,n2145);
and (n2212,n119,n70);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
or (n2215,n2216,n2219);
and (n2216,n2217,n2218);
xor (n2217,n2150,n2151);
and (n2218,n118,n70);
and (n2219,n2220,n2221);
xor (n2220,n2217,n2218);
or (n2221,n2222,n2225);
and (n2222,n2223,n2224);
xor (n2223,n2156,n2157);
and (n2224,n206,n70);
and (n2225,n2226,n2227);
xor (n2226,n2223,n2224);
or (n2227,n2228,n2231);
and (n2228,n2229,n2230);
xor (n2229,n2162,n2163);
and (n2230,n184,n70);
and (n2231,n2232,n2233);
xor (n2232,n2229,n2230);
and (n2233,n2234,n2235);
xor (n2234,n2168,n2169);
and (n2235,n186,n70);
and (n2236,n52,n76);
or (n2237,n2238,n2241);
and (n2238,n2239,n2240);
xor (n2239,n2173,n2174);
and (n2240,n61,n76);
and (n2241,n2242,n2243);
xor (n2242,n2239,n2240);
or (n2243,n2244,n2247);
and (n2244,n2245,n2246);
xor (n2245,n2179,n2180);
and (n2246,n38,n76);
and (n2247,n2248,n2249);
xor (n2248,n2245,n2246);
or (n2249,n2250,n2253);
and (n2250,n2251,n2252);
xor (n2251,n2185,n2186);
and (n2252,n33,n76);
and (n2253,n2254,n2255);
xor (n2254,n2251,n2252);
or (n2255,n2256,n2258);
and (n2256,n2257,n718);
xor (n2257,n2191,n2192);
and (n2258,n2259,n2260);
xor (n2259,n2257,n718);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2196,n2197);
and (n2263,n16,n76);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2202,n2203);
and (n2269,n24,n76);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2208,n2209);
and (n2275,n119,n76);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2281);
and (n2279,n2280,n214);
xor (n2280,n2214,n2215);
and (n2281,n2282,n2283);
xor (n2282,n2280,n214);
or (n2283,n2284,n2287);
and (n2284,n2285,n2286);
xor (n2285,n2220,n2221);
and (n2286,n206,n76);
and (n2287,n2288,n2289);
xor (n2288,n2285,n2286);
or (n2289,n2290,n2293);
and (n2290,n2291,n2292);
xor (n2291,n2226,n2227);
and (n2292,n184,n76);
and (n2293,n2294,n2295);
xor (n2294,n2291,n2292);
and (n2295,n2296,n2297);
xor (n2296,n2232,n2233);
and (n2297,n186,n76);
and (n2298,n61,n42);
or (n2299,n2300,n2303);
and (n2300,n2301,n2302);
xor (n2301,n2242,n2243);
and (n2302,n38,n42);
and (n2303,n2304,n2305);
xor (n2304,n2301,n2302);
or (n2305,n2306,n2309);
and (n2306,n2307,n2308);
xor (n2307,n2248,n2249);
and (n2308,n33,n42);
and (n2309,n2310,n2311);
xor (n2310,n2307,n2308);
or (n2311,n2312,n2315);
and (n2312,n2313,n2314);
xor (n2313,n2254,n2255);
and (n2314,n18,n42);
and (n2315,n2316,n2317);
xor (n2316,n2313,n2314);
or (n2317,n2318,n2321);
and (n2318,n2319,n2320);
xor (n2319,n2259,n2260);
and (n2320,n16,n42);
and (n2321,n2322,n2323);
xor (n2322,n2319,n2320);
or (n2323,n2324,n2327);
and (n2324,n2325,n2326);
xor (n2325,n2265,n2266);
and (n2326,n24,n42);
and (n2327,n2328,n2329);
xor (n2328,n2325,n2326);
or (n2329,n2330,n2333);
and (n2330,n2331,n2332);
xor (n2331,n2271,n2272);
and (n2332,n119,n42);
and (n2333,n2334,n2335);
xor (n2334,n2331,n2332);
or (n2335,n2336,n2338);
and (n2336,n2337,n303);
xor (n2337,n2277,n2278);
and (n2338,n2339,n2340);
xor (n2339,n2337,n303);
or (n2340,n2341,n2344);
and (n2341,n2342,n2343);
xor (n2342,n2282,n2283);
and (n2343,n206,n42);
and (n2344,n2345,n2346);
xor (n2345,n2342,n2343);
or (n2346,n2347,n2349);
and (n2347,n2348,n189);
xor (n2348,n2288,n2289);
and (n2349,n2350,n2351);
xor (n2350,n2348,n189);
and (n2351,n2352,n2353);
xor (n2352,n2294,n2295);
and (n2353,n186,n42);
and (n2354,n38,n48);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2304,n2305);
and (n2358,n33,n48);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2310,n2311);
and (n2364,n18,n48);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2316,n2317);
and (n2370,n16,n48);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2322,n2323);
and (n2376,n24,n48);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2328,n2329);
and (n2382,n119,n48);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2334,n2335);
and (n2388,n118,n48);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2339,n2340);
and (n2394,n206,n48);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2345,n2346);
and (n2400,n184,n48);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
and (n2403,n2404,n2405);
xor (n2404,n2350,n2351);
and (n2405,n186,n48);
endmodule
