module top (out,n13,n15,n22,n23,n32,n40,n42,n48,n58
        ,n67,n71,n93,n95,n103,n109,n132,n136,n141,n147
        ,n151,n157,n185,n262,n266,n328,n332,n364);
output out;
input n13;
input n15;
input n22;
input n23;
input n32;
input n40;
input n42;
input n48;
input n58;
input n67;
input n71;
input n93;
input n95;
input n103;
input n109;
input n132;
input n136;
input n141;
input n147;
input n151;
input n157;
input n185;
input n262;
input n266;
input n328;
input n332;
input n364;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n263;
wire n264;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n329;
wire n330;
wire n331;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
xor (out,n0,n377);
xor (n0,n1,n211);
and (n1,n2,n210);
nand (n2,n3,n177);
not (n3,n4);
xor (n4,n5,n123);
xor (n5,n6,n72);
xor (n6,n7,n60);
xor (n7,n8,n35);
nand (n8,n9,n26);
or (n9,n10,n17);
not (n10,n11);
nand (n11,n12,n16);
or (n12,n13,n14);
not (n14,n15);
nand (n16,n13,n14);
not (n17,n18);
nand (n18,n19,n24);
nand (n19,n20,n23);
nor (n20,n21,n13);
not (n21,n22);
nand (n24,n25,n13,n21);
not (n25,n23);
nand (n26,n27,n30);
nor (n27,n28,n29);
and (n28,n21,n25);
and (n29,n22,n23);
nand (n30,n31,n34);
or (n31,n32,n33);
not (n33,n13);
nand (n34,n33,n32);
nand (n35,n36,n51);
or (n36,n37,n44);
not (n37,n38);
nand (n38,n39,n43);
or (n39,n40,n41);
not (n41,n42);
nand (n43,n40,n41);
not (n44,n45);
nand (n45,n46,n49);
nand (n46,n33,n47,n40);
not (n47,n48);
nand (n49,n50,n48,n13);
not (n50,n40);
nand (n51,n52,n55);
nand (n52,n53,n54);
or (n53,n48,n33);
nand (n54,n33,n48);
nand (n55,n56,n59);
or (n56,n57,n40);
not (n57,n58);
nand (n59,n40,n57);
nor (n60,n61,n70);
not (n61,n62);
nor (n62,n63,n50);
and (n63,n64,n68);
nand (n64,n65,n33);
not (n65,n66);
and (n66,n67,n48);
nand (n68,n69,n47);
not (n69,n67);
not (n70,n71);
or (n72,n73,n122);
and (n73,n74,n106);
xor (n74,n75,n82);
nand (n75,n76,n81);
or (n76,n77,n44);
not (n77,n78);
nand (n78,n79,n80);
or (n79,n50,n67);
or (n80,n69,n40);
nand (n81,n52,n38);
nand (n82,n83,n97);
or (n83,n84,n89);
not (n84,n85);
nor (n85,n86,n87);
and (n86,n32,n23);
and (n87,n88,n25);
not (n88,n32);
not (n89,n90);
nand (n90,n91,n96);
nand (n91,n23,n92,n94);
not (n92,n93);
not (n94,n95);
nand (n96,n25,n93,n95);
nand (n97,n98,n101);
nand (n98,n99,n100);
or (n99,n92,n95);
nand (n100,n92,n95);
nor (n101,n102,n104);
and (n102,n103,n23);
and (n104,n105,n25);
not (n105,n103);
or (n106,n107,n121);
and (n107,n108,n111);
xor (n108,n109,n110);
and (n110,n52,n67);
nand (n111,n112,n117);
or (n112,n113,n17);
not (n113,n114);
nand (n114,n115,n116);
or (n115,n41,n13);
nand (n116,n13,n41);
nand (n117,n27,n118);
nand (n118,n119,n120);
or (n119,n57,n13);
nand (n120,n13,n57);
and (n121,n109,n110);
and (n122,n75,n82);
xor (n123,n124,n159);
xor (n124,n125,n134);
nand (n125,n126,n128);
or (n126,n127,n89);
not (n127,n101);
nand (n128,n98,n129);
nand (n129,n130,n133);
or (n130,n131,n23);
not (n131,n132);
nand (n133,n23,n131);
xor (n134,n135,n143);
xor (n135,n136,n137);
and (n137,n138,n67);
nand (n138,n139,n142);
or (n139,n140,n40);
not (n140,n141);
nand (n142,n40,n140);
nand (n143,n144,n153);
or (n144,n145,n148);
nand (n145,n146,n93);
not (n146,n147);
not (n148,n149);
nand (n149,n150,n152);
or (n150,n151,n92);
nand (n152,n92,n151);
nand (n153,n154,n147);
nand (n154,n155,n158);
or (n155,n156,n93);
not (n156,n157);
nand (n158,n93,n156);
or (n159,n160,n176);
and (n160,n161,n173);
xor (n161,n162,n169);
nand (n162,n163,n168);
or (n163,n145,n164);
not (n164,n165);
nand (n165,n166,n167);
or (n166,n131,n93);
nand (n167,n93,n131);
nand (n168,n149,n147);
nand (n169,n170,n172);
or (n170,n171,n17);
not (n171,n118);
nand (n172,n27,n11);
nand (n173,n174,n175);
or (n174,n71,n61);
nand (n175,n61,n71);
and (n176,n162,n169);
not (n177,n178);
or (n178,n179,n209);
and (n179,n180,n208);
xor (n180,n181,n207);
or (n181,n182,n206);
and (n182,n183,n199);
xor (n183,n184,n192);
and (n184,n185,n186);
nor (n186,n187,n33);
and (n187,n188,n191);
nand (n188,n189,n25);
not (n189,n190);
and (n190,n67,n22);
nand (n191,n21,n69);
nand (n192,n193,n198);
or (n193,n145,n194);
not (n194,n195);
nand (n195,n196,n197);
or (n196,n103,n92);
nand (n197,n92,n103);
nand (n198,n165,n147);
nand (n199,n200,n205);
or (n200,n201,n89);
not (n201,n202);
nor (n202,n203,n204);
and (n203,n15,n23);
and (n204,n14,n25);
nand (n205,n98,n85);
and (n206,n184,n192);
xor (n207,n161,n173);
xor (n208,n74,n106);
and (n209,n181,n207);
nand (n210,n4,n178);
nand (n211,n212,n376);
or (n212,n213,n241);
not (n213,n214);
or (n214,n215,n216);
xor (n215,n180,n208);
or (n216,n217,n240);
and (n217,n218,n239);
xor (n218,n219,n220);
xor (n219,n108,n111);
or (n220,n221,n238);
and (n221,n222,n231);
xor (n222,n223,n230);
nand (n223,n224,n229);
or (n224,n225,n17);
not (n225,n226);
nand (n226,n227,n228);
or (n227,n13,n69);
nand (n228,n69,n13);
nand (n229,n114,n27);
xor (n230,n185,n186);
nand (n231,n232,n237);
or (n232,n145,n233);
not (n233,n234);
nand (n234,n235,n236);
or (n235,n32,n92);
nand (n236,n92,n32);
nand (n237,n195,n147);
and (n238,n223,n230);
xor (n239,n183,n199);
and (n240,n219,n220);
not (n241,n242);
nand (n242,n243,n375);
or (n243,n244,n275);
not (n244,n245);
nand (n245,n246,n248);
not (n246,n247);
xor (n247,n218,n239);
not (n248,n249);
or (n249,n250,n274);
and (n250,n251,n273);
xor (n251,n252,n259);
nand (n252,n253,n258);
or (n253,n254,n89);
not (n254,n255);
nand (n255,n256,n257);
or (n256,n58,n25);
nand (n257,n25,n58);
nand (n258,n98,n202);
or (n259,n260,n272);
and (n260,n261,n264);
xor (n261,n262,n263);
and (n263,n27,n67);
nor (n264,n265,n267);
not (n265,n266);
nand (n267,n268,n23);
or (n268,n269,n271);
nor (n269,n270,n93);
and (n270,n67,n95);
nor (n271,n67,n95);
and (n272,n262,n263);
xor (n273,n222,n231);
and (n274,n252,n259);
not (n275,n276);
or (n276,n277,n374);
and (n277,n278,n298);
xor (n278,n279,n297);
or (n279,n280,n296);
and (n280,n281,n295);
xor (n281,n282,n289);
nand (n282,n283,n284);
or (n283,n146,n233);
nand (n284,n285,n286);
not (n285,n145);
nand (n286,n287,n288);
or (n287,n15,n92);
nand (n288,n92,n15);
nand (n289,n290,n294);
nand (n290,n90,n291);
nand (n291,n292,n293);
or (n292,n42,n25);
nand (n293,n25,n42);
nand (n294,n255,n98);
xor (n295,n261,n264);
and (n296,n282,n289);
xor (n297,n251,n273);
nand (n298,n299,n373);
or (n299,n300,n368);
nor (n300,n301,n367);
and (n301,n302,n337);
nand (n302,n303,n324);
not (n303,n304);
xor (n304,n305,n317);
xor (n305,n306,n313);
nand (n306,n307,n309);
or (n307,n146,n308);
not (n308,n286);
nand (n309,n310,n285);
nand (n310,n311,n312);
or (n311,n58,n92);
nand (n312,n92,n58);
nand (n313,n314,n316);
or (n314,n265,n315);
not (n315,n267);
nand (n316,n265,n315);
nand (n317,n318,n323);
or (n318,n319,n89);
not (n319,n320);
nand (n320,n321,n322);
or (n321,n25,n67);
nand (n322,n67,n25);
nand (n323,n98,n291);
not (n324,n325);
or (n325,n326,n336);
and (n326,n327,n330);
xor (n327,n328,n329);
and (n329,n98,n67);
nor (n330,n331,n333);
not (n331,n332);
nand (n333,n334,n93);
not (n334,n335);
and (n335,n67,n147);
and (n336,n328,n329);
nand (n337,n338,n366);
or (n338,n339,n349);
nor (n339,n340,n341);
xor (n340,n327,n330);
nand (n341,n342,n347);
or (n342,n343,n145);
not (n343,n344);
nor (n344,n345,n346);
and (n345,n41,n92);
and (n346,n42,n93);
or (n347,n348,n146);
not (n348,n310);
nor (n349,n350,n365);
and (n350,n351,n363);
nand (n351,n352,n356);
nor (n352,n353,n355);
and (n353,n354,n331);
not (n354,n333);
and (n355,n333,n332);
not (n356,n357);
nand (n357,n358,n359);
or (n358,n146,n343);
nand (n359,n360,n285);
nand (n360,n361,n362);
or (n361,n67,n92);
nand (n362,n92,n67);
and (n363,n335,n364);
nor (n365,n352,n356);
nand (n366,n340,n341);
nor (n367,n303,n324);
nor (n368,n369,n370);
xor (n369,n281,n295);
or (n370,n371,n372);
and (n371,n305,n317);
and (n372,n306,n313);
nand (n373,n369,n370);
and (n374,n279,n297);
nand (n375,n247,n249);
nand (n376,n215,n216);
xor (n377,n378,n543);
xor (n378,n379,n136);
xor (n379,n380,n542);
xor (n380,n381,n539);
xor (n381,n382,n538);
xor (n382,n383,n530);
xor (n383,n384,n529);
xor (n384,n385,n514);
xor (n385,n386,n513);
xor (n386,n387,n493);
xor (n387,n388,n492);
xor (n388,n389,n467);
xor (n389,n390,n102);
xor (n390,n391,n435);
xor (n391,n392,n434);
xor (n392,n393,n396);
xor (n393,n394,n395);
and (n394,n157,n147);
and (n395,n151,n93);
or (n396,n397,n400);
and (n397,n398,n399);
and (n398,n151,n147);
and (n399,n132,n93);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
and (n404,n132,n147);
and (n405,n103,n93);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
and (n410,n103,n147);
and (n411,n32,n93);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
and (n416,n32,n147);
and (n417,n15,n93);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
and (n422,n15,n147);
and (n423,n58,n93);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n429);
and (n427,n428,n346);
and (n428,n58,n147);
and (n429,n430,n431);
xor (n430,n428,n346);
and (n431,n432,n433);
and (n432,n42,n147);
and (n433,n67,n93);
and (n434,n132,n95);
or (n435,n436,n439);
and (n436,n437,n438);
xor (n437,n401,n402);
and (n438,n103,n95);
and (n439,n440,n441);
xor (n440,n437,n438);
or (n441,n442,n445);
and (n442,n443,n444);
xor (n443,n407,n408);
and (n444,n32,n95);
and (n445,n446,n447);
xor (n446,n443,n444);
or (n447,n448,n451);
and (n448,n449,n450);
xor (n449,n413,n414);
and (n450,n15,n95);
and (n451,n452,n453);
xor (n452,n449,n450);
or (n453,n454,n457);
and (n454,n455,n456);
xor (n455,n419,n420);
and (n456,n58,n95);
and (n457,n458,n459);
xor (n458,n455,n456);
or (n459,n460,n463);
and (n460,n461,n462);
xor (n461,n425,n426);
and (n462,n42,n95);
and (n463,n464,n465);
xor (n464,n461,n462);
and (n465,n466,n270);
xor (n466,n430,n431);
or (n467,n468,n470);
and (n468,n469,n86);
xor (n469,n440,n441);
and (n470,n471,n472);
xor (n471,n469,n86);
or (n472,n473,n475);
and (n473,n474,n203);
xor (n474,n446,n447);
and (n475,n476,n477);
xor (n476,n474,n203);
or (n477,n478,n481);
and (n478,n479,n480);
xor (n479,n452,n453);
and (n480,n58,n23);
and (n481,n482,n483);
xor (n482,n479,n480);
or (n483,n484,n487);
and (n484,n485,n486);
xor (n485,n458,n459);
and (n486,n42,n23);
and (n487,n488,n489);
xor (n488,n485,n486);
and (n489,n490,n491);
xor (n490,n464,n465);
and (n491,n67,n23);
and (n492,n32,n22);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n471,n472);
and (n496,n15,n22);
and (n497,n498,n499);
xor (n498,n495,n496);
or (n499,n500,n503);
and (n500,n501,n502);
xor (n501,n476,n477);
and (n502,n58,n22);
and (n503,n504,n505);
xor (n504,n501,n502);
or (n505,n506,n509);
and (n506,n507,n508);
xor (n507,n482,n483);
and (n508,n42,n22);
and (n509,n510,n511);
xor (n510,n507,n508);
and (n511,n512,n190);
xor (n512,n488,n489);
and (n513,n15,n13);
or (n514,n515,n518);
and (n515,n516,n517);
xor (n516,n498,n499);
and (n517,n58,n13);
and (n518,n519,n520);
xor (n519,n516,n517);
or (n520,n521,n524);
and (n521,n522,n523);
xor (n522,n504,n505);
and (n523,n42,n13);
and (n524,n525,n526);
xor (n525,n522,n523);
and (n526,n527,n528);
xor (n527,n510,n511);
and (n528,n67,n13);
and (n529,n58,n48);
or (n530,n531,n534);
and (n531,n532,n533);
xor (n532,n519,n520);
and (n533,n42,n48);
and (n534,n535,n536);
xor (n535,n532,n533);
and (n536,n537,n66);
xor (n537,n525,n526);
and (n538,n42,n40);
and (n539,n540,n541);
xor (n540,n535,n536);
and (n541,n67,n40);
and (n542,n67,n141);
or (n543,n544,n546,n577);
and (n544,n545,n71);
xor (n545,n540,n541);
and (n546,n71,n547);
or (n547,n548,n550,n576);
and (n548,n549,n109);
xor (n549,n537,n66);
and (n550,n109,n551);
or (n551,n552,n554,n575);
and (n552,n553,n185);
xor (n553,n527,n528);
and (n554,n185,n555);
or (n555,n556,n558,n574);
and (n556,n557,n262);
xor (n557,n512,n190);
and (n558,n262,n559);
or (n559,n560,n562,n573);
and (n560,n561,n266);
xor (n561,n490,n491);
and (n562,n266,n563);
or (n563,n564,n566,n572);
and (n564,n565,n328);
xor (n565,n466,n270);
and (n566,n328,n567);
or (n567,n568,n570,n571);
and (n568,n569,n332);
xor (n569,n432,n433);
and (n570,n332,n363);
and (n571,n569,n363);
and (n572,n565,n567);
and (n573,n561,n563);
and (n574,n557,n559);
and (n575,n553,n555);
and (n576,n549,n551);
and (n577,n545,n547);
endmodule
