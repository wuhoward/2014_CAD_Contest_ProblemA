module top (out,n18,n23,n25,n26,n28,n32,n35,n41,n59
        ,n73,n74,n75,n76,n77,n78,n79,n80,n84,n85
        ,n86,n90,n92,n94,n131,n133,n134,n135,n146,n147
        ,n148,n149,n161,n162,n163,n164,n177,n178,n179,n180
        ,n186,n188,n189,n192,n194,n197,n199,n200,n201,n281
        ,n387,n390,n392,n546,n548,n549,n552,n555,n556,n557
        ,n558,n561,n563,n567,n578,n579,n596,n599,n601,n602
        ,n604,n608,n614,n617,n619,n621,n625,n628,n630,n632
        ,n636,n639,n641,n643,n645,n653,n656,n658,n660,n664
        ,n667,n669,n671,n675,n678,n680,n682,n686,n689,n691
        ,n693,n701,n704,n706,n708,n712,n715,n717,n719,n723
        ,n726,n728,n730,n734,n737,n739,n741,n750,n753,n755
        ,n757,n771,n774,n776,n778,n797,n800,n802,n804,n813
        ,n816,n818,n820,n834,n837,n839,n841,n864,n867,n869
        ,n871,n887,n890,n892,n894,n939,n942,n944,n946,n950
        ,n953,n955,n957,n961,n964,n966,n968,n972,n975,n977
        ,n979,n987,n990,n992,n994,n998,n1001,n1003,n1005,n1009
        ,n1012,n1014,n1016,n1020,n1023,n1025,n1027,n1036,n1039,n1041
        ,n1043,n1048,n1051,n1053,n1055,n1065,n1068,n1070,n1072,n1090
        ,n1093,n1095,n1097,n1117,n1120,n1122,n1124,n1143,n1146,n1148
        ,n1150,n1172,n1175,n1177,n1179,n1191,n1194,n1196,n1198,n1230
        ,n1233,n1235,n1237,n1241,n1244,n1246,n1248,n1252,n1255,n1257
        ,n1259,n1263,n1266,n1268,n1270,n1291,n1294,n1296,n1298,n1305
        ,n1308,n1310,n1312,n1317,n1320,n1322,n1324,n1336,n1339,n1341
        ,n1343,n1352,n1355,n1357,n1359,n1369,n1372,n1374,n1376,n1384
        ,n1387,n1389,n1391,n1435,n1438,n1440,n1442,n1448,n1451,n1453
        ,n1455,n1465,n1468,n1470,n1472,n1501,n1504,n1506,n1508,n1620
        ,n1623,n1625,n1627,n1635,n1638,n1640,n1642,n1651,n1654,n1656
        ,n1658,n1667,n1670,n1672,n1674,n1682,n1685,n1687,n1689);
output out;
input n18;
input n23;
input n25;
input n26;
input n28;
input n32;
input n35;
input n41;
input n59;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n84;
input n85;
input n86;
input n90;
input n92;
input n94;
input n131;
input n133;
input n134;
input n135;
input n146;
input n147;
input n148;
input n149;
input n161;
input n162;
input n163;
input n164;
input n177;
input n178;
input n179;
input n180;
input n186;
input n188;
input n189;
input n192;
input n194;
input n197;
input n199;
input n200;
input n201;
input n281;
input n387;
input n390;
input n392;
input n546;
input n548;
input n549;
input n552;
input n555;
input n556;
input n557;
input n558;
input n561;
input n563;
input n567;
input n578;
input n579;
input n596;
input n599;
input n601;
input n602;
input n604;
input n608;
input n614;
input n617;
input n619;
input n621;
input n625;
input n628;
input n630;
input n632;
input n636;
input n639;
input n641;
input n643;
input n645;
input n653;
input n656;
input n658;
input n660;
input n664;
input n667;
input n669;
input n671;
input n675;
input n678;
input n680;
input n682;
input n686;
input n689;
input n691;
input n693;
input n701;
input n704;
input n706;
input n708;
input n712;
input n715;
input n717;
input n719;
input n723;
input n726;
input n728;
input n730;
input n734;
input n737;
input n739;
input n741;
input n750;
input n753;
input n755;
input n757;
input n771;
input n774;
input n776;
input n778;
input n797;
input n800;
input n802;
input n804;
input n813;
input n816;
input n818;
input n820;
input n834;
input n837;
input n839;
input n841;
input n864;
input n867;
input n869;
input n871;
input n887;
input n890;
input n892;
input n894;
input n939;
input n942;
input n944;
input n946;
input n950;
input n953;
input n955;
input n957;
input n961;
input n964;
input n966;
input n968;
input n972;
input n975;
input n977;
input n979;
input n987;
input n990;
input n992;
input n994;
input n998;
input n1001;
input n1003;
input n1005;
input n1009;
input n1012;
input n1014;
input n1016;
input n1020;
input n1023;
input n1025;
input n1027;
input n1036;
input n1039;
input n1041;
input n1043;
input n1048;
input n1051;
input n1053;
input n1055;
input n1065;
input n1068;
input n1070;
input n1072;
input n1090;
input n1093;
input n1095;
input n1097;
input n1117;
input n1120;
input n1122;
input n1124;
input n1143;
input n1146;
input n1148;
input n1150;
input n1172;
input n1175;
input n1177;
input n1179;
input n1191;
input n1194;
input n1196;
input n1198;
input n1230;
input n1233;
input n1235;
input n1237;
input n1241;
input n1244;
input n1246;
input n1248;
input n1252;
input n1255;
input n1257;
input n1259;
input n1263;
input n1266;
input n1268;
input n1270;
input n1291;
input n1294;
input n1296;
input n1298;
input n1305;
input n1308;
input n1310;
input n1312;
input n1317;
input n1320;
input n1322;
input n1324;
input n1336;
input n1339;
input n1341;
input n1343;
input n1352;
input n1355;
input n1357;
input n1359;
input n1369;
input n1372;
input n1374;
input n1376;
input n1384;
input n1387;
input n1389;
input n1391;
input n1435;
input n1438;
input n1440;
input n1442;
input n1448;
input n1451;
input n1453;
input n1455;
input n1465;
input n1468;
input n1470;
input n1472;
input n1501;
input n1504;
input n1506;
input n1508;
input n1620;
input n1623;
input n1625;
input n1627;
input n1635;
input n1638;
input n1640;
input n1642;
input n1651;
input n1654;
input n1656;
input n1658;
input n1667;
input n1670;
input n1672;
input n1674;
input n1682;
input n1685;
input n1687;
input n1689;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n20;
wire n21;
wire n22;
wire n24;
wire n27;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n81;
wire n82;
wire n83;
wire n87;
wire n88;
wire n89;
wire n91;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n190;
wire n191;
wire n193;
wire n195;
wire n196;
wire n198;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n388;
wire n389;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n547;
wire n550;
wire n551;
wire n553;
wire n554;
wire n559;
wire n560;
wire n562;
wire n564;
wire n565;
wire n566;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n597;
wire n598;
wire n600;
wire n603;
wire n605;
wire n606;
wire n607;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n615;
wire n616;
wire n618;
wire n620;
wire n622;
wire n623;
wire n624;
wire n626;
wire n627;
wire n629;
wire n631;
wire n633;
wire n634;
wire n635;
wire n637;
wire n638;
wire n640;
wire n642;
wire n644;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n654;
wire n655;
wire n657;
wire n659;
wire n661;
wire n662;
wire n663;
wire n665;
wire n666;
wire n668;
wire n670;
wire n672;
wire n673;
wire n674;
wire n676;
wire n677;
wire n679;
wire n681;
wire n683;
wire n684;
wire n685;
wire n687;
wire n688;
wire n690;
wire n692;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n702;
wire n703;
wire n705;
wire n707;
wire n709;
wire n710;
wire n711;
wire n713;
wire n714;
wire n716;
wire n718;
wire n720;
wire n721;
wire n722;
wire n724;
wire n725;
wire n727;
wire n729;
wire n731;
wire n732;
wire n733;
wire n735;
wire n736;
wire n738;
wire n740;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n751;
wire n752;
wire n754;
wire n756;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n772;
wire n773;
wire n775;
wire n777;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n798;
wire n799;
wire n801;
wire n803;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n814;
wire n815;
wire n817;
wire n819;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n835;
wire n836;
wire n838;
wire n840;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n868;
wire n870;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n888;
wire n889;
wire n891;
wire n893;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n940;
wire n941;
wire n943;
wire n945;
wire n947;
wire n948;
wire n949;
wire n951;
wire n952;
wire n954;
wire n956;
wire n958;
wire n959;
wire n960;
wire n962;
wire n963;
wire n965;
wire n967;
wire n969;
wire n970;
wire n971;
wire n973;
wire n974;
wire n976;
wire n978;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n988;
wire n989;
wire n991;
wire n993;
wire n995;
wire n996;
wire n997;
wire n999;
wire n1000;
wire n1002;
wire n1004;
wire n1006;
wire n1007;
wire n1008;
wire n1010;
wire n1011;
wire n1013;
wire n1015;
wire n1017;
wire n1018;
wire n1019;
wire n1021;
wire n1022;
wire n1024;
wire n1026;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1037;
wire n1038;
wire n1040;
wire n1042;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1049;
wire n1050;
wire n1052;
wire n1054;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1066;
wire n1067;
wire n1069;
wire n1071;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1091;
wire n1092;
wire n1094;
wire n1096;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1118;
wire n1119;
wire n1121;
wire n1123;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1144;
wire n1145;
wire n1147;
wire n1149;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1173;
wire n1174;
wire n1176;
wire n1178;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1192;
wire n1193;
wire n1195;
wire n1197;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1231;
wire n1232;
wire n1234;
wire n1236;
wire n1238;
wire n1239;
wire n1240;
wire n1242;
wire n1243;
wire n1245;
wire n1247;
wire n1249;
wire n1250;
wire n1251;
wire n1253;
wire n1254;
wire n1256;
wire n1258;
wire n1260;
wire n1261;
wire n1262;
wire n1264;
wire n1265;
wire n1267;
wire n1269;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1292;
wire n1293;
wire n1295;
wire n1297;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1306;
wire n1307;
wire n1309;
wire n1311;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1318;
wire n1319;
wire n1321;
wire n1323;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1337;
wire n1338;
wire n1340;
wire n1342;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1353;
wire n1354;
wire n1356;
wire n1358;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1370;
wire n1371;
wire n1373;
wire n1375;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1385;
wire n1386;
wire n1388;
wire n1390;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1436;
wire n1437;
wire n1439;
wire n1441;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1449;
wire n1450;
wire n1452;
wire n1454;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1466;
wire n1467;
wire n1469;
wire n1471;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1502;
wire n1503;
wire n1505;
wire n1507;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1621;
wire n1622;
wire n1624;
wire n1626;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1636;
wire n1637;
wire n1639;
wire n1641;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1652;
wire n1653;
wire n1655;
wire n1657;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1668;
wire n1669;
wire n1671;
wire n1673;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1683;
wire n1684;
wire n1686;
wire n1688;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
xnor (out,n0,n2743);
or (n0,n1,n2742);
and (n1,n2,n2286);
xor (n2,n3,n2215);
xor (n3,n4,n2153);
xor (n4,n5,n2122);
or (n5,n6,n2121);
and (n6,n7,n1946);
xor (n7,n8,n1902);
xor (n8,n9,n1779);
xor (n9,n10,n1277);
xor (n10,n11,n1272);
xor (n11,n12,n1029);
wire s0n12,s1n12,notn12;
or (n12,s0n12,s1n12);
not(notn12,n932);
and (s0n12,notn12,1'b0);
and (s1n12,n932,n14);
xor (n14,n15,n743);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n589);
and (s0n15,notn15,1'b0);
and (s1n15,n589,n16);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n572);
and (s0n16,notn16,n17);
and (s1n16,n572,n559);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n19);
and (s0n17,notn17,1'b0);
and (s1n17,n19,n18);
and (n19,n20,n553);
and (n20,n21,n37);
or (n21,n22,n27,n31,n34);
and (n22,n23,n24);
and (n24,n25,n26);
and (n27,n28,n29);
and (n29,n30,n26);
not (n30,n25);
and (n31,n32,n33);
nor (n33,n30,n26);
and (n34,n35,n36);
nor (n36,n25,n26);
and (n37,n38,n552);
not (n38,n39);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n551);
and (s0n39,notn39,n40);
and (s1n39,n551,1'b0);
wire s0n40,s1n40,notn40;
or (n40,s0n40,s1n40);
not(notn40,n181);
and (s0n40,notn40,n41);
and (s1n40,n181,n42);
wire s0n42,s1n42,notn42;
or (n42,s0n42,s1n42);
not(notn42,n544);
and (s0n42,notn42,n43);
and (s1n42,n544,n518);
or (n43,n44,n486,n517,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n44,n45,n485);
or (n45,n46,n484);
or (n46,n47,n483);
or (n47,n48,n481);
or (n48,n49,n480);
or (n49,n50,n478);
or (n50,n51,n476);
nor (n51,n52,n401,n410,n422,n434,n445,n456,n467);
or (n52,1'b0,n53,n395,n399);
and (n53,n54,n394);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n385);
and (s0n54,notn54,n55);
and (s1n54,n385,n293);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n252);
and (s0n55,notn55,1'b0);
and (s1n55,n252,n56);
or (n56,n57,n233,n237,n241,n244,n247,n249,1'b0);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n206,n217,n227);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n95);
and (s0n61,notn61,n62);
and (s1n61,n95,1'b0);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n93);
and (s0n62,notn62,n63);
and (s1n62,n93,n91);
wire s0n63,s1n63,notn63;
or (n63,s0n63,s1n63);
not(notn63,n87);
and (s0n63,notn63,n64);
and (s1n63,n87,n81);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n80);
and (s0n64,notn64,n65);
and (s1n64,n80,1'b0);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n79);
and (s0n65,notn65,n66);
and (s1n65,n79,1'b1);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n78);
and (s0n66,notn66,n67);
and (s1n66,n78,1'b0);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n77);
and (s0n67,notn67,n68);
and (s1n67,n77,1'b1);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n76);
and (s0n68,notn68,n69);
and (s1n68,n76,1'b0);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n75);
and (s0n69,notn69,n70);
and (s1n69,n75,1'b1);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n74);
and (s0n70,notn70,n71);
and (s1n70,n74,1'b0);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n73);
and (s0n71,notn71,n58);
and (s1n71,n73,1'b1);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n86);
and (s0n81,notn81,n82);
and (s1n81,n86,1'b0);
wire s0n82,s1n82,notn82;
or (n82,s0n82,s1n82);
not(notn82,n85);
and (s0n82,notn82,n83);
and (s1n82,n85,1'b1);
not (n83,n84);
or (n87,n88,n90);
or (n88,n89,n84);
or (n89,n86,n85);
not (n91,n92);
or (n93,n92,n94);
not (n95,n96);
or (n96,n97,n204);
or (n97,n98,n202);
or (n98,n99,n196);
or (n99,n100,n195);
or (n100,n101,n191);
or (n101,n102,n190);
or (n102,n103,n185);
or (n103,n104,n184);
or (n104,n105,n183);
or (n105,n106,n181);
or (n106,n107,n175);
or (n107,n108,n174);
or (n108,n109,n173);
or (n109,n110,n172);
or (n110,n111,n171);
or (n111,n112,n170);
or (n112,n113,n169);
or (n113,n114,n168);
or (n114,n115,n165);
or (n115,n116,n159);
or (n116,n117,n158);
or (n117,n118,n157);
or (n118,n119,n156);
or (n119,n120,n155);
or (n120,n121,n154);
or (n121,n122,n152);
or (n122,n123,n150);
or (n123,n124,n144);
or (n124,n125,n143);
or (n125,n126,n142);
or (n126,n127,n141);
or (n127,n128,n140);
or (n128,n129,n138);
or (n129,n130,n136);
nor (n130,n131,n132,n134,n135);
not (n132,n133);
nor (n136,n131,n132,n137,n135);
not (n137,n134);
and (n138,n131,n133,n134,n139);
not (n139,n135);
and (n140,n131,n132,n134,n139);
nor (n141,n131,n133,n137,n135);
and (n142,n131,n132,n134,n135);
and (n143,n131,n133,n134,n135);
nor (n144,n145,n147,n148,n149);
not (n145,n146);
nor (n150,n145,n151,n148,n149);
not (n151,n147);
and (n152,n145,n147,n148,n153);
not (n153,n149);
and (n154,n146,n147,n148,n153);
and (n155,n146,n151,n148,n153);
and (n156,n145,n151,n148,n149);
and (n157,n146,n151,n148,n149);
and (n158,n146,n147,n148,n149);
nor (n159,n160,n162,n163,n164);
not (n160,n161);
and (n165,n161,n162,n166,n167);
not (n166,n163);
not (n167,n164);
and (n168,n160,n162,n166,n167);
and (n169,n161,n162,n163,n167);
nor (n170,n161,n162,n166,n167);
and (n171,n160,n162,n163,n164);
and (n172,n160,n162,n166,n164);
and (n173,n161,n162,n166,n164);
nor (n174,n160,n162,n163,n167);
nor (n175,n176,n178,n179,n180);
not (n176,n177);
nor (n181,n177,n182,n179,n180);
not (n182,n178);
and (n183,n176,n182,n179,n180);
and (n184,n177,n182,n179,n180);
nor (n185,n186,n187,n189);
not (n187,n188);
and (n190,n186,n188,n189);
and (n191,n192,n193);
not (n193,n194);
nor (n195,n192,n193);
nor (n196,n197,n198,n200,n201);
not (n198,n199);
and (n202,n197,n199,n200,n203);
not (n203,n201);
and (n204,n205,n198,n200,n203);
not (n205,n197);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n95);
and (s0n206,notn206,n207);
and (s1n206,n95,1'b0);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n93);
and (s0n207,notn207,n208);
and (s1n207,n93,1'b0);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n87);
and (s0n208,notn208,n209);
and (s1n208,n87,n89);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n80);
and (s0n209,notn209,n210);
and (s1n209,n80,1'b1);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n79);
and (s0n210,notn210,n211);
and (s1n210,n79,1'b1);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n78);
and (s0n211,notn211,n212);
and (s1n211,n78,1'b0);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n77);
and (s0n212,notn212,n213);
and (s1n212,n77,1'b0);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n76);
and (s0n213,notn213,n214);
and (s1n213,n76,1'b1);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n75);
and (s0n214,notn214,n215);
and (s1n214,n75,1'b1);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n74);
and (s0n215,notn215,n216);
and (s1n215,n74,1'b0);
not (n216,n73);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n95);
and (s0n217,notn217,n218);
and (s1n217,n95,1'b0);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n93);
and (s0n218,notn218,n219);
and (s1n218,n93,1'b0);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n87);
and (s0n219,notn219,n220);
and (s1n219,n87,n226);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n80);
and (s0n220,notn220,n221);
and (s1n220,n80,1'b1);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n79);
and (s0n221,notn221,n222);
and (s1n221,n79,1'b1);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n78);
and (s0n222,notn222,n223);
and (s1n222,n78,1'b0);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n77);
and (s0n223,notn223,n224);
and (s1n223,n77,1'b0);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n76);
and (s0n224,notn224,n225);
and (s1n224,n76,1'b0);
not (n225,n75);
not (n226,n89);
not (n227,n228);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n95);
and (s0n228,notn228,n229);
and (s1n228,n95,1'b0);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n93);
and (s0n229,notn229,n230);
and (s1n229,n93,1'b0);
wire s0n230,s1n230,notn230;
or (n230,s0n230,s1n230);
not(notn230,n87);
and (s0n230,notn230,n231);
and (s1n230,n87,1'b0);
wire s0n231,s1n231,notn231;
or (n231,s0n231,s1n231);
not(notn231,n80);
and (s0n231,notn231,n232);
and (s1n231,n80,1'b0);
not (n232,n79);
and (n233,n234,n235);
not (n234,n74);
and (n235,n236,n206,n217,n227);
not (n236,n61);
and (n237,n238,n239);
not (n238,n76);
and (n239,n61,n240,n217,n227);
not (n240,n206);
and (n241,n242,n243);
not (n242,n78);
and (n243,n236,n240,n217,n227);
and (n244,n245,n246);
not (n245,n80);
nor (n246,n236,n240,n217,n228);
and (n247,n83,n248);
nor (n248,n61,n240,n217,n228);
and (n249,n250,n251);
not (n250,n86);
nor (n251,n236,n206,n217,n228);
or (n252,n253,n282);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n280);
and (s0n253,notn253,n254);
and (s1n253,n280,1'b0);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n279);
and (s0n254,notn254,n255);
and (s1n254,n279,n274);
wire s0n255,s1n255,notn255;
or (n255,s0n255,s1n255);
not(notn255,n273);
and (s0n255,notn255,n256);
and (s1n255,n273,n262);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n261);
and (s0n256,notn256,n257);
and (s1n256,n261,n124);
or (n257,n258,n155);
or (n258,n259,n154);
or (n259,n260,n152);
or (n260,n144,n150);
or (n261,n131,n133,n134,n135);
or (n262,1'b0,1'b0,n263,n269,n271);
and (n263,n264,n267);
or (n264,1'b0,1'b0,n265,n185);
and (n265,n266,n188,n189);
not (n266,n186);
and (n267,n176,n182,n179,n268);
not (n268,n180);
and (n269,n192,n270);
and (n270,n177,n182,n179,n268);
or (n271,n272,n183);
or (n272,n175,n181);
or (n273,n177,n178,n179,n180);
or (n274,n275,n174);
or (n275,n276,n172);
or (n276,n277,n169);
or (n277,n278,n168);
or (n278,n159,n165);
or (n279,n161,n162,n163,n164);
not (n280,n281);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n280);
and (s0n282,notn282,n283);
and (s1n282,n280,1'b0);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n279);
and (s0n283,notn283,n284);
and (s1n283,n279,n292);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n273);
and (s0n284,notn284,n285);
and (s1n284,n273,n288);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n261);
and (s0n285,notn285,n286);
and (s1n285,n261,1'b0);
or (n286,n287,n158);
or (n287,n156,n157);
or (n288,1'b0,n184,n289,n291,1'b0);
and (n289,n290,n267);
or (n290,1'b0,n190,n265,1'b0);
and (n291,n194,n270);
or (n292,n171,n173);
not (n293,n294);
nor (n294,n55,n295,n311,n331,n348,n362,n373,n381);
wire s0n295,s1n295,notn295;
or (n295,s0n295,s1n295);
not(notn295,n252);
and (s0n295,notn295,1'b0);
and (s1n295,n252,n296);
or (n296,n297,n299,n301,n303,n305,n307,n309,1'b0);
and (n297,n298,n60);
xnor (n298,n73,n59);
and (n299,n300,n235);
xnor (n300,n75,n74);
and (n301,n302,n239);
xnor (n302,n77,n76);
and (n303,n304,n243);
xnor (n304,n79,n78);
and (n305,n306,n246);
xnor (n306,n90,n80);
and (n307,n308,n248);
xnor (n308,n85,n84);
and (n309,n310,n251);
xnor (n310,n94,n86);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n252);
and (s0n311,notn311,1'b0);
and (s1n311,n252,n312);
or (n312,n313,n316,n319,n322,n325,n328,1'b0,1'b0);
and (n313,n314,n60);
xnor (n314,n74,n315);
or (n315,n73,n59);
and (n316,n317,n235);
xnor (n317,n76,n318);
or (n318,n75,n74);
and (n319,n320,n239);
xnor (n320,n78,n321);
or (n321,n77,n76);
and (n322,n323,n243);
xnor (n323,n80,n324);
or (n324,n79,n78);
and (n325,n326,n246);
xnor (n326,n84,n327);
or (n327,n90,n80);
and (n328,n329,n248);
xnor (n329,n86,n330);
or (n330,n85,n84);
wire s0n331,s1n331,notn331;
or (n331,s0n331,s1n331);
not(notn331,n252);
and (s0n331,notn331,1'b0);
and (s1n331,n252,n332);
or (n332,n333,n336,n339,n342,n345,1'b0,1'b0,1'b0);
and (n333,n334,n60);
xnor (n334,n75,n335);
or (n335,n74,n315);
and (n336,n337,n235);
xnor (n337,n77,n338);
or (n338,n76,n318);
and (n339,n340,n239);
xnor (n340,n79,n341);
or (n341,n78,n321);
and (n342,n343,n243);
xnor (n343,n90,n344);
or (n344,n80,n324);
and (n345,n346,n246);
xnor (n346,n85,n347);
or (n347,n84,n327);
wire s0n348,s1n348,notn348;
or (n348,s0n348,s1n348);
not(notn348,n252);
and (s0n348,notn348,1'b0);
and (s1n348,n252,n349);
or (n349,n350,n353,n356,n359,1'b0,1'b0,1'b0,1'b0);
and (n350,n351,n60);
xnor (n351,n76,n352);
or (n352,n75,n335);
and (n353,n354,n235);
xnor (n354,n78,n355);
or (n355,n77,n338);
and (n356,n357,n239);
xnor (n357,n80,n358);
or (n358,n79,n341);
and (n359,n360,n243);
xnor (n360,n84,n361);
or (n361,n90,n344);
wire s0n362,s1n362,notn362;
or (n362,s0n362,s1n362);
not(notn362,n252);
and (s0n362,notn362,1'b0);
and (s1n362,n252,n363);
or (n363,n364,n367,n370,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n364,n365,n60);
xnor (n365,n77,n366);
or (n366,n76,n352);
and (n367,n368,n235);
xnor (n368,n79,n369);
or (n369,n78,n355);
and (n370,n371,n239);
xnor (n371,n90,n372);
or (n372,n80,n358);
wire s0n373,s1n373,notn373;
or (n373,s0n373,s1n373);
not(notn373,n252);
and (s0n373,notn373,1'b0);
and (s1n373,n252,n374);
or (n374,n375,n378,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n375,n376,n60);
xnor (n376,n78,n377);
or (n377,n77,n366);
and (n378,n379,n235);
xnor (n379,n80,n380);
or (n380,n79,n369);
wire s0n381,s1n381,notn381;
or (n381,s0n381,s1n381);
not(notn381,n252);
and (s0n381,notn381,1'b0);
and (s1n381,n252,n382);
and (n382,n383,n60);
xnor (n383,n79,n384);
or (n384,n78,n377);
nor (n385,n386,n388,n391);
not (n386,n387);
not (n388,n389);
xor (n389,n390,n387);
xor (n391,n392,n393);
and (n393,n390,n387);
and (n394,n253,n282);
and (n395,n396,n397);
xor (n396,n295,n55);
nor (n397,n253,n398);
not (n398,n282);
and (n399,n55,n400);
and (n400,n253,n398);
not (n401,n402);
or (n402,1'b0,n403,n405,n409);
and (n403,n404,n394);
wire s0n404,s1n404,notn404;
or (n404,s0n404,s1n404);
not(notn404,n385);
and (s0n404,notn404,n295);
and (s1n404,n385,1'b0);
and (n405,n406,n397);
xor (n406,n407,n408);
not (n407,n311);
not (n408,n295);
and (n409,n295,n400);
or (n410,1'b0,n411,n413,n421);
and (n411,n412,n394);
wire s0n412,s1n412,notn412;
or (n412,s0n412,s1n412);
not(notn412,n385);
and (s0n412,notn412,n311);
and (s1n412,n385,1'b0);
and (n413,n414,n397);
wire s0n414,s1n414,notn414;
or (n414,s0n414,s1n414);
not(notn414,n55);
and (s0n414,notn414,n415);
and (s1n414,n55,n418);
xor (n415,n416,n417);
not (n416,n331);
and (n417,n407,n408);
xor (n418,n331,n419);
and (n419,n311,n420);
and (n420,n295,n55);
and (n421,n311,n400);
not (n422,n423);
or (n423,1'b0,n424,n426,n433);
and (n424,n425,n394);
wire s0n425,s1n425,notn425;
or (n425,s0n425,s1n425);
not(notn425,n385);
and (s0n425,notn425,n331);
and (s1n425,n385,1'b0);
and (n426,n427,n397);
wire s0n427,s1n427,notn427;
or (n427,s0n427,s1n427);
not(notn427,n55);
and (s0n427,notn427,n428);
and (s1n427,n55,n431);
xor (n428,n429,n430);
not (n429,n348);
and (n430,n416,n417);
xor (n431,n348,n432);
and (n432,n331,n419);
and (n433,n331,n400);
or (n434,1'b0,n435,n437,n444);
and (n435,n436,n394);
wire s0n436,s1n436,notn436;
or (n436,s0n436,s1n436);
not(notn436,n385);
and (s0n436,notn436,n348);
and (s1n436,n385,1'b0);
and (n437,n438,n397);
wire s0n438,s1n438,notn438;
or (n438,s0n438,s1n438);
not(notn438,n55);
and (s0n438,notn438,n439);
and (s1n438,n55,n442);
xor (n439,n440,n441);
not (n440,n362);
and (n441,n429,n430);
xor (n442,n362,n443);
and (n443,n348,n432);
and (n444,n348,n400);
or (n445,1'b0,n446,n448,n455);
and (n446,n447,n394);
wire s0n447,s1n447,notn447;
or (n447,s0n447,s1n447);
not(notn447,n385);
and (s0n447,notn447,n362);
and (s1n447,n385,1'b0);
and (n448,n449,n397);
wire s0n449,s1n449,notn449;
or (n449,s0n449,s1n449);
not(notn449,n55);
and (s0n449,notn449,n450);
and (s1n449,n55,n453);
xor (n450,n451,n452);
not (n451,n373);
and (n452,n440,n441);
xor (n453,n373,n454);
and (n454,n362,n443);
and (n455,n362,n400);
or (n456,1'b0,n457,n459,n466);
and (n457,n458,n394);
wire s0n458,s1n458,notn458;
or (n458,s0n458,s1n458);
not(notn458,n385);
and (s0n458,notn458,n373);
and (s1n458,n385,1'b0);
and (n459,n460,n397);
wire s0n460,s1n460,notn460;
or (n460,s0n460,s1n460);
not(notn460,n55);
and (s0n460,notn460,n461);
and (s1n460,n55,n464);
xor (n461,n462,n463);
not (n462,n381);
and (n463,n451,n452);
xor (n464,n381,n465);
and (n465,n373,n454);
and (n466,n373,n400);
or (n467,1'b0,n468,n470,n475);
and (n468,n469,n394);
wire s0n469,s1n469,notn469;
or (n469,s0n469,s1n469);
not(notn469,n385);
and (s0n469,notn469,n381);
and (s1n469,n385,1'b0);
and (n470,n471,n397);
wire s0n471,s1n471,notn471;
or (n471,s0n471,s1n471);
not(notn471,n55);
and (s0n471,notn471,n472);
and (s1n471,n55,n474);
not (n472,n473);
and (n473,n462,n463);
and (n474,n381,n465);
and (n475,n381,n400);
nor (n476,n477,n401,n410,n422,n434,n445,n456,n467);
not (n477,n52);
nor (n478,n52,n402,n479,n422,n434,n445,n456,n467);
not (n479,n410);
nor (n480,n477,n402,n479,n422,n434,n445,n456,n467);
nor (n481,n52,n401,n479,n423,n482,n445,n456,n467);
not (n482,n434);
nor (n483,n477,n401,n479,n423,n482,n445,n456,n467);
nor (n484,n52,n402,n410,n422,n482,n445,n456,n467);
nor (n485,n477,n402,n410,n422,n482,n445,n456,n467);
or (n486,n487,n502);
or (n487,n488,n501);
or (n488,n489,n500);
or (n489,n490,n499);
or (n490,n491,n498);
or (n491,n492,n497);
or (n492,n493,n496);
or (n493,n494,n495);
nor (n494,n52,n401,n479,n423,n434,n445,n456,n467);
nor (n495,n477,n401,n479,n423,n434,n445,n456,n467);
nor (n496,n52,n402,n410,n422,n434,n445,n456,n467);
nor (n497,n477,n402,n410,n422,n434,n445,n456,n467);
nor (n498,n52,n401,n410,n423,n482,n445,n456,n467);
nor (n499,n477,n401,n410,n423,n482,n445,n456,n467);
nor (n500,n52,n402,n479,n423,n482,n445,n456,n467);
nor (n501,n477,n402,n479,n423,n482,n445,n456,n467);
or (n502,n503,n516);
or (n503,n504,n515);
or (n504,n505,n514);
or (n505,n506,n513);
or (n506,n507,n512);
or (n507,n508,n511);
or (n508,n509,n510);
nor (n509,n52,n401,n479,n422,n434,n445,n456,n467);
nor (n510,n477,n401,n479,n422,n434,n445,n456,n467);
nor (n511,n52,n402,n410,n423,n482,n445,n456,n467);
nor (n512,n477,n402,n410,n423,n482,n445,n456,n467);
nor (n513,n52,n401,n410,n422,n482,n445,n456,n467);
nor (n514,n477,n401,n410,n422,n482,n445,n456,n467);
nor (n515,n52,n402,n479,n422,n482,n445,n456,n467);
nor (n516,n477,n402,n479,n422,n482,n445,n456,n467);
nor (n517,n477,n402,n479,n423,n434,n445,n456,n467);
or (n518,1'b0,n519,n526,n533,n294);
or (n519,n520,n484);
or (n520,n521,n483);
or (n521,n522,n481);
or (n522,n523,n501);
or (n523,n524,n478);
or (n524,n525,n476);
or (n525,n497,n51);
or (n526,n527,n500);
or (n527,n528,n499);
or (n528,n529,n498);
or (n529,n530,n512);
or (n530,n531,n496);
or (n531,n532,n495);
or (n532,n517,n494);
or (n533,n534,n511);
or (n534,n535,n510);
or (n535,n536,n509);
or (n536,n537,n480);
or (n537,n538,n543);
or (n538,n539,n542);
or (n539,n540,n541);
nor (n540,n477,n402,n410,n423,n434,n445,n456,n467);
nor (n541,n52,n401,n410,n423,n434,n445,n456,n467);
nor (n542,n477,n401,n410,n423,n434,n445,n456,n467);
nor (n543,n52,n402,n479,n423,n434,n445,n456,n467);
or (n544,n545,n550);
nor (n545,n546,n547,n549);
not (n547,n548);
and (n550,n546,n548,n549);
nor (n551,n176,n182,n179,n180);
nor (n553,n554,n556,n557,n558);
not (n554,n555);
or (n559,1'b0,n560,n562,n566,n569);
and (n560,n561,n553);
and (n562,n563,n564);
nor (n564,n555,n565,n557,n558);
not (n565,n556);
and (n566,n567,n568);
nor (n568,n554,n565,n557,n558);
and (n569,n18,n570);
and (n570,n554,n565,n557,n571);
not (n571,n558);
and (n572,n37,n573);
not (n573,n574);
wire s0n574,s1n574,notn574;
or (n574,s0n574,s1n574);
not(notn574,n587);
and (s0n574,notn574,n20);
and (s1n574,n587,n575);
or (n575,n576,n580,n583,n585);
and (n576,n23,n577);
and (n577,n578,n579);
and (n580,n28,n581);
and (n581,n582,n579);
not (n582,n578);
and (n583,n32,n584);
nor (n584,n582,n579);
and (n585,n35,n586);
nor (n586,n578,n579);
and (n587,n38,n588);
not (n588,n552);
and (n589,n590,n646);
not (n590,n591);
wire s0n591,s1n591,notn591;
or (n591,s0n591,s1n591);
not(notn591,n37);
and (s0n591,notn591,1'b0);
and (s1n591,n37,n592);
wire s0n592,s1n592,notn592;
or (n592,s0n592,s1n592);
not(notn592,n645);
and (s0n592,notn592,n593);
and (s1n592,n645,n636);
or (n593,n594,n612,n623,n634);
and (n594,n595,n24);
wire s0n595,s1n595,notn595;
or (n595,s0n595,s1n595);
not(notn595,n574);
and (s0n595,notn595,n596);
and (s1n595,n574,n597);
or (n597,n598,n603,n607,n610);
and (n598,n599,n600);
nor (n600,n601,n602);
and (n603,n604,n605);
nor (n605,n606,n602);
not (n606,n601);
and (n607,n608,n609);
and (n609,n606,n602);
and (n610,n596,n611);
and (n611,n601,n602);
and (n612,n613,n29);
wire s0n613,s1n613,notn613;
or (n613,s0n613,s1n613);
not(notn613,n574);
and (s0n613,notn613,n614);
and (s1n613,n574,n615);
or (n615,n616,n618,n620,n622);
and (n616,n617,n600);
and (n618,n619,n605);
and (n620,n621,n609);
and (n622,n614,n611);
and (n623,n624,n33);
wire s0n624,s1n624,notn624;
or (n624,s0n624,s1n624);
not(notn624,n574);
and (s0n624,notn624,n625);
and (s1n624,n574,n626);
or (n626,n627,n629,n631,n633);
and (n627,n628,n600);
and (n629,n630,n605);
and (n631,n632,n609);
and (n633,n625,n611);
and (n634,n635,n36);
wire s0n635,s1n635,notn635;
or (n635,s0n635,s1n635);
not(notn635,n574);
and (s0n635,notn635,n636);
and (s1n635,n574,n637);
or (n637,n638,n640,n642,n644);
and (n638,n639,n600);
and (n640,n641,n605);
and (n642,n643,n609);
and (n644,n636,n611);
and (n646,n647,n695);
not (n647,n648);
wire s0n648,s1n648,notn648;
or (n648,s0n648,s1n648);
not(notn648,n37);
and (s0n648,notn648,1'b0);
and (s1n648,n37,n649);
wire s0n649,s1n649,notn649;
or (n649,s0n649,s1n649);
not(notn649,n645);
and (s0n649,notn649,n650);
and (s1n649,n645,n686);
or (n650,n651,n662,n673,n684);
and (n651,n652,n24);
wire s0n652,s1n652,notn652;
or (n652,s0n652,s1n652);
not(notn652,n574);
and (s0n652,notn652,n653);
and (s1n652,n574,n654);
or (n654,n655,n657,n659,n661);
and (n655,n656,n600);
and (n657,n658,n605);
and (n659,n660,n609);
and (n661,n653,n611);
and (n662,n663,n29);
wire s0n663,s1n663,notn663;
or (n663,s0n663,s1n663);
not(notn663,n574);
and (s0n663,notn663,n664);
and (s1n663,n574,n665);
or (n665,n666,n668,n670,n672);
and (n666,n667,n600);
and (n668,n669,n605);
and (n670,n671,n609);
and (n672,n664,n611);
and (n673,n674,n33);
wire s0n674,s1n674,notn674;
or (n674,s0n674,s1n674);
not(notn674,n574);
and (s0n674,notn674,n675);
and (s1n674,n574,n676);
or (n676,n677,n679,n681,n683);
and (n677,n678,n600);
and (n679,n680,n605);
and (n681,n682,n609);
and (n683,n675,n611);
and (n684,n685,n36);
wire s0n685,s1n685,notn685;
or (n685,s0n685,s1n685);
not(notn685,n574);
and (s0n685,notn685,n686);
and (s1n685,n574,n687);
or (n687,n688,n690,n692,n694);
and (n688,n689,n600);
and (n690,n691,n605);
and (n692,n693,n609);
and (n694,n686,n611);
not (n695,n696);
wire s0n696,s1n696,notn696;
or (n696,s0n696,s1n696);
not(notn696,n37);
and (s0n696,notn696,1'b0);
and (s1n696,n37,n697);
wire s0n697,s1n697,notn697;
or (n697,s0n697,s1n697);
not(notn697,n645);
and (s0n697,notn697,n698);
and (s1n697,n645,n734);
or (n698,n699,n710,n721,n732);
and (n699,n700,n24);
wire s0n700,s1n700,notn700;
or (n700,s0n700,s1n700);
not(notn700,n574);
and (s0n700,notn700,n701);
and (s1n700,n574,n702);
or (n702,n703,n705,n707,n709);
and (n703,n704,n600);
and (n705,n706,n605);
and (n707,n708,n609);
and (n709,n701,n611);
and (n710,n711,n29);
wire s0n711,s1n711,notn711;
or (n711,s0n711,s1n711);
not(notn711,n574);
and (s0n711,notn711,n712);
and (s1n711,n574,n713);
or (n713,n714,n716,n718,n720);
and (n714,n715,n600);
and (n716,n717,n605);
and (n718,n719,n609);
and (n720,n712,n611);
and (n721,n722,n33);
wire s0n722,s1n722,notn722;
or (n722,s0n722,s1n722);
not(notn722,n574);
and (s0n722,notn722,n723);
and (s1n722,n574,n724);
or (n724,n725,n727,n729,n731);
and (n725,n726,n600);
and (n727,n728,n605);
and (n729,n730,n609);
and (n731,n723,n611);
and (n732,n733,n36);
wire s0n733,s1n733,notn733;
or (n733,s0n733,s1n733);
not(notn733,n574);
and (s0n733,notn733,n734);
and (s1n733,n574,n735);
or (n735,n736,n738,n740,n742);
and (n736,n737,n600);
and (n738,n739,n605);
and (n740,n741,n609);
and (n742,n734,n611);
or (n743,n744,n783);
and (n744,n745,n784);
xor (n745,n746,n761);
xor (n746,n747,n759);
wire s0n747,s1n747,notn747;
or (n747,s0n747,s1n747);
not(notn747,n589);
and (s0n747,notn747,1'b0);
and (s1n747,n589,n748);
wire s0n748,s1n748,notn748;
or (n748,s0n748,s1n748);
not(notn748,n572);
and (s0n748,notn748,n749);
and (s1n748,n572,n751);
wire s0n749,s1n749,notn749;
or (n749,s0n749,s1n749);
not(notn749,n19);
and (s0n749,notn749,1'b0);
and (s1n749,n19,n750);
or (n751,1'b0,n752,n754,n756,n758);
and (n752,n753,n553);
and (n754,n755,n564);
and (n756,n757,n568);
and (n758,n750,n570);
wire s0n759,s1n759,notn759;
or (n759,s0n759,s1n759);
not(notn759,n760);
and (s0n759,notn759,1'b0);
and (s1n759,n760,n16);
xor (n760,n590,n646);
or (n761,n762,n783);
and (n762,n763,n780);
xor (n763,n764,n765);
wire s0n764,s1n764,notn764;
or (n764,s0n764,s1n764);
not(notn764,n760);
and (s0n764,notn764,1'b0);
and (s1n764,n760,n748);
xor (n765,n766,n768);
wire s0n766,s1n766,notn766;
or (n766,s0n766,s1n766);
not(notn766,n767);
and (s0n766,notn766,1'b0);
and (s1n766,n767,n16);
xor (n767,n647,n695);
wire s0n768,s1n768,notn768;
or (n768,s0n768,s1n768);
not(notn768,n589);
and (s0n768,notn768,1'b0);
and (s1n768,n589,n769);
wire s0n769,s1n769,notn769;
or (n769,s0n769,s1n769);
not(notn769,n572);
and (s0n769,notn769,n770);
and (s1n769,n572,n772);
wire s0n770,s1n770,notn770;
or (n770,s0n770,s1n770);
not(notn770,n19);
and (s0n770,notn770,1'b0);
and (s1n770,n19,n771);
or (n772,1'b0,n773,n775,n777,n779);
and (n773,n774,n553);
and (n775,n776,n564);
and (n777,n778,n568);
and (n779,n771,n570);
and (n780,n781,n782);
wire s0n781,s1n781,notn781;
or (n781,s0n781,s1n781);
not(notn781,n767);
and (s0n781,notn781,1'b0);
and (s1n781,n767,n748);
wire s0n782,s1n782,notn782;
or (n782,s0n782,s1n782);
not(notn782,n696);
and (s0n782,notn782,1'b0);
and (s1n782,n696,n16);
and (n783,n764,n765);
nand (n784,n785,n931);
or (n785,n786,n926);
nor (n786,n787,n925);
and (n787,n788,n914);
nand (n788,n789,n913);
or (n789,n790,n847);
not (n790,n791);
or (n791,n792,n825);
xor (n792,n793,n822);
xor (n793,n794,n806);
wire s0n794,s1n794,notn794;
or (n794,s0n794,s1n794);
not(notn794,n760);
and (s0n794,notn794,1'b0);
and (s1n794,n760,n795);
wire s0n795,s1n795,notn795;
or (n795,s0n795,s1n795);
not(notn795,n572);
and (s0n795,notn795,n796);
and (s1n795,n572,n798);
wire s0n796,s1n796,notn796;
or (n796,s0n796,s1n796);
not(notn796,n19);
and (s0n796,notn796,1'b0);
and (s1n796,n19,n797);
or (n798,1'b0,n799,n801,n803,n805);
and (n799,n800,n553);
and (n801,n802,n564);
and (n803,n804,n568);
and (n805,n797,n570);
xor (n806,n807,n810);
xor (n807,n808,n809);
wire s0n808,s1n808,notn808;
or (n808,s0n808,s1n808);
not(notn808,n767);
and (s0n808,notn808,1'b0);
and (s1n808,n767,n769);
wire s0n809,s1n809,notn809;
or (n809,s0n809,s1n809);
not(notn809,n696);
and (s0n809,notn809,1'b0);
and (s1n809,n696,n748);
wire s0n810,s1n810,notn810;
or (n810,s0n810,s1n810);
not(notn810,n589);
and (s0n810,notn810,1'b0);
and (s1n810,n589,n811);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n572);
and (s0n811,notn811,n812);
and (s1n811,n572,n814);
wire s0n812,s1n812,notn812;
or (n812,s0n812,s1n812);
not(notn812,n19);
and (s0n812,notn812,1'b0);
and (s1n812,n19,n813);
or (n814,1'b0,n815,n817,n819,n821);
and (n815,n816,n553);
and (n817,n818,n564);
and (n819,n820,n568);
and (n821,n813,n570);
and (n822,n823,n824);
wire s0n823,s1n823,notn823;
or (n823,s0n823,s1n823);
not(notn823,n767);
and (s0n823,notn823,1'b0);
and (s1n823,n767,n795);
wire s0n824,s1n824,notn824;
or (n824,s0n824,s1n824);
not(notn824,n696);
and (s0n824,notn824,1'b0);
and (s1n824,n696,n769);
or (n825,n826,n846);
and (n826,n827,n843);
xor (n827,n828,n829);
wire s0n828,s1n828,notn828;
or (n828,s0n828,s1n828);
not(notn828,n760);
and (s0n828,notn828,1'b0);
and (s1n828,n760,n811);
xor (n829,n830,n831);
xor (n830,n823,n824);
wire s0n831,s1n831,notn831;
or (n831,s0n831,s1n831);
not(notn831,n589);
and (s0n831,notn831,1'b0);
and (s1n831,n589,n832);
wire s0n832,s1n832,notn832;
or (n832,s0n832,s1n832);
not(notn832,n572);
and (s0n832,notn832,n833);
and (s1n832,n572,n835);
wire s0n833,s1n833,notn833;
or (n833,s0n833,s1n833);
not(notn833,n19);
and (s0n833,notn833,1'b0);
and (s1n833,n19,n834);
or (n835,1'b0,n836,n838,n840,n842);
and (n836,n837,n553);
and (n838,n839,n564);
and (n840,n841,n568);
and (n842,n834,n570);
and (n843,n844,n845);
wire s0n844,s1n844,notn844;
or (n844,s0n844,s1n844);
not(notn844,n767);
and (s0n844,notn844,1'b0);
and (s1n844,n767,n811);
wire s0n845,s1n845,notn845;
or (n845,s0n845,s1n845);
not(notn845,n696);
and (s0n845,notn845,1'b0);
and (s1n845,n696,n795);
and (n846,n828,n829);
not (n847,n848);
nand (n848,n849,n909,n912);
nand (n849,n850,n874,n906);
or (n850,n851,n852);
xor (n851,n827,n843);
or (n852,n853,n873);
and (n853,n854,n859);
xor (n854,n855,n856);
wire s0n855,s1n855,notn855;
or (n855,s0n855,s1n855);
not(notn855,n760);
and (s0n855,notn855,1'b0);
and (s1n855,n760,n832);
and (n856,n857,n858);
wire s0n857,s1n857,notn857;
or (n857,s0n857,s1n857);
not(notn857,n767);
and (s0n857,notn857,1'b0);
and (s1n857,n767,n832);
wire s0n858,s1n858,notn858;
or (n858,s0n858,s1n858);
not(notn858,n696);
and (s0n858,notn858,1'b0);
and (s1n858,n696,n811);
xor (n859,n860,n861);
xor (n860,n844,n845);
wire s0n861,s1n861,notn861;
or (n861,s0n861,s1n861);
not(notn861,n589);
and (s0n861,notn861,1'b0);
and (s1n861,n589,n862);
wire s0n862,s1n862,notn862;
or (n862,s0n862,s1n862);
not(notn862,n572);
and (s0n862,notn862,n863);
and (s1n862,n572,n865);
wire s0n863,s1n863,notn863;
or (n863,s0n863,s1n863);
not(notn863,n19);
and (s0n863,notn863,1'b0);
and (s1n863,n19,n864);
or (n865,1'b0,n866,n868,n870,n872);
and (n866,n867,n553);
and (n868,n869,n564);
and (n870,n871,n568);
and (n872,n864,n570);
and (n873,n855,n856);
or (n874,n875,n905);
and (n875,n876,n900);
xor (n876,n877,n880);
and (n877,n878,n879);
wire s0n878,s1n878,notn878;
or (n878,s0n878,s1n878);
not(notn878,n767);
and (s0n878,notn878,1'b0);
and (s1n878,n767,n862);
wire s0n879,s1n879,notn879;
or (n879,s0n879,s1n879);
not(notn879,n696);
and (s0n879,notn879,1'b0);
and (s1n879,n696,n832);
or (n880,n881,n899);
and (n881,n882,n898);
xor (n882,n883,n897);
and (n883,n884,n896);
wire s0n884,s1n884,notn884;
or (n884,s0n884,s1n884);
not(notn884,n767);
and (s0n884,notn884,1'b0);
and (s1n884,n767,n885);
wire s0n885,s1n885,notn885;
or (n885,s0n885,s1n885);
not(notn885,n572);
and (s0n885,notn885,n886);
and (s1n885,n572,n888);
wire s0n886,s1n886,notn886;
or (n886,s0n886,s1n886);
not(notn886,n19);
and (s0n886,notn886,1'b0);
and (s1n886,n19,n887);
or (n888,1'b0,n889,n891,n893,n895);
and (n889,n890,n553);
and (n891,n892,n564);
and (n893,n894,n568);
and (n895,n887,n570);
wire s0n896,s1n896,notn896;
or (n896,s0n896,s1n896);
not(notn896,n696);
and (s0n896,notn896,1'b0);
and (s1n896,n696,n862);
wire s0n897,s1n897,notn897;
or (n897,s0n897,s1n897);
not(notn897,n760);
and (s0n897,notn897,1'b0);
and (s1n897,n760,n885);
xor (n898,n878,n879);
and (n899,n883,n897);
xor (n900,n901,n904);
xor (n901,n902,n903);
wire s0n902,s1n902,notn902;
or (n902,s0n902,s1n902);
not(notn902,n589);
and (s0n902,notn902,1'b0);
and (s1n902,n589,n885);
xor (n903,n857,n858);
wire s0n904,s1n904,notn904;
or (n904,s0n904,s1n904);
not(notn904,n760);
and (s0n904,notn904,1'b0);
and (s1n904,n760,n862);
and (n905,n877,n880);
or (n906,n907,n908);
xor (n907,n854,n859);
and (n908,n901,n904);
nand (n909,n910,n850);
not (n910,n911);
nand (n911,n907,n908);
nand (n912,n851,n852);
nand (n913,n792,n825);
or (n914,n915,n922);
xor (n915,n916,n921);
xor (n916,n917,n918);
wire s0n917,s1n917,notn917;
or (n917,s0n917,s1n917);
not(notn917,n760);
and (s0n917,notn917,1'b0);
and (s1n917,n760,n769);
xor (n918,n919,n920);
xor (n919,n781,n782);
wire s0n920,s1n920,notn920;
or (n920,s0n920,s1n920);
not(notn920,n589);
and (s0n920,notn920,1'b0);
and (s1n920,n589,n795);
and (n921,n808,n809);
or (n922,n923,n924);
and (n923,n793,n822);
and (n924,n794,n806);
and (n925,n915,n922);
nor (n926,n927,n930);
or (n927,n928,n929);
and (n928,n916,n921);
and (n929,n917,n918);
xor (n930,n763,n780);
nand (n931,n927,n930);
xor (n932,n933,n981);
not (n933,n934);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n37);
and (s0n934,notn934,1'b0);
and (s1n934,n37,n935);
wire s0n935,s1n935,notn935;
or (n935,s0n935,s1n935);
not(notn935,n645);
and (s0n935,notn935,n936);
and (s1n935,n645,n972);
or (n936,n937,n948,n959,n970);
and (n937,n938,n24);
wire s0n938,s1n938,notn938;
or (n938,s0n938,s1n938);
not(notn938,n574);
and (s0n938,notn938,n939);
and (s1n938,n574,n940);
or (n940,n941,n943,n945,n947);
and (n941,n942,n600);
and (n943,n944,n605);
and (n945,n946,n609);
and (n947,n939,n611);
and (n948,n949,n29);
wire s0n949,s1n949,notn949;
or (n949,s0n949,s1n949);
not(notn949,n574);
and (s0n949,notn949,n950);
and (s1n949,n574,n951);
or (n951,n952,n954,n956,n958);
and (n952,n953,n600);
and (n954,n955,n605);
and (n956,n957,n609);
and (n958,n950,n611);
and (n959,n960,n33);
wire s0n960,s1n960,notn960;
or (n960,s0n960,s1n960);
not(notn960,n574);
and (s0n960,notn960,n961);
and (s1n960,n574,n962);
or (n962,n963,n965,n967,n969);
and (n963,n964,n600);
and (n965,n966,n605);
and (n967,n968,n609);
and (n969,n961,n611);
and (n970,n971,n36);
wire s0n971,s1n971,notn971;
or (n971,s0n971,s1n971);
not(notn971,n574);
and (s0n971,notn971,n972);
and (s1n971,n574,n973);
or (n973,n974,n976,n978,n980);
and (n974,n975,n600);
and (n976,n977,n605);
and (n978,n979,n609);
and (n980,n972,n611);
not (n981,n982);
wire s0n982,s1n982,notn982;
or (n982,s0n982,s1n982);
not(notn982,n37);
and (s0n982,notn982,1'b0);
and (s1n982,n37,n983);
wire s0n983,s1n983,notn983;
or (n983,s0n983,s1n983);
not(notn983,n645);
and (s0n983,notn983,n984);
and (s1n983,n645,n1020);
or (n984,n985,n996,n1007,n1018);
and (n985,n986,n24);
wire s0n986,s1n986,notn986;
or (n986,s0n986,s1n986);
not(notn986,n574);
and (s0n986,notn986,n987);
and (s1n986,n574,n988);
or (n988,n989,n991,n993,n995);
and (n989,n990,n600);
and (n991,n992,n605);
and (n993,n994,n609);
and (n995,n987,n611);
and (n996,n997,n29);
wire s0n997,s1n997,notn997;
or (n997,s0n997,s1n997);
not(notn997,n574);
and (s0n997,notn997,n998);
and (s1n997,n574,n999);
or (n999,n1000,n1002,n1004,n1006);
and (n1000,n1001,n600);
and (n1002,n1003,n605);
and (n1004,n1005,n609);
and (n1006,n998,n611);
and (n1007,n1008,n33);
wire s0n1008,s1n1008,notn1008;
or (n1008,s0n1008,s1n1008);
not(notn1008,n574);
and (s0n1008,notn1008,n1009);
and (s1n1008,n574,n1010);
or (n1010,n1011,n1013,n1015,n1017);
and (n1011,n1012,n600);
and (n1013,n1014,n605);
and (n1015,n1016,n609);
and (n1017,n1009,n611);
and (n1018,n1019,n36);
wire s0n1019,s1n1019,notn1019;
or (n1019,s0n1019,s1n1019);
not(notn1019,n574);
and (s0n1019,notn1019,n1020);
and (s1n1019,n574,n1021);
or (n1021,n1022,n1024,n1026,n1028);
and (n1022,n1023,n600);
and (n1024,n1025,n605);
and (n1026,n1027,n609);
and (n1028,n1020,n611);
and (n1029,n1030,n1225);
xor (n1030,n1031,n1079);
xor (n1031,n1032,n1057);
xor (n1032,n1033,n1045);
and (n1033,n760,n1034);
wire s0n1034,s1n1034,notn1034;
or (n1034,s0n1034,s1n1034);
not(notn1034,n572);
and (s0n1034,notn1034,n1035);
and (s1n1034,n572,n1037);
wire s0n1035,s1n1035,notn1035;
or (n1035,s0n1035,s1n1035);
not(notn1035,n19);
and (s0n1035,notn1035,1'b0);
and (s1n1035,n19,n1036);
or (n1037,1'b0,n1038,n1040,n1042,n1044);
and (n1038,n1039,n553);
and (n1040,n1041,n564);
and (n1042,n1043,n568);
and (n1044,n1036,n570);
and (n1045,n589,n1046);
wire s0n1046,s1n1046,notn1046;
or (n1046,s0n1046,s1n1046);
not(notn1046,n572);
and (s0n1046,notn1046,n1047);
and (s1n1046,n572,n1049);
wire s0n1047,s1n1047,notn1047;
or (n1047,s0n1047,s1n1047);
not(notn1047,n19);
and (s0n1047,notn1047,1'b0);
and (s1n1047,n19,n1048);
or (n1049,1'b0,n1050,n1052,n1054,n1056);
and (n1050,n1051,n553);
and (n1052,n1053,n564);
and (n1054,n1055,n568);
and (n1056,n1048,n570);
or (n1057,n1058,n1078);
and (n1058,n1059,n1075);
xor (n1059,n1060,n1074);
xor (n1060,n1061,n1062);
and (n1061,n767,n1034);
and (n1062,n589,n1063);
wire s0n1063,s1n1063,notn1063;
or (n1063,s0n1063,s1n1063);
not(notn1063,n572);
and (s0n1063,notn1063,n1064);
and (s1n1063,n572,n1066);
wire s0n1064,s1n1064,notn1064;
or (n1064,s0n1064,s1n1064);
not(notn1064,n19);
and (s0n1064,notn1064,1'b0);
and (s1n1064,n19,n1065);
or (n1066,1'b0,n1067,n1069,n1071,n1073);
and (n1067,n1068,n553);
and (n1069,n1070,n564);
and (n1071,n1072,n568);
and (n1073,n1065,n570);
and (n1074,n760,n1046);
and (n1075,n1076,n1077);
and (n1076,n767,n1046);
wire s0n1077,s1n1077,notn1077;
or (n1077,s0n1077,s1n1077);
not(notn1077,n696);
and (s0n1077,notn1077,1'b0);
and (s1n1077,n696,n1034);
and (n1078,n1060,n1074);
or (n1079,n1080,n1224);
and (n1080,n1081,n1105);
xor (n1081,n1082,n1104);
or (n1082,n1083,n1103);
and (n1083,n1084,n1100);
xor (n1084,n1085,n1099);
xor (n1085,n1086,n1087);
xor (n1086,n1076,n1077);
and (n1087,n589,n1088);
wire s0n1088,s1n1088,notn1088;
or (n1088,s0n1088,s1n1088);
not(notn1088,n572);
and (s0n1088,notn1088,n1089);
and (s1n1088,n572,n1091);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n19);
and (s0n1089,notn1089,1'b0);
and (s1n1089,n19,n1090);
or (n1091,1'b0,n1092,n1094,n1096,n1098);
and (n1092,n1093,n553);
and (n1094,n1095,n564);
and (n1096,n1097,n568);
and (n1098,n1090,n570);
and (n1099,n760,n1063);
and (n1100,n1101,n1102);
wire s0n1101,s1n1101,notn1101;
or (n1101,s0n1101,s1n1101);
not(notn1101,n696);
and (s0n1101,notn1101,1'b0);
and (s1n1101,n696,n1046);
and (n1102,n767,n1063);
and (n1103,n1085,n1099);
xor (n1104,n1059,n1075);
or (n1105,n1106,n1223);
and (n1106,n1107,n1131);
xor (n1107,n1108,n1130);
or (n1108,n1109,n1129);
and (n1109,n1110,n1126);
xor (n1110,n1111,n1112);
and (n1111,n760,n1088);
xor (n1112,n1113,n1114);
xor (n1113,n1101,n1102);
and (n1114,n589,n1115);
wire s0n1115,s1n1115,notn1115;
or (n1115,s0n1115,s1n1115);
not(notn1115,n572);
and (s0n1115,notn1115,n1116);
and (s1n1115,n572,n1118);
wire s0n1116,s1n1116,notn1116;
or (n1116,s0n1116,s1n1116);
not(notn1116,n19);
and (s0n1116,notn1116,1'b0);
and (s1n1116,n19,n1117);
or (n1118,1'b0,n1119,n1121,n1123,n1125);
and (n1119,n1120,n553);
and (n1121,n1122,n564);
and (n1123,n1124,n568);
and (n1125,n1117,n570);
and (n1126,n1127,n1128);
wire s0n1127,s1n1127,notn1127;
or (n1127,s0n1127,s1n1127);
not(notn1127,n696);
and (s0n1127,notn1127,1'b0);
and (s1n1127,n696,n1063);
and (n1128,n767,n1088);
and (n1129,n1111,n1112);
xor (n1130,n1084,n1100);
or (n1131,n1132,n1222);
and (n1132,n1133,n1157);
xor (n1133,n1134,n1156);
or (n1134,n1135,n1155);
and (n1135,n1136,n1152);
xor (n1136,n1137,n1138);
and (n1137,n760,n1115);
xor (n1138,n1139,n1140);
xor (n1139,n1127,n1128);
and (n1140,n589,n1141);
wire s0n1141,s1n1141,notn1141;
or (n1141,s0n1141,s1n1141);
not(notn1141,n572);
and (s0n1141,notn1141,n1142);
and (s1n1141,n572,n1144);
wire s0n1142,s1n1142,notn1142;
or (n1142,s0n1142,s1n1142);
not(notn1142,n19);
and (s0n1142,notn1142,1'b0);
and (s1n1142,n19,n1143);
or (n1144,1'b0,n1145,n1147,n1149,n1151);
and (n1145,n1146,n553);
and (n1147,n1148,n564);
and (n1149,n1150,n568);
and (n1151,n1143,n570);
and (n1152,n1153,n1154);
and (n1153,n767,n1115);
wire s0n1154,s1n1154,notn1154;
or (n1154,s0n1154,s1n1154);
not(notn1154,n696);
and (s0n1154,notn1154,1'b0);
and (s1n1154,n696,n1088);
and (n1155,n1137,n1138);
xor (n1156,n1110,n1126);
or (n1157,n1158,n1221);
and (n1158,n1159,n1183);
xor (n1159,n1160,n1182);
or (n1160,n1161,n1181);
and (n1161,n1162,n1167);
xor (n1162,n1163,n1164);
and (n1163,n760,n1141);
and (n1164,n1165,n1166);
wire s0n1165,s1n1165,notn1165;
or (n1165,s0n1165,s1n1165);
not(notn1165,n696);
and (s0n1165,notn1165,1'b0);
and (s1n1165,n696,n1115);
and (n1166,n767,n1141);
xor (n1167,n1168,n1169);
xor (n1168,n1153,n1154);
and (n1169,n589,n1170);
wire s0n1170,s1n1170,notn1170;
or (n1170,s0n1170,s1n1170);
not(notn1170,n572);
and (s0n1170,notn1170,n1171);
and (s1n1170,n572,n1173);
wire s0n1171,s1n1171,notn1171;
or (n1171,s0n1171,s1n1171);
not(notn1171,n19);
and (s0n1171,notn1171,1'b0);
and (s1n1171,n19,n1172);
or (n1173,1'b0,n1174,n1176,n1178,n1180);
and (n1174,n1175,n553);
and (n1176,n1177,n564);
and (n1178,n1179,n568);
and (n1180,n1172,n570);
and (n1181,n1163,n1164);
xor (n1182,n1136,n1152);
or (n1183,n1184,n1220);
and (n1184,n1185,n1203);
xor (n1185,n1186,n1202);
and (n1186,n1187,n1201);
xor (n1187,n1188,n1200);
and (n1188,n589,n1189);
wire s0n1189,s1n1189,notn1189;
or (n1189,s0n1189,s1n1189);
not(notn1189,n572);
and (s0n1189,notn1189,n1190);
and (s1n1189,n572,n1192);
wire s0n1190,s1n1190,notn1190;
or (n1190,s0n1190,s1n1190);
not(notn1190,n19);
and (s0n1190,notn1190,1'b0);
and (s1n1190,n19,n1191);
or (n1192,1'b0,n1193,n1195,n1197,n1199);
and (n1193,n1194,n553);
and (n1195,n1196,n564);
and (n1197,n1198,n568);
and (n1199,n1191,n570);
and (n1200,n760,n1170);
xor (n1201,n1165,n1166);
xor (n1202,n1162,n1167);
or (n1203,n1204,n1219);
and (n1204,n1205,n1218);
xor (n1205,n1206,n1209);
and (n1206,n1207,n1208);
wire s0n1207,s1n1207,notn1207;
or (n1207,s0n1207,s1n1207);
not(notn1207,n696);
and (s0n1207,notn1207,1'b0);
and (s1n1207,n696,n1141);
and (n1208,n767,n1170);
or (n1209,n1210,n1217);
and (n1210,n1211,n1216);
xor (n1211,n1212,n1215);
and (n1212,n1213,n1214);
and (n1213,n767,n1189);
wire s0n1214,s1n1214,notn1214;
or (n1214,s0n1214,s1n1214);
not(notn1214,n696);
and (s0n1214,notn1214,1'b0);
and (s1n1214,n696,n1170);
xor (n1215,n1207,n1208);
and (n1216,n760,n1189);
and (n1217,n1212,n1215);
xor (n1218,n1187,n1201);
and (n1219,n1206,n1209);
and (n1220,n1186,n1202);
and (n1221,n1160,n1182);
and (n1222,n1134,n1156);
and (n1223,n1108,n1130);
and (n1224,n1082,n1104);
wire s0n1225,s1n1225,notn1225;
or (n1225,s0n1225,s1n1225);
not(notn1225,n37);
and (s0n1225,notn1225,1'b0);
and (s1n1225,n37,n1226);
wire s0n1226,s1n1226,notn1226;
or (n1226,s0n1226,s1n1226);
not(notn1226,n645);
and (s0n1226,notn1226,n1227);
and (s1n1226,n645,n1263);
or (n1227,n1228,n1239,n1250,n1261);
and (n1228,n1229,n24);
wire s0n1229,s1n1229,notn1229;
or (n1229,s0n1229,s1n1229);
not(notn1229,n574);
and (s0n1229,notn1229,n1230);
and (s1n1229,n574,n1231);
or (n1231,n1232,n1234,n1236,n1238);
and (n1232,n1233,n600);
and (n1234,n1235,n605);
and (n1236,n1237,n609);
and (n1238,n1230,n611);
and (n1239,n1240,n29);
wire s0n1240,s1n1240,notn1240;
or (n1240,s0n1240,s1n1240);
not(notn1240,n574);
and (s0n1240,notn1240,n1241);
and (s1n1240,n574,n1242);
or (n1242,n1243,n1245,n1247,n1249);
and (n1243,n1244,n600);
and (n1245,n1246,n605);
and (n1247,n1248,n609);
and (n1249,n1241,n611);
and (n1250,n1251,n33);
wire s0n1251,s1n1251,notn1251;
or (n1251,s0n1251,s1n1251);
not(notn1251,n574);
and (s0n1251,notn1251,n1252);
and (s1n1251,n574,n1253);
or (n1253,n1254,n1256,n1258,n1260);
and (n1254,n1255,n600);
and (n1256,n1257,n605);
and (n1258,n1259,n609);
and (n1260,n1252,n611);
and (n1261,n1262,n36);
wire s0n1262,s1n1262,notn1262;
or (n1262,s0n1262,s1n1262);
not(notn1262,n574);
and (s0n1262,notn1262,n1263);
and (s1n1262,n574,n1264);
or (n1264,n1265,n1267,n1269,n1271);
and (n1265,n1266,n600);
and (n1267,n1268,n605);
and (n1269,n1270,n609);
and (n1271,n1263,n611);
and (n1272,n1273,n1274);
xor (n1273,n745,n784);
xor (n1274,n1275,n1276);
not (n1275,n1225);
and (n1276,n933,n981);
xor (n1277,n1278,n1769);
xor (n1278,n1279,n1735);
or (n1279,n1280,n1734);
and (n1280,n1281,n1603);
xor (n1281,n1282,n1590);
and (n1282,n1283,n1516);
xor (n1283,n1284,n1426);
wire s0n1284,s1n1284,notn1284;
or (n1284,s0n1284,s1n1284);
not(notn1284,n1425);
and (s0n1284,notn1284,1'b0);
and (s1n1284,n1425,n1285);
xor (n1285,n1286,n1396);
xor (n1286,n1287,n1300);
not (n1287,n1288);
nand (n1288,n591,n1289);
wire s0n1289,s1n1289,notn1289;
or (n1289,s0n1289,s1n1289);
not(notn1289,n572);
and (s0n1289,notn1289,n1290);
and (s1n1289,n572,n1292);
wire s0n1290,s1n1290,notn1290;
or (n1290,s0n1290,s1n1290);
not(notn1290,n19);
and (s0n1290,notn1290,1'b0);
and (s1n1290,n19,n1291);
or (n1292,1'b0,n1293,n1295,n1297,n1299);
and (n1293,n1294,n553);
and (n1295,n1296,n564);
and (n1297,n1298,n568);
and (n1299,n1291,n570);
xor (n1300,n1301,n1326);
xor (n1301,n1302,n1314);
wire s0n1302,s1n1302,notn1302;
or (n1302,s0n1302,s1n1302);
not(notn1302,n648);
and (s0n1302,notn1302,1'b0);
and (s1n1302,n648,n1303);
wire s0n1303,s1n1303,notn1303;
or (n1303,s0n1303,s1n1303);
not(notn1303,n572);
and (s0n1303,notn1303,n1304);
and (s1n1303,n572,n1306);
wire s0n1304,s1n1304,notn1304;
or (n1304,s0n1304,s1n1304);
not(notn1304,n19);
and (s0n1304,notn1304,1'b0);
and (s1n1304,n19,n1305);
or (n1306,1'b0,n1307,n1309,n1311,n1313);
and (n1307,n1308,n553);
and (n1309,n1310,n564);
and (n1311,n1312,n568);
and (n1313,n1305,n570);
wire s0n1314,s1n1314,notn1314;
or (n1314,s0n1314,s1n1314);
not(notn1314,n696);
and (s0n1314,notn1314,1'b0);
and (s1n1314,n696,n1315);
wire s0n1315,s1n1315,notn1315;
or (n1315,s0n1315,s1n1315);
not(notn1315,n572);
and (s0n1315,notn1315,n1316);
and (s1n1315,n572,n1318);
wire s0n1316,s1n1316,notn1316;
or (n1316,s0n1316,s1n1316);
not(notn1316,n19);
and (s0n1316,notn1316,1'b0);
and (s1n1316,n19,n1317);
or (n1318,1'b0,n1319,n1321,n1323,n1325);
and (n1319,n1320,n553);
and (n1321,n1322,n564);
and (n1323,n1324,n568);
and (n1325,n1317,n570);
or (n1326,n1327,n1330,n1395);
and (n1327,n1328,n1329);
wire s0n1328,s1n1328,notn1328;
or (n1328,s0n1328,s1n1328);
not(notn1328,n648);
and (s0n1328,notn1328,1'b0);
and (s1n1328,n648,n1289);
wire s0n1329,s1n1329,notn1329;
or (n1329,s0n1329,s1n1329);
not(notn1329,n696);
and (s0n1329,notn1329,1'b0);
and (s1n1329,n696,n1303);
and (n1330,n1329,n1331);
or (n1331,n1332,n1346,n1394);
and (n1332,n1333,n1345);
wire s0n1333,s1n1333,notn1333;
or (n1333,s0n1333,s1n1333);
not(notn1333,n648);
and (s0n1333,notn1333,1'b0);
and (s1n1333,n648,n1334);
wire s0n1334,s1n1334,notn1334;
or (n1334,s0n1334,s1n1334);
not(notn1334,n572);
and (s0n1334,notn1334,n1335);
and (s1n1334,n572,n1337);
wire s0n1335,s1n1335,notn1335;
or (n1335,s0n1335,s1n1335);
not(notn1335,n19);
and (s0n1335,notn1335,1'b0);
and (s1n1335,n19,n1336);
or (n1337,1'b0,n1338,n1340,n1342,n1344);
and (n1338,n1339,n553);
and (n1340,n1341,n564);
and (n1342,n1343,n568);
and (n1344,n1336,n570);
wire s0n1345,s1n1345,notn1345;
or (n1345,s0n1345,s1n1345);
not(notn1345,n696);
and (s0n1345,notn1345,1'b0);
and (s1n1345,n696,n1289);
and (n1346,n1345,n1347);
or (n1347,n1348,n1362,n1364);
and (n1348,n1349,n1361);
wire s0n1349,s1n1349,notn1349;
or (n1349,s0n1349,s1n1349);
not(notn1349,n648);
and (s0n1349,notn1349,1'b0);
and (s1n1349,n648,n1350);
wire s0n1350,s1n1350,notn1350;
or (n1350,s0n1350,s1n1350);
not(notn1350,n572);
and (s0n1350,notn1350,n1351);
and (s1n1350,n572,n1353);
wire s0n1351,s1n1351,notn1351;
or (n1351,s0n1351,s1n1351);
not(notn1351,n19);
and (s0n1351,notn1351,1'b0);
and (s1n1351,n19,n1352);
or (n1353,1'b0,n1354,n1356,n1358,n1360);
and (n1354,n1355,n553);
and (n1356,n1357,n564);
and (n1358,n1359,n568);
and (n1360,n1352,n570);
wire s0n1361,s1n1361,notn1361;
or (n1361,s0n1361,s1n1361);
not(notn1361,n696);
and (s0n1361,notn1361,1'b0);
and (s1n1361,n696,n1334);
and (n1362,n1361,n1363);
or (n1363,n1364,n1379,n1380);
and (n1364,n1365,n1378);
not (n1365,n1366);
nand (n1366,n648,n1367);
wire s0n1367,s1n1367,notn1367;
or (n1367,s0n1367,s1n1367);
not(notn1367,n572);
and (s0n1367,notn1367,n1368);
and (s1n1367,n572,n1370);
wire s0n1368,s1n1368,notn1368;
or (n1368,s0n1368,s1n1368);
not(notn1368,n19);
and (s0n1368,notn1368,1'b0);
and (s1n1368,n19,n1369);
or (n1370,1'b0,n1371,n1373,n1375,n1377);
and (n1371,n1372,n553);
and (n1373,n1374,n564);
and (n1375,n1376,n568);
and (n1377,n1369,n570);
wire s0n1378,s1n1378,notn1378;
or (n1378,s0n1378,s1n1378);
not(notn1378,n696);
and (s0n1378,notn1378,1'b0);
and (s1n1378,n696,n1350);
and (n1379,n1378,n1380);
and (n1380,n1381,n1393);
wire s0n1381,s1n1381,notn1381;
or (n1381,s0n1381,s1n1381);
not(notn1381,n648);
and (s0n1381,notn1381,1'b0);
and (s1n1381,n648,n1382);
wire s0n1382,s1n1382,notn1382;
or (n1382,s0n1382,s1n1382);
not(notn1382,n572);
and (s0n1382,notn1382,n1383);
and (s1n1382,n572,n1385);
wire s0n1383,s1n1383,notn1383;
or (n1383,s0n1383,s1n1383);
not(notn1383,n19);
and (s0n1383,notn1383,1'b0);
and (s1n1383,n19,n1384);
or (n1385,1'b0,n1386,n1388,n1390,n1392);
and (n1386,n1387,n553);
and (n1388,n1389,n564);
and (n1390,n1391,n568);
and (n1392,n1384,n570);
wire s0n1393,s1n1393,notn1393;
or (n1393,s0n1393,s1n1393);
not(notn1393,n696);
and (s0n1393,notn1393,1'b0);
and (s1n1393,n696,n1367);
and (n1394,n1333,n1347);
and (n1395,n1328,n1331);
or (n1396,n1397,n1402,n1424);
and (n1397,n1398,n1400);
not (n1398,n1399);
nand (n1399,n591,n1334);
xor (n1400,n1401,n1331);
xor (n1401,n1328,n1329);
and (n1402,n1400,n1403);
or (n1403,n1404,n1409,n1423);
and (n1404,n1405,n1407);
not (n1405,n1406);
nand (n1406,n591,n1350);
xor (n1407,n1408,n1347);
xor (n1408,n1333,n1345);
and (n1409,n1407,n1410);
or (n1410,n1411,n1416,n1422);
and (n1411,n1412,n1414);
not (n1412,n1413);
nand (n1413,n591,n1367);
xor (n1414,n1415,n1363);
xor (n1415,n1349,n1361);
and (n1416,n1414,n1417);
and (n1417,n1418,n1420);
not (n1418,n1419);
nand (n1419,n591,n1382);
xor (n1420,n1421,n1380);
xor (n1421,n1365,n1378);
and (n1422,n1412,n1417);
and (n1423,n1405,n1410);
and (n1424,n1398,n1403);
and (n1425,n1275,n1276);
xor (n1426,n1427,n1474);
xor (n1427,n1428,n1459);
xor (n1428,n1429,n1457);
xor (n1429,n1430,n1444);
nor (n1430,n1431,n981);
not (n1431,n1432);
wire s0n1432,s1n1432,notn1432;
or (n1432,s0n1432,s1n1432);
not(notn1432,n591);
and (s0n1432,notn1432,1'b0);
and (s1n1432,n591,n1433);
wire s0n1433,s1n1433,notn1433;
or (n1433,s0n1433,s1n1433);
not(notn1433,n572);
and (s0n1433,notn1433,n1434);
and (s1n1433,n572,n1436);
wire s0n1434,s1n1434,notn1434;
or (n1434,s0n1434,s1n1434);
not(notn1434,n19);
and (s0n1434,notn1434,1'b0);
and (s1n1434,n19,n1435);
or (n1436,1'b0,n1437,n1439,n1441,n1443);
and (n1437,n1438,n553);
and (n1439,n1440,n564);
and (n1441,n1442,n568);
and (n1443,n1435,n570);
and (n1444,n1445,n982);
and (n1445,n591,n1446);
wire s0n1446,s1n1446,notn1446;
or (n1446,s0n1446,s1n1446);
not(notn1446,n572);
and (s0n1446,notn1446,n1447);
and (s1n1446,n572,n1449);
wire s0n1447,s1n1447,notn1447;
or (n1447,s0n1447,s1n1447);
not(notn1447,n19);
and (s0n1447,notn1447,1'b0);
and (s1n1447,n19,n1448);
or (n1449,1'b0,n1450,n1452,n1454,n1456);
and (n1450,n1451,n553);
and (n1452,n1453,n564);
and (n1454,n1455,n568);
and (n1456,n1448,n570);
and (n1457,n1444,n1458);
wire s0n1458,s1n1458,notn1458;
or (n1458,s0n1458,s1n1458);
not(notn1458,n648);
and (s0n1458,notn1458,1'b0);
and (s1n1458,n648,n1315);
and (n1459,n1430,n1460);
not (n1460,n1461);
not (n1461,n1462);
wire s0n1462,s1n1462,notn1462;
or (n1462,s0n1462,s1n1462);
not(notn1462,n648);
and (s0n1462,notn1462,1'b0);
and (s1n1462,n648,n1463);
wire s0n1463,s1n1463,notn1463;
or (n1463,s0n1463,s1n1463);
not(notn1463,n572);
and (s0n1463,notn1463,n1464);
and (s1n1463,n572,n1466);
wire s0n1464,s1n1464,notn1464;
or (n1464,s0n1464,s1n1464);
not(notn1464,n19);
and (s0n1464,notn1464,1'b0);
and (s1n1464,n19,n1465);
or (n1466,1'b0,n1467,n1469,n1471,n1473);
and (n1467,n1468,n553);
and (n1469,n1470,n564);
and (n1471,n1472,n568);
and (n1473,n1465,n570);
or (n1474,n1475,n1515);
and (n1475,n1476,n1493);
xor (n1476,n1477,n1484);
nor (n1477,n1478,n981);
xnor (n1478,n1479,n1482);
not (n1479,n1480);
not (n1480,n1481);
nand (n1481,n591,n1315);
not (n1482,n1483);
wire s0n1483,s1n1483,notn1483;
or (n1483,s0n1483,s1n1483);
not(notn1483,n648);
and (s0n1483,notn1483,1'b0);
and (s1n1483,n648,n1446);
and (n1484,n1485,n982);
nand (n1485,n1486,n1492);
or (n1486,n1487,n1489);
not (n1487,n1488);
wire s0n1488,s1n1488,notn1488;
or (n1488,s0n1488,s1n1488);
not(notn1488,n648);
and (s0n1488,notn1488,1'b0);
and (s1n1488,n648,n1433);
not (n1489,n1490);
not (n1490,n1491);
wire s0n1491,s1n1491,notn1491;
or (n1491,s0n1491,s1n1491);
not(notn1491,n591);
and (s0n1491,notn1491,1'b0);
and (s1n1491,n591,n1463);
or (n1492,n1490,n1488);
and (n1493,n1494,n982);
or (n1494,n1495,n1512);
nor (n1495,n1496,n1461);
and (n1496,n1497,n1510);
not (n1497,n1498);
wire s0n1498,s1n1498,notn1498;
or (n1498,s0n1498,s1n1498);
not(notn1498,n591);
and (s0n1498,notn1498,1'b0);
and (s1n1498,n591,n1499);
wire s0n1499,s1n1499,notn1499;
or (n1499,s0n1499,s1n1499);
not(notn1499,n572);
and (s0n1499,notn1499,n1500);
and (s1n1499,n572,n1502);
wire s0n1500,s1n1500,notn1500;
or (n1500,s0n1500,s1n1500);
not(notn1500,n19);
and (s0n1500,notn1500,1'b0);
and (s1n1500,n19,n1501);
or (n1502,1'b0,n1503,n1505,n1507,n1509);
and (n1503,n1504,n553);
and (n1505,n1506,n564);
and (n1507,n1508,n568);
and (n1509,n1501,n570);
not (n1510,n1511);
wire s0n1511,s1n1511,notn1511;
or (n1511,s0n1511,s1n1511);
not(notn1511,n696);
and (s0n1511,notn1511,1'b0);
and (s1n1511,n696,n1433);
nor (n1512,n1513,n1431);
not (n1513,n1514);
wire s0n1514,s1n1514,notn1514;
or (n1514,s0n1514,s1n1514);
not(notn1514,n696);
and (s0n1514,notn1514,1'b0);
and (s1n1514,n696,n1499);
and (n1515,n1477,n1484);
and (n1516,n1517,n1274);
xor (n1517,n1518,n1535);
xor (n1518,n1519,n1528);
nor (n1519,n1520,n1525);
and (n1520,n1521,n1458);
xor (n1521,n1522,n1524);
not (n1522,n1523);
wire s0n1523,s1n1523,notn1523;
or (n1523,s0n1523,s1n1523);
not(notn1523,n696);
and (s0n1523,notn1523,1'b0);
and (s1n1523,n696,n1446);
nand (n1524,n591,n1303);
and (n1525,n1526,n1527);
not (n1526,n1521);
not (n1527,n1458);
nand (n1528,n1529,n1531,n1533);
or (n1529,n1524,n1530);
not (n1530,n1328);
or (n1531,n1288,n1532);
not (n1532,n1314);
not (n1533,n1534);
and (n1534,n1302,n1314);
nand (n1535,n1536,n1589);
or (n1536,n1537,n1550);
not (n1537,n1538);
nand (n1538,n1539,n1541);
xor (n1539,n1301,n1540);
not (n1540,n1287);
not (n1541,n1542);
nand (n1542,n1543,n1547,n1549);
or (n1543,n1544,n1545);
not (n1544,n1361);
not (n1545,n1546);
not (n1546,n1524);
or (n1547,n1540,n1548);
not (n1548,n1333);
not (n1549,n1327);
not (n1550,n1551);
or (n1551,n1552,n1588);
and (n1552,n1553,n1563);
xor (n1553,n1554,n1560);
nand (n1554,n1555,n1557,n1559);
or (n1555,n1288,n1556);
not (n1556,n1378);
or (n1557,n1399,n1558);
not (n1558,n1349);
not (n1559,n1332);
nand (n1560,n1561,n1562);
or (n1561,n1399,n1401);
nand (n1562,n1401,n1399);
or (n1563,n1564,n1587);
and (n1564,n1565,n1574);
xor (n1565,n1566,n1572);
nand (n1566,n1567,n1569,n1571);
not (n1567,n1568);
and (n1568,n1405,n1365);
or (n1569,n1399,n1570);
not (n1570,n1393);
not (n1571,n1348);
xnor (n1572,n1573,n1408);
not (n1573,n1405);
or (n1574,n1575,n1586);
and (n1575,n1576,n1582);
xor (n1576,n1577,n1578);
nor (n1577,n1419,n1556);
xnor (n1578,n1579,n1558);
nand (n1579,n1580,n1581);
or (n1580,n1412,n1544);
nand (n1581,n1412,n1544);
nand (n1582,n1583,n1585);
or (n1583,n1584,n1366);
xnor (n1584,n1556,n1419);
not (n1585,n1380);
and (n1586,n1577,n1578);
and (n1587,n1566,n1572);
and (n1588,n1554,n1560);
or (n1589,n1539,n1541);
and (n1590,n1591,n1274);
xor (n1591,n1592,n1600);
xor (n1592,n1593,n1599);
nand (n1593,n1594,n1596);
or (n1594,n1595,n1527);
and (n1595,n1522,n1524);
or (n1596,n1597,n1598);
not (n1597,n1329);
not (n1598,n1445);
not (n1599,n1478);
or (n1600,n1601,n1602);
and (n1601,n1518,n1535);
and (n1602,n1519,n1528);
wire s0n1603,s1n1603,notn1603;
or (n1603,s0n1603,s1n1603);
not(notn1603,n1225);
and (s0n1603,notn1603,1'b0);
and (s1n1603,n1225,n1604);
xor (n1604,n1605,n1696);
xor (n1605,n1491,n1606);
xor (n1606,n1488,n1607);
or (n1607,n1608,n1609,n1695);
and (n1608,n1462,n1511);
and (n1609,n1511,n1610);
or (n1610,n1611,n1614,n1694);
and (n1611,n1612,n1613);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n648);
and (s0n1612,notn1612,1'b0);
and (s1n1612,n648,n1499);
wire s0n1613,s1n1613,notn1613;
or (n1613,s0n1613,s1n1613);
not(notn1613,n696);
and (s0n1613,notn1613,1'b0);
and (s1n1613,n696,n1463);
and (n1614,n1613,n1615);
or (n1615,n1616,n1629,n1693);
and (n1616,n1617,n1514);
wire s0n1617,s1n1617,notn1617;
or (n1617,s0n1617,s1n1617);
not(notn1617,n648);
and (s0n1617,notn1617,1'b0);
and (s1n1617,n648,n1618);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n572);
and (s0n1618,notn1618,n1619);
and (s1n1618,n572,n1621);
wire s0n1619,s1n1619,notn1619;
or (n1619,s0n1619,s1n1619);
not(notn1619,n19);
and (s0n1619,notn1619,1'b0);
and (s1n1619,n19,n1620);
or (n1621,1'b0,n1622,n1624,n1626,n1628);
and (n1622,n1623,n553);
and (n1624,n1625,n564);
and (n1626,n1627,n568);
and (n1628,n1620,n570);
and (n1629,n1514,n1630);
or (n1630,n1631,n1645,n1692);
and (n1631,n1632,n1644);
wire s0n1632,s1n1632,notn1632;
or (n1632,s0n1632,s1n1632);
not(notn1632,n648);
and (s0n1632,notn1632,1'b0);
and (s1n1632,n648,n1633);
wire s0n1633,s1n1633,notn1633;
or (n1633,s0n1633,s1n1633);
not(notn1633,n572);
and (s0n1633,notn1633,n1634);
and (s1n1633,n572,n1636);
wire s0n1634,s1n1634,notn1634;
or (n1634,s0n1634,s1n1634);
not(notn1634,n19);
and (s0n1634,notn1634,1'b0);
and (s1n1634,n19,n1635);
or (n1636,1'b0,n1637,n1639,n1641,n1643);
and (n1637,n1638,n553);
and (n1639,n1640,n564);
and (n1641,n1642,n568);
and (n1643,n1635,n570);
wire s0n1644,s1n1644,notn1644;
or (n1644,s0n1644,s1n1644);
not(notn1644,n696);
and (s0n1644,notn1644,1'b0);
and (s1n1644,n696,n1618);
and (n1645,n1644,n1646);
or (n1646,n1647,n1661,n1663);
and (n1647,n1648,n1660);
wire s0n1648,s1n1648,notn1648;
or (n1648,s0n1648,s1n1648);
not(notn1648,n648);
and (s0n1648,notn1648,1'b0);
and (s1n1648,n648,n1649);
wire s0n1649,s1n1649,notn1649;
or (n1649,s0n1649,s1n1649);
not(notn1649,n572);
and (s0n1649,notn1649,n1650);
and (s1n1649,n572,n1652);
wire s0n1650,s1n1650,notn1650;
or (n1650,s0n1650,s1n1650);
not(notn1650,n19);
and (s0n1650,notn1650,1'b0);
and (s1n1650,n19,n1651);
or (n1652,1'b0,n1653,n1655,n1657,n1659);
and (n1653,n1654,n553);
and (n1655,n1656,n564);
and (n1657,n1658,n568);
and (n1659,n1651,n570);
wire s0n1660,s1n1660,notn1660;
or (n1660,s0n1660,s1n1660);
not(notn1660,n696);
and (s0n1660,notn1660,1'b0);
and (s1n1660,n696,n1633);
and (n1661,n1660,n1662);
or (n1662,n1663,n1677,n1678);
and (n1663,n1664,n1676);
wire s0n1664,s1n1664,notn1664;
or (n1664,s0n1664,s1n1664);
not(notn1664,n648);
and (s0n1664,notn1664,1'b0);
and (s1n1664,n648,n1665);
wire s0n1665,s1n1665,notn1665;
or (n1665,s0n1665,s1n1665);
not(notn1665,n572);
and (s0n1665,notn1665,n1666);
and (s1n1665,n572,n1668);
wire s0n1666,s1n1666,notn1666;
or (n1666,s0n1666,s1n1666);
not(notn1666,n19);
and (s0n1666,notn1666,1'b0);
and (s1n1666,n19,n1667);
or (n1668,1'b0,n1669,n1671,n1673,n1675);
and (n1669,n1670,n553);
and (n1671,n1672,n564);
and (n1673,n1674,n568);
and (n1675,n1667,n570);
wire s0n1676,s1n1676,notn1676;
or (n1676,s0n1676,s1n1676);
not(notn1676,n696);
and (s0n1676,notn1676,1'b0);
and (s1n1676,n696,n1649);
and (n1677,n1676,n1678);
and (n1678,n1679,n1691);
wire s0n1679,s1n1679,notn1679;
or (n1679,s0n1679,s1n1679);
not(notn1679,n648);
and (s0n1679,notn1679,1'b0);
and (s1n1679,n648,n1680);
wire s0n1680,s1n1680,notn1680;
or (n1680,s0n1680,s1n1680);
not(notn1680,n572);
and (s0n1680,notn1680,n1681);
and (s1n1680,n572,n1683);
wire s0n1681,s1n1681,notn1681;
or (n1681,s0n1681,s1n1681);
not(notn1681,n19);
and (s0n1681,notn1681,1'b0);
and (s1n1681,n19,n1682);
or (n1683,1'b0,n1684,n1686,n1688,n1690);
and (n1684,n1685,n553);
and (n1686,n1687,n564);
and (n1688,n1689,n568);
and (n1690,n1682,n570);
wire s0n1691,s1n1691,notn1691;
or (n1691,s0n1691,s1n1691);
not(notn1691,n696);
and (s0n1691,notn1691,1'b0);
and (s1n1691,n696,n1665);
and (n1692,n1632,n1646);
and (n1693,n1617,n1630);
and (n1694,n1612,n1615);
and (n1695,n1462,n1610);
or (n1696,n1697,n1700,n1733);
and (n1697,n1498,n1698);
xor (n1698,n1699,n1610);
xor (n1699,n1462,n1511);
and (n1700,n1698,n1701);
or (n1701,n1702,n1706,n1732);
and (n1702,n1703,n1704);
wire s0n1703,s1n1703,notn1703;
or (n1703,s0n1703,s1n1703);
not(notn1703,n591);
and (s0n1703,notn1703,1'b0);
and (s1n1703,n591,n1618);
xor (n1704,n1705,n1615);
xor (n1705,n1612,n1613);
and (n1706,n1704,n1707);
or (n1707,n1708,n1712,n1731);
and (n1708,n1709,n1710);
wire s0n1709,s1n1709,notn1709;
or (n1709,s0n1709,s1n1709);
not(notn1709,n591);
and (s0n1709,notn1709,1'b0);
and (s1n1709,n591,n1633);
xor (n1710,n1711,n1630);
xor (n1711,n1617,n1514);
and (n1712,n1710,n1713);
or (n1713,n1714,n1718,n1730);
and (n1714,n1715,n1716);
wire s0n1715,s1n1715,notn1715;
or (n1715,s0n1715,s1n1715);
not(notn1715,n591);
and (s0n1715,notn1715,1'b0);
and (s1n1715,n591,n1649);
xor (n1716,n1717,n1646);
xor (n1717,n1632,n1644);
and (n1718,n1716,n1719);
or (n1719,n1720,n1724,n1729);
and (n1720,n1721,n1722);
wire s0n1721,s1n1721,notn1721;
or (n1721,s0n1721,s1n1721);
not(notn1721,n591);
and (s0n1721,notn1721,1'b0);
and (s1n1721,n591,n1665);
xor (n1722,n1723,n1662);
xor (n1723,n1648,n1660);
and (n1724,n1722,n1725);
and (n1725,n1726,n1727);
wire s0n1726,s1n1726,notn1726;
or (n1726,s0n1726,s1n1726);
not(notn1726,n591);
and (s0n1726,notn1726,1'b0);
and (s1n1726,n591,n1680);
xor (n1727,n1728,n1678);
xor (n1728,n1664,n1676);
and (n1729,n1721,n1725);
and (n1730,n1715,n1719);
and (n1731,n1709,n1713);
and (n1732,n1703,n1707);
and (n1733,n1498,n1701);
and (n1734,n1282,n1590);
xor (n1735,n1736,n1766);
xor (n1736,n1737,n1765);
wire s0n1737,s1n1737,notn1737;
or (n1737,s0n1737,s1n1737);
not(notn1737,n932);
and (s0n1737,notn1737,1'b0);
and (s1n1737,n932,n1738);
or (n1738,n1739,n1748,n1764);
and (n1739,n1445,n1740);
and (n1740,n1483,n1741);
or (n1741,n1742,n1743,n1747);
and (n1742,n1458,n1523);
and (n1743,n1523,n1744);
or (n1744,n1534,n1745,n1746);
and (n1745,n1314,n1326);
and (n1746,n1302,n1326);
and (n1747,n1458,n1744);
and (n1748,n1740,n1749);
or (n1749,n1750,n1752,n1763);
and (n1750,n1480,n1751);
xor (n1751,n1483,n1741);
and (n1752,n1751,n1753);
or (n1753,n1754,n1757,n1762);
and (n1754,n1546,n1755);
xor (n1755,n1756,n1744);
xor (n1756,n1458,n1523);
and (n1757,n1755,n1758);
or (n1758,n1759,n1760,n1761);
and (n1759,n1287,n1300);
and (n1760,n1300,n1396);
and (n1761,n1287,n1396);
and (n1762,n1546,n1758);
and (n1763,n1480,n1753);
and (n1764,n1445,n1749);
and (n1765,n1591,n1425);
wire s0n1766,s1n1766,notn1766;
or (n1766,s0n1766,s1n1766);
not(notn1766,n1274);
and (s0n1766,notn1766,1'b0);
and (s1n1766,n1274,n1767);
xor (n1767,n1768,n1749);
xor (n1768,n1445,n1740);
wire s0n1769,s1n1769,notn1769;
or (n1769,s0n1769,s1n1769);
not(notn1769,n934);
and (s0n1769,notn1769,1'b0);
and (s1n1769,n934,n1770);
or (n1770,n1771,n1773,n1778);
and (n1771,n1432,n1772);
and (n1772,n1488,n1607);
and (n1773,n1772,n1774);
or (n1774,n1775,n1776,n1777);
and (n1775,n1491,n1606);
and (n1776,n1606,n1696);
and (n1777,n1491,n1696);
and (n1778,n1432,n1774);
or (n1779,n1780,n1901);
and (n1780,n1781,n1795);
xor (n1781,n1782,n1794);
or (n1782,n1783,n1793);
and (n1783,n1784,n1789);
xor (n1784,n1785,n1787);
and (n1785,n1786,n1225);
xor (n1786,n1107,n1131);
and (n1787,n1788,n934);
xor (n1788,n1081,n1105);
and (n1789,n1790,n1274);
xor (n1790,n1791,n788);
nor (n1791,n1792,n925);
not (n1792,n914);
and (n1793,n1785,n1787);
xor (n1794,n1281,n1603);
and (n1795,n1796,n1848);
xor (n1796,n1797,n1800);
and (n1797,n1798,n1425);
xnor (n1798,n848,n1799);
nand (n1799,n791,n913);
or (n1800,n1801,n1847);
and (n1801,n1802,n1827);
xor (n1802,n1803,n1806);
wire s0n1803,s1n1803,notn1803;
or (n1803,s0n1803,s1n1803);
not(notn1803,n1225);
and (s0n1803,notn1803,1'b0);
and (s1n1803,n1225,n1804);
xor (n1804,n1805,n1707);
xor (n1805,n1703,n1704);
and (n1806,n1807,n1821);
or (n1807,n1808,n1820);
and (n1808,n1809,n1819);
xor (n1809,n1810,n1818);
and (n1810,n1811,n982);
nand (n1811,n1812,n1814,n1817);
or (n1812,n1813,n1497);
not (n1813,n1660);
or (n1814,n1815,n1816);
not (n1815,n1703);
not (n1816,n1632);
not (n1817,n1616);
and (n1818,n1542,n982);
nor (n1819,n1539,n981);
and (n1820,n1810,n1818);
and (n1821,n1822,n982);
nor (n1822,n1823,n1825);
and (n1823,n1824,n1460);
xor (n1824,n1497,n1510);
and (n1825,n1826,n1461);
not (n1826,n1824);
or (n1827,n1828,n1846);
and (n1828,n1829,n1843);
xor (n1829,n1830,n1832);
and (n1830,n1831,n1274);
xor (n1831,n1553,n1563);
xor (n1832,n1833,n1842);
xor (n1833,n1834,n1835);
and (n1834,n1528,n982);
and (n1835,n1836,n982);
nand (n1836,n1837,n1841);
or (n1837,n1838,n1815);
and (n1838,n1839,n1840);
not (n1839,n1612);
not (n1840,n1613);
not (n1841,n1611);
and (n1842,n1519,n982);
wire s0n1843,s1n1843,notn1843;
or (n1843,s0n1843,s1n1843);
not(notn1843,n1225);
and (s0n1843,notn1843,1'b0);
and (s1n1843,n1225,n1844);
xor (n1844,n1845,n1713);
xor (n1845,n1709,n1710);
and (n1846,n1830,n1832);
and (n1847,n1803,n1806);
wire s0n1848,s1n1848,notn1848;
or (n1848,s0n1848,s1n1848);
not(notn1848,n932);
and (s0n1848,notn1848,1'b0);
and (s1n1848,n932,n1849);
xor (n1849,n1850,n1869);
xor (n1850,n1851,n1852);
xor (n1851,n768,n764);
xor (n1852,n766,n1853);
or (n1853,n780,n1854,n1868);
and (n1854,n782,n1855);
or (n1855,n921,n1856,n1867);
and (n1856,n809,n1857);
or (n1857,n822,n1858,n1866);
and (n1858,n824,n1859);
or (n1859,n843,n1860,n1865);
and (n1860,n845,n1861);
or (n1861,n856,n1862,n877);
and (n1862,n858,n1863);
or (n1863,n877,n1864,n883);
and (n1864,n879,n883);
and (n1865,n844,n1861);
and (n1866,n823,n1859);
and (n1867,n808,n1857);
and (n1868,n781,n1855);
or (n1869,n1870,n1873,n1900);
and (n1870,n1871,n1872);
xor (n1871,n920,n917);
xor (n1872,n919,n1855);
and (n1873,n1872,n1874);
or (n1874,n1875,n1878,n1899);
and (n1875,n1876,n1877);
xor (n1876,n810,n794);
xor (n1877,n807,n1857);
and (n1878,n1877,n1879);
or (n1879,n1880,n1883,n1898);
and (n1880,n1881,n1882);
xor (n1881,n831,n828);
xor (n1882,n830,n1859);
and (n1883,n1882,n1884);
or (n1884,n1885,n1888,n1897);
and (n1885,n1886,n1887);
xor (n1886,n861,n855);
xor (n1887,n860,n1861);
and (n1888,n1887,n1889);
or (n1889,n1890,n1893,n1896);
and (n1890,n1891,n1892);
xor (n1891,n902,n904);
xor (n1892,n903,n1863);
and (n1893,n1892,n1894);
and (n1894,n897,n1895);
xor (n1895,n898,n883);
and (n1896,n1891,n1894);
and (n1897,n1886,n1889);
and (n1898,n1881,n1884);
and (n1899,n1876,n1879);
and (n1900,n1871,n1874);
and (n1901,n1782,n1794);
xor (n1902,n1903,n1934);
xor (n1903,n1904,n1917);
xor (n1904,n1905,n1914);
xor (n1905,n1906,n1907);
wire s0n1906,s1n1906,notn1906;
or (n1906,s0n1906,s1n1906);
not(notn1906,n1425);
and (s0n1906,notn1906,1'b0);
and (s1n1906,n1425,n1849);
and (n1907,n1908,n1911);
or (n1908,n1909,n1910);
and (n1909,n1427,n1474);
and (n1910,n1428,n1459);
or (n1911,n1912,n1913);
and (n1912,n1429,n1457);
and (n1913,n1430,n1444);
wire s0n1914,s1n1914,notn1914;
or (n1914,s0n1914,s1n1914);
not(notn1914,n1225);
and (s0n1914,notn1914,1'b0);
and (s1n1914,n1225,n1915);
xor (n1915,n1916,n1774);
xor (n1916,n1432,n1772);
or (n1917,n1918,n1933);
and (n1918,n1919,n1932);
xor (n1919,n1920,n1931);
or (n1920,n1921,n1930);
and (n1921,n1922,n1929);
xor (n1922,n1923,n1924);
xor (n1923,n1283,n1516);
and (n1924,n1925,n1928);
xor (n1925,n1926,n1927);
and (n1926,n1831,n1425);
wire s0n1927,s1n1927,notn1927;
or (n1927,s0n1927,s1n1927);
not(notn1927,n1274);
and (s0n1927,notn1927,1'b0);
and (s1n1927,n1274,n1285);
and (n1928,n1517,n932);
wire s0n1929,s1n1929,notn1929;
or (n1929,s0n1929,s1n1929);
not(notn1929,n934);
and (s0n1929,notn1929,1'b0);
and (s1n1929,n934,n1604);
and (n1930,n1923,n1924);
and (n1931,n1788,n1225);
wire s0n1932,s1n1932,notn1932;
or (n1932,s0n1932,s1n1932);
not(notn1932,n1274);
and (s0n1932,notn1932,1'b0);
and (s1n1932,n1274,n1849);
and (n1933,n1920,n1931);
or (n1934,n1935,n1945);
and (n1935,n1936,n1944);
xor (n1936,n1937,n1938);
wire s0n1937,s1n1937,notn1937;
or (n1937,s0n1937,s1n1937);
not(notn1937,n982);
and (s0n1937,notn1937,1'b0);
and (s1n1937,n982,n14);
and (n1938,n1939,n982);
xnor (n1939,n1940,n1942);
not (n1940,n1941);
and (n1941,n589,n1034);
or (n1942,n1943,n1078);
and (n1943,n1031,n1079);
and (n1944,n1273,n932);
and (n1945,n1937,n1938);
or (n1946,n1947,n2120);
and (n1947,n1948,n1987);
xor (n1948,n1949,n1950);
xor (n1949,n1781,n1795);
or (n1950,n1951,n1986);
and (n1951,n1952,n1961);
xor (n1952,n1953,n1960);
or (n1953,n1954,n1959);
and (n1954,n1955,n1958);
xor (n1955,n1956,n1957);
and (n1956,n1798,n1274);
xor (n1957,n1802,n1827);
and (n1958,n1788,n982);
and (n1959,n1956,n1957);
xor (n1960,n1796,n1848);
or (n1961,n1962,n1985);
and (n1962,n1963,n1984);
xor (n1963,n1964,n1965);
and (n1964,n1786,n934);
or (n1965,n1966,n1983);
and (n1966,n1967,n1980);
xor (n1967,n1968,n1972);
xor (n1968,n1969,n1970);
xor (n1969,n1807,n1821);
and (n1970,n1971,n1425);
xor (n1971,n1565,n1574);
and (n1972,n1973,n1977);
xor (n1973,n1974,n1975);
xor (n1974,n1809,n1819);
and (n1975,n1976,n1425);
xor (n1976,n1576,n1582);
wire s0n1977,s1n1977,notn1977;
or (n1977,s0n1977,s1n1977);
not(notn1977,n1225);
and (s0n1977,notn1977,1'b0);
and (s1n1977,n1225,n1978);
xor (n1978,n1979,n1719);
xor (n1979,n1715,n1716);
wire s0n1980,s1n1980,notn1980;
or (n1980,s0n1980,s1n1980);
not(notn1980,n1425);
and (s0n1980,notn1980,1'b0);
and (s1n1980,n1425,n1981);
xor (n1981,n1982,n1889);
xor (n1982,n1886,n1887);
and (n1983,n1968,n1972);
and (n1984,n1790,n932);
and (n1985,n1964,n1965);
and (n1986,n1953,n1960);
or (n1987,n1988,n2119);
and (n1988,n1989,n2100);
xor (n1989,n1990,n2099);
or (n1990,n1991,n2098);
and (n1991,n1992,n2097);
xor (n1992,n1993,n2068);
or (n1993,n1994,n2067);
and (n1994,n1995,n2064);
xor (n1995,n1996,n2019);
xor (n1996,n1997,n2018);
xor (n1997,n1998,n1999);
wire s0n1998,s1n1998,notn1998;
or (n1998,s0n1998,s1n1998);
not(notn1998,n932);
and (s0n1998,notn1998,1'b0);
and (s1n1998,n932,n1285);
or (n1999,n2000,n2017);
and (n2000,n2001,n2016);
xor (n2001,n2002,n2014);
or (n2002,n2003,n2004);
and (n2003,n1554,n982);
and (n2004,n2005,n982);
nand (n2005,n2006,n2007);
not (n2006,n1631);
nand (n2007,n2008,n2012);
or (n2008,n2009,n2010);
not (n2009,n1816);
not (n2010,n2011);
not (n2011,n1644);
not (n2012,n2013);
not (n2013,n1715);
nor (n2014,n981,n2015);
xor (n2015,n1705,n1815);
and (n2016,n1971,n1274);
and (n2017,n2002,n2014);
wire s0n2018,s1n2018,notn2018;
or (n2018,s0n2018,s1n2018);
not(notn2018,n934);
and (s0n2018,notn2018,1'b0);
and (s1n2018,n934,n1804);
and (n2019,n2020,n2063);
xor (n2020,n2021,n2057);
or (n2021,n2022,n2056);
and (n2022,n2023,n2053);
xor (n2023,n2024,n2038);
and (n2024,n2025,n2030);
xor (n2025,n2026,n2028);
and (n2026,n2027,n982);
xnor (n2027,n2013,n1717);
and (n2028,n1425,n2029);
xor (n2029,n1381,n1393);
and (n2030,n2031,n2034);
and (n2031,n2032,n2012);
wire s0n2032,s1n2032,notn2032;
or (n2032,s0n2032,s1n2032);
not(notn2032,n982);
and (s0n2032,notn2032,1'b0);
and (s1n2032,n982,n2033);
wire s0n2033,s1n2033,notn2033;
or (n2033,s0n2033,s1n2033);
not(notn2033,n696);
and (s0n2033,notn2033,1'b0);
and (s1n2033,n696,n1680);
nor (n2034,n2035,n1573);
not (n2035,n2036);
wire s0n2036,s1n2036,notn2036;
or (n2036,s0n2036,s1n2036);
not(notn2036,n982);
and (s0n2036,notn2036,1'b0);
and (s1n2036,n982,n2037);
wire s0n2037,s1n2037,notn2037;
or (n2037,s0n2037,s1n2037);
not(notn2037,n696);
and (s0n2037,notn2037,1'b0);
and (s1n2037,n696,n1382);
or (n2038,n2039,n2052);
and (n2039,n2040,n2051);
xor (n2040,n2041,n2050);
and (n2041,n2042,n982);
not (n2042,n2043);
nor (n2043,n2044,n2045);
and (n2044,n2012,n1664);
and (n2045,n2046,n2049);
nand (n2046,n2047,n2048);
not (n2047,n1721);
not (n2048,n1648);
not (n2049,n1813);
and (n2050,n1566,n982);
and (n2051,n1572,n982);
and (n2052,n2041,n2050);
wire s0n2053,s1n2053,notn2053;
or (n2053,s0n2053,s1n2053);
not(notn2053,n1225);
and (s0n2053,notn2053,1'b0);
and (s1n2053,n1225,n2054);
xor (n2054,n2055,n1725);
xor (n2055,n1721,n1722);
and (n2056,n2024,n2038);
and (n2057,n2058,n2062);
xor (n2058,n2059,n2060);
wire s0n2059,s1n2059,notn2059;
or (n2059,s0n2059,s1n2059);
not(notn2059,n934);
and (s0n2059,notn2059,1'b0);
and (s1n2059,n934,n1978);
wire s0n2060,s1n2060,notn2060;
or (n2060,s0n2060,s1n2060);
not(notn2060,n1425);
and (s0n2060,notn2060,1'b0);
and (s1n2060,n1425,n2061);
xor (n2061,n1418,n1420);
and (n2062,n1971,n932);
xor (n2063,n1973,n1977);
wire s0n2064,s1n2064,notn2064;
or (n2064,s0n2064,s1n2064);
not(notn2064,n1274);
and (s0n2064,notn2064,1'b0);
and (s1n2064,n1274,n2065);
xor (n2065,n2066,n1884);
xor (n2066,n1881,n1882);
and (n2067,n1996,n2019);
or (n2068,n2069,n2096);
and (n2069,n2070,n2094);
xor (n2070,n2071,n2072);
xor (n2071,n1829,n1843);
or (n2072,n2073,n2093);
and (n2073,n2074,n2092);
xor (n2074,n2075,n2076);
and (n2075,n1831,n932);
or (n2076,n2077,n2091);
and (n2077,n2078,n2090);
xor (n2078,n2079,n2089);
and (n2079,n2080,n982);
not (n2080,n2081);
nor (n2081,n2082,n2088);
and (n2082,n2083,n2086);
not (n2083,n2084);
xor (n2084,n1513,n2085);
not (n2085,n1709);
not (n2086,n2087);
not (n2087,n1617);
and (n2088,n2084,n2087);
and (n2089,n1560,n982);
and (n2090,n1976,n1274);
and (n2091,n2079,n2089);
wire s0n2092,s1n2092,notn2092;
or (n2092,s0n2092,s1n2092);
not(notn2092,n934);
and (s0n2092,notn2092,1'b0);
and (s1n2092,n934,n1844);
and (n2093,n2075,n2076);
and (n2094,n2095,n1225);
xor (n2095,n1159,n1183);
and (n2096,n2071,n2072);
wire s0n2097,s1n2097,notn2097;
or (n2097,s0n2097,s1n2097);
not(notn2097,n982);
and (s0n2097,notn2097,1'b0);
and (s1n2097,n982,n1849);
and (n2098,n1993,n2068);
xor (n2099,n1784,n1789);
xor (n2100,n2101,n2118);
xor (n2101,n2102,n2103);
and (n2102,n1030,n982);
xor (n2103,n2104,n2115);
xor (n2104,n2105,n2106);
and (n2105,n1591,n932);
or (n2106,n2107,n2114);
and (n2107,n2108,n2111);
xor (n2108,n2109,n2110);
xor (n2109,n1476,n1493);
and (n2110,n1593,n982);
or (n2111,n2112,n2113);
and (n2112,n1833,n1842);
and (n2113,n1834,n1835);
and (n2114,n2109,n2110);
wire s0n2115,s1n2115,notn2115;
or (n2115,s0n2115,s1n2115);
not(notn2115,n1225);
and (s0n2115,notn2115,1'b0);
and (s1n2115,n1225,n2116);
xor (n2116,n2117,n1701);
xor (n2117,n1498,n1698);
and (n2118,n1273,n982);
and (n2119,n1990,n2099);
and (n2120,n1949,n1950);
and (n2121,n8,n1902);
xor (n2122,n2123,n2150);
xor (n2123,n2124,n2131);
xor (n2124,n2125,n2128);
xor (n2125,n2126,n2127);
and (n2126,n1905,n1914);
and (n2127,n1736,n1766);
or (n2128,n2129,n2130);
and (n2129,n11,n1272);
and (n2130,n12,n1029);
and (n2131,n2132,n2143);
xor (n2132,n2133,n2142);
or (n2133,n2134,n2141);
and (n2134,n2135,n2140);
xor (n2135,n2136,n2137);
wire s0n2136,s1n2136,notn2136;
or (n2136,s0n2136,s1n2136);
not(notn2136,n932);
and (s0n2136,notn2136,1'b0);
and (s1n2136,n932,n1767);
xor (n2137,n2138,n2139);
xor (n2138,n1908,n1911);
and (n2139,n1517,n1425);
and (n2140,n1030,n934);
and (n2141,n2136,n2137);
and (n2142,n1939,n934);
and (n2143,n2144,n2149);
xor (n2144,n2145,n2146);
and (n2145,n1790,n1425);
or (n2146,n2147,n2148);
and (n2147,n2104,n2115);
and (n2148,n2105,n2106);
wire s0n2149,s1n2149,notn2149;
or (n2149,s0n2149,s1n2149);
not(notn2149,n934);
and (s0n2149,notn2149,1'b0);
and (s1n2149,n934,n1915);
or (n2150,n2151,n2152);
and (n2151,n1903,n1934);
and (n2152,n1904,n1917);
xor (n2153,n2154,n2173);
xor (n2154,n2155,n2158);
or (n2155,n2156,n2157);
and (n2156,n9,n1779);
and (n2157,n10,n1277);
xor (n2158,n2159,n2168);
xor (n2159,n2160,n2163);
or (n2160,n2161,n2162);
and (n2161,n1278,n1769);
and (n2162,n1279,n1735);
xor (n2163,n2164,n2167);
xor (n2164,n2165,n2166);
wire s0n2165,s1n2165,notn2165;
or (n2165,s0n2165,s1n2165);
not(notn2165,n1425);
and (s0n2165,notn2165,1'b0);
and (s1n2165,n1425,n1767);
wire s0n2166,s1n2166,notn2166;
or (n2166,s0n2166,s1n2166);
not(notn2166,n1274);
and (s0n2166,notn2166,1'b0);
and (s1n2166,n1274,n1738);
and (n2167,n1273,n1425);
xor (n2168,n2169,n2172);
xor (n2169,n2170,n2171);
and (n2170,n1939,n1225);
wire s0n2171,s1n2171,notn2171;
or (n2171,s0n2171,s1n2171);
not(notn2171,n1225);
and (s0n2171,notn2171,1'b0);
and (s1n2171,n1225,n1770);
wire s0n2172,s1n2172,notn2172;
or (n2172,s0n2172,s1n2172);
not(notn2172,n1274);
and (s0n2172,notn2172,1'b0);
and (s1n2172,n1274,n14);
or (n2173,n2174,n2214);
and (n2174,n2175,n2186);
xor (n2175,n2176,n2185);
or (n2176,n2177,n2184);
and (n2177,n2178,n2183);
xor (n2178,n2179,n2182);
or (n2179,n2180,n2181);
and (n2180,n2101,n2118);
and (n2181,n2102,n2103);
xor (n2182,n2135,n2140);
xor (n2183,n1919,n1932);
and (n2184,n2179,n2182);
xor (n2185,n2132,n2143);
or (n2186,n2187,n2213);
and (n2187,n2188,n2212);
xor (n2188,n2189,n2190);
xor (n2189,n2144,n2149);
or (n2190,n2191,n2211);
and (n2191,n2192,n2203);
xor (n2192,n2193,n2194);
xor (n2193,n1922,n1929);
or (n2194,n2195,n2202);
and (n2195,n2196,n2201);
xor (n2196,n2197,n2200);
or (n2197,n2198,n2199);
and (n2198,n1997,n2018);
and (n2199,n1998,n1999);
xor (n2200,n2108,n2111);
wire s0n2201,s1n2201,notn2201;
or (n2201,s0n2201,s1n2201);
not(notn2201,n934);
and (s0n2201,notn2201,1'b0);
and (s1n2201,n934,n2116);
and (n2202,n2197,n2200);
or (n2203,n2204,n2210);
and (n2204,n2205,n2208);
xor (n2205,n2206,n2207);
wire s0n2206,s1n2206,notn2206;
or (n2206,s0n2206,s1n2206);
not(notn2206,n1425);
and (s0n2206,notn2206,1'b0);
and (s1n2206,n1425,n2065);
xor (n2207,n1925,n1928);
and (n2208,n2209,n1225);
xor (n2209,n1133,n1157);
and (n2210,n2206,n2207);
and (n2211,n2193,n2194);
xor (n2212,n1936,n1944);
and (n2213,n2189,n2190);
and (n2214,n2176,n2185);
or (n2215,n2216,n2285);
and (n2216,n2217,n2284);
xor (n2217,n2218,n2283);
or (n2218,n2219,n2282);
and (n2219,n2220,n2223);
xor (n2220,n2221,n2222);
xor (n2221,n2188,n2212);
xor (n2222,n2178,n2183);
or (n2223,n2224,n2281);
and (n2224,n2225,n2268);
xor (n2225,n2226,n2267);
or (n2226,n2227,n2266);
and (n2227,n2228,n2231);
xor (n2228,n2229,n2230);
xor (n2229,n2205,n2208);
xor (n2230,n2196,n2201);
or (n2231,n2232,n2265);
and (n2232,n2233,n2264);
xor (n2233,n2234,n2241);
and (n2234,n2235,n2239);
xor (n2235,n2236,n2238);
and (n2236,n2237,n1425);
xor (n2237,n876,n900);
xor (n2238,n2001,n2016);
and (n2239,n2240,n1225);
xor (n2240,n1185,n1203);
or (n2241,n2242,n2263);
and (n2242,n2243,n2262);
xor (n2243,n2244,n2245);
xor (n2244,n2074,n2092);
or (n2245,n2246,n2261);
and (n2246,n2247,n2253);
xor (n2247,n2248,n2249);
xor (n2248,n2078,n2090);
nand (n2249,n2250,n2002);
or (n2250,n2251,n2252);
not (n2251,n2004);
not (n2252,n2003);
or (n2253,n2254,n2260);
and (n2254,n2255,n2259);
xor (n2255,n2256,n2257);
wire s0n2256,s1n2256,notn2256;
or (n2256,s0n2256,s1n2256);
not(notn2256,n1274);
and (s0n2256,notn2256,1'b0);
and (s1n2256,n1274,n2061);
wire s0n2257,s1n2257,notn2257;
or (n2257,s0n2257,s1n2257);
not(notn2257,n1225);
and (s0n2257,notn2257,1'b0);
and (s1n2257,n1225,n2258);
xor (n2258,n1726,n1727);
and (n2259,n1976,n932);
and (n2260,n2256,n2257);
and (n2261,n2248,n2249);
wire s0n2262,s1n2262,notn2262;
or (n2262,s0n2262,s1n2262);
not(notn2262,n1274);
and (s0n2262,notn2262,1'b0);
and (s1n2262,n1274,n1981);
and (n2263,n2244,n2245);
and (n2264,n1786,n982);
and (n2265,n2234,n2241);
and (n2266,n2229,n2230);
xor (n2267,n2192,n2203);
or (n2268,n2269,n2280);
and (n2269,n2270,n2279);
xor (n2270,n2271,n2272);
xor (n2271,n1955,n1958);
or (n2272,n2273,n2278);
and (n2273,n2274,n2277);
xor (n2274,n2275,n2276);
and (n2275,n1798,n932);
and (n2276,n2209,n934);
and (n2277,n1790,n982);
and (n2278,n2275,n2276);
xor (n2279,n1963,n1984);
and (n2280,n2271,n2272);
and (n2281,n2226,n2267);
and (n2282,n2221,n2222);
xor (n2283,n2175,n2186);
xor (n2284,n7,n1946);
and (n2285,n2218,n2283);
or (n2286,n2287,n2741);
and (n2287,n2288,n2373);
xor (n2288,n2289,n2290);
xor (n2289,n2217,n2284);
or (n2290,n2291,n2372);
and (n2291,n2292,n2371);
xor (n2292,n2293,n2370);
or (n2293,n2294,n2369);
and (n2294,n2295,n2368);
xor (n2295,n2296,n2297);
xor (n2296,n1952,n1961);
or (n2297,n2298,n2367);
and (n2298,n2299,n2336);
xor (n2299,n2300,n2301);
xor (n2300,n1992,n2097);
or (n2301,n2302,n2335);
and (n2302,n2303,n2306);
xor (n2303,n2304,n2305);
xor (n2304,n1967,n1980);
xor (n2305,n2070,n2094);
or (n2306,n2307,n2334);
and (n2307,n2308,n2333);
xor (n2308,n2309,n2332);
and (n2309,n2310,n2331);
and (n2310,n2311,n2318);
or (n2311,n2312,n2317);
and (n2312,n2313,n2316);
xor (n2313,n2314,n2315);
and (n2314,n1274,n2029);
xor (n2315,n2031,n2034);
wire s0n2316,s1n2316,notn2316;
or (n2316,s0n2316,s1n2316);
not(notn2316,n934);
and (s0n2316,notn2316,1'b0);
and (s1n2316,n934,n2258);
and (n2317,n2314,n2315);
and (n2318,n2319,n2330);
xor (n2319,n2320,n2328);
and (n2320,n2321,n982);
nand (n2321,n2322,n2327);
or (n2322,n2048,n2323);
nand (n2323,n2324,n2326);
or (n2324,n2325,n1813);
not (n2325,n2047);
nand (n2326,n2325,n1813);
nand (n2327,n2323,n2048);
wire s0n2328,s1n2328,notn2328;
or (n2328,s0n2328,s1n2328);
not(notn2328,n1425);
and (s0n2328,notn2328,1'b0);
and (s1n2328,n1425,n2329);
wire s0n2329,s1n2329,notn2329;
or (n2329,s0n2329,s1n2329);
not(notn2329,n696);
and (s0n2329,notn2329,1'b0);
and (s1n2329,n696,n885);
and (n2330,n1578,n982);
xor (n2331,n2023,n2053);
wire s0n2332,s1n2332,notn2332;
or (n2332,s0n2332,s1n2332);
not(notn2332,n932);
and (s0n2332,notn2332,1'b0);
and (s1n2332,n932,n2065);
and (n2333,n2095,n934);
and (n2334,n2309,n2332);
and (n2335,n2304,n2305);
or (n2336,n2337,n2366);
and (n2337,n2338,n2365);
xor (n2338,n2339,n2364);
or (n2339,n2340,n2363);
and (n2340,n2341,n2362);
xor (n2341,n2342,n2361);
or (n2342,n2343,n2360);
and (n2343,n2344,n2359);
xor (n2344,n2345,n2346);
xor (n2345,n2058,n2062);
or (n2346,n2347,n2358);
and (n2347,n2348,n2357);
xor (n2348,n2349,n2350);
xor (n2349,n2040,n2051);
and (n2350,n2351,n2353);
wire s0n2351,s1n2351,notn2351;
or (n2351,s0n2351,s1n2351);
not(notn2351,n1225);
and (s0n2351,notn2351,1'b0);
and (s1n2351,n1225,n2352);
xor (n2352,n1679,n1691);
and (n2353,n2354,n2355);
wire s0n2354,s1n2354,notn2354;
or (n2354,s0n2354,s1n2354);
not(notn2354,n1225);
and (s0n2354,notn2354,1'b0);
and (s1n2354,n1225,n2033);
wire s0n2355,s1n2355,notn2355;
or (n2355,s0n2355,s1n2355);
not(notn2355,n1225);
and (s0n2355,notn2355,1'b0);
and (s1n2355,n1225,n2356);
wire s0n2356,s1n2356,notn2356;
or (n2356,s0n2356,s1n2356);
not(notn2356,n696);
and (s0n2356,notn2356,1'b0);
and (s1n2356,n696,n1189);
wire s0n2357,s1n2357,notn2357;
or (n2357,s0n2357,s1n2357);
not(notn2357,n934);
and (s0n2357,notn2357,1'b0);
and (s1n2357,n934,n2054);
and (n2358,n2349,n2350);
and (n2359,n2237,n1274);
and (n2360,n2345,n2346);
xor (n2361,n2020,n2063);
and (n2362,n1798,n982);
and (n2363,n2342,n2361);
xor (n2364,n1995,n2064);
xor (n2365,n2274,n2277);
and (n2366,n2339,n2364);
and (n2367,n2300,n2301);
xor (n2368,n1989,n2100);
and (n2369,n2296,n2297);
xor (n2370,n1948,n1987);
xor (n2371,n2220,n2223);
and (n2372,n2293,n2370);
or (n2373,n2374,n2740);
and (n2374,n2375,n2483);
xor (n2375,n2376,n2377);
xor (n2376,n2292,n2371);
or (n2377,n2378,n2482);
and (n2378,n2379,n2481);
xor (n2379,n2380,n2381);
xor (n2380,n2225,n2268);
or (n2381,n2382,n2480);
and (n2382,n2383,n2479);
xor (n2383,n2384,n2385);
xor (n2384,n2228,n2231);
or (n2385,n2386,n2478);
and (n2386,n2387,n2411);
xor (n2387,n2388,n2410);
or (n2388,n2389,n2409);
and (n2389,n2390,n2393);
xor (n2390,n2391,n2392);
and (n2391,n2209,n982);
xor (n2392,n2235,n2239);
or (n2393,n2394,n2408);
and (n2394,n2395,n2407);
xor (n2395,n2396,n2405);
or (n2396,n2397,n2404);
and (n2397,n2398,n2402);
xor (n2398,n2399,n2401);
and (n2399,n2400,n1225);
xor (n2400,n1211,n1216);
xor (n2401,n2025,n2030);
and (n2402,n2403,n1274);
xor (n2403,n882,n898);
and (n2404,n2399,n2401);
and (n2405,n2406,n1225);
xor (n2406,n1205,n1218);
wire s0n2407,s1n2407,notn2407;
or (n2407,s0n2407,s1n2407);
not(notn2407,n932);
and (s0n2407,notn2407,1'b0);
and (s1n2407,n932,n1981);
and (n2408,n2396,n2405);
and (n2409,n2391,n2392);
xor (n2410,n2233,n2264);
or (n2411,n2412,n2477);
and (n2412,n2413,n2476);
xor (n2413,n2414,n2415);
xor (n2414,n2243,n2262);
or (n2415,n2416,n2475);
and (n2416,n2417,n2474);
xor (n2417,n2418,n2419);
and (n2418,n2240,n934);
or (n2419,n2420,n2473);
and (n2420,n2421,n2446);
xor (n2421,n2422,n2423);
xor (n2422,n2255,n2259);
or (n2423,n2424,n2445);
and (n2424,n2425,n2444);
xor (n2425,n2426,n2434);
or (n2426,n2427,n2433);
and (n2427,n2428,n2431);
xor (n2428,n2429,n2430);
xor (n2429,n2354,n2355);
wire s0n2430,s1n2430,notn2430;
or (n2430,s0n2430,s1n2430);
not(notn2430,n934);
and (s0n2430,notn2430,1'b0);
and (s1n2430,n934,n2352);
and (n2431,n2432,n982);
not (n2432,n1584);
and (n2433,n2429,n2430);
or (n2434,n2435,n2443);
and (n2435,n2436,n2439);
xor (n2436,n2437,n2438);
and (n2437,n1365,n982);
and (n2438,n1664,n982);
and (n2439,n2440,n982);
xor (n2440,n2441,n2442);
not (n2441,n1676);
not (n2442,n1726);
and (n2443,n2437,n2438);
wire s0n2444,s1n2444,notn2444;
or (n2444,s0n2444,s1n2444);
not(notn2444,n932);
and (s0n2444,notn2444,1'b0);
and (s1n2444,n932,n2061);
and (n2445,n2426,n2434);
or (n2446,n2447,n2472);
and (n2447,n2448,n2470);
xor (n2448,n2449,n2467);
or (n2449,n2450,n2466);
and (n2450,n2451,n2465);
xor (n2451,n2452,n2460);
or (n2452,n2453,n2459);
and (n2453,n2454,n2457);
xor (n2454,n2455,n2456);
nor (n2455,n1570,n981);
wire s0n2456,s1n2456,notn2456;
or (n2456,s0n2456,s1n2456);
not(notn2456,n934);
and (s0n2456,notn2456,1'b0);
and (s1n2456,n934,n2033);
nor (n2457,n2458,n981);
not (n2458,n1691);
and (n2459,n2455,n2456);
and (n2460,n2461,n2463);
nor (n2461,n2462,n981);
not (n2462,n1381);
nor (n2463,n2464,n981);
not (n2464,n1679);
wire s0n2465,s1n2465,notn2465;
or (n2465,s0n2465,s1n2465);
not(notn2465,n1274);
and (s0n2465,notn2465,1'b0);
and (s1n2465,n1274,n2329);
and (n2466,n2452,n2460);
xor (n2467,n2468,n2469);
xor (n2468,n2351,n2353);
wire s0n2469,s1n2469,notn2469;
or (n2469,s0n2469,s1n2469);
not(notn2469,n1425);
and (s0n2469,notn2469,1'b0);
and (s1n2469,n1425,n2037);
and (n2470,n2471,n1225);
xor (n2471,n1213,n1214);
and (n2472,n2449,n2467);
and (n2473,n2422,n2423);
and (n2474,n2095,n982);
and (n2475,n2418,n2419);
xor (n2476,n2308,n2333);
and (n2477,n2414,n2415);
and (n2478,n2388,n2410);
xor (n2479,n2270,n2279);
and (n2480,n2384,n2385);
xor (n2481,n2295,n2368);
and (n2482,n2380,n2381);
or (n2483,n2484,n2739);
and (n2484,n2485,n2547);
xor (n2485,n2486,n2546);
or (n2486,n2487,n2545);
and (n2487,n2488,n2544);
xor (n2488,n2489,n2543);
or (n2489,n2490,n2542);
and (n2490,n2491,n2541);
xor (n2491,n2492,n2540);
or (n2492,n2493,n2539);
and (n2493,n2494,n2538);
xor (n2494,n2495,n2531);
or (n2495,n2496,n2530);
and (n2496,n2497,n2523);
xor (n2497,n2498,n2501);
xor (n2498,n2499,n2500);
xor (n2499,n2310,n2331);
and (n2500,n2403,n1425);
or (n2501,n2502,n2522);
and (n2502,n2503,n2521);
xor (n2503,n2504,n2518);
or (n2504,n2505,n2517);
and (n2505,n2506,n2516);
xor (n2506,n2507,n2509);
wire s0n2507,s1n2507,notn2507;
or (n2507,s0n2507,s1n2507);
not(notn2507,n1274);
and (s0n2507,notn2507,1'b0);
and (s1n2507,n1274,n2508);
xor (n2508,n884,n896);
or (n2509,n2510,n2515);
and (n2510,n2511,n2514);
xor (n2511,n2512,n2513);
xor (n2512,n2436,n2439);
wire s0n2513,s1n2513,notn2513;
or (n2513,s0n2513,s1n2513);
not(notn2513,n932);
and (s0n2513,notn2513,1'b0);
and (s1n2513,n932,n2029);
wire s0n2514,s1n2514,notn2514;
or (n2514,s0n2514,s1n2514);
not(notn2514,n1274);
and (s0n2514,notn2514,1'b0);
and (s1n2514,n1274,n2037);
and (n2515,n2512,n2513);
xor (n2516,n2313,n2316);
and (n2517,n2507,n2509);
xor (n2518,n2519,n2520);
xor (n2519,n2311,n2318);
wire s0n2520,s1n2520,notn2520;
or (n2520,s0n2520,s1n2520);
not(notn2520,n1425);
and (s0n2520,notn2520,1'b0);
and (s1n2520,n1425,n2508);
and (n2521,n2237,n932);
and (n2522,n2504,n2518);
or (n2523,n2524,n2529);
and (n2524,n2525,n2528);
xor (n2525,n2526,n2527);
and (n2526,n2406,n934);
xor (n2527,n2348,n2357);
wire s0n2528,s1n2528,notn2528;
or (n2528,s0n2528,s1n2528);
not(notn2528,n982);
and (s0n2528,notn2528,1'b0);
and (s1n2528,n982,n1981);
and (n2529,n2526,n2527);
and (n2530,n2498,n2501);
or (n2531,n2532,n2537);
and (n2532,n2533,n2536);
xor (n2533,n2534,n2535);
xor (n2534,n2247,n2253);
xor (n2535,n2344,n2359);
wire s0n2536,s1n2536,notn2536;
or (n2536,s0n2536,s1n2536);
not(notn2536,n982);
and (s0n2536,notn2536,1'b0);
and (s1n2536,n982,n2065);
and (n2537,n2534,n2535);
xor (n2538,n2341,n2362);
and (n2539,n2495,n2531);
xor (n2540,n2303,n2306);
xor (n2541,n2338,n2365);
and (n2542,n2492,n2540);
xor (n2543,n2299,n2336);
xor (n2544,n2383,n2479);
and (n2545,n2489,n2543);
xor (n2546,n2379,n2481);
or (n2547,n2548,n2738);
and (n2548,n2549,n2625);
xor (n2549,n2550,n2624);
or (n2550,n2551,n2623);
and (n2551,n2552,n2622);
xor (n2552,n2553,n2554);
xor (n2553,n2387,n2411);
or (n2554,n2555,n2621);
and (n2555,n2556,n2620);
xor (n2556,n2557,n2558);
xor (n2557,n2390,n2393);
or (n2558,n2559,n2619);
and (n2559,n2560,n2575);
xor (n2560,n2561,n2562);
xor (n2561,n2395,n2407);
or (n2562,n2563,n2574);
and (n2563,n2564,n2573);
xor (n2564,n2565,n2566);
xor (n2565,n2398,n2402);
or (n2566,n2567,n2572);
and (n2567,n2568,n2571);
xor (n2568,n2569,n2570);
and (n2569,n2400,n934);
xor (n2570,n2319,n2330);
and (n2571,n2403,n932);
and (n2572,n2569,n2570);
and (n2573,n2240,n982);
and (n2574,n2565,n2566);
or (n2575,n2576,n2618);
and (n2576,n2577,n2599);
xor (n2577,n2578,n2579);
xor (n2578,n2421,n2446);
or (n2579,n2580,n2598);
and (n2580,n2581,n2597);
xor (n2581,n2582,n2596);
or (n2582,n2583,n2595);
and (n2583,n2584,n2594);
xor (n2584,n2585,n2586);
xor (n2585,n2428,n2431);
or (n2586,n2587,n2593);
and (n2587,n2588,n2592);
xor (n2588,n2589,n2591);
and (n2589,n2036,n2590);
wire s0n2590,s1n2590,notn2590;
or (n2590,s0n2590,s1n2590);
not(notn2590,n982);
and (s0n2590,notn2590,1'b0);
and (s1n2590,n982,n2356);
wire s0n2591,s1n2591,notn2591;
or (n2591,s0n2591,s1n2591);
not(notn2591,n934);
and (s0n2591,notn2591,1'b0);
and (s1n2591,n934,n2356);
xor (n2592,n2461,n2463);
and (n2593,n2589,n2591);
wire s0n2594,s1n2594,notn2594;
or (n2594,s0n2594,s1n2594);
not(notn2594,n932);
and (s0n2594,notn2594,1'b0);
and (s1n2594,n932,n2508);
and (n2595,n2585,n2586);
xor (n2596,n2425,n2444);
and (n2597,n2406,n982);
and (n2598,n2582,n2596);
or (n2599,n2600,n2617);
and (n2600,n2601,n2616);
xor (n2601,n2602,n2603);
xor (n2602,n2448,n2470);
or (n2603,n2604,n2615);
and (n2604,n2605,n2614);
xor (n2605,n2606,n2607);
xor (n2606,n2511,n2514);
or (n2607,n2608,n2613);
and (n2608,n2609,n2612);
xor (n2609,n2610,n2611);
wire s0n2610,s1n2610,notn2610;
or (n2610,s0n2610,s1n2610);
not(notn2610,n932);
and (s0n2610,notn2610,1'b0);
and (s1n2610,n932,n2329);
xor (n2611,n2454,n2457);
wire s0n2612,s1n2612,notn2612;
or (n2612,s0n2612,s1n2612);
not(notn2612,n932);
and (s0n2612,notn2612,1'b0);
and (s1n2612,n932,n2037);
and (n2613,n2610,n2611);
and (n2614,n2471,n934);
and (n2615,n2606,n2607);
and (n2616,n2237,n982);
and (n2617,n2602,n2603);
and (n2618,n2578,n2579);
and (n2619,n2561,n2562);
xor (n2620,n2413,n2476);
and (n2621,n2557,n2558);
xor (n2622,n2491,n2541);
and (n2623,n2553,n2554);
xor (n2624,n2488,n2544);
nand (n2625,n2626,n2737);
or (n2626,n2627,n2642);
nor (n2627,n2628,n2629);
xor (n2628,n2552,n2622);
or (n2629,n2630,n2641);
and (n2630,n2631,n2640);
xor (n2631,n2632,n2633);
xor (n2632,n2494,n2538);
or (n2633,n2634,n2639);
and (n2634,n2635,n2638);
xor (n2635,n2636,n2637);
xor (n2636,n2417,n2474);
xor (n2637,n2533,n2536);
xor (n2638,n2497,n2523);
and (n2639,n2636,n2637);
xor (n2640,n2556,n2620);
and (n2641,n2632,n2633);
and (n2642,n2643,n2736);
nand (n2643,n2644,n2659);
or (n2644,n2645,n2646);
xor (n2645,n2631,n2640);
or (n2646,n2647,n2658);
and (n2647,n2648,n2657);
xor (n2648,n2649,n2656);
or (n2649,n2650,n2655);
and (n2650,n2651,n2654);
xor (n2651,n2652,n2653);
xor (n2652,n2525,n2528);
xor (n2653,n2503,n2521);
xor (n2654,n2564,n2573);
and (n2655,n2652,n2653);
xor (n2656,n2560,n2575);
xor (n2657,n2635,n2638);
and (n2658,n2649,n2656);
nand (n2659,n2660,n2729);
nand (n2660,n2661,n2700,n2703);
or (n2661,n2662,n2699);
or (n2662,n2663,n2698);
and (n2663,n2664,n2697);
xor (n2664,n2665,n2684);
or (n2665,n2666,n2683);
and (n2666,n2667,n2682);
xor (n2667,n2668,n2669);
xor (n2668,n2581,n2597);
or (n2669,n2670,n2681);
and (n2670,n2671,n2680);
xor (n2671,n2672,n2673);
xor (n2672,n2584,n2594);
or (n2673,n2674,n2679);
and (n2674,n2675,n2678);
xor (n2675,n2676,n2677);
xor (n2676,n2588,n2592);
wire s0n2677,s1n2677,notn2677;
or (n2677,s0n2677,s1n2677);
not(notn2677,n982);
and (s0n2677,notn2677,1'b0);
and (s1n2677,n982,n2508);
and (n2678,n2471,n982);
and (n2679,n2676,n2677);
xor (n2680,n2605,n2614);
and (n2681,n2672,n2673);
xor (n2682,n2601,n2616);
and (n2683,n2668,n2669);
or (n2684,n2685,n2696);
and (n2685,n2686,n2695);
xor (n2686,n2687,n2694);
or (n2687,n2688,n2693);
and (n2688,n2689,n2692);
xor (n2689,n2690,n2691);
and (n2690,n2400,n982);
xor (n2691,n2451,n2465);
and (n2692,n2403,n982);
and (n2693,n2690,n2691);
xor (n2694,n2506,n2516);
xor (n2695,n2568,n2571);
and (n2696,n2687,n2694);
xor (n2697,n2577,n2599);
and (n2698,n2665,n2684);
xor (n2699,n2648,n2657);
or (n2700,n2701,n2702);
xor (n2701,n2664,n2697);
xor (n2702,n2651,n2654);
nand (n2703,n2704,n2725);
or (n2704,n2705,n2708);
nor (n2705,n2706,n2707);
xor (n2706,n2667,n2682);
xor (n2707,n2686,n2695);
nand (n2708,n2709,n2712,n2715);
or (n2709,n2710,n2711);
xor (n2710,n2689,n2692);
xor (n2711,n2671,n2680);
or (n2712,n2713,n2714);
xor (n2713,n2609,n2612);
xor (n2714,n2675,n2678);
nand (n2715,n2716,n2719);
or (n2716,n2717,n2718);
not (n2717,n2713);
not (n2718,n2714);
nor (n2719,n2720,n2724);
and (n2720,n2721,n2722);
xor (n2721,n2036,n2590);
or (n2722,n2723,n2032);
wire s0n2723,s1n2723,notn2723;
or (n2723,s0n2723,s1n2723);
not(notn2723,n982);
and (s0n2723,notn2723,1'b0);
and (s1n2723,n982,n2329);
and (n2724,n2723,n2032);
nor (n2725,n2726,n2728);
and (n2726,n2727,n2710,n2711);
not (n2727,n2705);
and (n2728,n2706,n2707);
nor (n2729,n2730,n2734);
and (n2730,n2699,n2731);
nand (n2731,n2732,n2733);
not (n2732,n2662);
nand (n2733,n2701,n2702);
and (n2734,n2735,n2662);
not (n2735,n2733);
nand (n2736,n2645,n2646);
nand (n2737,n2628,n2629);
and (n2738,n2550,n2624);
and (n2739,n2486,n2546);
and (n2740,n2376,n2377);
and (n2741,n2289,n2290);
and (n2742,n3,n2215);
or (n2743,n2744,n2775);
not (n2744,n2745);
nand (n2745,n2746,n2774);
or (n2746,n2747,n2770);
not (n2747,n2748);
nand (n2748,n2749,n2753);
not (n2749,n2750);
or (n2750,n2751,n2752);
and (n2751,n2154,n2173);
and (n2752,n2155,n2158);
nor (n2753,n2754,n2769);
not (n2754,n2755);
nor (n2755,n2756,n2766);
not (n2756,n2757);
nor (n2757,n2758,n2759);
and (n2758,n2169,n2172);
not (n2759,n2760);
nor (n2760,n2761,n2762);
and (n2761,n2164,n2167);
not (n2762,n2763);
xnor (n2763,n2764,n2765);
wire s0n2764,s1n2764,notn2764;
or (n2764,s0n2764,s1n2764);
not(notn2764,n1425);
and (s0n2764,notn2764,1'b0);
and (s1n2764,n1425,n14);
wire s0n2765,s1n2765,notn2765;
or (n2765,s0n2765,s1n2765);
not(notn2765,n1425);
and (s0n2765,notn2765,1'b0);
and (s1n2765,n1425,n1738);
or (n2766,n2767,n2768);
and (n2767,n2159,n2168);
and (n2768,n2160,n2163);
and (n2769,n2123,n2150);
not (n2770,n2771);
or (n2771,n2772,n2773);
and (n2772,n4,n2153);
and (n2773,n5,n2122);
or (n2774,n2771,n2748);
not (n2775,n0);
endmodule
