module top (out,n6,n8,n9,n13,n21,n22,n29,n43,n62
        ,n64,n73,n74,n98,n99,n111,n164,n165,n169,n174
        ,n194,n196,n212,n266,n298,n427,n441,n442,n514,n523
        ,n524,n560,n632,n662,n663,n853,n857,n859,n885,n886
        ,n993,n1010,n1011,n1197,n1201,n1203,n1214,n1226,n1240);
output out;
input n6;
input n8;
input n9;
input n13;
input n21;
input n22;
input n29;
input n43;
input n62;
input n64;
input n73;
input n74;
input n98;
input n99;
input n111;
input n164;
input n165;
input n169;
input n174;
input n194;
input n196;
input n212;
input n266;
input n298;
input n427;
input n441;
input n442;
input n514;
input n523;
input n524;
input n560;
input n632;
input n662;
input n663;
input n853;
input n857;
input n859;
input n885;
input n886;
input n993;
input n1010;
input n1011;
input n1197;
input n1201;
input n1203;
input n1214;
input n1226;
input n1240;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n7;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n166;
wire n167;
wire n168;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n854;
wire n855;
wire n856;
wire n858;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1198;
wire n1199;
wire n1200;
wire n1202;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
xnor (out,n0,n3142);
nand (n0,n1,n46);
nand (n1,n2,n32);
xor (n2,n3,n14);
not (n3,n4);
or (n4,n5,n10);
and (n5,n6,n7);
xor (n7,n8,n9);
and (n10,n6,n11);
nor (n11,n7,n12);
xnor (n12,n13,n8);
nand (n14,n15,n30,n31);
nand (n15,n16,n26);
not (n16,n17);
xor (n17,n18,n9);
or (n18,n19,n23);
and (n19,n6,n20);
xor (n20,n21,n22);
and (n23,n6,n24);
nor (n24,n20,n25);
xnor (n25,n9,n21);
xor (n26,n27,n13);
or (n27,n5,n28);
and (n28,n29,n11);
nand (n30,n13,n26);
nand (n31,n16,n13);
nand (n32,n33,n36,n45);
nand (n33,n17,n34);
xor (n34,n35,n13);
xor (n35,n16,n26);
nand (n36,n37,n34);
nand (n37,n38,n31,n44);
nand (n38,n39,n13);
xor (n39,n40,n13);
or (n40,n41,n42);
and (n41,n29,n7);
and (n42,n43,n11);
nand (n44,n39,n16);
nand (n45,n17,n37);
nand (n46,n47,n3140);
nand (n47,n48,n144);
nor (n48,n49,n142);
nor (n49,n50,n135);
nand (n50,n51,n124);
nand (n51,n52,n88,n123);
nand (n52,n53,n67);
nand (n53,n54,n65,n66);
nand (n54,n55,n59);
xor (n55,n56,n9);
or (n56,n57,n58);
and (n57,n29,n20);
and (n58,n43,n24);
xor (n59,n60,n13);
or (n60,n61,n63);
and (n61,n62,n7);
and (n63,n64,n11);
nand (n65,n13,n59);
nand (n66,n55,n13);
xor (n67,n68,n78);
xor (n68,n13,n69);
xor (n69,n70,n22);
or (n70,n71,n75);
and (n71,n6,n72);
xor (n72,n73,n74);
and (n75,n6,n76);
nor (n76,n72,n77);
xnor (n77,n22,n73);
xor (n78,n79,n84);
xor (n79,n80,n81);
not (n80,n69);
xor (n81,n82,n9);
or (n82,n19,n83);
and (n83,n29,n24);
xor (n84,n85,n13);
or (n85,n86,n87);
and (n86,n43,n7);
and (n87,n62,n11);
nand (n88,n89,n67);
nand (n89,n90,n113,n122);
nand (n90,n80,n91);
nand (n91,n92,n106,n112);
nand (n92,n93,n103);
not (n93,n94);
xor (n94,n95,n74);
or (n95,n96,n100);
and (n96,n6,n97);
xor (n97,n98,n99);
and (n100,n6,n101);
nor (n101,n97,n102);
xnor (n102,n74,n98);
xor (n103,n104,n22);
or (n104,n71,n105);
and (n105,n29,n76);
nand (n106,n107,n103);
xor (n107,n108,n13);
or (n108,n109,n110);
and (n109,n64,n7);
and (n110,n111,n11);
nand (n112,n93,n107);
nand (n113,n114,n91);
nand (n114,n115,n120,n121);
nand (n115,n116,n13);
xor (n116,n117,n9);
or (n117,n118,n119);
and (n118,n43,n20);
and (n119,n62,n24);
nand (n120,n94,n13);
nand (n121,n116,n94);
nand (n122,n80,n114);
nand (n123,n53,n89);
xor (n124,n125,n131);
xor (n125,n126,n130);
nand (n126,n127,n128,n129);
nand (n127,n80,n81);
nand (n128,n84,n81);
nand (n129,n80,n84);
xor (n130,n40,n16);
nand (n131,n132,n133,n134);
nand (n132,n13,n69);
nand (n133,n78,n69);
nand (n134,n13,n78);
nor (n135,n136,n138);
xor (n136,n137,n37);
not (n137,n27);
nand (n138,n139,n140,n141);
nand (n139,n126,n130);
nand (n140,n131,n130);
nand (n141,n126,n131);
not (n142,n143);
nand (n143,n136,n138);
nand (n144,n145,n147);
nor (n145,n146,n135);
nor (n146,n51,n124);
nand (n147,n148,n402);
nor (n148,n149,n396);
nor (n149,n150,n372);
nor (n150,n151,n370);
nor (n151,n152,n345);
nand (n152,n153,n309);
nand (n153,n154,n255,n308);
nand (n154,n155,n214);
nand (n155,n156,n198,n213);
nand (n156,n157,n184);
nand (n157,n158,n178,n183);
nand (n158,n159,n170);
not (n159,n160);
xor (n160,n161,n169);
or (n161,n162,n166);
and (n162,n6,n163);
xor (n163,n164,n165);
and (n166,n6,n167);
nor (n167,n163,n168);
xnor (n168,n169,n164);
xor (n170,n171,n99);
or (n171,n172,n175);
and (n172,n6,n173);
xor (n173,n174,n169);
and (n175,n29,n176);
nor (n176,n173,n177);
xnor (n177,n99,n174);
nand (n178,n179,n170);
xor (n179,n180,n74);
or (n180,n181,n182);
and (n181,n43,n97);
and (n182,n62,n101);
nand (n183,n159,n179);
nand (n184,n185,n190,n197);
nand (n185,n186,n160);
xor (n186,n187,n22);
or (n187,n188,n189);
and (n188,n64,n72);
and (n189,n111,n76);
nand (n190,n191,n160);
xor (n191,n192,n9);
or (n192,n193,n195);
and (n193,n194,n20);
and (n195,n196,n24);
nand (n197,n186,n191);
nand (n198,n199,n184);
xor (n199,n200,n208);
xor (n200,n201,n204);
xor (n201,n202,n99);
or (n202,n172,n203);
and (n203,n6,n176);
xor (n204,n205,n9);
or (n205,n206,n207);
and (n206,n111,n20);
and (n207,n194,n24);
xor (n208,n209,n13);
or (n209,n210,n211);
and (n210,n196,n7);
and (n211,n212,n11);
nand (n213,n157,n199);
xor (n214,n215,n239);
xor (n215,n216,n229);
nand (n216,n217,n227,n228);
nand (n217,n218,n222);
xor (n218,n219,n22);
or (n219,n220,n221);
and (n220,n62,n72);
and (n221,n64,n76);
not (n222,n223);
xor (n223,n224,n74);
or (n224,n225,n226);
and (n225,n29,n97);
and (n226,n43,n101);
nand (n227,n13,n222);
nand (n228,n218,n13);
xor (n229,n230,n13);
xor (n230,n231,n235);
xor (n231,n232,n13);
or (n232,n233,n234);
and (n233,n194,n7);
and (n234,n196,n11);
xor (n235,n236,n22);
or (n236,n237,n238);
and (n237,n43,n72);
and (n238,n62,n76);
xor (n239,n240,n245);
xor (n240,n223,n241);
nand (n241,n242,n243,n244);
nand (n242,n201,n204);
nand (n243,n208,n204);
nand (n244,n201,n208);
xor (n245,n246,n251);
xor (n246,n247,n248);
not (n247,n201);
xor (n248,n249,n74);
or (n249,n96,n250);
and (n250,n29,n101);
xor (n251,n252,n9);
or (n252,n253,n254);
and (n253,n64,n20);
and (n254,n111,n24);
nand (n255,n256,n214);
nand (n256,n257,n285,n307);
nand (n257,n258,n260);
xor (n258,n259,n13);
xor (n259,n218,n222);
nand (n260,n261,n267,n284);
nand (n261,n262,n13);
xor (n262,n263,n13);
or (n263,n264,n265);
and (n264,n212,n7);
and (n265,n266,n11);
nand (n267,n268,n13);
nand (n268,n269,n278,n283);
nand (n269,n270,n274);
xor (n270,n271,n99);
or (n271,n272,n273);
and (n272,n29,n173);
and (n273,n43,n176);
xor (n274,n275,n74);
or (n275,n276,n277);
and (n276,n62,n97);
and (n277,n64,n101);
nand (n278,n279,n274);
xor (n279,n280,n22);
or (n280,n281,n282);
and (n281,n111,n72);
and (n282,n194,n76);
nand (n283,n270,n279);
nand (n284,n262,n268);
nand (n285,n286,n260);
nand (n286,n287,n303,n306);
nand (n287,n288,n301);
nand (n288,n289,n299,n300);
nand (n289,n290,n294);
xor (n290,n291,n9);
or (n291,n292,n293);
and (n292,n196,n20);
and (n293,n212,n24);
xor (n294,n295,n13);
or (n295,n296,n297);
and (n296,n266,n7);
and (n297,n298,n11);
nand (n299,n159,n294);
nand (n300,n290,n159);
xor (n301,n302,n179);
xor (n302,n159,n170);
nand (n303,n304,n301);
xor (n304,n305,n191);
xor (n305,n186,n160);
nand (n306,n288,n304);
nand (n307,n258,n286);
nand (n308,n155,n256);
xor (n309,n310,n341);
xor (n310,n311,n315);
nand (n311,n312,n313,n314);
nand (n312,n223,n241);
nand (n313,n245,n241);
nand (n314,n223,n245);
xor (n315,n316,n335);
xor (n316,n317,n331);
xor (n317,n318,n327);
xor (n318,n319,n323);
xor (n319,n320,n22);
or (n320,n321,n322);
and (n321,n29,n72);
and (n322,n43,n76);
xor (n323,n324,n13);
or (n324,n325,n326);
and (n325,n111,n7);
and (n326,n194,n11);
xor (n327,n328,n9);
or (n328,n329,n330);
and (n329,n62,n20);
and (n330,n64,n24);
nand (n331,n332,n333,n334);
nand (n332,n231,n235);
nand (n333,n13,n235);
nand (n334,n231,n13);
xor (n335,n336,n337);
xor (n336,n93,n13);
nand (n337,n338,n339,n340);
nand (n338,n247,n248);
nand (n339,n251,n248);
nand (n340,n247,n251);
nand (n341,n342,n343,n344);
nand (n342,n216,n229);
nand (n343,n239,n229);
nand (n344,n216,n239);
nor (n345,n346,n366);
xor (n346,n347,n362);
xor (n347,n348,n352);
nand (n348,n349,n350,n351);
nand (n349,n93,n13);
nand (n350,n337,n13);
nand (n351,n93,n337);
xor (n352,n353,n360);
xor (n353,n354,n358);
nand (n354,n355,n356,n357);
nand (n355,n319,n323);
nand (n356,n327,n323);
nand (n357,n319,n327);
xor (n358,n359,n107);
xor (n359,n93,n103);
xor (n360,n361,n94);
xor (n361,n116,n13);
nand (n362,n363,n364,n365);
nand (n363,n317,n331);
nand (n364,n335,n331);
nand (n365,n317,n335);
nand (n366,n367,n368,n369);
nand (n367,n311,n315);
nand (n368,n341,n315);
nand (n369,n311,n341);
not (n370,n371);
nand (n371,n346,n366);
not (n372,n373);
nor (n373,n374,n389);
nor (n374,n375,n385);
xor (n375,n376,n381);
xor (n376,n377,n379);
xor (n377,n378,n13);
xor (n378,n55,n59);
xor (n379,n380,n114);
xor (n380,n80,n91);
nand (n381,n382,n383,n384);
nand (n382,n354,n358);
nand (n383,n360,n358);
nand (n384,n354,n360);
nand (n385,n386,n387,n388);
nand (n386,n348,n352);
nand (n387,n362,n352);
nand (n388,n348,n362);
nor (n389,n390,n394);
nand (n390,n391,n392,n393);
nand (n391,n377,n379);
nand (n392,n381,n379);
nand (n393,n377,n381);
xor (n394,n395,n89);
xor (n395,n53,n67);
not (n396,n397);
nor (n397,n398,n400);
nor (n398,n399,n389);
nand (n399,n375,n385);
not (n400,n401);
nand (n401,n390,n394);
nand (n402,n403,n3136);
nand (n403,n404,n1174);
nor (n404,n405,n1159);
nor (n405,n406,n752);
nand (n406,n407,n729);
nor (n407,n408,n705);
nor (n408,n409,n582);
xor (n409,n410,n539);
xor (n410,n411,n430);
xor (n411,n412,n417);
xor (n412,n413,n415);
xor (n413,n414,n279);
xor (n414,n270,n274);
xor (n415,n416,n159);
xor (n416,n290,n294);
nand (n417,n418,n428,n429);
nand (n418,n419,n423);
xor (n419,n420,n9);
or (n420,n421,n422);
and (n421,n212,n20);
and (n422,n266,n24);
xor (n423,n424,n13);
or (n424,n425,n426);
and (n425,n298,n7);
and (n426,n427,n11);
nand (n428,n13,n423);
nand (n429,n419,n13);
xor (n430,n431,n501);
xor (n431,n432,n467);
xor (n432,n433,n455);
xor (n433,n13,n434);
nand (n434,n435,n449,n454);
nand (n435,n436,n446);
not (n436,n437);
xor (n437,n438,n165);
or (n438,n439,n443);
and (n439,n6,n440);
xor (n440,n441,n442);
and (n443,n6,n444);
nor (n444,n440,n445);
xnor (n445,n165,n441);
xor (n446,n447,n169);
or (n447,n162,n448);
and (n448,n29,n167);
nand (n449,n450,n446);
xor (n450,n451,n74);
or (n451,n452,n453);
and (n452,n64,n97);
and (n453,n111,n101);
nand (n454,n436,n450);
nand (n455,n456,n461,n466);
nand (n456,n457,n437);
xor (n457,n458,n99);
or (n458,n459,n460);
and (n459,n43,n173);
and (n460,n62,n176);
nand (n461,n462,n437);
xor (n462,n463,n22);
or (n463,n464,n465);
and (n464,n194,n72);
and (n465,n196,n76);
nand (n466,n457,n462);
nand (n467,n468,n487,n500);
nand (n468,n469,n471);
xor (n469,n470,n450);
xor (n470,n436,n446);
nand (n471,n472,n481,n486);
nand (n472,n473,n477);
xor (n473,n474,n169);
or (n474,n475,n476);
and (n475,n29,n163);
and (n476,n43,n167);
xor (n477,n478,n74);
or (n478,n479,n480);
and (n479,n111,n97);
and (n480,n194,n101);
nand (n481,n482,n477);
xor (n482,n483,n99);
or (n483,n484,n485);
and (n484,n62,n173);
and (n485,n64,n176);
nand (n486,n473,n482);
nand (n487,n488,n471);
nand (n488,n489,n494,n499);
nand (n489,n436,n490);
xor (n490,n491,n22);
or (n491,n492,n493);
and (n492,n196,n72);
and (n493,n212,n76);
nand (n494,n495,n490);
xor (n495,n496,n9);
or (n496,n497,n498);
and (n497,n266,n20);
and (n498,n298,n24);
nand (n499,n436,n495);
nand (n500,n469,n488);
nand (n501,n502,n507,n538);
nand (n502,n503,n505);
xor (n503,n504,n13);
xor (n504,n419,n423);
xor (n505,n506,n462);
xor (n506,n457,n437);
nand (n507,n508,n505);
nand (n508,n509,n515,n537);
nand (n509,n510,n13);
xor (n510,n511,n13);
or (n511,n512,n513);
and (n512,n427,n7);
and (n513,n514,n11);
nand (n515,n516,n13);
nand (n516,n517,n531,n536);
nand (n517,n518,n528);
not (n518,n519);
xor (n519,n520,n442);
or (n520,n521,n525);
and (n521,n6,n522);
xor (n522,n523,n524);
and (n525,n6,n526);
nor (n526,n522,n527);
xnor (n527,n442,n523);
xor (n528,n529,n165);
or (n529,n439,n530);
and (n530,n29,n444);
nand (n531,n532,n528);
xor (n532,n533,n169);
or (n533,n534,n535);
and (n534,n43,n163);
and (n535,n62,n167);
nand (n536,n518,n532);
nand (n537,n510,n516);
nand (n538,n503,n508);
nand (n539,n540,n578,n581);
nand (n540,n541,n576);
nand (n541,n542,n562,n575);
nand (n542,n543,n545);
xor (n543,n544,n482);
xor (n544,n473,n477);
nand (n545,n546,n555,n561);
nand (n546,n547,n551);
xor (n547,n548,n99);
or (n548,n549,n550);
and (n549,n64,n173);
and (n550,n111,n176);
xor (n551,n552,n74);
or (n552,n553,n554);
and (n553,n194,n97);
and (n554,n196,n101);
nand (n555,n556,n551);
xor (n556,n557,n13);
or (n557,n558,n559);
and (n558,n514,n7);
and (n559,n560,n11);
nand (n561,n547,n556);
nand (n562,n563,n545);
nand (n563,n564,n569,n574);
nand (n564,n519,n565);
xor (n565,n566,n22);
or (n566,n567,n568);
and (n567,n212,n72);
and (n568,n266,n76);
nand (n569,n570,n565);
xor (n570,n571,n9);
or (n571,n572,n573);
and (n572,n298,n20);
and (n573,n427,n24);
nand (n574,n519,n570);
nand (n575,n543,n563);
xor (n576,n577,n488);
xor (n577,n469,n471);
nand (n578,n579,n576);
xor (n579,n580,n508);
xor (n580,n503,n505);
nand (n581,n541,n579);
nand (n582,n583,n615,n704);
nand (n583,n584,n613);
nand (n584,n585,n589,n612);
nand (n585,n586,n588);
xor (n586,n587,n495);
xor (n587,n436,n490);
xor (n588,n511,n516);
nand (n589,n590,n588);
nand (n590,n591,n594,n611);
nand (n591,n13,n592);
xor (n592,n593,n532);
xor (n593,n518,n528);
nand (n594,n595,n592);
nand (n595,n596,n605,n610);
nand (n596,n597,n601);
xor (n597,n598,n165);
or (n598,n599,n600);
and (n599,n29,n440);
and (n600,n43,n444);
xor (n601,n602,n169);
or (n602,n603,n604);
and (n603,n62,n163);
and (n604,n64,n167);
nand (n605,n606,n601);
xor (n606,n607,n99);
or (n607,n608,n609);
and (n608,n111,n173);
and (n609,n194,n176);
nand (n610,n597,n606);
nand (n611,n13,n595);
nand (n612,n586,n590);
xor (n613,n614,n579);
xor (n614,n541,n576);
nand (n615,n616,n613);
nand (n616,n617,n641,n703);
nand (n617,n618,n620);
xor (n618,n619,n563);
xor (n619,n543,n545);
nand (n620,n621,n637,n640);
nand (n621,n622,n635);
nand (n622,n623,n633,n634);
nand (n623,n624,n628);
xor (n624,n625,n74);
or (n625,n626,n627);
and (n626,n196,n97);
and (n627,n212,n101);
xor (n628,n629,n13);
or (n629,n630,n631);
and (n630,n560,n7);
and (n631,n632,n11);
nand (n633,n518,n628);
nand (n634,n624,n518);
xor (n635,n636,n556);
xor (n636,n547,n551);
nand (n637,n638,n635);
xor (n638,n639,n570);
xor (n639,n519,n565);
nand (n640,n622,n638);
nand (n641,n642,n620);
nand (n642,n643,n699,n702);
nand (n643,n644,n677);
nand (n644,n645,n654,n676);
nand (n645,n646,n650);
xor (n646,n647,n22);
or (n647,n648,n649);
and (n648,n266,n72);
and (n649,n298,n76);
xor (n650,n651,n9);
or (n651,n652,n653);
and (n652,n427,n20);
and (n653,n514,n24);
nand (n654,n655,n650);
nand (n655,n656,n670,n675);
nand (n656,n657,n667);
not (n657,n658);
xor (n658,n659,n524);
or (n659,n660,n664);
and (n660,n6,n661);
xor (n661,n662,n663);
and (n664,n6,n665);
nor (n665,n661,n666);
xnor (n666,n524,n662);
xor (n667,n668,n442);
or (n668,n521,n669);
and (n669,n29,n526);
nand (n670,n671,n667);
xor (n671,n672,n169);
or (n672,n673,n674);
and (n673,n64,n163);
and (n674,n111,n167);
nand (n675,n657,n671);
nand (n676,n646,n655);
nand (n677,n678,n681,n698);
nand (n678,n13,n679);
xor (n679,n680,n606);
xor (n680,n597,n601);
nand (n681,n682,n679);
nand (n682,n683,n692,n697);
nand (n683,n684,n688);
xor (n684,n685,n165);
or (n685,n686,n687);
and (n686,n43,n440);
and (n687,n62,n444);
xor (n688,n689,n99);
or (n689,n690,n691);
and (n690,n194,n173);
and (n691,n196,n176);
nand (n692,n693,n688);
xor (n693,n694,n74);
or (n694,n695,n696);
and (n695,n212,n97);
and (n696,n266,n101);
nand (n697,n684,n693);
nand (n698,n13,n682);
nand (n699,n700,n677);
xor (n700,n701,n595);
xor (n701,n13,n592);
nand (n702,n644,n700);
nand (n703,n618,n642);
nand (n704,n584,n616);
nor (n705,n706,n710);
nand (n706,n707,n708,n709);
nand (n707,n411,n430);
nand (n708,n539,n430);
nand (n709,n411,n539);
xor (n710,n711,n725);
xor (n711,n712,n716);
nand (n712,n713,n714,n715);
nand (n713,n413,n415);
nand (n714,n417,n415);
nand (n715,n413,n417);
xor (n716,n717,n723);
xor (n717,n718,n722);
nand (n718,n719,n720,n721);
nand (n719,n13,n434);
nand (n720,n455,n434);
nand (n721,n13,n455);
xor (n722,n263,n268);
xor (n723,n724,n304);
xor (n724,n288,n301);
nand (n725,n726,n727,n728);
nand (n726,n432,n467);
nand (n727,n501,n467);
nand (n728,n432,n501);
nor (n729,n730,n745);
nor (n730,n731,n735);
nand (n731,n732,n733,n734);
nand (n732,n712,n716);
nand (n733,n725,n716);
nand (n734,n712,n725);
xor (n735,n736,n741);
xor (n736,n737,n739);
xor (n737,n738,n199);
xor (n738,n157,n184);
xor (n739,n740,n286);
xor (n740,n258,n260);
nand (n741,n742,n743,n744);
nand (n742,n718,n722);
nand (n743,n723,n722);
nand (n744,n718,n723);
nor (n745,n746,n750);
nand (n746,n747,n748,n749);
nand (n747,n737,n739);
nand (n748,n741,n739);
nand (n749,n737,n741);
xor (n750,n751,n256);
xor (n751,n155,n214);
nor (n752,n753,n1153);
nor (n753,n754,n1129);
nor (n754,n755,n1127);
nor (n755,n756,n1102);
nand (n756,n757,n1064);
nand (n757,n758,n980,n1063);
nand (n758,n759,n843);
xor (n759,n760,n833);
xor (n760,n761,n783);
xor (n761,n762,n767);
xor (n762,n763,n13);
xor (n763,n764,n22);
or (n764,n765,n766);
and (n765,n298,n72);
and (n766,n427,n76);
nand (n767,n768,n777,n782);
nand (n768,n769,n773);
xor (n769,n770,n169);
or (n770,n771,n772);
and (n771,n111,n163);
and (n772,n194,n167);
xor (n773,n774,n442);
or (n774,n775,n776);
and (n775,n29,n522);
and (n776,n43,n526);
nand (n777,n778,n773);
xor (n778,n779,n165);
or (n779,n780,n781);
and (n780,n62,n440);
and (n781,n64,n444);
nand (n782,n769,n778);
nand (n783,n784,n815,n832);
nand (n784,n785,n801);
nand (n785,n786,n795,n800);
nand (n786,n787,n791);
xor (n787,n788,n169);
or (n788,n789,n790);
and (n789,n194,n163);
and (n790,n196,n167);
xor (n791,n792,n442);
or (n792,n793,n794);
and (n793,n43,n522);
and (n794,n62,n526);
nand (n795,n796,n791);
xor (n796,n797,n99);
or (n797,n798,n799);
and (n798,n212,n173);
and (n799,n266,n176);
nand (n800,n787,n796);
xor (n801,n802,n811);
xor (n802,n803,n807);
xor (n803,n804,n99);
or (n804,n805,n806);
and (n805,n196,n173);
and (n806,n212,n176);
xor (n807,n808,n74);
or (n808,n809,n810);
and (n809,n266,n97);
and (n810,n298,n101);
xor (n811,n812,n9);
or (n812,n813,n814);
and (n813,n560,n20);
and (n814,n632,n24);
nand (n815,n816,n801);
nand (n816,n817,n826,n831);
nand (n817,n818,n822);
xor (n818,n819,n524);
or (n819,n820,n821);
and (n820,n29,n661);
and (n821,n43,n665);
xor (n822,n823,n74);
or (n823,n824,n825);
and (n824,n298,n97);
and (n825,n427,n101);
nand (n826,n827,n822);
xor (n827,n828,n22);
or (n828,n829,n830);
and (n829,n514,n72);
and (n830,n560,n76);
nand (n831,n818,n827);
nand (n832,n785,n816);
xor (n833,n834,n839);
xor (n834,n835,n837);
xor (n835,n836,n671);
xor (n836,n657,n667);
xor (n837,n838,n693);
xor (n838,n684,n688);
nand (n839,n840,n841,n842);
nand (n840,n803,n807);
nand (n841,n811,n807);
nand (n842,n803,n811);
xor (n843,n844,n919);
xor (n844,n845,n899);
nand (n845,n846,n872,n898);
nand (n846,n847,n862);
nand (n847,n848,n860,n861);
nand (n848,n849,n854);
xor (n849,n850,n9);
or (n850,n851,n852);
and (n851,n632,n20);
and (n852,n853,n24);
xor (n854,n855,n13);
or (n855,n856,n858);
and (n856,n857,n7);
and (n858,n859,n11);
nand (n860,n13,n854);
nand (n861,n849,n13);
xor (n862,n863,n868);
xor (n863,n864,n657);
xor (n864,n865,n13);
or (n865,n866,n867);
and (n866,n853,n7);
and (n867,n857,n11);
xor (n868,n869,n22);
or (n869,n870,n871);
and (n870,n427,n72);
and (n871,n514,n76);
nand (n872,n873,n862);
xor (n873,n874,n896);
xor (n874,n13,n875);
nand (n875,n876,n890,n895);
nand (n876,n877,n880);
xor (n877,n878,n524);
or (n878,n660,n879);
and (n879,n29,n665);
not (n880,n881);
xor (n881,n882,n663);
or (n882,n883,n887);
and (n883,n6,n884);
xor (n884,n885,n886);
and (n887,n6,n888);
nor (n888,n884,n889);
xnor (n889,n663,n885);
nand (n890,n891,n880);
xor (n891,n892,n165);
or (n892,n893,n894);
and (n893,n64,n440);
and (n894,n111,n444);
nand (n895,n877,n891);
xor (n896,n897,n778);
xor (n897,n769,n773);
nand (n898,n847,n873);
xor (n899,n900,n915);
xor (n900,n901,n905);
nand (n901,n902,n903,n904);
nand (n902,n864,n657);
nand (n903,n868,n657);
nand (n904,n864,n868);
xor (n905,n906,n658);
xor (n906,n907,n911);
xor (n907,n908,n9);
or (n908,n909,n910);
and (n909,n514,n20);
and (n910,n560,n24);
xor (n911,n912,n13);
or (n912,n913,n914);
and (n913,n632,n7);
and (n914,n853,n11);
nand (n915,n916,n917,n918);
nand (n916,n13,n875);
nand (n917,n896,n875);
nand (n918,n13,n896);
nand (n919,n920,n976,n979);
nand (n920,n921,n941);
nand (n921,n922,n937,n940);
nand (n922,n923,n935);
nand (n923,n924,n929,n934);
nand (n924,n881,n925);
xor (n925,n926,n165);
or (n926,n927,n928);
and (n927,n111,n440);
and (n928,n194,n444);
nand (n929,n930,n925);
xor (n930,n931,n169);
or (n931,n932,n933);
and (n932,n196,n163);
and (n933,n212,n167);
nand (n934,n881,n930);
xor (n935,n936,n796);
xor (n936,n787,n791);
nand (n937,n938,n935);
xor (n938,n939,n891);
xor (n939,n877,n880);
nand (n940,n923,n938);
nand (n941,n942,n972,n975);
nand (n942,n943,n956);
nand (n943,n944,n950,n955);
nand (n944,n945,n949);
xor (n945,n946,n442);
or (n946,n947,n948);
and (n947,n62,n522);
and (n948,n64,n526);
not (n949,n818);
nand (n950,n951,n949);
xor (n951,n952,n99);
or (n952,n953,n954);
and (n953,n266,n173);
and (n954,n298,n176);
nand (n955,n945,n951);
nand (n956,n957,n966,n971);
nand (n957,n958,n962);
xor (n958,n959,n74);
or (n959,n960,n961);
and (n960,n427,n97);
and (n961,n514,n101);
xor (n962,n963,n22);
or (n963,n964,n965);
and (n964,n560,n72);
and (n965,n632,n76);
nand (n966,n967,n962);
xor (n967,n968,n9);
or (n968,n969,n970);
and (n969,n853,n20);
and (n970,n857,n24);
nand (n971,n958,n967);
nand (n972,n973,n956);
xor (n973,n974,n827);
xor (n974,n818,n822);
nand (n975,n943,n973);
nand (n976,n977,n941);
xor (n977,n978,n816);
xor (n978,n785,n801);
nand (n979,n921,n977);
nand (n980,n981,n843);
nand (n981,n982,n1059,n1062);
nand (n982,n983,n985);
xor (n983,n984,n873);
xor (n984,n847,n862);
nand (n985,n986,n1019,n1058);
nand (n986,n987,n1017);
nand (n987,n988,n994,n1016);
nand (n988,n989,n13);
xor (n989,n990,n13);
or (n990,n991,n992);
and (n991,n859,n7);
and (n992,n993,n11);
nand (n994,n995,n13);
nand (n995,n996,n1004,n1015);
nand (n996,n997,n1000);
xor (n997,n998,n663);
or (n998,n883,n999);
and (n999,n29,n888);
xor (n1000,n1001,n524);
or (n1001,n1002,n1003);
and (n1002,n43,n661);
and (n1003,n62,n665);
nand (n1004,n1005,n1000);
not (n1005,n1006);
xor (n1006,n1007,n886);
or (n1007,n1008,n1012);
and (n1008,n6,n1009);
xor (n1009,n1010,n1011);
and (n1012,n6,n1013);
nor (n1013,n1009,n1014);
xnor (n1014,n886,n1010);
nand (n1015,n997,n1005);
nand (n1016,n989,n995);
xor (n1017,n1018,n13);
xor (n1018,n849,n854);
nand (n1019,n1020,n1017);
nand (n1020,n1021,n1040,n1057);
nand (n1021,n1022,n1038);
nand (n1022,n1023,n1032,n1037);
nand (n1023,n1024,n1028);
xor (n1024,n1025,n442);
or (n1025,n1026,n1027);
and (n1026,n64,n522);
and (n1027,n111,n526);
xor (n1028,n1029,n165);
or (n1029,n1030,n1031);
and (n1030,n194,n440);
and (n1031,n196,n444);
nand (n1032,n1033,n1028);
xor (n1033,n1034,n169);
or (n1034,n1035,n1036);
and (n1035,n212,n163);
and (n1036,n266,n167);
nand (n1037,n1024,n1033);
xor (n1038,n1039,n930);
xor (n1039,n881,n925);
nand (n1040,n1041,n1038);
nand (n1041,n1042,n1051,n1056);
nand (n1042,n1043,n1047);
xor (n1043,n1044,n74);
or (n1044,n1045,n1046);
and (n1045,n514,n97);
and (n1046,n560,n101);
xor (n1047,n1048,n663);
or (n1048,n1049,n1050);
and (n1049,n29,n884);
and (n1050,n43,n888);
nand (n1051,n1052,n1047);
xor (n1052,n1053,n99);
or (n1053,n1054,n1055);
and (n1054,n298,n173);
and (n1055,n427,n176);
nand (n1056,n1043,n1052);
nand (n1057,n1022,n1041);
nand (n1058,n987,n1020);
nand (n1059,n1060,n985);
xor (n1060,n1061,n977);
xor (n1061,n921,n941);
nand (n1062,n983,n1060);
nand (n1063,n759,n981);
xor (n1064,n1065,n1098);
xor (n1065,n1066,n1070);
nand (n1066,n1067,n1068,n1069);
nand (n1067,n761,n783);
nand (n1068,n833,n783);
nand (n1069,n761,n833);
xor (n1070,n1071,n1086);
xor (n1071,n1072,n1076);
nand (n1072,n1073,n1074,n1075);
nand (n1073,n901,n905);
nand (n1074,n915,n905);
nand (n1075,n901,n915);
xor (n1076,n1077,n1084);
xor (n1077,n1078,n1082);
nand (n1078,n1079,n1080,n1081);
nand (n1079,n907,n911);
nand (n1080,n658,n911);
nand (n1081,n907,n658);
xor (n1082,n1083,n655);
xor (n1083,n646,n650);
xor (n1084,n1085,n518);
xor (n1085,n624,n628);
xor (n1086,n1087,n1094);
xor (n1087,n1088,n1092);
nand (n1088,n1089,n1090,n1091);
nand (n1089,n763,n13);
nand (n1090,n767,n13);
nand (n1091,n763,n767);
xor (n1092,n1093,n682);
xor (n1093,n13,n679);
nand (n1094,n1095,n1096,n1097);
nand (n1095,n835,n837);
nand (n1096,n839,n837);
nand (n1097,n835,n839);
nand (n1098,n1099,n1100,n1101);
nand (n1099,n845,n899);
nand (n1100,n919,n899);
nand (n1101,n845,n919);
nor (n1102,n1103,n1107);
nand (n1103,n1104,n1105,n1106);
nand (n1104,n1066,n1070);
nand (n1105,n1098,n1070);
nand (n1106,n1066,n1098);
xor (n1107,n1108,n1123);
xor (n1108,n1109,n1111);
xor (n1109,n1110,n700);
xor (n1110,n644,n677);
xor (n1111,n1112,n1119);
xor (n1112,n1113,n1115);
xor (n1113,n1114,n638);
xor (n1114,n622,n635);
nand (n1115,n1116,n1117,n1118);
nand (n1116,n1078,n1082);
nand (n1117,n1084,n1082);
nand (n1118,n1078,n1084);
nand (n1119,n1120,n1121,n1122);
nand (n1120,n1088,n1092);
nand (n1121,n1094,n1092);
nand (n1122,n1088,n1094);
nand (n1123,n1124,n1125,n1126);
nand (n1124,n1072,n1076);
nand (n1125,n1086,n1076);
nand (n1126,n1072,n1086);
not (n1127,n1128);
nand (n1128,n1103,n1107);
not (n1129,n1130);
nor (n1130,n1131,n1146);
nor (n1131,n1132,n1136);
nand (n1132,n1133,n1134,n1135);
nand (n1133,n1109,n1111);
nand (n1134,n1123,n1111);
nand (n1135,n1109,n1123);
xor (n1136,n1137,n1142);
xor (n1137,n1138,n1140);
xor (n1138,n1139,n590);
xor (n1139,n586,n588);
xor (n1140,n1141,n642);
xor (n1141,n618,n620);
nand (n1142,n1143,n1144,n1145);
nand (n1143,n1113,n1115);
nand (n1144,n1119,n1115);
nand (n1145,n1113,n1119);
nor (n1146,n1147,n1151);
nand (n1147,n1148,n1149,n1150);
nand (n1148,n1138,n1140);
nand (n1149,n1142,n1140);
nand (n1150,n1138,n1142);
xor (n1151,n1152,n616);
xor (n1152,n584,n613);
not (n1153,n1154);
nor (n1154,n1155,n1157);
nor (n1155,n1156,n1146);
nand (n1156,n1132,n1136);
not (n1157,n1158);
nand (n1158,n1147,n1151);
not (n1159,n1160);
nor (n1160,n1161,n1168);
nor (n1161,n1162,n1167);
nor (n1162,n1163,n1165);
nor (n1163,n1164,n705);
nand (n1164,n409,n582);
not (n1165,n1166);
nand (n1166,n706,n710);
not (n1167,n729);
not (n1168,n1169);
nor (n1169,n1170,n1172);
nor (n1170,n1171,n745);
nand (n1171,n731,n735);
not (n1172,n1173);
nand (n1173,n746,n750);
nand (n1174,n1175,n1179);
nor (n1175,n1176,n406);
nand (n1176,n1177,n1130);
nor (n1177,n1178,n1102);
nor (n1178,n757,n1064);
nand (n1179,n1180,n2710);
nor (n1180,n1181,n2678);
nor (n1181,n1182,n2151);
nor (n1182,n1183,n2136);
nor (n1183,n1184,n1857);
nand (n1184,n1185,n1640);
nor (n1185,n1186,n1539);
nor (n1186,n1187,n1449);
nand (n1187,n1188,n1364,n1448);
nand (n1188,n1189,n1266);
xor (n1189,n1190,n1242);
xor (n1190,n1191,n1216);
xor (n1191,n1192,n1204);
xor (n1192,n1193,n1198);
xor (n1193,n1194,n99);
or (n1194,n1195,n1196);
and (n1195,n993,n173);
and (n1196,n1197,n176);
xor (n1198,n1199,n74);
or (n1199,n1200,n1202);
and (n1200,n1201,n97);
and (n1202,n1203,n101);
xor (n1204,n1205,n1209);
xor (n1205,n1206,n886);
or (n1206,n1207,n1208);
and (n1207,n194,n1009);
and (n1208,n196,n1013);
xnor (n1209,n1210,n1011);
nor (n1210,n1211,n1215);
and (n1211,n111,n1212);
and (n1212,n1213,n1011);
not (n1213,n1214);
and (n1215,n64,n1214);
nand (n1216,n1217,n1227,n1241);
nand (n1217,n1218,n1222);
xor (n1218,n1219,n99);
or (n1219,n1220,n1221);
and (n1220,n1197,n173);
and (n1221,n1201,n176);
xor (n1222,n1223,n74);
or (n1223,n1224,n1225);
and (n1224,n1203,n97);
and (n1225,n1226,n101);
nand (n1227,n1228,n1222);
xor (n1228,n1229,n1238);
xor (n1229,n1230,n1234);
xor (n1230,n1231,n886);
or (n1231,n1232,n1233);
and (n1232,n196,n1009);
and (n1233,n212,n1013);
xor (n1234,n1235,n524);
or (n1235,n1236,n1237);
and (n1236,n427,n661);
and (n1237,n514,n665);
xnor (n1238,n1239,n22);
nand (n1239,n1240,n72);
nand (n1241,n1218,n1228);
xor (n1242,n1243,n1252);
xor (n1243,n1244,n1248);
xor (n1244,n1245,n22);
or (n1245,n1246,n1247);
and (n1246,n1226,n72);
and (n1247,n1240,n76);
nand (n1248,n1249,n1250,n1251);
nand (n1249,n1230,n1234);
nand (n1250,n1238,n1234);
nand (n1251,n1230,n1238);
xor (n1252,n1253,n1262);
xor (n1253,n1254,n1258);
xor (n1254,n1255,n524);
or (n1255,n1256,n1257);
and (n1256,n298,n661);
and (n1257,n427,n665);
xor (n1258,n1259,n663);
or (n1259,n1260,n1261);
and (n1260,n212,n884);
and (n1261,n266,n888);
xor (n1262,n1263,n442);
or (n1263,n1264,n1265);
and (n1264,n514,n522);
and (n1265,n560,n526);
nand (n1266,n1267,n1321,n1363);
nand (n1267,n1268,n1270);
xor (n1268,n1269,n1228);
xor (n1269,n1218,n1222);
xor (n1270,n1271,n1310);
xor (n1271,n1272,n1288);
nand (n1272,n1273,n1282,n1287);
nand (n1273,n1274,n1278);
xor (n1274,n1275,n524);
or (n1275,n1276,n1277);
and (n1276,n514,n661);
and (n1277,n560,n665);
xor (n1278,n1279,n663);
or (n1279,n1280,n1281);
and (n1280,n298,n884);
and (n1281,n427,n888);
nand (n1282,n1283,n1278);
xor (n1283,n1284,n442);
or (n1284,n1285,n1286);
and (n1285,n632,n522);
and (n1286,n853,n526);
nand (n1287,n1274,n1283);
nand (n1288,n1289,n1304,n1309);
nand (n1289,n1290,n1299);
xor (n1290,n1291,n1295);
xnor (n1291,n1292,n1011);
nor (n1292,n1293,n1294);
and (n1293,n196,n1212);
and (n1294,n194,n1214);
xor (n1295,n1296,n886);
or (n1296,n1297,n1298);
and (n1297,n212,n1009);
and (n1298,n266,n1013);
and (n1299,n1300,n74);
xnor (n1300,n1301,n1011);
nor (n1301,n1302,n1303);
and (n1302,n212,n1212);
and (n1303,n196,n1214);
nand (n1304,n1305,n1299);
xor (n1305,n1306,n165);
or (n1306,n1307,n1308);
and (n1307,n857,n440);
and (n1308,n859,n444);
nand (n1309,n1290,n1305);
xor (n1310,n1311,n1317);
xor (n1311,n1312,n1316);
xor (n1312,n1313,n165);
or (n1313,n1314,n1315);
and (n1314,n853,n440);
and (n1315,n857,n444);
and (n1316,n1291,n1295);
xor (n1317,n1318,n169);
or (n1318,n1319,n1320);
and (n1319,n859,n163);
and (n1320,n993,n167);
nand (n1321,n1322,n1270);
nand (n1322,n1323,n1347,n1362);
nand (n1323,n1324,n1345);
nand (n1324,n1325,n1339,n1344);
nand (n1325,n1326,n1335);
and (n1326,n1327,n1331);
xnor (n1327,n1328,n1011);
nor (n1328,n1329,n1330);
and (n1329,n266,n1212);
and (n1330,n212,n1214);
xor (n1331,n1332,n886);
or (n1332,n1333,n1334);
and (n1333,n298,n1009);
and (n1334,n427,n1013);
xor (n1335,n1336,n165);
or (n1336,n1337,n1338);
and (n1337,n859,n440);
and (n1338,n993,n444);
nand (n1339,n1340,n1335);
xor (n1340,n1341,n169);
or (n1341,n1342,n1343);
and (n1342,n1197,n163);
and (n1343,n1201,n167);
nand (n1344,n1326,n1340);
xor (n1345,n1346,n1305);
xor (n1346,n1290,n1299);
nand (n1347,n1348,n1345);
xor (n1348,n1349,n1358);
xor (n1349,n1350,n1354);
xor (n1350,n1351,n169);
or (n1351,n1352,n1353);
and (n1352,n993,n163);
and (n1353,n1197,n167);
xor (n1354,n1355,n99);
or (n1355,n1356,n1357);
and (n1356,n1201,n173);
and (n1357,n1203,n176);
xor (n1358,n1359,n74);
or (n1359,n1360,n1361);
and (n1360,n1226,n97);
and (n1361,n1240,n101);
nand (n1362,n1324,n1348);
nand (n1363,n1268,n1322);
nand (n1364,n1365,n1266);
xor (n1365,n1366,n1405);
xor (n1366,n1367,n1371);
nand (n1367,n1368,n1369,n1370);
nand (n1368,n1272,n1288);
nand (n1369,n1310,n1288);
nand (n1370,n1272,n1310);
xor (n1371,n1372,n1394);
xor (n1372,n1373,n1390);
nand (n1373,n1374,n1384,n1389);
nand (n1374,n1375,n1379);
xor (n1375,n1376,n663);
or (n1376,n1377,n1378);
and (n1377,n266,n884);
and (n1378,n298,n888);
xor (n1379,n1380,n22);
xnor (n1380,n1381,n1011);
nor (n1381,n1382,n1383);
and (n1382,n194,n1212);
and (n1383,n111,n1214);
nand (n1384,n1385,n1379);
xor (n1385,n1386,n442);
or (n1386,n1387,n1388);
and (n1387,n560,n522);
and (n1388,n632,n526);
nand (n1389,n1375,n1385);
nand (n1390,n1391,n1392,n1393);
nand (n1391,n1312,n1316);
nand (n1392,n1317,n1316);
nand (n1393,n1312,n1317);
xor (n1394,n1395,n1401);
xor (n1395,n1396,n1397);
and (n1396,n1380,n22);
xor (n1397,n1398,n165);
or (n1398,n1399,n1400);
and (n1399,n632,n440);
and (n1400,n853,n444);
xor (n1401,n1402,n169);
or (n1402,n1403,n1404);
and (n1403,n857,n163);
and (n1404,n859,n167);
nand (n1405,n1406,n1413,n1447);
nand (n1406,n1407,n1411);
nand (n1407,n1408,n1409,n1410);
nand (n1408,n1350,n1354);
nand (n1409,n1358,n1354);
nand (n1410,n1350,n1358);
xor (n1411,n1412,n1385);
xor (n1412,n1375,n1379);
nand (n1413,n1414,n1411);
nand (n1414,n1415,n1432,n1446);
nand (n1415,n1416,n1430);
nand (n1416,n1417,n1426,n1429);
nand (n1417,n1418,n1422);
xor (n1418,n1419,n886);
or (n1419,n1420,n1421);
and (n1420,n266,n1009);
and (n1421,n298,n1013);
xor (n1422,n1423,n524);
or (n1423,n1424,n1425);
and (n1424,n560,n661);
and (n1425,n632,n665);
nand (n1426,n1427,n1422);
xnor (n1427,n1428,n74);
nand (n1428,n1240,n97);
nand (n1429,n1418,n1427);
xor (n1430,n1431,n1283);
xor (n1431,n1274,n1278);
nand (n1432,n1433,n1430);
nand (n1433,n1434,n1440,n1445);
nand (n1434,n1435,n1439);
xor (n1435,n1436,n663);
or (n1436,n1437,n1438);
and (n1437,n427,n884);
and (n1438,n514,n888);
xor (n1439,n1300,n74);
nand (n1440,n1441,n1439);
xor (n1441,n1442,n442);
or (n1442,n1443,n1444);
and (n1443,n853,n522);
and (n1444,n857,n526);
nand (n1445,n1435,n1441);
nand (n1446,n1416,n1433);
nand (n1447,n1407,n1414);
nand (n1448,n1189,n1365);
xor (n1449,n1450,n1535);
xor (n1450,n1451,n1472);
xor (n1451,n1452,n1468);
xor (n1452,n1453,n1464);
xor (n1453,n1454,n1460);
xor (n1454,n1455,n1459);
xor (n1455,n1456,n74);
or (n1456,n1457,n1458);
and (n1457,n1197,n97);
and (n1458,n1201,n101);
and (n1459,n1205,n1209);
xor (n1460,n1461,n22);
or (n1461,n1462,n1463);
and (n1462,n1203,n72);
and (n1463,n1226,n76);
nand (n1464,n1465,n1466,n1467);
nand (n1465,n1244,n1248);
nand (n1466,n1252,n1248);
nand (n1467,n1244,n1252);
nand (n1468,n1469,n1470,n1471);
nand (n1469,n1373,n1390);
nand (n1470,n1394,n1390);
nand (n1471,n1373,n1394);
xor (n1472,n1473,n1531);
xor (n1473,n1474,n1498);
xor (n1474,n1475,n1494);
xor (n1475,n1476,n1480);
nand (n1476,n1477,n1478,n1479);
nand (n1477,n1396,n1397);
nand (n1478,n1401,n1397);
nand (n1479,n1396,n1401);
xor (n1480,n1481,n1490);
xor (n1481,n1482,n1486);
xnor (n1482,n1483,n1011);
nor (n1483,n1484,n1485);
and (n1484,n64,n1212);
and (n1485,n62,n1214);
xor (n1486,n1487,n524);
or (n1487,n1488,n1489);
and (n1488,n266,n661);
and (n1489,n298,n665);
xor (n1490,n1491,n663);
or (n1491,n1492,n1493);
and (n1492,n196,n884);
and (n1493,n212,n888);
nand (n1494,n1495,n1496,n1497);
nand (n1495,n1254,n1258);
nand (n1496,n1262,n1258);
nand (n1497,n1254,n1262);
xor (n1498,n1499,n1517);
xor (n1499,n1500,n1504);
nand (n1500,n1501,n1502,n1503);
nand (n1501,n1193,n1198);
nand (n1502,n1204,n1198);
nand (n1503,n1193,n1204);
xor (n1504,n1505,n1515);
xor (n1505,n1506,n1510);
xor (n1506,n1507,n442);
or (n1507,n1508,n1509);
and (n1508,n427,n522);
and (n1509,n514,n526);
xor (n1510,n9,n1511);
xor (n1511,n1512,n886);
or (n1512,n1513,n1514);
and (n1513,n111,n1009);
and (n1514,n194,n1013);
xnor (n1515,n1516,n9);
nand (n1516,n1240,n20);
xor (n1517,n1518,n1527);
xor (n1518,n1519,n1523);
xor (n1519,n1520,n165);
or (n1520,n1521,n1522);
and (n1521,n560,n440);
and (n1522,n632,n444);
xor (n1523,n1524,n169);
or (n1524,n1525,n1526);
and (n1525,n853,n163);
and (n1526,n857,n167);
xor (n1527,n1528,n99);
or (n1528,n1529,n1530);
and (n1529,n859,n173);
and (n1530,n993,n176);
nand (n1531,n1532,n1533,n1534);
nand (n1532,n1191,n1216);
nand (n1533,n1242,n1216);
nand (n1534,n1191,n1242);
nand (n1535,n1536,n1537,n1538);
nand (n1536,n1367,n1371);
nand (n1537,n1405,n1371);
nand (n1538,n1367,n1405);
nor (n1539,n1540,n1544);
nand (n1540,n1541,n1542,n1543);
nand (n1541,n1451,n1472);
nand (n1542,n1535,n1472);
nand (n1543,n1451,n1535);
xor (n1544,n1545,n1554);
xor (n1545,n1546,n1550);
nand (n1546,n1547,n1548,n1549);
nand (n1547,n1453,n1464);
nand (n1548,n1468,n1464);
nand (n1549,n1453,n1468);
nand (n1550,n1551,n1552,n1553);
nand (n1551,n1474,n1498);
nand (n1552,n1531,n1498);
nand (n1553,n1474,n1531);
xor (n1554,n1555,n1616);
xor (n1555,n1556,n1587);
xor (n1556,n1557,n1576);
xor (n1557,n1558,n1572);
xor (n1558,n1559,n1568);
xor (n1559,n1560,n1564);
xor (n1560,n1561,n524);
or (n1561,n1562,n1563);
and (n1562,n212,n661);
and (n1563,n266,n665);
xor (n1564,n1565,n663);
or (n1565,n1566,n1567);
and (n1566,n194,n884);
and (n1567,n196,n888);
xor (n1568,n1569,n442);
or (n1569,n1570,n1571);
and (n1570,n298,n522);
and (n1571,n427,n526);
nand (n1572,n1573,n1574,n1575);
nand (n1573,n1506,n1510);
nand (n1574,n1515,n1510);
nand (n1575,n1506,n1515);
xor (n1576,n1577,n1583);
xor (n1577,n1578,n1582);
xor (n1578,n1579,n165);
or (n1579,n1580,n1581);
and (n1580,n514,n440);
and (n1581,n560,n444);
and (n1582,n9,n1511);
xor (n1583,n1584,n169);
or (n1584,n1585,n1586);
and (n1585,n632,n163);
and (n1586,n853,n167);
xor (n1587,n1588,n1612);
xor (n1588,n1589,n1593);
nand (n1589,n1590,n1591,n1592);
nand (n1590,n1519,n1523);
nand (n1591,n1527,n1523);
nand (n1592,n1519,n1527);
xor (n1593,n1594,n1603);
xor (n1594,n1595,n1599);
xor (n1595,n1596,n99);
or (n1596,n1597,n1598);
and (n1597,n857,n173);
and (n1598,n859,n176);
xor (n1599,n1600,n74);
or (n1600,n1601,n1602);
and (n1601,n993,n97);
and (n1602,n1197,n101);
xor (n1603,n1604,n1608);
xnor (n1604,n1605,n1011);
nor (n1605,n1606,n1607);
and (n1606,n62,n1212);
and (n1607,n43,n1214);
xor (n1608,n1609,n886);
or (n1609,n1610,n1611);
and (n1610,n64,n1009);
and (n1611,n111,n1013);
nand (n1612,n1613,n1614,n1615);
nand (n1613,n1455,n1459);
nand (n1614,n1460,n1459);
nand (n1615,n1455,n1460);
xor (n1616,n1617,n1636);
xor (n1617,n1618,n1632);
xor (n1618,n1619,n1628);
xor (n1619,n1620,n1624);
xor (n1620,n1621,n22);
or (n1621,n1622,n1623);
and (n1622,n1201,n72);
and (n1623,n1203,n76);
xor (n1624,n1625,n9);
or (n1625,n1626,n1627);
and (n1626,n1226,n20);
and (n1627,n1240,n24);
nand (n1628,n1629,n1630,n1631);
nand (n1629,n1482,n1486);
nand (n1630,n1490,n1486);
nand (n1631,n1482,n1490);
nand (n1632,n1633,n1634,n1635);
nand (n1633,n1476,n1480);
nand (n1634,n1494,n1480);
nand (n1635,n1476,n1494);
nand (n1636,n1637,n1638,n1639);
nand (n1637,n1500,n1504);
nand (n1638,n1517,n1504);
nand (n1639,n1500,n1517);
nor (n1640,n1641,n1746);
nor (n1641,n1642,n1646);
nand (n1642,n1643,n1644,n1645);
nand (n1643,n1546,n1550);
nand (n1644,n1554,n1550);
nand (n1645,n1546,n1554);
xor (n1646,n1647,n1742);
xor (n1647,n1648,n1682);
xor (n1648,n1649,n1678);
xor (n1649,n1650,n1654);
nand (n1650,n1651,n1652,n1653);
nand (n1651,n1558,n1572);
nand (n1652,n1576,n1572);
nand (n1653,n1558,n1576);
xor (n1654,n1655,n1664);
xor (n1655,n1656,n1660);
xor (n1656,n1657,n9);
or (n1657,n1658,n1659);
and (n1658,n1203,n20);
and (n1659,n1226,n24);
nand (n1660,n1661,n1662,n1663);
nand (n1661,n1578,n1582);
nand (n1662,n1583,n1582);
nand (n1663,n1578,n1583);
xor (n1664,n1665,n1674);
xor (n1665,n1666,n1670);
xor (n1666,n1667,n524);
or (n1667,n1668,n1669);
and (n1668,n196,n661);
and (n1669,n212,n665);
xnor (n1670,n1671,n1011);
nor (n1671,n1672,n1673);
and (n1672,n43,n1212);
and (n1673,n29,n1214);
xor (n1674,n1675,n663);
or (n1675,n1676,n1677);
and (n1676,n111,n884);
and (n1677,n194,n888);
nand (n1678,n1679,n1680,n1681);
nand (n1679,n1589,n1593);
nand (n1680,n1612,n1593);
nand (n1681,n1589,n1612);
xor (n1682,n1683,n1738);
xor (n1683,n1684,n1706);
xor (n1684,n1685,n1694);
xor (n1685,n1686,n1690);
nand (n1686,n1687,n1688,n1689);
nand (n1687,n1560,n1564);
nand (n1688,n1568,n1564);
nand (n1689,n1560,n1568);
nand (n1690,n1691,n1692,n1693);
nand (n1691,n1595,n1599);
nand (n1692,n1603,n1599);
nand (n1693,n1595,n1603);
xor (n1694,n1695,n1702);
xor (n1695,n1696,n1700);
xor (n1696,n1697,n442);
or (n1697,n1698,n1699);
and (n1698,n266,n522);
and (n1699,n298,n526);
xnor (n1700,n1701,n13);
nand (n1701,n1240,n7);
xor (n1702,n1703,n165);
or (n1703,n1704,n1705);
and (n1704,n427,n440);
and (n1705,n514,n444);
xor (n1706,n1707,n1726);
xor (n1707,n1708,n1712);
nand (n1708,n1709,n1710,n1711);
nand (n1709,n1620,n1624);
nand (n1710,n1628,n1624);
nand (n1711,n1620,n1628);
xor (n1712,n1713,n1722);
xor (n1713,n1714,n1718);
xor (n1714,n1715,n169);
or (n1715,n1716,n1717);
and (n1716,n560,n163);
and (n1717,n632,n167);
xor (n1718,n1719,n99);
or (n1719,n1720,n1721);
and (n1720,n853,n173);
and (n1721,n857,n176);
xor (n1722,n1723,n74);
or (n1723,n1724,n1725);
and (n1724,n859,n97);
and (n1725,n993,n101);
xor (n1726,n1727,n1734);
xor (n1727,n1728,n1733);
xor (n1728,n13,n1729);
xor (n1729,n1730,n886);
or (n1730,n1731,n1732);
and (n1731,n62,n1009);
and (n1732,n64,n1013);
and (n1733,n1604,n1608);
xor (n1734,n1735,n22);
or (n1735,n1736,n1737);
and (n1736,n1197,n72);
and (n1737,n1201,n76);
nand (n1738,n1739,n1740,n1741);
nand (n1739,n1618,n1632);
nand (n1740,n1636,n1632);
nand (n1741,n1618,n1636);
nand (n1742,n1743,n1744,n1745);
nand (n1743,n1556,n1587);
nand (n1744,n1616,n1587);
nand (n1745,n1556,n1616);
nor (n1746,n1747,n1751);
nand (n1747,n1748,n1749,n1750);
nand (n1748,n1648,n1682);
nand (n1749,n1742,n1682);
nand (n1750,n1648,n1742);
xor (n1751,n1752,n1761);
xor (n1752,n1753,n1757);
nand (n1753,n1754,n1755,n1756);
nand (n1754,n1650,n1654);
nand (n1755,n1678,n1654);
nand (n1756,n1650,n1678);
nand (n1757,n1758,n1759,n1760);
nand (n1758,n1684,n1706);
nand (n1759,n1738,n1706);
nand (n1760,n1684,n1738);
xor (n1761,n1762,n1823);
xor (n1762,n1763,n1787);
xor (n1763,n1764,n1783);
xor (n1764,n1765,n1769);
nand (n1765,n1766,n1767,n1768);
nand (n1766,n1714,n1718);
nand (n1767,n1722,n1718);
nand (n1768,n1714,n1722);
xor (n1769,n1770,n1779);
xor (n1770,n1771,n1775);
xor (n1771,n1772,n165);
or (n1772,n1773,n1774);
and (n1773,n298,n440);
and (n1774,n427,n444);
xor (n1775,n1776,n169);
or (n1776,n1777,n1778);
and (n1777,n514,n163);
and (n1778,n560,n167);
xor (n1779,n1780,n99);
or (n1780,n1781,n1782);
and (n1781,n632,n173);
and (n1782,n853,n176);
nand (n1783,n1784,n1785,n1786);
nand (n1784,n1728,n1733);
nand (n1785,n1734,n1733);
nand (n1786,n1728,n1734);
xor (n1787,n1788,n1809);
xor (n1788,n1789,n1805);
xor (n1789,n1790,n1804);
xor (n1790,n1791,n1795);
xor (n1791,n1792,n74);
or (n1792,n1793,n1794);
and (n1793,n857,n97);
and (n1794,n859,n101);
xor (n1795,n1796,n1800);
xnor (n1796,n1797,n1011);
nor (n1797,n1798,n1799);
and (n1798,n29,n1212);
and (n1799,n6,n1214);
xor (n1800,n1801,n886);
or (n1801,n1802,n1803);
and (n1802,n43,n1009);
and (n1803,n62,n1013);
and (n1804,n13,n1729);
nand (n1805,n1806,n1807,n1808);
nand (n1806,n1656,n1660);
nand (n1807,n1664,n1660);
nand (n1808,n1656,n1664);
xor (n1809,n1810,n1819);
xor (n1810,n1811,n1815);
xor (n1811,n1812,n22);
or (n1812,n1813,n1814);
and (n1813,n993,n72);
and (n1814,n1197,n76);
xor (n1815,n1816,n13);
or (n1816,n1817,n1818);
and (n1817,n1226,n7);
and (n1818,n1240,n11);
xor (n1819,n1820,n9);
or (n1820,n1821,n1822);
and (n1821,n1201,n20);
and (n1822,n1203,n24);
xor (n1823,n1824,n1853);
xor (n1824,n1825,n1849);
xor (n1825,n1826,n1845);
xor (n1826,n1827,n1831);
nand (n1827,n1828,n1829,n1830);
nand (n1828,n1666,n1670);
nand (n1829,n1674,n1670);
nand (n1830,n1666,n1674);
xor (n1831,n1832,n1841);
xor (n1832,n1833,n1837);
xor (n1833,n1834,n524);
or (n1834,n1835,n1836);
and (n1835,n194,n661);
and (n1836,n196,n665);
xor (n1837,n1838,n663);
or (n1838,n1839,n1840);
and (n1839,n64,n884);
and (n1840,n111,n888);
xor (n1841,n1842,n442);
or (n1842,n1843,n1844);
and (n1843,n212,n522);
and (n1844,n266,n526);
nand (n1845,n1846,n1847,n1848);
nand (n1846,n1696,n1700);
nand (n1847,n1702,n1700);
nand (n1848,n1696,n1702);
nand (n1849,n1850,n1851,n1852);
nand (n1850,n1686,n1690);
nand (n1851,n1694,n1690);
nand (n1852,n1686,n1694);
nand (n1853,n1854,n1855,n1856);
nand (n1854,n1708,n1712);
nand (n1855,n1726,n1712);
nand (n1856,n1708,n1726);
nor (n1857,n1858,n2130);
nor (n1858,n1859,n2106);
nor (n1859,n1860,n2104);
nor (n1860,n1861,n2079);
nand (n1861,n1862,n2041);
nand (n1862,n1863,n1988,n2040);
nand (n1863,n1864,n1915);
xor (n1864,n1865,n1902);
xor (n1865,n1866,n1887);
nand (n1866,n1867,n1881,n1886);
nand (n1867,n1868,n1877);
and (n1868,n1869,n1873);
xnor (n1869,n1870,n1011);
nor (n1870,n1871,n1872);
and (n1871,n427,n1212);
and (n1872,n298,n1214);
xor (n1873,n1874,n886);
or (n1874,n1875,n1876);
and (n1875,n514,n1009);
and (n1876,n560,n1013);
xor (n1877,n1878,n165);
or (n1878,n1879,n1880);
and (n1879,n1197,n440);
and (n1880,n1201,n444);
nand (n1881,n1882,n1877);
xor (n1882,n1883,n169);
or (n1883,n1884,n1885);
and (n1884,n1203,n163);
and (n1885,n1226,n167);
nand (n1886,n1868,n1882);
xor (n1887,n1888,n1897);
xor (n1888,n1889,n1893);
xor (n1889,n1890,n524);
or (n1890,n1891,n1892);
and (n1891,n632,n661);
and (n1892,n853,n665);
xor (n1893,n1894,n663);
or (n1894,n1895,n1896);
and (n1895,n514,n884);
and (n1896,n560,n888);
and (n1897,n1898,n99);
xnor (n1898,n1899,n1011);
nor (n1899,n1900,n1901);
and (n1900,n298,n1212);
and (n1901,n266,n1214);
nand (n1902,n1903,n1909,n1914);
nand (n1903,n1904,n1908);
xor (n1904,n1905,n663);
or (n1905,n1906,n1907);
and (n1906,n560,n884);
and (n1907,n632,n888);
xor (n1908,n1898,n99);
nand (n1909,n1910,n1908);
xor (n1910,n1911,n442);
or (n1911,n1912,n1913);
and (n1912,n859,n522);
and (n1913,n993,n526);
nand (n1914,n1904,n1910);
xor (n1915,n1916,n1952);
xor (n1916,n1917,n1928);
xor (n1917,n1918,n1924);
xor (n1918,n1919,n1923);
xor (n1919,n1920,n442);
or (n1920,n1921,n1922);
and (n1921,n857,n522);
and (n1922,n859,n526);
xor (n1923,n1327,n1331);
xor (n1924,n1925,n165);
or (n1925,n1926,n1927);
and (n1926,n993,n440);
and (n1927,n1197,n444);
xor (n1928,n1929,n1938);
xor (n1929,n1930,n1934);
xor (n1930,n1931,n169);
or (n1931,n1932,n1933);
and (n1932,n1201,n163);
and (n1933,n1203,n167);
xor (n1934,n1935,n99);
or (n1935,n1936,n1937);
and (n1936,n1226,n173);
and (n1937,n1240,n176);
nand (n1938,n1939,n1946,n1951);
nand (n1939,n1940,n1944);
xor (n1940,n1941,n886);
or (n1941,n1942,n1943);
and (n1942,n427,n1009);
and (n1943,n514,n1013);
xnor (n1944,n1945,n99);
nand (n1945,n1240,n173);
nand (n1946,n1947,n1944);
xor (n1947,n1948,n524);
or (n1948,n1949,n1950);
and (n1949,n853,n661);
and (n1950,n857,n665);
nand (n1951,n1940,n1947);
nand (n1952,n1953,n1973,n1987);
nand (n1953,n1954,n1956);
xor (n1954,n1955,n1947);
xor (n1955,n1940,n1944);
nand (n1956,n1957,n1966,n1972);
nand (n1957,n1958,n1962);
xor (n1958,n1959,n524);
or (n1959,n1960,n1961);
and (n1960,n857,n661);
and (n1961,n859,n665);
xor (n1962,n1963,n663);
or (n1963,n1964,n1965);
and (n1964,n632,n884);
and (n1965,n853,n888);
nand (n1966,n1967,n1962);
and (n1967,n1968,n169);
xnor (n1968,n1969,n1011);
nor (n1969,n1970,n1971);
and (n1970,n514,n1212);
and (n1971,n427,n1214);
nand (n1972,n1958,n1967);
nand (n1973,n1974,n1956);
nand (n1974,n1975,n1981,n1986);
nand (n1975,n1976,n1980);
xor (n1976,n1977,n442);
or (n1977,n1978,n1979);
and (n1978,n993,n522);
and (n1979,n1197,n526);
xor (n1980,n1869,n1873);
nand (n1981,n1982,n1980);
xor (n1982,n1983,n165);
or (n1983,n1984,n1985);
and (n1984,n1201,n440);
and (n1985,n1203,n444);
nand (n1986,n1976,n1982);
nand (n1987,n1954,n1974);
nand (n1988,n1989,n1915);
nand (n1989,n1990,n1995,n2039);
nand (n1990,n1991,n1993);
xor (n1991,n1992,n1882);
xor (n1992,n1868,n1877);
xor (n1993,n1994,n1910);
xor (n1994,n1904,n1908);
nand (n1995,n1996,n1993);
nand (n1996,n1997,n2016,n2038);
nand (n1997,n1998,n2002);
xor (n1998,n1999,n169);
or (n1999,n2000,n2001);
and (n2000,n1226,n163);
and (n2001,n1240,n167);
nand (n2002,n2003,n2010,n2015);
nand (n2003,n2004,n2008);
xor (n2004,n2005,n886);
or (n2005,n2006,n2007);
and (n2006,n560,n1009);
and (n2007,n632,n1013);
xnor (n2008,n2009,n169);
nand (n2009,n1240,n163);
nand (n2010,n2011,n2008);
xor (n2011,n2012,n524);
or (n2012,n2013,n2014);
and (n2013,n859,n661);
and (n2014,n993,n665);
nand (n2015,n2004,n2011);
nand (n2016,n2017,n2002);
nand (n2017,n2018,n2032,n2037);
nand (n2018,n2019,n2023);
xor (n2019,n2020,n663);
or (n2020,n2021,n2022);
and (n2021,n853,n884);
and (n2022,n857,n888);
and (n2023,n2024,n2028);
xnor (n2024,n2025,n1011);
nor (n2025,n2026,n2027);
and (n2026,n560,n1212);
and (n2027,n514,n1214);
xor (n2028,n2029,n886);
or (n2029,n2030,n2031);
and (n2030,n632,n1009);
and (n2031,n853,n1013);
nand (n2032,n2033,n2023);
xor (n2033,n2034,n442);
or (n2034,n2035,n2036);
and (n2035,n1197,n522);
and (n2036,n1201,n526);
nand (n2037,n2019,n2033);
nand (n2038,n1998,n2017);
nand (n2039,n1991,n1996);
nand (n2040,n1864,n1989);
xor (n2041,n2042,n2057);
xor (n2042,n2043,n2053);
xor (n2043,n2044,n2051);
xor (n2044,n2045,n2049);
nand (n2045,n2046,n2047,n2048);
nand (n2046,n1889,n1893);
nand (n2047,n1897,n1893);
nand (n2048,n1889,n1897);
xor (n2049,n2050,n1340);
xor (n2050,n1326,n1335);
xor (n2051,n2052,n1441);
xor (n2052,n1435,n1439);
nand (n2053,n2054,n2055,n2056);
nand (n2054,n1917,n1928);
nand (n2055,n1952,n1928);
nand (n2056,n1917,n1952);
xor (n2057,n2058,n2067);
xor (n2058,n2059,n2063);
nand (n2059,n2060,n2061,n2062);
nand (n2060,n1930,n1934);
nand (n2061,n1938,n1934);
nand (n2062,n1930,n1938);
nand (n2063,n2064,n2065,n2066);
nand (n2064,n1866,n1887);
nand (n2065,n1902,n1887);
nand (n2066,n1866,n1902);
xor (n2067,n2068,n2077);
xor (n2068,n2069,n2073);
xor (n2069,n2070,n99);
or (n2070,n2071,n2072);
and (n2071,n1203,n173);
and (n2072,n1226,n176);
nand (n2073,n2074,n2075,n2076);
nand (n2074,n1919,n1923);
nand (n2075,n1924,n1923);
nand (n2076,n1919,n1924);
xor (n2077,n2078,n1427);
xor (n2078,n1418,n1422);
nor (n2079,n2080,n2084);
nand (n2080,n2081,n2082,n2083);
nand (n2081,n2043,n2053);
nand (n2082,n2057,n2053);
nand (n2083,n2043,n2057);
xor (n2084,n2085,n2092);
xor (n2085,n2086,n2088);
xor (n2086,n2087,n1348);
xor (n2087,n1324,n1345);
nand (n2088,n2089,n2090,n2091);
nand (n2089,n2059,n2063);
nand (n2090,n2067,n2063);
nand (n2091,n2059,n2067);
xor (n2092,n2093,n2102);
xor (n2093,n2094,n2098);
nand (n2094,n2095,n2096,n2097);
nand (n2095,n2069,n2073);
nand (n2096,n2077,n2073);
nand (n2097,n2069,n2077);
nand (n2098,n2099,n2100,n2101);
nand (n2099,n2045,n2049);
nand (n2100,n2051,n2049);
nand (n2101,n2045,n2051);
xor (n2102,n2103,n1433);
xor (n2103,n1416,n1430);
not (n2104,n2105);
nand (n2105,n2080,n2084);
not (n2106,n2107);
nor (n2107,n2108,n2123);
nor (n2108,n2109,n2113);
nand (n2109,n2110,n2111,n2112);
nand (n2110,n2086,n2088);
nand (n2111,n2092,n2088);
nand (n2112,n2086,n2092);
xor (n2113,n2114,n2121);
xor (n2114,n2115,n2117);
xor (n2115,n2116,n1414);
xor (n2116,n1407,n1411);
nand (n2117,n2118,n2119,n2120);
nand (n2118,n2094,n2098);
nand (n2119,n2102,n2098);
nand (n2120,n2094,n2102);
xor (n2121,n2122,n1322);
xor (n2122,n1268,n1270);
nor (n2123,n2124,n2128);
nand (n2124,n2125,n2126,n2127);
nand (n2125,n2115,n2117);
nand (n2126,n2121,n2117);
nand (n2127,n2115,n2121);
xor (n2128,n2129,n1365);
xor (n2129,n1189,n1266);
not (n2130,n2131);
nor (n2131,n2132,n2134);
nor (n2132,n2133,n2123);
nand (n2133,n2109,n2113);
not (n2134,n2135);
nand (n2135,n2124,n2128);
not (n2136,n2137);
nor (n2137,n2138,n2145);
nor (n2138,n2139,n2144);
nor (n2139,n2140,n2142);
nor (n2140,n2141,n1539);
nand (n2141,n1187,n1449);
not (n2142,n2143);
nand (n2143,n1540,n1544);
not (n2144,n1640);
not (n2145,n2146);
nor (n2146,n2147,n2149);
nor (n2147,n2148,n1746);
nand (n2148,n1642,n1646);
not (n2149,n2150);
nand (n2150,n1747,n1751);
not (n2151,n2152);
nor (n2152,n2153,n2568);
nand (n2153,n2154,n2381);
nor (n2154,n2155,n2267);
nor (n2155,n2156,n2160);
nand (n2156,n2157,n2158,n2159);
nand (n2157,n1753,n1757);
nand (n2158,n1761,n1757);
nand (n2159,n1753,n1761);
xor (n2160,n2161,n2263);
xor (n2161,n2162,n2195);
xor (n2162,n2163,n2191);
xor (n2163,n2164,n2187);
xor (n2164,n2165,n2183);
xor (n2165,n2166,n2179);
xor (n2166,n2167,n2176);
xor (n2167,n2168,n2172);
xor (n2168,n2169,n886);
or (n2169,n2170,n2171);
and (n2170,n29,n1009);
and (n2171,n43,n1013);
xor (n2172,n2173,n663);
or (n2173,n2174,n2175);
and (n2174,n62,n884);
and (n2175,n64,n888);
xnor (n2176,n2177,n1011);
nor (n2177,n2178,n1799);
and (n2178,n6,n1212);
nand (n2179,n2180,n2181,n2182);
nand (n2180,n1771,n1775);
nand (n2181,n1779,n1775);
nand (n2182,n1771,n1779);
nand (n2183,n2184,n2185,n2186);
nand (n2184,n1791,n1795);
nand (n2185,n1804,n1795);
nand (n2186,n1791,n1804);
nand (n2187,n2188,n2189,n2190);
nand (n2188,n1765,n1769);
nand (n2189,n1783,n1769);
nand (n2190,n1765,n1783);
nand (n2191,n2192,n2193,n2194);
nand (n2192,n1789,n1805);
nand (n2193,n1809,n1805);
nand (n2194,n1789,n1809);
xor (n2195,n2196,n2259);
xor (n2196,n2197,n2235);
xor (n2197,n2198,n2220);
xor (n2198,n2199,n2213);
xor (n2199,n2200,n2209);
xor (n2200,n2201,n2205);
xor (n2201,n2202,n442);
or (n2202,n2203,n2204);
and (n2203,n196,n522);
and (n2204,n212,n526);
xor (n2205,n2206,n165);
or (n2206,n2207,n2208);
and (n2207,n266,n440);
and (n2208,n298,n444);
xor (n2209,n2210,n169);
or (n2210,n2211,n2212);
and (n2211,n427,n163);
and (n2212,n514,n167);
xor (n2213,n2214,n2216);
xor (n2214,n13,n2215);
and (n2215,n1796,n1800);
xor (n2216,n2217,n22);
or (n2217,n2218,n2219);
and (n2218,n859,n72);
and (n2219,n993,n76);
xor (n2220,n2221,n2230);
xor (n2221,n2222,n2226);
xor (n2222,n2223,n99);
or (n2223,n2224,n2225);
and (n2224,n560,n173);
and (n2225,n632,n176);
xor (n2226,n2227,n74);
or (n2227,n2228,n2229);
and (n2228,n853,n97);
and (n2229,n857,n101);
xor (n2230,n13,n2231);
xor (n2231,n2232,n524);
or (n2232,n2233,n2234);
and (n2233,n111,n661);
and (n2234,n194,n665);
xor (n2235,n2236,n2245);
xor (n2236,n2237,n2241);
nand (n2237,n2238,n2239,n2240);
nand (n2238,n1811,n1815);
nand (n2239,n1819,n1815);
nand (n2240,n1811,n1819);
nand (n2241,n2242,n2243,n2244);
nand (n2242,n1827,n1831);
nand (n2243,n1845,n1831);
nand (n2244,n1827,n1845);
xor (n2245,n2246,n2255);
xor (n2246,n2247,n2251);
xor (n2247,n2248,n9);
or (n2248,n2249,n2250);
and (n2249,n1197,n20);
and (n2250,n1201,n24);
xor (n2251,n2252,n13);
or (n2252,n2253,n2254);
and (n2253,n1203,n7);
and (n2254,n1226,n11);
nand (n2255,n2256,n2257,n2258);
nand (n2256,n1833,n1837);
nand (n2257,n1841,n1837);
nand (n2258,n1833,n1841);
nand (n2259,n2260,n2261,n2262);
nand (n2260,n1825,n1849);
nand (n2261,n1853,n1849);
nand (n2262,n1825,n1853);
nand (n2263,n2264,n2265,n2266);
nand (n2264,n1763,n1787);
nand (n2265,n1823,n1787);
nand (n2266,n1763,n1823);
nor (n2267,n2268,n2272);
nand (n2268,n2269,n2270,n2271);
nand (n2269,n2162,n2195);
nand (n2270,n2263,n2195);
nand (n2271,n2162,n2263);
xor (n2272,n2273,n2282);
xor (n2273,n2274,n2278);
nand (n2274,n2275,n2276,n2277);
nand (n2275,n2164,n2187);
nand (n2276,n2191,n2187);
nand (n2277,n2164,n2191);
nand (n2278,n2279,n2280,n2281);
nand (n2279,n2197,n2235);
nand (n2280,n2259,n2235);
nand (n2281,n2197,n2259);
xor (n2282,n2283,n2340);
xor (n2283,n2284,n2315);
xor (n2284,n2285,n2301);
xor (n2285,n2286,n2290);
nand (n2286,n2287,n2288,n2289);
nand (n2287,n13,n2215);
nand (n2288,n2216,n2215);
nand (n2289,n13,n2216);
xor (n2290,n2291,n2297);
xor (n2291,n2292,n2296);
xor (n2292,n2293,n74);
or (n2293,n2294,n2295);
and (n2294,n632,n97);
and (n2295,n853,n101);
and (n2296,n13,n2231);
xor (n2297,n2298,n22);
or (n2298,n2299,n2300);
and (n2299,n857,n72);
and (n2300,n859,n76);
xor (n2301,n2302,n2311);
xor (n2302,n2303,n2307);
xor (n2303,n2304,n9);
or (n2304,n2305,n2306);
and (n2305,n993,n20);
and (n2306,n1197,n24);
xor (n2307,n2308,n13);
or (n2308,n2309,n2310);
and (n2309,n1201,n7);
and (n2310,n1203,n11);
nand (n2311,n2312,n2313,n2314);
nand (n2312,n2168,n2172);
nand (n2313,n2176,n2172);
nand (n2314,n2168,n2176);
xor (n2315,n2316,n2325);
xor (n2316,n2317,n2321);
nand (n2317,n2318,n2319,n2320);
nand (n2318,n2247,n2251);
nand (n2319,n2255,n2251);
nand (n2320,n2247,n2255);
nand (n2321,n2322,n2323,n2324);
nand (n2322,n2166,n2179);
nand (n2323,n2183,n2179);
nand (n2324,n2166,n2183);
xor (n2325,n2326,n13);
xor (n2326,n2327,n2331);
nand (n2327,n2328,n2329,n2330);
nand (n2328,n2201,n2205);
nand (n2329,n2209,n2205);
nand (n2330,n2201,n2209);
xor (n2331,n2332,n2337);
not (n2332,n2333);
xor (n2333,n2334,n524);
or (n2334,n2335,n2336);
and (n2335,n64,n661);
and (n2336,n111,n665);
xor (n2337,n2338,n886);
or (n2338,n1008,n2339);
and (n2339,n29,n1013);
xor (n2340,n2341,n2377);
xor (n2341,n2342,n2346);
nand (n2342,n2343,n2344,n2345);
nand (n2343,n2199,n2213);
nand (n2344,n2220,n2213);
nand (n2345,n2199,n2220);
xor (n2346,n2347,n2366);
xor (n2347,n2348,n2352);
nand (n2348,n2349,n2350,n2351);
nand (n2349,n2222,n2226);
nand (n2350,n2230,n2226);
nand (n2351,n2222,n2230);
xor (n2352,n2353,n2362);
xor (n2353,n2354,n2358);
xor (n2354,n2355,n165);
or (n2355,n2356,n2357);
and (n2356,n212,n440);
and (n2357,n266,n444);
xor (n2358,n2359,n169);
or (n2359,n2360,n2361);
and (n2360,n298,n163);
and (n2361,n427,n167);
xor (n2362,n2363,n99);
or (n2363,n2364,n2365);
and (n2364,n514,n173);
and (n2365,n560,n176);
xor (n2366,n2367,n2373);
xor (n2367,n2368,n2372);
xor (n2368,n2369,n663);
or (n2369,n2370,n2371);
and (n2370,n43,n884);
and (n2371,n62,n888);
not (n2372,n2176);
xor (n2373,n2374,n442);
or (n2374,n2375,n2376);
and (n2375,n194,n522);
and (n2376,n196,n526);
nand (n2377,n2378,n2379,n2380);
nand (n2378,n2237,n2241);
nand (n2379,n2245,n2241);
nand (n2380,n2237,n2245);
nor (n2381,n2382,n2489);
nor (n2382,n2383,n2387);
nand (n2383,n2384,n2385,n2386);
nand (n2384,n2274,n2278);
nand (n2385,n2282,n2278);
nand (n2386,n2274,n2282);
xor (n2387,n2388,n2485);
xor (n2388,n2389,n2429);
xor (n2389,n2390,n2425);
xor (n2390,n2391,n2421);
xor (n2391,n2392,n2417);
xor (n2392,n2393,n2407);
xor (n2393,n2394,n2403);
xor (n2394,n2395,n2399);
xor (n2395,n2396,n165);
or (n2396,n2397,n2398);
and (n2397,n196,n440);
and (n2398,n212,n444);
xor (n2399,n2400,n169);
or (n2400,n2401,n2402);
and (n2401,n266,n163);
and (n2402,n298,n167);
xor (n2403,n2404,n74);
or (n2404,n2405,n2406);
and (n2405,n560,n97);
and (n2406,n632,n101);
xor (n2407,n2408,n2413);
xor (n2408,n2409,n1006);
xor (n2409,n2410,n524);
or (n2410,n2411,n2412);
and (n2411,n62,n661);
and (n2412,n64,n665);
xor (n2413,n2414,n442);
or (n2414,n2415,n2416);
and (n2415,n111,n522);
and (n2416,n194,n526);
nand (n2417,n2418,n2419,n2420);
nand (n2418,n2292,n2296);
nand (n2419,n2297,n2296);
nand (n2420,n2292,n2297);
nand (n2421,n2422,n2423,n2424);
nand (n2422,n2286,n2290);
nand (n2423,n2301,n2290);
nand (n2424,n2286,n2301);
nand (n2425,n2426,n2427,n2428);
nand (n2426,n2317,n2321);
nand (n2427,n2325,n2321);
nand (n2428,n2317,n2325);
xor (n2429,n2430,n2481);
xor (n2430,n2431,n2452);
xor (n2431,n2432,n2448);
xor (n2432,n2433,n2444);
xor (n2433,n2434,n2440);
xor (n2434,n2435,n2436);
not (n2435,n1047);
xor (n2436,n2437,n99);
or (n2437,n2438,n2439);
and (n2438,n427,n173);
and (n2439,n514,n176);
xor (n2440,n2441,n22);
or (n2441,n2442,n2443);
and (n2442,n853,n72);
and (n2443,n857,n76);
nand (n2444,n2445,n2446,n2447);
nand (n2445,n2303,n2307);
nand (n2446,n2311,n2307);
nand (n2447,n2303,n2311);
nand (n2448,n2449,n2450,n2451);
nand (n2449,n2327,n2331);
nand (n2450,n13,n2331);
nand (n2451,n2327,n13);
xor (n2452,n2453,n2477);
xor (n2453,n2454,n2467);
xor (n2454,n2455,n2464);
xor (n2455,n2456,n2460);
xor (n2456,n2457,n9);
or (n2457,n2458,n2459);
and (n2458,n859,n20);
and (n2459,n993,n24);
xor (n2460,n2461,n13);
or (n2461,n2462,n2463);
and (n2462,n1197,n7);
and (n2463,n1201,n11);
nand (n2464,n2332,n2465,n2466);
nand (n2465,n2337,n2333);
not (n2466,n2337);
xor (n2467,n2468,n2473);
xor (n2468,n13,n2469);
nand (n2469,n2470,n2471,n2472);
nand (n2470,n2368,n2372);
nand (n2471,n2373,n2372);
nand (n2472,n2368,n2373);
nand (n2473,n2474,n2475,n2476);
nand (n2474,n2354,n2358);
nand (n2475,n2362,n2358);
nand (n2476,n2354,n2362);
nand (n2477,n2478,n2479,n2480);
nand (n2478,n2348,n2352);
nand (n2479,n2366,n2352);
nand (n2480,n2348,n2366);
nand (n2481,n2482,n2483,n2484);
nand (n2482,n2342,n2346);
nand (n2483,n2377,n2346);
nand (n2484,n2342,n2377);
nand (n2485,n2486,n2487,n2488);
nand (n2486,n2284,n2315);
nand (n2487,n2340,n2315);
nand (n2488,n2284,n2340);
nor (n2489,n2490,n2494);
nand (n2490,n2491,n2492,n2493);
nand (n2491,n2389,n2429);
nand (n2492,n2485,n2429);
nand (n2493,n2389,n2485);
xor (n2494,n2495,n2504);
xor (n2495,n2496,n2500);
nand (n2496,n2497,n2498,n2499);
nand (n2497,n2391,n2421);
nand (n2498,n2425,n2421);
nand (n2499,n2391,n2425);
nand (n2500,n2501,n2502,n2503);
nand (n2501,n2431,n2452);
nand (n2502,n2481,n2452);
nand (n2503,n2431,n2481);
xor (n2504,n2505,n2536);
xor (n2505,n2506,n2510);
nand (n2506,n2507,n2508,n2509);
nand (n2507,n2454,n2467);
nand (n2508,n2477,n2467);
nand (n2509,n2454,n2477);
xor (n2510,n2511,n2524);
xor (n2511,n2512,n2516);
nand (n2512,n2513,n2514,n2515);
nand (n2513,n13,n2469);
nand (n2514,n2473,n2469);
nand (n2515,n13,n2473);
xor (n2516,n2517,n2520);
xor (n2517,n2518,n13);
xor (n2518,n2519,n1005);
xor (n2519,n997,n1000);
nand (n2520,n2521,n2522,n2523);
nand (n2521,n2409,n1006);
nand (n2522,n2413,n1006);
nand (n2523,n2409,n2413);
xor (n2524,n2525,n2532);
xor (n2525,n2526,n2528);
xor (n2526,n2527,n1033);
xor (n2527,n1024,n1028);
nand (n2528,n2529,n2530,n2531);
nand (n2529,n2395,n2399);
nand (n2530,n2403,n2399);
nand (n2531,n2395,n2403);
nand (n2532,n2533,n2534,n2535);
nand (n2533,n2456,n2460);
nand (n2534,n2464,n2460);
nand (n2535,n2456,n2464);
xor (n2536,n2537,n2546);
xor (n2537,n2538,n2542);
nand (n2538,n2539,n2540,n2541);
nand (n2539,n2393,n2407);
nand (n2540,n2417,n2407);
nand (n2541,n2393,n2417);
nand (n2542,n2543,n2544,n2545);
nand (n2543,n2433,n2444);
nand (n2544,n2448,n2444);
nand (n2545,n2433,n2448);
xor (n2546,n2547,n2554);
xor (n2547,n2548,n2552);
nand (n2548,n2549,n2550,n2551);
nand (n2549,n2435,n2436);
nand (n2550,n2440,n2436);
nand (n2551,n2435,n2440);
xor (n2552,n2553,n1052);
xor (n2553,n1043,n1047);
xor (n2554,n2555,n2564);
xor (n2555,n2556,n2560);
xor (n2556,n2557,n22);
or (n2557,n2558,n2559);
and (n2558,n632,n72);
and (n2559,n853,n76);
xor (n2560,n2561,n9);
or (n2561,n2562,n2563);
and (n2562,n857,n20);
and (n2563,n859,n24);
xor (n2564,n2565,n13);
or (n2565,n2566,n2567);
and (n2566,n993,n7);
and (n2567,n1197,n11);
nand (n2568,n2569,n2653);
nor (n2569,n2570,n2620);
nor (n2570,n2571,n2575);
nand (n2571,n2572,n2573,n2574);
nand (n2572,n2496,n2500);
nand (n2573,n2504,n2500);
nand (n2574,n2496,n2504);
xor (n2575,n2576,n2616);
xor (n2576,n2577,n2597);
xor (n2577,n2578,n2585);
xor (n2578,n2579,n2581);
xor (n2579,n2580,n1041);
xor (n2580,n1022,n1038);
nand (n2581,n2582,n2583,n2584);
nand (n2582,n2548,n2552);
nand (n2583,n2554,n2552);
nand (n2584,n2548,n2554);
xor (n2585,n2586,n2593);
xor (n2586,n2587,n2591);
nand (n2587,n2588,n2589,n2590);
nand (n2588,n2556,n2560);
nand (n2589,n2564,n2560);
nand (n2590,n2556,n2564);
xor (n2591,n2592,n951);
xor (n2592,n945,n949);
nand (n2593,n2594,n2595,n2596);
nand (n2594,n2518,n13);
nand (n2595,n2520,n13);
nand (n2596,n2518,n2520);
xor (n2597,n2598,n2612);
xor (n2598,n2599,n2603);
nand (n2599,n2600,n2601,n2602);
nand (n2600,n2512,n2516);
nand (n2601,n2524,n2516);
nand (n2602,n2512,n2524);
xor (n2603,n2604,n2608);
xor (n2604,n2605,n2607);
xor (n2605,n2606,n967);
xor (n2606,n958,n962);
xor (n2607,n990,n995);
nand (n2608,n2609,n2610,n2611);
nand (n2609,n2526,n2528);
nand (n2610,n2532,n2528);
nand (n2611,n2526,n2532);
nand (n2612,n2613,n2614,n2615);
nand (n2613,n2538,n2542);
nand (n2614,n2546,n2542);
nand (n2615,n2538,n2546);
nand (n2616,n2617,n2618,n2619);
nand (n2617,n2506,n2510);
nand (n2618,n2536,n2510);
nand (n2619,n2506,n2536);
nor (n2620,n2621,n2625);
nand (n2621,n2622,n2623,n2624);
nand (n2622,n2577,n2597);
nand (n2623,n2616,n2597);
nand (n2624,n2577,n2616);
xor (n2625,n2626,n2649);
xor (n2626,n2627,n2637);
xor (n2627,n2628,n2635);
xor (n2628,n2629,n2631);
xor (n2629,n2630,n938);
xor (n2630,n923,n935);
nand (n2631,n2632,n2633,n2634);
nand (n2632,n2587,n2591);
nand (n2633,n2593,n2591);
nand (n2634,n2587,n2593);
xor (n2635,n2636,n973);
xor (n2636,n943,n956);
xor (n2637,n2638,n2645);
xor (n2638,n2639,n2641);
xor (n2639,n2640,n1020);
xor (n2640,n987,n1017);
nand (n2641,n2642,n2643,n2644);
nand (n2642,n2605,n2607);
nand (n2643,n2608,n2607);
nand (n2644,n2605,n2608);
nand (n2645,n2646,n2647,n2648);
nand (n2646,n2579,n2581);
nand (n2647,n2585,n2581);
nand (n2648,n2579,n2585);
nand (n2649,n2650,n2651,n2652);
nand (n2650,n2599,n2603);
nand (n2651,n2612,n2603);
nand (n2652,n2599,n2612);
nor (n2653,n2654,n2671);
nor (n2654,n2655,n2659);
nand (n2655,n2656,n2657,n2658);
nand (n2656,n2627,n2637);
nand (n2657,n2649,n2637);
nand (n2658,n2627,n2649);
xor (n2659,n2660,n2667);
xor (n2660,n2661,n2665);
nand (n2661,n2662,n2663,n2664);
nand (n2662,n2629,n2631);
nand (n2663,n2635,n2631);
nand (n2664,n2629,n2635);
xor (n2665,n2666,n1060);
xor (n2666,n983,n985);
nand (n2667,n2668,n2669,n2670);
nand (n2668,n2639,n2641);
nand (n2669,n2645,n2641);
nand (n2670,n2639,n2645);
nor (n2671,n2672,n2676);
nand (n2672,n2673,n2674,n2675);
nand (n2673,n2661,n2665);
nand (n2674,n2667,n2665);
nand (n2675,n2661,n2667);
xor (n2676,n2677,n981);
xor (n2677,n759,n843);
not (n2678,n2679);
nor (n2679,n2680,n2695);
nor (n2680,n2568,n2681);
nor (n2681,n2682,n2689);
nor (n2682,n2683,n2688);
nor (n2683,n2684,n2686);
nor (n2684,n2685,n2267);
nand (n2685,n2156,n2160);
not (n2686,n2687);
nand (n2687,n2268,n2272);
not (n2688,n2381);
not (n2689,n2690);
nor (n2690,n2691,n2693);
nor (n2691,n2692,n2489);
nand (n2692,n2383,n2387);
not (n2693,n2694);
nand (n2694,n2490,n2494);
not (n2695,n2696);
nor (n2696,n2697,n2704);
nor (n2697,n2698,n2703);
nor (n2698,n2699,n2701);
nor (n2699,n2700,n2620);
nand (n2700,n2571,n2575);
not (n2701,n2702);
nand (n2702,n2621,n2625);
not (n2703,n2653);
not (n2704,n2705);
nor (n2705,n2706,n2708);
nor (n2706,n2707,n2671);
nand (n2707,n2655,n2659);
not (n2708,n2709);
nand (n2709,n2672,n2676);
nand (n2710,n2711,n3130);
nand (n2711,n2712,n3023);
nor (n2712,n2713,n3008);
nor (n2713,n2714,n2879);
nand (n2714,n2715,n2856);
nor (n2715,n2716,n2833);
nor (n2716,n2717,n2806);
nand (n2717,n2718,n2763,n2805);
nand (n2718,n2719,n2731);
xor (n2719,n2720,n2726);
xor (n2720,n2721,n2722);
xor (n2721,n2024,n2028);
xor (n2722,n2723,n165);
or (n2723,n2724,n2725);
and (n2724,n1226,n440);
and (n2725,n1240,n444);
and (n2726,n165,n2727);
xor (n2727,n2728,n886);
or (n2728,n2729,n2730);
and (n2729,n853,n1009);
and (n2730,n857,n1013);
nand (n2731,n2732,n2749,n2762);
nand (n2732,n2733,n2734);
xor (n2733,n165,n2727);
nand (n2734,n2735,n2744,n2748);
nand (n2735,n2736,n2740);
xor (n2736,n2737,n524);
or (n2737,n2738,n2739);
and (n2738,n1201,n661);
and (n2739,n1203,n665);
xor (n2740,n2741,n663);
or (n2741,n2742,n2743);
and (n2742,n993,n884);
and (n2743,n1197,n888);
nand (n2744,n2745,n2740);
and (n2745,n442,n2746);
xnor (n2746,n2747,n442);
nand (n2747,n1240,n522);
nand (n2748,n2736,n2745);
nand (n2749,n2750,n2734);
xor (n2750,n2751,n2758);
xor (n2751,n2752,n2756);
xnor (n2752,n2753,n1011);
nor (n2753,n2754,n2755);
and (n2754,n632,n1212);
and (n2755,n560,n1214);
xnor (n2756,n2757,n165);
nand (n2757,n1240,n440);
xor (n2758,n2759,n524);
or (n2759,n2760,n2761);
and (n2760,n1197,n661);
and (n2761,n1201,n665);
nand (n2762,n2733,n2750);
nand (n2763,n2764,n2731);
xor (n2764,n2765,n2784);
xor (n2765,n2766,n2770);
nand (n2766,n2767,n2768,n2769);
nand (n2767,n2752,n2756);
nand (n2768,n2758,n2756);
nand (n2769,n2752,n2758);
xor (n2770,n2771,n2780);
xor (n2771,n2772,n2776);
xor (n2772,n2773,n524);
or (n2773,n2774,n2775);
and (n2774,n993,n661);
and (n2775,n1197,n665);
xor (n2776,n2777,n663);
or (n2777,n2778,n2779);
and (n2778,n857,n884);
and (n2779,n859,n888);
xor (n2780,n2781,n442);
or (n2781,n2782,n2783);
and (n2782,n1201,n522);
and (n2783,n1203,n526);
nand (n2784,n2785,n2799,n2804);
nand (n2785,n2786,n2790);
xor (n2786,n2787,n663);
or (n2787,n2788,n2789);
and (n2788,n859,n884);
and (n2789,n993,n888);
and (n2790,n2791,n2795);
xnor (n2791,n2792,n1011);
nor (n2792,n2793,n2794);
and (n2793,n853,n1212);
and (n2794,n632,n1214);
xor (n2795,n2796,n886);
or (n2796,n2797,n2798);
and (n2797,n857,n1009);
and (n2798,n859,n1013);
nand (n2799,n2800,n2790);
xor (n2800,n2801,n442);
or (n2801,n2802,n2803);
and (n2802,n1203,n522);
and (n2803,n1226,n526);
nand (n2804,n2786,n2800);
nand (n2805,n2719,n2764);
xor (n2806,n2807,n2821);
xor (n2807,n2808,n2817);
xor (n2808,n2809,n2815);
xor (n2809,n2810,n2814);
xor (n2810,n2811,n165);
or (n2811,n2812,n2813);
and (n2812,n1203,n440);
and (n2813,n1226,n444);
xor (n2814,n1968,n169);
xor (n2815,n2816,n2011);
xor (n2816,n2004,n2008);
nand (n2817,n2818,n2819,n2820);
nand (n2818,n2766,n2770);
nand (n2819,n2784,n2770);
nand (n2820,n2766,n2784);
xor (n2821,n2822,n2831);
xor (n2822,n2823,n2827);
nand (n2823,n2824,n2825,n2826);
nand (n2824,n2721,n2722);
nand (n2825,n2726,n2722);
nand (n2826,n2721,n2726);
nand (n2827,n2828,n2829,n2830);
nand (n2828,n2772,n2776);
nand (n2829,n2780,n2776);
nand (n2830,n2772,n2780);
xor (n2831,n2832,n2033);
xor (n2832,n2019,n2023);
nor (n2833,n2834,n2838);
nand (n2834,n2835,n2836,n2837);
nand (n2835,n2808,n2817);
nand (n2836,n2821,n2817);
nand (n2837,n2808,n2821);
xor (n2838,n2839,n2846);
xor (n2839,n2840,n2842);
xor (n2840,n2841,n2017);
xor (n2841,n1998,n2002);
nand (n2842,n2843,n2844,n2845);
nand (n2843,n2823,n2827);
nand (n2844,n2831,n2827);
nand (n2845,n2823,n2831);
xor (n2846,n2847,n2852);
xor (n2847,n2848,n2850);
xor (n2848,n2849,n1967);
xor (n2849,n1958,n1962);
xor (n2850,n2851,n1982);
xor (n2851,n1976,n1980);
nand (n2852,n2853,n2854,n2855);
nand (n2853,n2810,n2814);
nand (n2854,n2815,n2814);
nand (n2855,n2810,n2815);
nor (n2856,n2857,n2872);
nor (n2857,n2858,n2862);
nand (n2858,n2859,n2860,n2861);
nand (n2859,n2840,n2842);
nand (n2860,n2846,n2842);
nand (n2861,n2840,n2846);
xor (n2862,n2863,n2870);
xor (n2863,n2864,n2866);
xor (n2864,n2865,n1974);
xor (n2865,n1954,n1956);
nand (n2866,n2867,n2868,n2869);
nand (n2867,n2848,n2850);
nand (n2868,n2852,n2850);
nand (n2869,n2848,n2852);
xor (n2870,n2871,n1996);
xor (n2871,n1991,n1993);
nor (n2872,n2873,n2877);
nand (n2873,n2874,n2875,n2876);
nand (n2874,n2864,n2866);
nand (n2875,n2870,n2866);
nand (n2876,n2864,n2870);
xor (n2877,n2878,n1989);
xor (n2878,n1864,n1915);
nor (n2879,n2880,n3002);
nor (n2880,n2881,n2978);
nor (n2881,n2882,n2975);
nor (n2882,n2883,n2951);
nand (n2883,n2884,n2923);
or (n2884,n2885,n2909,n2922);
and (n2885,n2886,n2895);
xor (n2886,n2887,n2891);
xnor (n2887,n2888,n1011);
nor (n2888,n2889,n2890);
and (n2889,n859,n1212);
and (n2890,n857,n1214);
xnor (n2891,n2892,n886);
nor (n2892,n2893,n2894);
and (n2893,n1197,n1013);
and (n2894,n993,n1009);
or (n2895,n2896,n2903,n2908);
and (n2896,n2897,n2899);
not (n2897,n2898);
nand (n2898,n1240,n661);
xnor (n2899,n2900,n1011);
nor (n2900,n2901,n2902);
and (n2901,n993,n1212);
and (n2902,n859,n1214);
and (n2903,n2899,n2904);
xnor (n2904,n2905,n886);
nor (n2905,n2906,n2907);
and (n2906,n1201,n1013);
and (n2907,n1197,n1009);
and (n2908,n2897,n2904);
and (n2909,n2895,n2910);
xor (n2910,n2911,n2918);
xor (n2911,n2912,n2914);
and (n2912,n524,n2913);
xnor (n2913,n2898,n524);
xnor (n2914,n2915,n663);
nor (n2915,n2916,n2917);
and (n2916,n1203,n888);
and (n2917,n1201,n884);
xnor (n2918,n2919,n524);
nor (n2919,n2920,n2921);
and (n2920,n1240,n665);
and (n2921,n1226,n661);
and (n2922,n2886,n2910);
xor (n2923,n2924,n2940);
xor (n2924,n2925,n2929);
or (n2925,n2926,n2927,n2928);
and (n2926,n2912,n2914);
and (n2927,n2914,n2918);
and (n2928,n2912,n2918);
xor (n2929,n2930,n2936);
xor (n2930,n2931,n2932);
and (n2931,n2887,n2891);
xnor (n2932,n2933,n663);
nor (n2933,n2934,n2935);
and (n2934,n1201,n888);
and (n2935,n1197,n884);
xnor (n2936,n2937,n524);
nor (n2937,n2938,n2939);
and (n2938,n1226,n665);
and (n2939,n1203,n661);
xor (n2940,n2941,n2947);
xor (n2941,n2942,n2943);
not (n2942,n2747);
xnor (n2943,n2944,n1011);
nor (n2944,n2945,n2946);
and (n2945,n857,n1212);
and (n2946,n853,n1214);
xnor (n2947,n2948,n886);
nor (n2948,n2949,n2950);
and (n2949,n993,n1013);
and (n2950,n859,n1009);
nor (n2951,n2952,n2956);
or (n2952,n2953,n2954,n2955);
and (n2953,n2925,n2929);
and (n2954,n2929,n2940);
and (n2955,n2925,n2940);
xor (n2956,n2957,n2964);
xor (n2957,n2958,n2962);
or (n2958,n2959,n2960,n2961);
and (n2959,n2931,n2932);
and (n2960,n2932,n2936);
and (n2961,n2931,n2936);
xor (n2962,n2963,n2745);
xor (n2963,n2736,n2740);
xor (n2964,n2965,n2971);
xor (n2965,n2966,n2970);
xor (n2966,n2967,n442);
or (n2967,n2968,n2969);
and (n2968,n1226,n522);
and (n2969,n1240,n526);
xor (n2970,n2791,n2795);
or (n2971,n2972,n2973,n2974);
and (n2972,n2942,n2943);
and (n2973,n2943,n2947);
and (n2974,n2942,n2947);
not (n2975,n2976);
not (n2976,n2977);
and (n2977,n2952,n2956);
not (n2978,n2979);
nor (n2979,n2980,n2995);
nor (n2980,n2981,n2985);
nand (n2981,n2982,n2983,n2984);
nand (n2982,n2958,n2962);
nand (n2983,n2964,n2962);
nand (n2984,n2958,n2964);
xor (n2985,n2986,n2993);
xor (n2986,n2987,n2989);
xor (n2987,n2988,n2800);
xor (n2988,n2786,n2790);
nand (n2989,n2990,n2991,n2992);
nand (n2990,n2966,n2970);
nand (n2991,n2971,n2970);
nand (n2992,n2966,n2971);
xor (n2993,n2994,n2750);
xor (n2994,n2733,n2734);
nor (n2995,n2996,n3000);
nand (n2996,n2997,n2998,n2999);
nand (n2997,n2987,n2989);
nand (n2998,n2993,n2989);
nand (n2999,n2987,n2993);
xor (n3000,n3001,n2764);
xor (n3001,n2719,n2731);
not (n3002,n3003);
nor (n3003,n3004,n3006);
nor (n3004,n3005,n2995);
nand (n3005,n2981,n2985);
not (n3006,n3007);
nand (n3007,n2996,n3000);
not (n3008,n3009);
nor (n3009,n3010,n3017);
nor (n3010,n3011,n3016);
nor (n3011,n3012,n3014);
nor (n3012,n3013,n2833);
nand (n3013,n2717,n2806);
not (n3014,n3015);
nand (n3015,n2834,n2838);
not (n3016,n2856);
not (n3017,n3018);
nor (n3018,n3019,n3021);
nor (n3019,n3020,n2872);
nand (n3020,n2858,n2862);
not (n3021,n3022);
nand (n3022,n2873,n2877);
nand (n3023,n3024,n3028);
nor (n3024,n3025,n2714);
nand (n3025,n3026,n2979);
nor (n3026,n3027,n2951);
nor (n3027,n2884,n2923);
or (n3028,n3029,n3051);
and (n3029,n3030,n3032);
xor (n3030,n3031,n2910);
xor (n3031,n2886,n2895);
or (n3032,n3033,n3047,n3050);
and (n3033,n3034,n3043);
and (n3034,n3035,n3039);
xnor (n3035,n3036,n1011);
nor (n3036,n3037,n3038);
and (n3037,n1197,n1212);
and (n3038,n993,n1214);
xnor (n3039,n3040,n886);
nor (n3040,n3041,n3042);
and (n3041,n1203,n1013);
and (n3042,n1201,n1009);
xnor (n3043,n3044,n663);
nor (n3044,n3045,n3046);
and (n3045,n1226,n888);
and (n3046,n1203,n884);
and (n3047,n3043,n3048);
xor (n3048,n3049,n2904);
xor (n3049,n2897,n2899);
and (n3050,n3034,n3048);
and (n3051,n3052,n3053);
xor (n3052,n3030,n3032);
or (n3053,n3054,n3069);
and (n3054,n3055,n3067);
or (n3055,n3056,n3061,n3066);
and (n3056,n3057,n3058);
xor (n3057,n3035,n3039);
and (n3058,n663,n3059);
xnor (n3059,n3060,n663);
nand (n3060,n1240,n884);
and (n3061,n3058,n3062);
xnor (n3062,n3063,n663);
nor (n3063,n3064,n3065);
and (n3064,n1240,n888);
and (n3065,n1226,n884);
and (n3066,n3057,n3062);
xor (n3067,n3068,n3048);
xor (n3068,n3034,n3043);
and (n3069,n3070,n3071);
xor (n3070,n3055,n3067);
or (n3071,n3072,n3088);
and (n3072,n3073,n3075);
xor (n3073,n3074,n3062);
xor (n3074,n3057,n3058);
or (n3075,n3076,n3082,n3087);
and (n3076,n3077,n3078);
not (n3077,n3060);
xnor (n3078,n3079,n1011);
nor (n3079,n3080,n3081);
and (n3080,n1201,n1212);
and (n3081,n1197,n1214);
and (n3082,n3078,n3083);
xnor (n3083,n3084,n886);
nor (n3084,n3085,n3086);
and (n3085,n1226,n1013);
and (n3086,n1203,n1009);
and (n3087,n3077,n3083);
and (n3088,n3089,n3090);
xor (n3089,n3073,n3075);
or (n3090,n3091,n3102);
and (n3091,n3092,n3094);
xor (n3092,n3093,n3083);
xor (n3093,n3077,n3078);
and (n3094,n3095,n3098);
and (n3095,n886,n3096);
xnor (n3096,n3097,n886);
nand (n3097,n1240,n1009);
xnor (n3098,n3099,n1011);
nor (n3099,n3100,n3101);
and (n3100,n1203,n1212);
and (n3101,n1201,n1214);
and (n3102,n3103,n3104);
xor (n3103,n3092,n3094);
or (n3104,n3105,n3111);
and (n3105,n3106,n3110);
xnor (n3106,n3107,n886);
nor (n3107,n3108,n3109);
and (n3108,n1240,n1013);
and (n3109,n1226,n1009);
xor (n3110,n3095,n3098);
and (n3111,n3112,n3113);
xor (n3112,n3106,n3110);
or (n3113,n3114,n3120);
and (n3114,n3115,n3119);
xnor (n3115,n3116,n1011);
nor (n3116,n3117,n3118);
and (n3117,n1226,n1212);
and (n3118,n1203,n1214);
not (n3119,n3097);
and (n3120,n3121,n3122);
xor (n3121,n3115,n3119);
and (n3122,n3123,n3127);
xnor (n3123,n3124,n1011);
nor (n3124,n3125,n3126);
and (n3125,n1240,n1212);
and (n3126,n1226,n1214);
and (n3127,n3128,n1011);
xnor (n3128,n3129,n1011);
nand (n3129,n1240,n1214);
not (n3130,n3131);
nand (n3131,n3132,n2152);
nor (n3132,n3133,n1184);
nand (n3133,n3134,n2107);
nor (n3134,n3135,n2079);
nor (n3135,n1862,n2041);
not (n3136,n3137);
nand (n3137,n3138,n373);
nor (n3138,n3139,n345);
nor (n3139,n153,n309);
not (n3140,n3141);
nor (n3141,n2,n32);
xor (n3142,n3143,n3155);
xor (n3143,n3144,n3146);
not (n3144,n3145);
xnor (n3145,n3,n13);
or (n3146,n3145,n3147);
or (n3147,n3148,n3149,n3154);
not (n3148,n15);
and (n3149,n26,n3150);
or (n3150,n3151,n3152,n3153);
and (n3151,n17,n39);
and (n3152,n39,n126);
and (n3153,n17,n126);
and (n3154,n16,n3150);
and (n3155,n3156,n3157);
xnor (n3156,n3145,n3147);
or (n3157,n3158,n3462);
and (n3158,n3159,n3160);
xor (n3159,n35,n3150);
or (n3160,n3161,n3177,n3461);
and (n3161,n3162,n3164);
xor (n3162,n3163,n126);
xor (n3163,n17,n39);
or (n3164,n3165,n3167,n3176);
and (n3165,n3166,n78);
not (n3166,n54);
and (n3167,n78,n3168);
or (n3168,n3169,n3170,n3175);
and (n3169,n69,n378);
and (n3170,n378,n3171);
or (n3171,n3172,n3173,n3174);
not (n3172,n92);
and (n3173,n103,n116);
and (n3174,n93,n116);
and (n3175,n69,n3171);
and (n3176,n3166,n3168);
and (n3177,n3164,n3178);
or (n3178,n3179,n3219,n3460);
and (n3179,n3180,n3182);
xor (n3180,n3181,n3168);
xor (n3181,n3166,n78);
or (n3182,n3183,n3191,n3218);
and (n3183,n3184,n3189);
or (n3184,n3185,n3186,n3188);
and (n3185,n107,n354);
and (n3186,n354,n3187);
xor (n3187,n359,n116);
and (n3188,n107,n3187);
xor (n3189,n3190,n3171);
xor (n3190,n69,n378);
and (n3191,n3189,n3192);
or (n3192,n3193,n3201,n3217);
and (n3193,n3194,n3199);
or (n3194,n3195,n3196,n3198);
and (n3195,n94,n317);
and (n3196,n317,n3197);
not (n3197,n332);
and (n3198,n94,n3197);
xor (n3199,n3200,n3187);
xor (n3200,n107,n354);
and (n3201,n3199,n3202);
or (n3202,n3203,n3213,n3216);
and (n3203,n3204,n3208);
or (n3204,n3205,n3206,n3207);
and (n3205,n201,n248);
not (n3206,n339);
and (n3207,n201,n251);
or (n3208,n3209,n3210,n3212);
and (n3209,n247,n230);
and (n3210,n230,n3211);
not (n3211,n217);
and (n3212,n247,n3211);
and (n3213,n3208,n3214);
xor (n3214,n3215,n3197);
xor (n3215,n94,n317);
and (n3216,n3204,n3214);
and (n3217,n3194,n3202);
and (n3218,n3184,n3192);
and (n3219,n3182,n3220);
or (n3220,n3221,n3223);
xor (n3221,n3222,n3192);
xor (n3222,n3184,n3189);
or (n3223,n3224,n3255,n3459);
and (n3224,n3225,n3227);
xor (n3225,n3226,n3202);
xor (n3226,n3194,n3199);
or (n3227,n3228,n3240,n3254);
and (n3228,n3229,n3238);
or (n3229,n3230,n3235,n3237);
and (n3230,n3231,n223);
or (n3231,n3232,n3233,n3234);
and (n3232,n247,n204);
not (n3233,n243);
and (n3234,n247,n208);
and (n3235,n223,n3236);
not (n3236,n245);
and (n3237,n3231,n3236);
xor (n3238,n3239,n3214);
xor (n3239,n3204,n3208);
and (n3240,n3238,n3241);
or (n3241,n3242,n3250,n3253);
and (n3242,n3243,n3248);
or (n3243,n3244,n3246,n3247);
and (n3244,n3245,n259);
not (n3245,n199);
and (n3246,n259,n157);
and (n3247,n3245,n157);
xor (n3248,n3249,n3211);
xor (n3249,n247,n230);
and (n3250,n3248,n3251);
xor (n3251,n3252,n3236);
xor (n3252,n3231,n223);
and (n3253,n3243,n3251);
and (n3254,n3229,n3241);
and (n3255,n3227,n3256);
or (n3256,n3257,n3345,n3458);
and (n3257,n3258,n3260);
xor (n3258,n3259,n3241);
xor (n3259,n3229,n3238);
or (n3260,n3261,n3282,n3344);
and (n3261,n3262,n3280);
or (n3262,n3263,n3276,n3279);
and (n3263,n3264,n3268);
or (n3264,n3265,n3266,n3267);
not (n3265,n197);
and (n3266,n191,n262);
and (n3267,n186,n262);
or (n3268,n3269,n3274,n3275);
and (n3269,n268,n3270);
or (n3270,n3271,n3272,n3273);
and (n3271,n160,n290);
not (n3272,n289);
and (n3273,n160,n294);
and (n3274,n3270,n301);
and (n3275,n268,n301);
and (n3276,n3268,n3277);
xor (n3277,n3278,n157);
xor (n3278,n3245,n259);
and (n3279,n3264,n3277);
xor (n3280,n3281,n3251);
xor (n3281,n3243,n3248);
and (n3282,n3280,n3283);
or (n3283,n3284,n3297,n3343);
and (n3284,n3285,n3295);
or (n3285,n3286,n3291,n3294);
and (n3286,n3287,n3289);
xor (n3287,n3288,n262);
xor (n3288,n186,n191);
and (n3289,n413,n3290);
not (n3290,n415);
and (n3291,n3289,n3292);
xor (n3292,n3293,n301);
xor (n3293,n268,n3270);
and (n3294,n3287,n3292);
xor (n3295,n3296,n3277);
xor (n3296,n3264,n3268);
and (n3297,n3295,n3298);
or (n3298,n3299,n3312,n3342);
and (n3299,n3300,n3310);
or (n3300,n3301,n3307,n3309);
and (n3301,n3302,n3303);
not (n3302,n418);
or (n3303,n3304,n3305,n3306);
not (n3304,n435);
and (n3305,n446,n457);
and (n3306,n436,n457);
and (n3307,n3303,n3308);
not (n3308,n412);
and (n3309,n3302,n3308);
xor (n3310,n3311,n3292);
xor (n3311,n3287,n3289);
and (n3312,n3310,n3313);
or (n3313,n3314,n3328,n3341);
and (n3314,n3315,n3319);
or (n3315,n3316,n3317,n3318);
and (n3316,n450,n462);
and (n3317,n462,n504);
and (n3318,n450,n504);
or (n3319,n3320,n3325,n3327);
and (n3320,n471,n3321);
or (n3321,n3322,n3323,n3324);
and (n3322,n437,n490);
not (n3323,n494);
and (n3324,n437,n495);
and (n3325,n3321,n3326);
xor (n3326,n470,n457);
and (n3327,n471,n3326);
and (n3328,n3319,n3329);
or (n3329,n3330,n3337,n3340);
and (n3330,n3331,n3332);
not (n3331,n542);
or (n3332,n3333,n3335,n3336);
and (n3333,n510,n3334);
not (n3334,n586);
and (n3335,n3334,n516);
not (n3336,n537);
and (n3337,n3332,n3338);
xor (n3338,n3339,n504);
xor (n3339,n450,n462);
and (n3340,n3331,n3338);
and (n3341,n3315,n3329);
and (n3342,n3300,n3313);
and (n3343,n3285,n3298);
and (n3344,n3262,n3283);
and (n3345,n3260,n3346);
or (n3346,n3347,n3349);
xor (n3347,n3348,n3283);
xor (n3348,n3262,n3280);
or (n3349,n3350,n3352);
xor (n3350,n3351,n3298);
xor (n3351,n3285,n3295);
or (n3352,n3353,n3385,n3457);
and (n3353,n3354,n3383);
or (n3354,n3355,n3379,n3382);
and (n3355,n3356,n3358);
xor (n3356,n3357,n3308);
xor (n3357,n3302,n3303);
or (n3358,n3359,n3375,n3378);
and (n3359,n3360,n3362);
xor (n3360,n3361,n3326);
xor (n3361,n471,n3321);
or (n3362,n3363,n3369,n3374);
and (n3363,n619,n3364);
and (n3364,n3365,n635);
or (n3365,n3366,n3367,n3368);
and (n3366,n519,n624);
not (n3367,n623);
and (n3368,n519,n628);
and (n3369,n3364,n3370);
or (n3370,n3371,n3372,n3373);
not (n3371,n569);
and (n3372,n570,n595);
and (n3373,n565,n595);
and (n3374,n619,n3370);
and (n3375,n3362,n3376);
xor (n3376,n3377,n3338);
xor (n3377,n3331,n3332);
and (n3378,n3360,n3376);
and (n3379,n3358,n3380);
xor (n3380,n3381,n3329);
xor (n3381,n3315,n3319);
and (n3382,n3356,n3380);
xor (n3383,n3384,n3313);
xor (n3384,n3300,n3310);
and (n3385,n3383,n3386);
or (n3386,n3387,n3389);
xor (n3387,n3388,n3380);
xor (n3388,n3356,n3358);
or (n3389,n3390,n3421,n3456);
and (n3390,n3391,n3419);
or (n3391,n3392,n3401,n3418);
and (n3392,n3393,n3395);
xor (n3393,n3394,n516);
xor (n3394,n510,n3334);
or (n3395,n3396,n3398,n3400);
and (n3396,n3397,n592);
not (n3397,n645);
and (n3398,n592,n3399);
xor (n3399,n3365,n635);
and (n3400,n3397,n3399);
and (n3401,n3395,n3402);
or (n3402,n3403,n3414,n3417);
and (n3403,n3404,n3409);
or (n3404,n3405,n3407,n3408);
and (n3405,n679,n3406);
not (n3406,n1084);
and (n3407,n3406,n1083);
and (n3408,n679,n1083);
or (n3409,n3410,n3412,n3413);
and (n3410,n682,n3411);
not (n3411,n1079);
and (n3412,n3411,n655);
and (n3413,n682,n655);
and (n3414,n3409,n3415);
xor (n3415,n3416,n595);
xor (n3416,n565,n570);
and (n3417,n3404,n3415);
and (n3418,n3393,n3402);
xor (n3419,n3420,n3376);
xor (n3420,n3360,n3362);
and (n3421,n3419,n3422);
or (n3422,n3423,n3452,n3455);
and (n3423,n3424,n3426);
xor (n3424,n3425,n3370);
xor (n3425,n619,n3364);
or (n3426,n3427,n3448,n3451);
and (n3427,n3428,n3446);
or (n3428,n3429,n3442,n3445);
and (n3429,n3430,n3434);
or (n3430,n3431,n3432,n3433);
and (n3431,n763,n837);
and (n3432,n837,n906);
and (n3433,n763,n906);
or (n3434,n3435,n3436,n3441);
and (n3435,n767,n839);
and (n3436,n839,n3437);
or (n3437,n3438,n3439,n3440);
and (n3438,n658,n868);
not (n3439,n904);
and (n3440,n658,n864);
and (n3441,n767,n3437);
and (n3442,n3434,n3443);
xor (n3443,n3444,n1083);
xor (n3444,n679,n3406);
and (n3445,n3430,n3443);
xor (n3446,n3447,n3399);
xor (n3447,n3397,n592);
and (n3448,n3446,n3449);
xor (n3449,n3450,n3415);
xor (n3450,n3404,n3409);
and (n3451,n3428,n3449);
and (n3452,n3426,n3453);
xor (n3453,n3454,n3402);
xor (n3454,n3393,n3395);
and (n3455,n3424,n3453);
and (n3456,n3391,n3422);
and (n3457,n3354,n3386);
and (n3458,n3258,n3346);
and (n3459,n3225,n3256);
and (n3460,n3180,n3220);
and (n3461,n3162,n3178);
and (n3462,n3463,n3464);
xor (n3463,n3159,n3160);
or (n3464,n3465,n3467);
xor (n3465,n3466,n3178);
xor (n3466,n3162,n3164);
and (n3467,n3468,n3469);
not (n3468,n3465);
and (n3469,n3470,n3472);
xor (n3470,n3471,n3220);
xor (n3471,n3180,n3182);
and (n3472,n3473,n3474);
xnor (n3473,n3221,n3223);
and (n3474,n3475,n3477);
xor (n3475,n3476,n3256);
xor (n3476,n3225,n3227);
and (n3477,n3478,n3480);
xor (n3478,n3479,n3346);
xor (n3479,n3258,n3260);
and (n3480,n3481,n3482);
xnor (n3481,n3347,n3349);
and (n3482,n3483,n3484);
xnor (n3483,n3350,n3352);
and (n3484,n3485,n3487);
xor (n3485,n3486,n3386);
xor (n3486,n3354,n3383);
and (n3487,n3488,n3489);
xnor (n3488,n3387,n3389);
or (n3489,n3490,n3570);
and (n3490,n3491,n3493);
xor (n3491,n3492,n3422);
xor (n3492,n3391,n3419);
or (n3493,n3494,n3496);
xor (n3494,n3495,n3453);
xor (n3495,n3424,n3426);
or (n3496,n3497,n3520,n3569);
and (n3497,n3498,n3518);
or (n3498,n3499,n3514,n3517);
and (n3499,n3500,n3502);
xor (n3500,n3501,n655);
xor (n3501,n682,n3411);
or (n3502,n3503,n3510,n3513);
and (n3503,n835,n3504);
or (n3504,n3505,n3507,n3509);
and (n3505,n896,n3506);
not (n3506,n862);
and (n3507,n3506,n3508);
not (n3508,n848);
and (n3509,n896,n3508);
and (n3510,n3504,n3511);
xor (n3511,n3512,n906);
xor (n3512,n763,n837);
and (n3513,n835,n3511);
and (n3514,n3502,n3515);
xor (n3515,n3516,n3443);
xor (n3516,n3430,n3434);
and (n3517,n3500,n3515);
xor (n3518,n3519,n3449);
xor (n3519,n3428,n3446);
and (n3520,n3518,n3521);
or (n3521,n3522,n3533,n3568);
and (n3522,n3523,n3531);
or (n3523,n3524,n3527,n3530);
and (n3524,n3525,n783);
xor (n3525,n3526,n3437);
xor (n3526,n767,n839);
and (n3527,n783,n3528);
xor (n3528,n3529,n3511);
xor (n3529,n835,n3504);
and (n3530,n3525,n3528);
xor (n3531,n3532,n3515);
xor (n3532,n3500,n3502);
and (n3533,n3531,n3534);
or (n3534,n3535,n3564,n3567);
and (n3535,n3536,n3549);
or (n3536,n3537,n3547,n3548);
and (n3537,n3538,n941);
or (n3538,n3539,n3544,n3546);
and (n3539,n3540,n935);
or (n3540,n3541,n3542,n3543);
and (n3541,n880,n925);
not (n3542,n929);
and (n3543,n880,n930);
and (n3544,n935,n3545);
not (n3545,n938);
and (n3546,n3540,n3545);
not (n3547,n976);
and (n3548,n3538,n977);
or (n3549,n3550,n3557,n3563);
and (n3550,n3551,n3555);
or (n3551,n3552,n3553,n3554);
and (n3552,n881,n877);
not (n3553,n895);
and (n3554,n881,n891);
xor (n3555,n3556,n3508);
xor (n3556,n896,n3506);
and (n3557,n3555,n3558);
or (n3558,n3559,n3560,n3562);
and (n3559,n880,n1018);
and (n3560,n1018,n3561);
not (n3561,n2632);
and (n3562,n880,n3561);
and (n3563,n3551,n3558);
and (n3564,n3549,n3565);
xor (n3565,n3566,n3528);
xor (n3566,n3525,n783);
and (n3567,n3536,n3565);
and (n3568,n3523,n3534);
and (n3569,n3498,n3521);
and (n3570,n3571,n3572);
xor (n3571,n3491,n3493);
and (n3572,n3573,n3574);
xnor (n3573,n3494,n3496);
or (n3574,n3575,n3660);
and (n3575,n3576,n3578);
xor (n3576,n3577,n3521);
xor (n3577,n3498,n3518);
or (n3578,n3579,n3581);
xor (n3579,n3580,n3534);
xor (n3580,n3523,n3531);
or (n3581,n3582,n3604,n3659);
and (n3582,n3583,n3602);
or (n3583,n3584,n3598,n3601);
and (n3584,n3585,n3587);
xor (n3585,n3586,n977);
xor (n3586,n3538,n941);
or (n3587,n3588,n3591,n3597);
and (n3588,n3589,n2635);
xor (n3589,n3590,n3545);
xor (n3590,n3540,n935);
and (n3591,n2635,n3592);
or (n3592,n3593,n3594,n3596);
not (n3593,n1057);
and (n3594,n1041,n3595);
not (n3595,n1038);
and (n3596,n1022,n3595);
and (n3597,n3589,n3592);
and (n3598,n3587,n3599);
xor (n3599,n3600,n3558);
xor (n3600,n3551,n3555);
and (n3601,n3585,n3599);
xor (n3602,n3603,n3565);
xor (n3603,n3536,n3549);
and (n3604,n3602,n3605);
or (n3605,n3606,n3621,n3658);
and (n3606,n3607,n3619);
or (n3607,n3608,n3615,n3618);
and (n3608,n3609,n3613);
or (n3609,n3610,n3611,n3612);
and (n3610,n989,n2605);
and (n3611,n2605,n2586);
and (n3612,n989,n2586);
xor (n3613,n3614,n3561);
xor (n3614,n880,n1018);
and (n3615,n3613,n3616);
and (n3616,n2581,n3617);
not (n3617,n2579);
and (n3618,n3609,n3616);
xor (n3619,n3620,n3599);
xor (n3620,n3585,n3587);
and (n3621,n3619,n3622);
or (n3622,n3623,n3643,n3657);
and (n3623,n3624,n3641);
or (n3624,n3625,n3630,n3640);
and (n3625,n3626,n2608);
or (n3626,n3627,n3628,n3629);
and (n3627,n1006,n997);
not (n3628,n996);
and (n3629,n1006,n1000);
and (n3630,n2608,n3631);
or (n3631,n3632,n3637,n3639);
and (n3632,n1005,n3633);
or (n3633,n3634,n3635,n3636);
and (n3634,n1005,n2409);
not (n3635,n2523);
and (n3636,n1005,n2413);
and (n3637,n3633,n3638);
not (n3638,n2518);
and (n3639,n1005,n3638);
and (n3640,n3626,n3631);
xor (n3641,n3642,n3592);
xor (n3642,n3589,n2635);
and (n3643,n3641,n3644);
or (n3644,n3645,n3649,n3656);
and (n3645,n3646,n3648);
xor (n3646,n3647,n2586);
xor (n3647,n989,n2605);
not (n3648,n2578);
and (n3649,n3648,n3650);
or (n3650,n3651,n3654,n3655);
and (n3651,n3652,n2524);
and (n3652,n2393,n3653);
not (n3653,n2407);
and (n3654,n2524,n2546);
and (n3655,n3652,n2546);
and (n3656,n3646,n3650);
and (n3657,n3624,n3644);
and (n3658,n3607,n3622);
and (n3659,n3583,n3605);
and (n3660,n3661,n3662);
xor (n3661,n3576,n3578);
and (n3662,n3663,n3664);
xnor (n3663,n3579,n3581);
or (n3664,n3665,n3869);
and (n3665,n3666,n3668);
xor (n3666,n3667,n3605);
xor (n3667,n3583,n3602);
or (n3668,n3669,n3744,n3868);
and (n3669,n3670,n3742);
or (n3670,n3671,n3738,n3741);
and (n3671,n3672,n3674);
xor (n3672,n3673,n3616);
xor (n3673,n3609,n3613);
or (n3674,n3675,n3709,n3737);
and (n3675,n3676,n3707);
or (n3676,n3677,n3695,n3706);
and (n3677,n3678,n3687);
and (n3678,n3679,n2433);
or (n3679,n3680,n3685,n3686);
and (n3680,n3681,n2303);
or (n3681,n3682,n3683,n3684);
and (n3682,n2372,n2168);
not (n3683,n2312);
and (n3684,n2372,n2172);
not (n3685,n2445);
and (n3686,n3681,n2307);
or (n3687,n3688,n3693,n3694);
and (n3688,n2473,n3689);
or (n3689,n3690,n3691,n3692);
and (n3690,n2372,n2292);
not (n3691,n2420);
and (n3692,n2372,n2297);
and (n3693,n3689,n2454);
and (n3694,n2473,n2454);
and (n3695,n3687,n3696);
or (n3696,n3697,n3703,n3705);
and (n3697,n3698,n3699);
not (n3698,n2392);
or (n3699,n3700,n3701,n3702);
and (n3700,n2176,n2368);
not (n3701,n2472);
and (n3702,n2176,n2373);
and (n3703,n3699,n3704);
not (n3704,n2449);
and (n3705,n3698,n3704);
and (n3706,n3678,n3696);
xor (n3707,n3708,n3631);
xor (n3708,n3626,n2608);
and (n3709,n3707,n3710);
or (n3710,n3711,n3733,n3736);
and (n3711,n3712,n3714);
xor (n3712,n3713,n3638);
xor (n3713,n1005,n3633);
or (n3714,n3715,n3724,n3732);
and (n3715,n3716,n3723);
or (n3716,n3717,n3719,n3722);
and (n3717,n2352,n3718);
not (n3718,n2349);
and (n3719,n3718,n3720);
xor (n3720,n3721,n2297);
xor (n3721,n2372,n2292);
and (n3722,n2352,n3720);
xor (n3723,n3679,n2433);
and (n3724,n3723,n3725);
or (n3725,n3726,n3730,n3731);
and (n3726,n3727,n3728);
not (n3727,n2366);
xor (n3728,n3729,n2307);
xor (n3729,n3681,n2303);
and (n3730,n3728,n2326);
and (n3731,n3727,n2326);
and (n3732,n3716,n3725);
and (n3733,n3714,n3734);
xor (n3734,n3735,n2546);
xor (n3735,n3652,n2524);
and (n3736,n3712,n3734);
and (n3737,n3676,n3710);
and (n3738,n3674,n3739);
xor (n3739,n3740,n3644);
xor (n3740,n3624,n3641);
and (n3741,n3672,n3739);
xor (n3742,n3743,n3622);
xor (n3743,n3607,n3619);
and (n3744,n3742,n3745);
or (n3745,n3746,n3779,n3867);
and (n3746,n3747,n3777);
or (n3747,n3748,n3773,n3776);
and (n3748,n3749,n3751);
xor (n3749,n3750,n3650);
xor (n3750,n3646,n3648);
or (n3751,n3752,n3769,n3772);
and (n3752,n3753,n3755);
xor (n3753,n3754,n3696);
xor (n3754,n3678,n3687);
or (n3755,n3756,n3761,n3768);
and (n3756,n3757,n3759);
xor (n3757,n3758,n2454);
xor (n3758,n2473,n3689);
xor (n3759,n3760,n3704);
xor (n3760,n3698,n3699);
and (n3761,n3759,n3762);
and (n3762,n2317,n3763);
or (n3763,n3764,n3765,n3767);
not (n3764,n2323);
and (n3765,n2183,n3766);
not (n3766,n2166);
and (n3767,n2179,n3766);
and (n3768,n3757,n3762);
and (n3769,n3755,n3770);
xor (n3770,n3771,n3734);
xor (n3771,n3712,n3714);
and (n3772,n3753,n3770);
and (n3773,n3751,n3774);
xor (n3774,n3775,n3710);
xor (n3775,n3676,n3707);
and (n3776,n3749,n3774);
xor (n3777,n3778,n3739);
xor (n3778,n3672,n3674);
and (n3779,n3777,n3780);
or (n3780,n3781,n3838,n3866);
and (n3781,n3782,n3784);
xor (n3782,n3783,n3774);
xor (n3783,n3749,n3751);
or (n3784,n3785,n3817,n3837);
and (n3785,n3786,n3815);
or (n3786,n3787,n3800,n3814);
and (n3787,n3788,n3798);
or (n3788,n3789,n3796,n3797);
and (n3789,n3790,n3794);
or (n3790,n3791,n3792,n3793);
and (n3791,n2231,n2216);
and (n3792,n2216,n2199);
and (n3793,n2231,n2199);
xor (n3794,n3795,n3720);
xor (n3795,n2352,n3718);
and (n3796,n3794,n2377);
and (n3797,n3790,n2377);
xor (n3798,n3799,n3725);
xor (n3799,n3716,n3723);
and (n3800,n3798,n3801);
or (n3801,n3802,n3811,n3813);
and (n3802,n3803,n3809);
or (n3803,n3804,n3805,n3808);
and (n3804,n2221,n2215);
and (n3805,n2215,n3806);
xor (n3806,n3807,n2199);
xor (n3807,n2231,n2216);
and (n3808,n2221,n3806);
xor (n3809,n3810,n2326);
xor (n3810,n3727,n3728);
and (n3811,n3809,n3812);
xor (n3812,n2317,n3763);
and (n3813,n3803,n3812);
and (n3814,n3788,n3801);
xor (n3815,n3816,n3770);
xor (n3816,n3753,n3755);
and (n3817,n3815,n3818);
or (n3818,n3819,n3833,n3836);
and (n3819,n3820,n3822);
xor (n3820,n3821,n3762);
xor (n3821,n3757,n3759);
or (n3822,n3823,n3831,n3832);
and (n3823,n3824,n3826);
xor (n3824,n3825,n2377);
xor (n3825,n3790,n3794);
or (n3826,n3827,n3828,n3830);
not (n3827,n2276);
and (n3828,n2191,n3829);
not (n3829,n2164);
and (n3830,n2187,n3829);
and (n3831,n3826,n2278);
and (n3832,n3824,n2278);
and (n3833,n3822,n3834);
xor (n3834,n3835,n3801);
xor (n3835,n3788,n3798);
and (n3836,n3820,n3834);
and (n3837,n3786,n3818);
and (n3838,n3784,n3839);
or (n3839,n3840,n3842);
xor (n3840,n3841,n3818);
xor (n3841,n3786,n3815);
or (n3842,n3843,n3859,n3865);
and (n3843,n3844,n3857);
or (n3844,n3845,n3853,n3856);
and (n3845,n3846,n3848);
xor (n3846,n3847,n3812);
xor (n3847,n3803,n3809);
or (n3848,n3849,n3851,n3852);
and (n3849,n3850,n2263);
not (n3850,n2162);
not (n3851,n2270);
and (n3852,n3850,n2195);
and (n3853,n3848,n3854);
xor (n3854,n3855,n2278);
xor (n3855,n3824,n3826);
and (n3856,n3846,n3854);
xor (n3857,n3858,n3834);
xor (n3858,n3820,n3822);
and (n3859,n3857,n3860);
or (n3860,n3861,n3863);
or (n3861,n2156,n3862);
not (n3862,n2160);
xor (n3863,n3864,n3854);
xor (n3864,n3846,n3848);
and (n3865,n3844,n3860);
and (n3866,n3782,n3839);
and (n3867,n3747,n3780);
and (n3868,n3670,n3745);
and (n3869,n3870,n3871);
xor (n3870,n3666,n3668);
and (n3871,n3872,n3874);
xor (n3872,n3873,n3745);
xor (n3873,n3670,n3742);
or (n3874,n3875,n3877);
xor (n3875,n3876,n3780);
xor (n3876,n3747,n3777);
and (n3877,n3878,n3879);
not (n3878,n3875);
and (n3879,n3880,n3882);
xor (n3880,n3881,n3839);
xor (n3881,n3782,n3784);
and (n3882,n3883,n3884);
xnor (n3883,n3840,n3842);
and (n3884,n3885,n3887);
xor (n3885,n3886,n3860);
xor (n3886,n3844,n3857);
and (n3887,n3888,n3889);
xnor (n3888,n3861,n3863);
and (n3889,n3890,n3893);
not (n3890,n3891);
nand (n3891,n3892,n2685);
not (n3892,n2155);
nand (n3893,n1182,n3894);
nand (n3894,n3132,n2711);
endmodule
