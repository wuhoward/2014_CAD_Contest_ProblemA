module top (out,n3,n4,n5,n19,n20,n28,n29,n38,n46
        ,n48,n54,n61,n72,n73,n77,n83,n94,n96,n104
        ,n113,n122,n135,n155,n210,n235);
output out;
input n3;
input n4;
input n5;
input n19;
input n20;
input n28;
input n29;
input n38;
input n46;
input n48;
input n54;
input n61;
input n72;
input n73;
input n77;
input n83;
input n94;
input n96;
input n104;
input n113;
input n122;
input n135;
input n155;
input n210;
input n235;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
xnor (out,n0,n461);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n458);
xor (n7,n8,n251);
xor (n8,n9,n194);
or (n9,n10,n193);
and (n10,n11,n158);
xor (n11,n12,n86);
xor (n12,n13,n68);
xor (n13,n14,n41);
nand (n14,n15,n34);
or (n15,n16,n23);
nor (n16,n17,n21);
and (n17,n18,n20);
not (n18,n19);
and (n21,n19,n22);
not (n22,n20);
nand (n23,n24,n31);
not (n24,n25);
nand (n25,n26,n30);
or (n26,n27,n29);
not (n27,n28);
nand (n30,n29,n27);
nand (n31,n32,n33);
or (n32,n29,n18);
nand (n33,n18,n29);
nand (n34,n35,n25);
not (n35,n36);
nor (n36,n37,n39);
and (n37,n18,n38);
and (n39,n19,n40);
not (n40,n38);
nand (n41,n42,n56);
or (n42,n43,n51);
not (n43,n44);
nand (n44,n45,n49);
or (n45,n46,n47);
not (n47,n48);
or (n49,n50,n48);
not (n50,n46);
not (n51,n52);
nand (n52,n53,n55);
or (n53,n18,n54);
nand (n55,n54,n18);
nand (n56,n57,n63);
not (n57,n58);
nor (n58,n59,n62);
and (n59,n60,n46);
not (n60,n61);
and (n62,n50,n61);
nor (n63,n52,n64);
nor (n64,n65,n66);
and (n65,n50,n54);
and (n66,n46,n67);
not (n67,n54);
nand (n68,n69,n80);
or (n69,n70,n74);
nand (n70,n71,n73);
not (n71,n72);
nor (n74,n75,n78);
and (n75,n76,n77);
not (n76,n73);
and (n78,n73,n79);
not (n79,n77);
or (n80,n81,n71);
nor (n81,n82,n84);
and (n82,n76,n83);
and (n84,n73,n85);
not (n85,n83);
or (n86,n87,n157);
and (n87,n88,n138);
xor (n88,n89,n116);
nand (n89,n90,n109);
or (n90,n91,n99);
not (n91,n92);
nand (n92,n93,n97);
or (n93,n94,n95);
not (n95,n96);
or (n97,n98,n96);
not (n98,n94);
nand (n99,n100,n106);
not (n100,n101);
nand (n101,n102,n105);
or (n102,n103,n73);
not (n103,n104);
nand (n105,n73,n103);
nand (n106,n107,n108);
or (n107,n103,n94);
nand (n108,n103,n94);
nand (n109,n110,n101);
not (n110,n111);
nor (n111,n112,n114);
and (n112,n98,n113);
and (n114,n94,n115);
not (n115,n113);
nand (n116,n117,n131);
or (n117,n118,n128);
not (n118,n119);
nor (n119,n120,n124);
nand (n120,n121,n123);
or (n121,n98,n122);
nand (n123,n122,n98);
nor (n124,n125,n127);
and (n125,n126,n28);
not (n126,n122);
and (n127,n122,n27);
nor (n128,n129,n130);
and (n129,n27,n38);
and (n130,n28,n40);
or (n131,n132,n133);
not (n132,n120);
nor (n133,n134,n136);
and (n134,n27,n135);
and (n136,n28,n137);
not (n137,n135);
and (n138,n139,n145);
nor (n139,n140,n18);
nor (n140,n141,n143);
and (n141,n60,n142);
not (n142,n29);
nor (n143,n144,n28);
and (n144,n61,n29);
nand (n145,n146,n151);
or (n146,n70,n147);
not (n147,n148);
nor (n148,n149,n150);
and (n149,n115,n76);
and (n150,n113,n73);
or (n151,n152,n71);
nor (n152,n153,n156);
and (n153,n154,n73);
not (n154,n155);
and (n156,n155,n76);
and (n157,n89,n116);
xor (n158,n159,n179);
xor (n159,n160,n166);
nand (n160,n161,n162);
or (n161,n118,n133);
or (n162,n132,n163);
nor (n163,n164,n165);
and (n164,n27,n96);
and (n165,n28,n95);
xor (n166,n167,n173);
and (n167,n168,n46);
nand (n168,n169,n170);
or (n169,n61,n54);
nand (n170,n171,n18);
not (n171,n172);
and (n172,n61,n54);
nand (n173,n174,n175);
or (n174,n99,n111);
or (n175,n100,n176);
nor (n176,n177,n178);
and (n177,n98,n155);
and (n178,n94,n154);
or (n179,n180,n192);
and (n180,n181,n186);
xor (n181,n182,n183);
nor (n182,n51,n60);
nand (n183,n184,n185);
or (n184,n152,n70);
or (n185,n74,n71);
nand (n186,n187,n191);
or (n187,n23,n188);
nor (n188,n189,n190);
and (n189,n18,n48);
and (n190,n19,n47);
or (n191,n24,n16);
and (n192,n182,n183);
and (n193,n12,n86);
xor (n194,n195,n222);
xor (n195,n196,n219);
xor (n196,n197,n213);
xor (n197,n198,n205);
nand (n198,n199,n201);
or (n199,n43,n200);
not (n200,n63);
nand (n201,n52,n202);
nand (n202,n203,n204);
or (n203,n46,n22);
or (n204,n50,n20);
nand (n205,n206,n207);
or (n206,n81,n70);
or (n207,n208,n71);
nor (n208,n209,n211);
and (n209,n76,n210);
and (n211,n73,n212);
not (n212,n210);
nand (n213,n214,n215);
or (n214,n118,n163);
or (n215,n132,n216);
nor (n216,n217,n218);
and (n217,n27,n113);
and (n218,n28,n115);
or (n219,n220,n221);
and (n220,n159,n179);
and (n221,n160,n166);
xor (n222,n223,n228);
xor (n223,n224,n225);
and (n224,n167,n173);
or (n225,n226,n227);
and (n226,n13,n68);
and (n227,n14,n41);
xor (n228,n229,n244);
xor (n229,n230,n237);
nor (n230,n231,n60);
not (n231,n232);
nand (n232,n233,n236);
or (n233,n234,n46);
not (n234,n235);
nand (n236,n46,n234);
nand (n237,n238,n239);
or (n238,n176,n99);
nand (n239,n240,n101);
not (n240,n241);
nor (n241,n242,n243);
and (n242,n77,n98);
and (n243,n79,n94);
nand (n244,n245,n250);
or (n245,n246,n24);
not (n246,n247);
nand (n247,n248,n249);
or (n248,n19,n137);
or (n249,n18,n135);
or (n250,n23,n36);
nand (n251,n252,n455,n457);
nand (n252,n253,n288,n448);
nand (n253,n254,n256);
not (n254,n255);
xor (n255,n11,n158);
not (n256,n257);
or (n257,n258,n287);
and (n258,n259,n286);
xor (n259,n260,n285);
or (n260,n261,n284);
and (n261,n262,n278);
xor (n262,n263,n271);
nand (n263,n264,n269);
or (n264,n265,n23);
not (n265,n266);
nand (n266,n267,n268);
or (n267,n18,n61);
or (n268,n60,n19);
nand (n269,n270,n25);
not (n270,n188);
nand (n271,n272,n277);
or (n272,n273,n99);
not (n273,n274);
nand (n274,n275,n276);
or (n275,n94,n137);
or (n276,n98,n135);
nand (n277,n101,n92);
nand (n278,n279,n283);
or (n279,n118,n280);
nor (n280,n281,n282);
and (n281,n27,n20);
and (n282,n28,n22);
or (n283,n132,n128);
and (n284,n263,n271);
xor (n285,n181,n186);
xor (n286,n88,n138);
and (n287,n260,n285);
nand (n288,n289,n447);
or (n289,n290,n340);
not (n290,n291);
nand (n291,n292,n316);
not (n292,n293);
xor (n293,n294,n315);
xor (n294,n295,n296);
xor (n295,n139,n145);
or (n296,n297,n314);
and (n297,n298,n307);
xor (n298,n299,n300);
and (n299,n25,n61);
nand (n300,n301,n306);
or (n301,n70,n302);
not (n302,n303);
nor (n303,n304,n305);
and (n304,n95,n76);
and (n305,n96,n73);
nand (n306,n148,n72);
nand (n307,n308,n313);
or (n308,n309,n99);
not (n309,n310);
nor (n310,n311,n312);
and (n311,n40,n98);
and (n312,n38,n94);
nand (n313,n101,n274);
and (n314,n299,n300);
xor (n315,n262,n278);
not (n316,n317);
or (n317,n318,n339);
and (n318,n319,n338);
xor (n319,n320,n326);
nand (n320,n321,n325);
or (n321,n118,n322);
nor (n322,n323,n324);
and (n323,n47,n28);
and (n324,n48,n27);
or (n325,n132,n280);
and (n326,n327,n332);
and (n327,n328,n28);
nand (n328,n329,n331);
or (n329,n330,n94);
and (n330,n61,n122);
or (n331,n61,n122);
nand (n332,n333,n334);
or (n333,n71,n302);
or (n334,n335,n70);
nor (n335,n336,n337);
and (n336,n76,n135);
and (n337,n73,n137);
xor (n338,n298,n307);
and (n339,n320,n326);
not (n340,n341);
nand (n341,n342,n446);
or (n342,n343,n366);
not (n343,n344);
nand (n344,n345,n347);
not (n345,n346);
xor (n346,n319,n338);
not (n347,n348);
or (n348,n349,n365);
and (n349,n350,n364);
xor (n350,n351,n358);
nand (n351,n352,n357);
or (n352,n353,n99);
not (n353,n354);
nor (n354,n355,n356);
and (n355,n22,n98);
and (n356,n20,n94);
nand (n357,n310,n101);
nand (n358,n359,n360);
or (n359,n132,n322);
nand (n360,n119,n361);
nand (n361,n362,n363);
or (n362,n61,n27);
or (n363,n60,n28);
xor (n364,n327,n332);
and (n365,n351,n358);
not (n366,n367);
or (n367,n368,n445);
and (n368,n369,n390);
xor (n369,n370,n389);
or (n370,n371,n388);
and (n371,n372,n381);
xor (n372,n373,n374);
and (n373,n120,n61);
nand (n374,n375,n380);
or (n375,n376,n99);
not (n376,n377);
nor (n377,n378,n379);
and (n378,n47,n98);
and (n379,n48,n94);
nand (n380,n354,n101);
nand (n381,n382,n387);
or (n382,n70,n383);
not (n383,n384);
nor (n384,n385,n386);
and (n385,n40,n76);
and (n386,n38,n73);
or (n387,n335,n71);
and (n388,n373,n374);
xor (n389,n350,n364);
nand (n390,n391,n444);
or (n391,n392,n408);
nor (n392,n393,n394);
xor (n393,n372,n381);
nor (n394,n395,n403);
not (n395,n396);
nand (n396,n397,n398);
or (n397,n71,n383);
nand (n398,n399,n402);
nand (n399,n400,n401);
or (n400,n20,n76);
nand (n401,n76,n20);
not (n402,n70);
nand (n403,n404,n94);
nand (n404,n405,n407);
or (n405,n406,n73);
and (n406,n61,n104);
or (n407,n61,n104);
nor (n408,n409,n443);
and (n409,n410,n422);
nand (n410,n411,n418);
not (n411,n412);
nand (n412,n413,n417);
or (n413,n99,n414);
nor (n414,n415,n416);
and (n415,n94,n60);
and (n416,n61,n98);
or (n417,n100,n376);
nor (n418,n419,n420);
and (n419,n403,n396);
and (n420,n421,n395);
not (n421,n403);
or (n422,n423,n442);
and (n423,n424,n433);
xor (n424,n425,n426);
nor (n425,n100,n60);
nand (n426,n427,n432);
or (n427,n70,n428);
not (n428,n429);
nand (n429,n430,n431);
or (n430,n47,n73);
nand (n431,n73,n47);
nand (n432,n399,n72);
nor (n433,n434,n440);
nor (n434,n435,n436);
and (n435,n429,n72);
nor (n436,n437,n70);
nor (n437,n438,n439);
and (n438,n60,n73);
and (n439,n61,n76);
or (n440,n441,n76);
and (n441,n61,n72);
and (n442,n425,n426);
nor (n443,n411,n418);
nand (n444,n393,n394);
and (n445,n370,n389);
nand (n446,n346,n348);
nand (n447,n293,n317);
nand (n448,n449,n453);
not (n449,n450);
or (n450,n451,n452);
and (n451,n294,n315);
and (n452,n295,n296);
not (n453,n454);
xor (n454,n259,n286);
nand (n455,n253,n456);
and (n456,n454,n450);
nand (n457,n257,n255);
not (n458,n459);
nand (n459,n460,n3);
not (n460,n4);
wire s0n461,s1n461,notn461;
or (n461,s0n461,s1n461);
not(notn461,n4);
and (s0n461,notn461,n462);
and (s1n461,n4,1'b0);
wire s0n462,s1n462,notn462;
or (n462,s0n462,s1n462);
not(notn462,n3);
and (s0n462,notn462,n5);
and (s1n462,n3,n463);
xor (n463,n464,n725);
xor (n464,n465,n722);
xor (n465,n466,n721);
xor (n466,n467,n713);
xor (n467,n468,n712);
xor (n468,n469,n697);
xor (n469,n470,n696);
xor (n470,n471,n676);
xor (n471,n472,n675);
xor (n472,n473,n648);
xor (n473,n474,n647);
xor (n474,n475,n615);
xor (n475,n476,n614);
xor (n476,n477,n578);
xor (n477,n478,n577);
xor (n478,n479,n533);
xor (n479,n480,n532);
xor (n480,n481,n484);
xor (n481,n482,n483);
and (n482,n210,n72);
and (n483,n83,n73);
or (n484,n485,n488);
and (n485,n486,n487);
and (n486,n83,n72);
and (n487,n77,n73);
and (n488,n489,n490);
xor (n489,n486,n487);
or (n490,n491,n494);
and (n491,n492,n493);
and (n492,n77,n72);
and (n493,n155,n73);
and (n494,n495,n496);
xor (n495,n492,n493);
or (n496,n497,n499);
and (n497,n498,n150);
and (n498,n155,n72);
and (n499,n500,n501);
xor (n500,n498,n150);
or (n501,n502,n504);
and (n502,n503,n305);
and (n503,n113,n72);
and (n504,n505,n506);
xor (n505,n503,n305);
or (n506,n507,n510);
and (n507,n508,n509);
and (n508,n96,n72);
and (n509,n135,n73);
and (n510,n511,n512);
xor (n511,n508,n509);
or (n512,n513,n515);
and (n513,n514,n386);
and (n514,n135,n72);
and (n515,n516,n517);
xor (n516,n514,n386);
or (n517,n518,n521);
and (n518,n519,n520);
and (n519,n38,n72);
and (n520,n20,n73);
and (n521,n522,n523);
xor (n522,n519,n520);
or (n523,n524,n527);
and (n524,n525,n526);
and (n525,n20,n72);
and (n526,n48,n73);
and (n527,n528,n529);
xor (n528,n525,n526);
and (n529,n530,n531);
and (n530,n48,n72);
and (n531,n61,n73);
and (n532,n77,n104);
or (n533,n534,n537);
and (n534,n535,n536);
xor (n535,n489,n490);
and (n536,n155,n104);
and (n537,n538,n539);
xor (n538,n535,n536);
or (n539,n540,n543);
and (n540,n541,n542);
xor (n541,n495,n496);
and (n542,n113,n104);
and (n543,n544,n545);
xor (n544,n541,n542);
or (n545,n546,n549);
and (n546,n547,n548);
xor (n547,n500,n501);
and (n548,n96,n104);
and (n549,n550,n551);
xor (n550,n547,n548);
or (n551,n552,n555);
and (n552,n553,n554);
xor (n553,n505,n506);
and (n554,n135,n104);
and (n555,n556,n557);
xor (n556,n553,n554);
or (n557,n558,n561);
and (n558,n559,n560);
xor (n559,n511,n512);
and (n560,n38,n104);
and (n561,n562,n563);
xor (n562,n559,n560);
or (n563,n564,n567);
and (n564,n565,n566);
xor (n565,n516,n517);
and (n566,n20,n104);
and (n567,n568,n569);
xor (n568,n565,n566);
or (n569,n570,n573);
and (n570,n571,n572);
xor (n571,n522,n523);
and (n572,n48,n104);
and (n573,n574,n575);
xor (n574,n571,n572);
and (n575,n576,n406);
xor (n576,n528,n529);
and (n577,n155,n94);
or (n578,n579,n582);
and (n579,n580,n581);
xor (n580,n538,n539);
and (n581,n113,n94);
and (n582,n583,n584);
xor (n583,n580,n581);
or (n584,n585,n588);
and (n585,n586,n587);
xor (n586,n544,n545);
and (n587,n96,n94);
and (n588,n589,n590);
xor (n589,n586,n587);
or (n590,n591,n594);
and (n591,n592,n593);
xor (n592,n550,n551);
and (n593,n135,n94);
and (n594,n595,n596);
xor (n595,n592,n593);
or (n596,n597,n599);
and (n597,n598,n312);
xor (n598,n556,n557);
and (n599,n600,n601);
xor (n600,n598,n312);
or (n601,n602,n604);
and (n602,n603,n356);
xor (n603,n562,n563);
and (n604,n605,n606);
xor (n605,n603,n356);
or (n606,n607,n609);
and (n607,n608,n379);
xor (n608,n568,n569);
and (n609,n610,n611);
xor (n610,n608,n379);
and (n611,n612,n613);
xor (n612,n574,n575);
and (n613,n61,n94);
and (n614,n113,n122);
or (n615,n616,n619);
and (n616,n617,n618);
xor (n617,n583,n584);
and (n618,n96,n122);
and (n619,n620,n621);
xor (n620,n617,n618);
or (n621,n622,n625);
and (n622,n623,n624);
xor (n623,n589,n590);
and (n624,n135,n122);
and (n625,n626,n627);
xor (n626,n623,n624);
or (n627,n628,n631);
and (n628,n629,n630);
xor (n629,n595,n596);
and (n630,n38,n122);
and (n631,n632,n633);
xor (n632,n629,n630);
or (n633,n634,n637);
and (n634,n635,n636);
xor (n635,n600,n601);
and (n636,n20,n122);
and (n637,n638,n639);
xor (n638,n635,n636);
or (n639,n640,n643);
and (n640,n641,n642);
xor (n641,n605,n606);
and (n642,n48,n122);
and (n643,n644,n645);
xor (n644,n641,n642);
and (n645,n646,n330);
xor (n646,n610,n611);
and (n647,n96,n28);
or (n648,n649,n652);
and (n649,n650,n651);
xor (n650,n620,n621);
and (n651,n135,n28);
and (n652,n653,n654);
xor (n653,n650,n651);
or (n654,n655,n658);
and (n655,n656,n657);
xor (n656,n626,n627);
and (n657,n38,n28);
and (n658,n659,n660);
xor (n659,n656,n657);
or (n660,n661,n664);
and (n661,n662,n663);
xor (n662,n632,n633);
and (n663,n20,n28);
and (n664,n665,n666);
xor (n665,n662,n663);
or (n666,n667,n670);
and (n667,n668,n669);
xor (n668,n638,n639);
and (n669,n48,n28);
and (n670,n671,n672);
xor (n671,n668,n669);
and (n672,n673,n674);
xor (n673,n644,n645);
and (n674,n61,n28);
and (n675,n135,n29);
or (n676,n677,n680);
and (n677,n678,n679);
xor (n678,n653,n654);
and (n679,n38,n29);
and (n680,n681,n682);
xor (n681,n678,n679);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n659,n660);
and (n685,n20,n29);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n665,n666);
and (n691,n48,n29);
and (n692,n693,n694);
xor (n693,n690,n691);
and (n694,n695,n144);
xor (n695,n671,n672);
and (n696,n38,n19);
or (n697,n698,n701);
and (n698,n699,n700);
xor (n699,n681,n682);
and (n700,n20,n19);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n687,n688);
and (n706,n48,n19);
and (n707,n708,n709);
xor (n708,n705,n706);
and (n709,n710,n711);
xor (n710,n693,n694);
and (n711,n61,n19);
and (n712,n20,n54);
or (n713,n714,n717);
and (n714,n715,n716);
xor (n715,n702,n703);
and (n716,n48,n54);
and (n717,n718,n719);
xor (n718,n715,n716);
and (n719,n720,n172);
xor (n720,n708,n709);
and (n721,n48,n46);
and (n722,n723,n724);
xor (n723,n718,n719);
and (n724,n61,n46);
and (n725,n61,n235);
endmodule
