module top (out,n27,n40,n43,n45,n46,n48,n52,n61,n63
        ,n64,n66,n71,n74,n76,n81,n85,n93,n97,n98
        ,n99,n111,n115,n116,n117,n132,n133,n134,n135,n136
        ,n140,n141,n142,n147,n149,n151,n188,n190,n191,n192
        ,n203,n204,n205,n206,n218,n219,n220,n221,n235,n241
        ,n243,n244,n248,n249,n252,n254,n255,n256,n329,n384
        ,n387,n389,n477,n479,n480,n594,n597,n599,n601,n605
        ,n608,n610,n612,n616,n619,n621,n623,n625,n684,n687
        ,n689,n691,n695,n698,n700,n702,n706,n709,n711,n713
        ,n717,n720,n722,n724,n758,n761,n763,n765,n769,n772
        ,n774,n776,n780,n783,n785,n787,n791,n794,n796,n798
        ,n831,n834,n836,n838,n842,n845,n847,n849,n853,n856
        ,n858,n860,n864,n867,n869,n871,n901,n902,n904,n905
        ,n920,n924,n926,n931,n933,n975,n987,n992,n997,n1002
        ,n1010,n1013,n1022,n1026,n1032,n1034,n1036,n1038,n1040,n1048
        ,n1051,n1053,n1055,n1057,n1064,n1065,n1075,n1078,n1082,n1087
        ,n1090,n1093,n1096,n1101,n1103,n1105,n1107,n1109,n1114,n1116
        ,n1123,n1126,n1128,n1138,n1140,n1142,n1144,n1146,n1151,n1153
        ,n1156,n1158,n1160,n1164,n1166,n1169,n1172,n1176,n1178,n1181
        ,n1183,n1184,n1192,n1197,n1201,n1205,n1209,n1214,n1216,n1219
        ,n1221,n1223,n1227,n1229,n1232,n1235,n1239,n1243,n1248,n1252
        ,n1253,n1263,n1265,n1267,n1269,n1271,n1277,n1279,n1281,n1283
        ,n1288,n1289,n1292,n1295,n1298,n1303,n1306,n1309,n1312,n1313
        ,n1320,n1321,n1324,n1327,n1330,n1335,n1338,n1341,n1344,n1349
        ,n1351,n1354,n1358,n1360,n1365,n1367,n1373,n1376,n1377,n1387
        ,n1389,n1391,n1393,n1395,n1398,n1400,n1406,n1408,n1410,n1412
        ,n1414,n1419,n1422,n1424,n1426,n1429,n1431,n1432,n1439,n1440
        ,n1443,n1446,n1449,n1454,n1457,n1460,n1463,n1468,n1470,n1472
        ,n1474,n1476,n1481,n1483,n1489,n1491,n1492,n1502,n1504,n1506
        ,n1508,n1510,n1516,n1518,n1520,n1522,n1527,n1528,n1531,n1534
        ,n1537,n1542,n1545,n1548,n1551,n1552,n1559,n1560,n1563,n1566
        ,n1569,n1574,n1577,n1580,n1583,n1588,n1590,n1593,n1597,n1599
        ,n1604,n1606,n1612,n1615,n1616,n1626,n1628,n1630,n1632,n1634
        ,n1640,n1642,n1644,n1646,n1651,n1652,n1655,n1658,n1661,n1666
        ,n1669,n1672,n1675,n1676,n1683,n1684,n1687,n1690,n1693,n1698
        ,n1701,n1704,n1707,n1712,n1714,n1717,n1721,n1723,n1728,n1730
        ,n1733,n1738,n1739,n1748,n1750,n1753,n1755,n1757,n1761,n1763
        ,n1767,n1769,n1774,n1775,n1778,n1781,n1784,n1789,n1792,n1795
        ,n1798,n1799,n1806,n1807,n1810,n1813,n1816,n1821,n1824,n1827
        ,n1830,n1836,n1838,n1840,n1842,n1844,n1853,n1855,n1857,n1859
        ,n1860,n1869,n1871,n1873,n1875,n1877,n1882,n1885,n1887,n1889
        ,n1894,n1895,n1898,n1901,n1904,n1909,n1912,n1915,n1918,n1919
        ,n1926,n1927,n1930,n1933,n1936,n1941,n1944,n1947,n1950,n1955
        ,n1957,n1960,n1964,n1966,n1971,n1973,n1976,n1981,n1982,n1998
        ,n2000,n2010,n2012,n2014,n2016,n2018,n2023,n2026,n2028,n2030
        ,n2033,n2036,n2038,n2040,n2042,n2045,n2047,n2050,n2052,n2053
        ,n2060,n2062,n2064,n2066,n2068,n2074,n2076,n2078,n2080,n2082
        ,n2087,n2090,n2092,n2094,n2097,n2099,n2102,n2104,n2105,n2116
        ,n2118,n2120,n2122,n2124,n2129,n2132,n2134,n2136,n2139,n2143
        ,n2145,n2147,n2149,n2152,n2154,n2157,n2159,n2160,n2167,n2169
        ,n2174,n2176,n2179,n2184,n2186,n2192,n2195,n2200,n2201,n2204
        ,n2207,n2210,n2215,n2218,n2221,n2224,n2225,n2233,n2237,n2240
        ,n2242,n2244,n2249,n2251,n2254,n2256,n2258,n2262,n2264,n2267
        ,n2270,n2273,n2275,n2278,n2280,n2281,n2286,n2289,n2292,n2294
        ,n2296,n2302,n2304,n2306,n2308,n2310,n2312,n2319,n2321,n2323
        ,n2325,n2327,n2330,n2332,n2333,n2343,n2345,n2350,n2352,n2355
        ,n2360,n2362,n2368,n2371,n2376,n2377,n2380,n2383,n2386,n2391
        ,n2394,n2397,n2400,n2401,n2408,n2410,n2412,n2414,n2416,n2421
        ,n2423,n2429,n2431,n2436,n2437,n2440,n2443,n2446,n2451,n2454
        ,n2457,n2460,n2461,n2471,n2473,n2478,n2480,n2483,n2488,n2490
        ,n2496,n2499,n2504,n2505,n2508,n2511,n2514,n2519,n2522,n2525
        ,n2528,n2529,n2535,n2537,n2540,n2542,n2544,n2548,n2550,n2554
        ,n2556,n2561,n2562,n2565,n2568,n2571,n2576,n2579,n2582,n2585
        ,n2586,n2596,n2598,n2600,n2602,n2604,n2610,n2612,n2614,n2616
        ,n2621,n2622,n2625,n2628,n2631,n2636,n2639,n2642,n2645,n2646
        ,n2653,n2655,n2657,n2659,n2661,n2666,n2669,n2671,n2673,n2678
        ,n2679,n2682,n2685,n2688,n2693,n2696,n2699,n2702,n2703,n2713
        ,n2714,n2717,n2720,n2723,n2728,n2730,n2734,n2736,n2741,n2742
        ,n2745,n2748,n2751,n2756,n2759,n2762,n2765,n2766,n2776,n2778
        ,n2780,n2782,n2784,n2791,n2793,n2795,n2797,n2802,n2803,n2806
        ,n2809,n2812,n2817,n2820,n2823,n2826,n2827,n2837,n2839,n2842
        ,n2844,n2846,n2851,n2853,n2857,n2859,n2864,n2865,n2868,n2871
        ,n2874,n2879,n2882,n2885,n2888,n2889,n2896,n2898,n2901,n2905
        ,n2907,n2912,n2914,n2917,n2922,n2927,n2928,n2931,n2934,n2937
        ,n2942,n2945,n2948,n2951,n2952,n2966,n2968,n2988,n2989,n2992
        ,n2995,n2998,n3003,n3006,n3009,n3012,n3013,n3016,n3021,n3023
        ,n3026,n3028,n3030,n3036,n3038,n3042,n3044,n3056,n3057,n3060
        ,n3063,n3066,n3071,n3074,n3077,n3080,n3081,n3091,n3093,n3095
        ,n3097,n3099,n3105,n3107,n3109,n3111,n3112,n3122,n3124,n3127
        ,n3129,n3146,n3147,n3150,n3153,n3156,n3161,n3164,n3167,n3170
        ,n3171,n3175,n3182,n3184,n3186,n3188,n3190,n3196,n3199,n3201
        ,n3203,n3213,n3214,n3217,n3220,n3223,n3228,n3231,n3234,n3237
        ,n3238,n3245,n3247,n3250,n3252,n3254,n3260,n3262,n3266,n3268
        ,n3270,n3282,n3283,n3286,n3289,n3292,n3297,n3300,n3303,n3306
        ,n3307,n3314,n3316,n3321,n3323,n3326,n3333,n3336,n3338,n3340
        ,n3341,n3355,n3356,n3359,n3362,n3365,n3370,n3373,n3376,n3379
        ,n3380,n3383,n3389,n3391,n3393,n3395,n3397,n3405,n3407,n3409
        ,n3411,n3428,n3429,n3432,n3435,n3438,n3443,n3446,n3449,n3452
        ,n3453,n3461,n3463,n3465,n3467,n3469,n3477,n3479,n3481,n3483
        ,n3484,n3495,n3496,n3499,n3502,n3505,n3510,n3513,n3516,n3519
        ,n3520,n3525,n3534,n3536,n3538,n3540,n3542,n3549,n3551,n3553
        ,n3555,n3851,n3853,n3857,n3859,n3864,n3866,n3884,n3886,n3892
        ,n3894,n3909,n3911,n3977,n3979,n3991,n3993,n4011,n4013,n4032
        ,n4038,n4054,n4061,n4080,n4087,n4093,n4095,n4520,n4522,n5454
        ,n5455,n5458,n5459,n5466,n5467,n5470,n5471,n5505,n5506,n5511
        ,n5512,n5549,n5550,n5553,n5554,n5582,n5583,n5587,n5588,n5619
        ,n5620,n5623,n5624,n5661,n5662,n5666,n5667,n5709,n5710,n5713
        ,n5714,n5745,n5746,n5749,n5750,n5788,n5789,n5792,n5793,n5824
        ,n5825,n5828,n5829,n5866,n5867,n5870,n5871,n5891,n5892,n5897
        ,n5898,n5927,n5928,n5931,n5932,n5963,n5964,n5969,n5970,n5999
        ,n6000,n6003,n6004,n6163,n6166,n6182,n6186,n6196,n6207,n6211
        ,n6215,n6227,n6237,n6240,n6242,n6246,n6248,n6262,n6264,n6276
        ,n6286,n6289,n6291,n6295,n6297,n6311,n6313,n6327,n6335,n6338
        ,n6340,n6356,n6358,n6361,n6363,n6378,n6389,n6392,n6394,n6400
        ,n6415,n6417,n6419,n6431,n6441,n6444,n6446,n6462,n6464,n6467
        ,n6469,n6484,n6494,n6497,n6499,n6505,n6520,n6522,n6524,n6541
        ,n6543,n6545,n6555,n6576,n6578,n6581,n6583,n6761,n6764,n6877
        ,n6880,n6971,n6974,n7099,n7102,n7357,n7360,n7376,n7379,n7510
        ,n7513,n7619,n7622,n7733,n7743,n7746,n7748,n7750,n7754,n7757
        ,n7759,n7761,n7765,n7768,n7770,n7772,n7776,n7779,n7781,n7783
        ,n7791,n7794,n7796,n7798,n7802,n7805,n7807,n7809,n7813,n7816
        ,n7818,n7820,n7824,n7827,n7829,n7831,n7875,n7902,n7917,n7932
        ,n7947,n7962,n7981,n8059,n8070,n8090,n8105,n8120,n8140,n8155
        ,n8164,n8259,n8272,n8278,n8296,n8316,n8326,n8340,n8392,n8399
        ,n8418,n8449,n8510,n8524,n8534,n8554,n8568);
output out;
input n27;
input n40;
input n43;
input n45;
input n46;
input n48;
input n52;
input n61;
input n63;
input n64;
input n66;
input n71;
input n74;
input n76;
input n81;
input n85;
input n93;
input n97;
input n98;
input n99;
input n111;
input n115;
input n116;
input n117;
input n132;
input n133;
input n134;
input n135;
input n136;
input n140;
input n141;
input n142;
input n147;
input n149;
input n151;
input n188;
input n190;
input n191;
input n192;
input n203;
input n204;
input n205;
input n206;
input n218;
input n219;
input n220;
input n221;
input n235;
input n241;
input n243;
input n244;
input n248;
input n249;
input n252;
input n254;
input n255;
input n256;
input n329;
input n384;
input n387;
input n389;
input n477;
input n479;
input n480;
input n594;
input n597;
input n599;
input n601;
input n605;
input n608;
input n610;
input n612;
input n616;
input n619;
input n621;
input n623;
input n625;
input n684;
input n687;
input n689;
input n691;
input n695;
input n698;
input n700;
input n702;
input n706;
input n709;
input n711;
input n713;
input n717;
input n720;
input n722;
input n724;
input n758;
input n761;
input n763;
input n765;
input n769;
input n772;
input n774;
input n776;
input n780;
input n783;
input n785;
input n787;
input n791;
input n794;
input n796;
input n798;
input n831;
input n834;
input n836;
input n838;
input n842;
input n845;
input n847;
input n849;
input n853;
input n856;
input n858;
input n860;
input n864;
input n867;
input n869;
input n871;
input n901;
input n902;
input n904;
input n905;
input n920;
input n924;
input n926;
input n931;
input n933;
input n975;
input n987;
input n992;
input n997;
input n1002;
input n1010;
input n1013;
input n1022;
input n1026;
input n1032;
input n1034;
input n1036;
input n1038;
input n1040;
input n1048;
input n1051;
input n1053;
input n1055;
input n1057;
input n1064;
input n1065;
input n1075;
input n1078;
input n1082;
input n1087;
input n1090;
input n1093;
input n1096;
input n1101;
input n1103;
input n1105;
input n1107;
input n1109;
input n1114;
input n1116;
input n1123;
input n1126;
input n1128;
input n1138;
input n1140;
input n1142;
input n1144;
input n1146;
input n1151;
input n1153;
input n1156;
input n1158;
input n1160;
input n1164;
input n1166;
input n1169;
input n1172;
input n1176;
input n1178;
input n1181;
input n1183;
input n1184;
input n1192;
input n1197;
input n1201;
input n1205;
input n1209;
input n1214;
input n1216;
input n1219;
input n1221;
input n1223;
input n1227;
input n1229;
input n1232;
input n1235;
input n1239;
input n1243;
input n1248;
input n1252;
input n1253;
input n1263;
input n1265;
input n1267;
input n1269;
input n1271;
input n1277;
input n1279;
input n1281;
input n1283;
input n1288;
input n1289;
input n1292;
input n1295;
input n1298;
input n1303;
input n1306;
input n1309;
input n1312;
input n1313;
input n1320;
input n1321;
input n1324;
input n1327;
input n1330;
input n1335;
input n1338;
input n1341;
input n1344;
input n1349;
input n1351;
input n1354;
input n1358;
input n1360;
input n1365;
input n1367;
input n1373;
input n1376;
input n1377;
input n1387;
input n1389;
input n1391;
input n1393;
input n1395;
input n1398;
input n1400;
input n1406;
input n1408;
input n1410;
input n1412;
input n1414;
input n1419;
input n1422;
input n1424;
input n1426;
input n1429;
input n1431;
input n1432;
input n1439;
input n1440;
input n1443;
input n1446;
input n1449;
input n1454;
input n1457;
input n1460;
input n1463;
input n1468;
input n1470;
input n1472;
input n1474;
input n1476;
input n1481;
input n1483;
input n1489;
input n1491;
input n1492;
input n1502;
input n1504;
input n1506;
input n1508;
input n1510;
input n1516;
input n1518;
input n1520;
input n1522;
input n1527;
input n1528;
input n1531;
input n1534;
input n1537;
input n1542;
input n1545;
input n1548;
input n1551;
input n1552;
input n1559;
input n1560;
input n1563;
input n1566;
input n1569;
input n1574;
input n1577;
input n1580;
input n1583;
input n1588;
input n1590;
input n1593;
input n1597;
input n1599;
input n1604;
input n1606;
input n1612;
input n1615;
input n1616;
input n1626;
input n1628;
input n1630;
input n1632;
input n1634;
input n1640;
input n1642;
input n1644;
input n1646;
input n1651;
input n1652;
input n1655;
input n1658;
input n1661;
input n1666;
input n1669;
input n1672;
input n1675;
input n1676;
input n1683;
input n1684;
input n1687;
input n1690;
input n1693;
input n1698;
input n1701;
input n1704;
input n1707;
input n1712;
input n1714;
input n1717;
input n1721;
input n1723;
input n1728;
input n1730;
input n1733;
input n1738;
input n1739;
input n1748;
input n1750;
input n1753;
input n1755;
input n1757;
input n1761;
input n1763;
input n1767;
input n1769;
input n1774;
input n1775;
input n1778;
input n1781;
input n1784;
input n1789;
input n1792;
input n1795;
input n1798;
input n1799;
input n1806;
input n1807;
input n1810;
input n1813;
input n1816;
input n1821;
input n1824;
input n1827;
input n1830;
input n1836;
input n1838;
input n1840;
input n1842;
input n1844;
input n1853;
input n1855;
input n1857;
input n1859;
input n1860;
input n1869;
input n1871;
input n1873;
input n1875;
input n1877;
input n1882;
input n1885;
input n1887;
input n1889;
input n1894;
input n1895;
input n1898;
input n1901;
input n1904;
input n1909;
input n1912;
input n1915;
input n1918;
input n1919;
input n1926;
input n1927;
input n1930;
input n1933;
input n1936;
input n1941;
input n1944;
input n1947;
input n1950;
input n1955;
input n1957;
input n1960;
input n1964;
input n1966;
input n1971;
input n1973;
input n1976;
input n1981;
input n1982;
input n1998;
input n2000;
input n2010;
input n2012;
input n2014;
input n2016;
input n2018;
input n2023;
input n2026;
input n2028;
input n2030;
input n2033;
input n2036;
input n2038;
input n2040;
input n2042;
input n2045;
input n2047;
input n2050;
input n2052;
input n2053;
input n2060;
input n2062;
input n2064;
input n2066;
input n2068;
input n2074;
input n2076;
input n2078;
input n2080;
input n2082;
input n2087;
input n2090;
input n2092;
input n2094;
input n2097;
input n2099;
input n2102;
input n2104;
input n2105;
input n2116;
input n2118;
input n2120;
input n2122;
input n2124;
input n2129;
input n2132;
input n2134;
input n2136;
input n2139;
input n2143;
input n2145;
input n2147;
input n2149;
input n2152;
input n2154;
input n2157;
input n2159;
input n2160;
input n2167;
input n2169;
input n2174;
input n2176;
input n2179;
input n2184;
input n2186;
input n2192;
input n2195;
input n2200;
input n2201;
input n2204;
input n2207;
input n2210;
input n2215;
input n2218;
input n2221;
input n2224;
input n2225;
input n2233;
input n2237;
input n2240;
input n2242;
input n2244;
input n2249;
input n2251;
input n2254;
input n2256;
input n2258;
input n2262;
input n2264;
input n2267;
input n2270;
input n2273;
input n2275;
input n2278;
input n2280;
input n2281;
input n2286;
input n2289;
input n2292;
input n2294;
input n2296;
input n2302;
input n2304;
input n2306;
input n2308;
input n2310;
input n2312;
input n2319;
input n2321;
input n2323;
input n2325;
input n2327;
input n2330;
input n2332;
input n2333;
input n2343;
input n2345;
input n2350;
input n2352;
input n2355;
input n2360;
input n2362;
input n2368;
input n2371;
input n2376;
input n2377;
input n2380;
input n2383;
input n2386;
input n2391;
input n2394;
input n2397;
input n2400;
input n2401;
input n2408;
input n2410;
input n2412;
input n2414;
input n2416;
input n2421;
input n2423;
input n2429;
input n2431;
input n2436;
input n2437;
input n2440;
input n2443;
input n2446;
input n2451;
input n2454;
input n2457;
input n2460;
input n2461;
input n2471;
input n2473;
input n2478;
input n2480;
input n2483;
input n2488;
input n2490;
input n2496;
input n2499;
input n2504;
input n2505;
input n2508;
input n2511;
input n2514;
input n2519;
input n2522;
input n2525;
input n2528;
input n2529;
input n2535;
input n2537;
input n2540;
input n2542;
input n2544;
input n2548;
input n2550;
input n2554;
input n2556;
input n2561;
input n2562;
input n2565;
input n2568;
input n2571;
input n2576;
input n2579;
input n2582;
input n2585;
input n2586;
input n2596;
input n2598;
input n2600;
input n2602;
input n2604;
input n2610;
input n2612;
input n2614;
input n2616;
input n2621;
input n2622;
input n2625;
input n2628;
input n2631;
input n2636;
input n2639;
input n2642;
input n2645;
input n2646;
input n2653;
input n2655;
input n2657;
input n2659;
input n2661;
input n2666;
input n2669;
input n2671;
input n2673;
input n2678;
input n2679;
input n2682;
input n2685;
input n2688;
input n2693;
input n2696;
input n2699;
input n2702;
input n2703;
input n2713;
input n2714;
input n2717;
input n2720;
input n2723;
input n2728;
input n2730;
input n2734;
input n2736;
input n2741;
input n2742;
input n2745;
input n2748;
input n2751;
input n2756;
input n2759;
input n2762;
input n2765;
input n2766;
input n2776;
input n2778;
input n2780;
input n2782;
input n2784;
input n2791;
input n2793;
input n2795;
input n2797;
input n2802;
input n2803;
input n2806;
input n2809;
input n2812;
input n2817;
input n2820;
input n2823;
input n2826;
input n2827;
input n2837;
input n2839;
input n2842;
input n2844;
input n2846;
input n2851;
input n2853;
input n2857;
input n2859;
input n2864;
input n2865;
input n2868;
input n2871;
input n2874;
input n2879;
input n2882;
input n2885;
input n2888;
input n2889;
input n2896;
input n2898;
input n2901;
input n2905;
input n2907;
input n2912;
input n2914;
input n2917;
input n2922;
input n2927;
input n2928;
input n2931;
input n2934;
input n2937;
input n2942;
input n2945;
input n2948;
input n2951;
input n2952;
input n2966;
input n2968;
input n2988;
input n2989;
input n2992;
input n2995;
input n2998;
input n3003;
input n3006;
input n3009;
input n3012;
input n3013;
input n3016;
input n3021;
input n3023;
input n3026;
input n3028;
input n3030;
input n3036;
input n3038;
input n3042;
input n3044;
input n3056;
input n3057;
input n3060;
input n3063;
input n3066;
input n3071;
input n3074;
input n3077;
input n3080;
input n3081;
input n3091;
input n3093;
input n3095;
input n3097;
input n3099;
input n3105;
input n3107;
input n3109;
input n3111;
input n3112;
input n3122;
input n3124;
input n3127;
input n3129;
input n3146;
input n3147;
input n3150;
input n3153;
input n3156;
input n3161;
input n3164;
input n3167;
input n3170;
input n3171;
input n3175;
input n3182;
input n3184;
input n3186;
input n3188;
input n3190;
input n3196;
input n3199;
input n3201;
input n3203;
input n3213;
input n3214;
input n3217;
input n3220;
input n3223;
input n3228;
input n3231;
input n3234;
input n3237;
input n3238;
input n3245;
input n3247;
input n3250;
input n3252;
input n3254;
input n3260;
input n3262;
input n3266;
input n3268;
input n3270;
input n3282;
input n3283;
input n3286;
input n3289;
input n3292;
input n3297;
input n3300;
input n3303;
input n3306;
input n3307;
input n3314;
input n3316;
input n3321;
input n3323;
input n3326;
input n3333;
input n3336;
input n3338;
input n3340;
input n3341;
input n3355;
input n3356;
input n3359;
input n3362;
input n3365;
input n3370;
input n3373;
input n3376;
input n3379;
input n3380;
input n3383;
input n3389;
input n3391;
input n3393;
input n3395;
input n3397;
input n3405;
input n3407;
input n3409;
input n3411;
input n3428;
input n3429;
input n3432;
input n3435;
input n3438;
input n3443;
input n3446;
input n3449;
input n3452;
input n3453;
input n3461;
input n3463;
input n3465;
input n3467;
input n3469;
input n3477;
input n3479;
input n3481;
input n3483;
input n3484;
input n3495;
input n3496;
input n3499;
input n3502;
input n3505;
input n3510;
input n3513;
input n3516;
input n3519;
input n3520;
input n3525;
input n3534;
input n3536;
input n3538;
input n3540;
input n3542;
input n3549;
input n3551;
input n3553;
input n3555;
input n3851;
input n3853;
input n3857;
input n3859;
input n3864;
input n3866;
input n3884;
input n3886;
input n3892;
input n3894;
input n3909;
input n3911;
input n3977;
input n3979;
input n3991;
input n3993;
input n4011;
input n4013;
input n4032;
input n4038;
input n4054;
input n4061;
input n4080;
input n4087;
input n4093;
input n4095;
input n4520;
input n4522;
input n5454;
input n5455;
input n5458;
input n5459;
input n5466;
input n5467;
input n5470;
input n5471;
input n5505;
input n5506;
input n5511;
input n5512;
input n5549;
input n5550;
input n5553;
input n5554;
input n5582;
input n5583;
input n5587;
input n5588;
input n5619;
input n5620;
input n5623;
input n5624;
input n5661;
input n5662;
input n5666;
input n5667;
input n5709;
input n5710;
input n5713;
input n5714;
input n5745;
input n5746;
input n5749;
input n5750;
input n5788;
input n5789;
input n5792;
input n5793;
input n5824;
input n5825;
input n5828;
input n5829;
input n5866;
input n5867;
input n5870;
input n5871;
input n5891;
input n5892;
input n5897;
input n5898;
input n5927;
input n5928;
input n5931;
input n5932;
input n5963;
input n5964;
input n5969;
input n5970;
input n5999;
input n6000;
input n6003;
input n6004;
input n6163;
input n6166;
input n6182;
input n6186;
input n6196;
input n6207;
input n6211;
input n6215;
input n6227;
input n6237;
input n6240;
input n6242;
input n6246;
input n6248;
input n6262;
input n6264;
input n6276;
input n6286;
input n6289;
input n6291;
input n6295;
input n6297;
input n6311;
input n6313;
input n6327;
input n6335;
input n6338;
input n6340;
input n6356;
input n6358;
input n6361;
input n6363;
input n6378;
input n6389;
input n6392;
input n6394;
input n6400;
input n6415;
input n6417;
input n6419;
input n6431;
input n6441;
input n6444;
input n6446;
input n6462;
input n6464;
input n6467;
input n6469;
input n6484;
input n6494;
input n6497;
input n6499;
input n6505;
input n6520;
input n6522;
input n6524;
input n6541;
input n6543;
input n6545;
input n6555;
input n6576;
input n6578;
input n6581;
input n6583;
input n6761;
input n6764;
input n6877;
input n6880;
input n6971;
input n6974;
input n7099;
input n7102;
input n7357;
input n7360;
input n7376;
input n7379;
input n7510;
input n7513;
input n7619;
input n7622;
input n7733;
input n7743;
input n7746;
input n7748;
input n7750;
input n7754;
input n7757;
input n7759;
input n7761;
input n7765;
input n7768;
input n7770;
input n7772;
input n7776;
input n7779;
input n7781;
input n7783;
input n7791;
input n7794;
input n7796;
input n7798;
input n7802;
input n7805;
input n7807;
input n7809;
input n7813;
input n7816;
input n7818;
input n7820;
input n7824;
input n7827;
input n7829;
input n7831;
input n7875;
input n7902;
input n7917;
input n7932;
input n7947;
input n7962;
input n7981;
input n8059;
input n8070;
input n8090;
input n8105;
input n8120;
input n8140;
input n8155;
input n8164;
input n8259;
input n8272;
input n8278;
input n8296;
input n8316;
input n8326;
input n8340;
input n8392;
input n8399;
input n8418;
input n8449;
input n8510;
input n8524;
input n8534;
input n8554;
input n8568;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n44;
wire n47;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n137;
wire n138;
wire n139;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n242;
wire n245;
wire n246;
wire n247;
wire n250;
wire n251;
wire n253;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n385;
wire n386;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n478;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n595;
wire n596;
wire n598;
wire n600;
wire n602;
wire n603;
wire n604;
wire n606;
wire n607;
wire n609;
wire n611;
wire n613;
wire n614;
wire n615;
wire n617;
wire n618;
wire n620;
wire n622;
wire n624;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n685;
wire n686;
wire n688;
wire n690;
wire n692;
wire n693;
wire n694;
wire n696;
wire n697;
wire n699;
wire n701;
wire n703;
wire n704;
wire n705;
wire n707;
wire n708;
wire n710;
wire n712;
wire n714;
wire n715;
wire n716;
wire n718;
wire n719;
wire n721;
wire n723;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n759;
wire n760;
wire n762;
wire n764;
wire n766;
wire n767;
wire n768;
wire n770;
wire n771;
wire n773;
wire n775;
wire n777;
wire n778;
wire n779;
wire n781;
wire n782;
wire n784;
wire n786;
wire n788;
wire n789;
wire n790;
wire n792;
wire n793;
wire n795;
wire n797;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n832;
wire n833;
wire n835;
wire n837;
wire n839;
wire n840;
wire n841;
wire n843;
wire n844;
wire n846;
wire n848;
wire n850;
wire n851;
wire n852;
wire n854;
wire n855;
wire n857;
wire n859;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n868;
wire n870;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n903;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n921;
wire n922;
wire n923;
wire n925;
wire n927;
wire n928;
wire n929;
wire n930;
wire n932;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n988;
wire n989;
wire n990;
wire n991;
wire n993;
wire n994;
wire n995;
wire n996;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1011;
wire n1012;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1023;
wire n1024;
wire n1025;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1033;
wire n1035;
wire n1037;
wire n1039;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1049;
wire n1050;
wire n1052;
wire n1054;
wire n1056;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1076;
wire n1077;
wire n1079;
wire n1080;
wire n1081;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1088;
wire n1089;
wire n1091;
wire n1092;
wire n1094;
wire n1095;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1102;
wire n1104;
wire n1106;
wire n1108;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1115;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1124;
wire n1125;
wire n1127;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1139;
wire n1141;
wire n1143;
wire n1145;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1152;
wire n1154;
wire n1155;
wire n1157;
wire n1159;
wire n1161;
wire n1162;
wire n1163;
wire n1165;
wire n1167;
wire n1168;
wire n1170;
wire n1171;
wire n1173;
wire n1174;
wire n1175;
wire n1177;
wire n1179;
wire n1180;
wire n1182;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1198;
wire n1199;
wire n1200;
wire n1202;
wire n1203;
wire n1204;
wire n1206;
wire n1207;
wire n1208;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1215;
wire n1217;
wire n1218;
wire n1220;
wire n1222;
wire n1224;
wire n1225;
wire n1226;
wire n1228;
wire n1230;
wire n1231;
wire n1233;
wire n1234;
wire n1236;
wire n1237;
wire n1238;
wire n1240;
wire n1241;
wire n1242;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1249;
wire n1250;
wire n1251;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1264;
wire n1266;
wire n1268;
wire n1270;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1278;
wire n1280;
wire n1282;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1290;
wire n1291;
wire n1293;
wire n1294;
wire n1296;
wire n1297;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1304;
wire n1305;
wire n1307;
wire n1308;
wire n1310;
wire n1311;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1322;
wire n1323;
wire n1325;
wire n1326;
wire n1328;
wire n1329;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1336;
wire n1337;
wire n1339;
wire n1340;
wire n1342;
wire n1343;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1350;
wire n1352;
wire n1353;
wire n1355;
wire n1356;
wire n1357;
wire n1359;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1366;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1374;
wire n1375;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1388;
wire n1390;
wire n1392;
wire n1394;
wire n1396;
wire n1397;
wire n1399;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1407;
wire n1409;
wire n1411;
wire n1413;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1420;
wire n1421;
wire n1423;
wire n1425;
wire n1427;
wire n1428;
wire n1430;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1441;
wire n1442;
wire n1444;
wire n1445;
wire n1447;
wire n1448;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1455;
wire n1456;
wire n1458;
wire n1459;
wire n1461;
wire n1462;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1469;
wire n1471;
wire n1473;
wire n1475;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1482;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1490;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1503;
wire n1505;
wire n1507;
wire n1509;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1517;
wire n1519;
wire n1521;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1529;
wire n1530;
wire n1532;
wire n1533;
wire n1535;
wire n1536;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1543;
wire n1544;
wire n1546;
wire n1547;
wire n1549;
wire n1550;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1561;
wire n1562;
wire n1564;
wire n1565;
wire n1567;
wire n1568;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1575;
wire n1576;
wire n1578;
wire n1579;
wire n1581;
wire n1582;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1589;
wire n1591;
wire n1592;
wire n1594;
wire n1595;
wire n1596;
wire n1598;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1605;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1613;
wire n1614;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1627;
wire n1629;
wire n1631;
wire n1633;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1641;
wire n1643;
wire n1645;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1653;
wire n1654;
wire n1656;
wire n1657;
wire n1659;
wire n1660;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1667;
wire n1668;
wire n1670;
wire n1671;
wire n1673;
wire n1674;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1685;
wire n1686;
wire n1688;
wire n1689;
wire n1691;
wire n1692;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1699;
wire n1700;
wire n1702;
wire n1703;
wire n1705;
wire n1706;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1713;
wire n1715;
wire n1716;
wire n1718;
wire n1719;
wire n1720;
wire n1722;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1729;
wire n1731;
wire n1732;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1749;
wire n1751;
wire n1752;
wire n1754;
wire n1756;
wire n1758;
wire n1759;
wire n1760;
wire n1762;
wire n1764;
wire n1765;
wire n1766;
wire n1768;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1776;
wire n1777;
wire n1779;
wire n1780;
wire n1782;
wire n1783;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1790;
wire n1791;
wire n1793;
wire n1794;
wire n1796;
wire n1797;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1808;
wire n1809;
wire n1811;
wire n1812;
wire n1814;
wire n1815;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1822;
wire n1823;
wire n1825;
wire n1826;
wire n1828;
wire n1829;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1837;
wire n1839;
wire n1841;
wire n1843;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1854;
wire n1856;
wire n1858;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1870;
wire n1872;
wire n1874;
wire n1876;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1883;
wire n1884;
wire n1886;
wire n1888;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1896;
wire n1897;
wire n1899;
wire n1900;
wire n1902;
wire n1903;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1910;
wire n1911;
wire n1913;
wire n1914;
wire n1916;
wire n1917;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1928;
wire n1929;
wire n1931;
wire n1932;
wire n1934;
wire n1935;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1942;
wire n1943;
wire n1945;
wire n1946;
wire n1948;
wire n1949;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1956;
wire n1958;
wire n1959;
wire n1961;
wire n1962;
wire n1963;
wire n1965;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1972;
wire n1974;
wire n1975;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1999;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2011;
wire n2013;
wire n2015;
wire n2017;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2024;
wire n2025;
wire n2027;
wire n2029;
wire n2031;
wire n2032;
wire n2034;
wire n2035;
wire n2037;
wire n2039;
wire n2041;
wire n2043;
wire n2044;
wire n2046;
wire n2048;
wire n2049;
wire n2051;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2061;
wire n2063;
wire n2065;
wire n2067;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2075;
wire n2077;
wire n2079;
wire n2081;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2088;
wire n2089;
wire n2091;
wire n2093;
wire n2095;
wire n2096;
wire n2098;
wire n2100;
wire n2101;
wire n2103;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2117;
wire n2119;
wire n2121;
wire n2123;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2130;
wire n2131;
wire n2133;
wire n2135;
wire n2137;
wire n2138;
wire n2140;
wire n2141;
wire n2142;
wire n2144;
wire n2146;
wire n2148;
wire n2150;
wire n2151;
wire n2153;
wire n2155;
wire n2156;
wire n2158;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2168;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2175;
wire n2177;
wire n2178;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2185;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2193;
wire n2194;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2202;
wire n2203;
wire n2205;
wire n2206;
wire n2208;
wire n2209;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2216;
wire n2217;
wire n2219;
wire n2220;
wire n2222;
wire n2223;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2234;
wire n2235;
wire n2236;
wire n2238;
wire n2239;
wire n2241;
wire n2243;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2250;
wire n2252;
wire n2253;
wire n2255;
wire n2257;
wire n2259;
wire n2260;
wire n2261;
wire n2263;
wire n2265;
wire n2266;
wire n2268;
wire n2269;
wire n2271;
wire n2272;
wire n2274;
wire n2276;
wire n2277;
wire n2279;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2287;
wire n2288;
wire n2290;
wire n2291;
wire n2293;
wire n2295;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2303;
wire n2305;
wire n2307;
wire n2309;
wire n2311;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2320;
wire n2322;
wire n2324;
wire n2326;
wire n2328;
wire n2329;
wire n2331;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2344;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2351;
wire n2353;
wire n2354;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2361;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2369;
wire n2370;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2378;
wire n2379;
wire n2381;
wire n2382;
wire n2384;
wire n2385;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2392;
wire n2393;
wire n2395;
wire n2396;
wire n2398;
wire n2399;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2409;
wire n2411;
wire n2413;
wire n2415;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2422;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2430;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2438;
wire n2439;
wire n2441;
wire n2442;
wire n2444;
wire n2445;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2452;
wire n2453;
wire n2455;
wire n2456;
wire n2458;
wire n2459;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2472;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2479;
wire n2481;
wire n2482;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2489;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2497;
wire n2498;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2506;
wire n2507;
wire n2509;
wire n2510;
wire n2512;
wire n2513;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2520;
wire n2521;
wire n2523;
wire n2524;
wire n2526;
wire n2527;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2536;
wire n2538;
wire n2539;
wire n2541;
wire n2543;
wire n2545;
wire n2546;
wire n2547;
wire n2549;
wire n2551;
wire n2552;
wire n2553;
wire n2555;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2563;
wire n2564;
wire n2566;
wire n2567;
wire n2569;
wire n2570;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2577;
wire n2578;
wire n2580;
wire n2581;
wire n2583;
wire n2584;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2597;
wire n2599;
wire n2601;
wire n2603;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2611;
wire n2613;
wire n2615;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2623;
wire n2624;
wire n2626;
wire n2627;
wire n2629;
wire n2630;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2637;
wire n2638;
wire n2640;
wire n2641;
wire n2643;
wire n2644;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2654;
wire n2656;
wire n2658;
wire n2660;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2667;
wire n2668;
wire n2670;
wire n2672;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2680;
wire n2681;
wire n2683;
wire n2684;
wire n2686;
wire n2687;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2694;
wire n2695;
wire n2697;
wire n2698;
wire n2700;
wire n2701;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2715;
wire n2716;
wire n2718;
wire n2719;
wire n2721;
wire n2722;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2729;
wire n2731;
wire n2732;
wire n2733;
wire n2735;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2743;
wire n2744;
wire n2746;
wire n2747;
wire n2749;
wire n2750;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2757;
wire n2758;
wire n2760;
wire n2761;
wire n2763;
wire n2764;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2777;
wire n2779;
wire n2781;
wire n2783;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2792;
wire n2794;
wire n2796;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2804;
wire n2805;
wire n2807;
wire n2808;
wire n2810;
wire n2811;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2818;
wire n2819;
wire n2821;
wire n2822;
wire n2824;
wire n2825;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2838;
wire n2840;
wire n2841;
wire n2843;
wire n2845;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2852;
wire n2854;
wire n2855;
wire n2856;
wire n2858;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2866;
wire n2867;
wire n2869;
wire n2870;
wire n2872;
wire n2873;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2880;
wire n2881;
wire n2883;
wire n2884;
wire n2886;
wire n2887;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2897;
wire n2899;
wire n2900;
wire n2902;
wire n2903;
wire n2904;
wire n2906;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2913;
wire n2915;
wire n2916;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2929;
wire n2930;
wire n2932;
wire n2933;
wire n2935;
wire n2936;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2943;
wire n2944;
wire n2946;
wire n2947;
wire n2949;
wire n2950;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2967;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2990;
wire n2991;
wire n2993;
wire n2994;
wire n2996;
wire n2997;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3004;
wire n3005;
wire n3007;
wire n3008;
wire n3010;
wire n3011;
wire n3014;
wire n3015;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3022;
wire n3024;
wire n3025;
wire n3027;
wire n3029;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3037;
wire n3039;
wire n3040;
wire n3041;
wire n3043;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3058;
wire n3059;
wire n3061;
wire n3062;
wire n3064;
wire n3065;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3072;
wire n3073;
wire n3075;
wire n3076;
wire n3078;
wire n3079;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3092;
wire n3094;
wire n3096;
wire n3098;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3106;
wire n3108;
wire n3110;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3123;
wire n3125;
wire n3126;
wire n3128;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3148;
wire n3149;
wire n3151;
wire n3152;
wire n3154;
wire n3155;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3162;
wire n3163;
wire n3165;
wire n3166;
wire n3168;
wire n3169;
wire n3172;
wire n3173;
wire n3174;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3183;
wire n3185;
wire n3187;
wire n3189;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3197;
wire n3198;
wire n3200;
wire n3202;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3215;
wire n3216;
wire n3218;
wire n3219;
wire n3221;
wire n3222;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3229;
wire n3230;
wire n3232;
wire n3233;
wire n3235;
wire n3236;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3246;
wire n3248;
wire n3249;
wire n3251;
wire n3253;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3261;
wire n3263;
wire n3264;
wire n3265;
wire n3267;
wire n3269;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3284;
wire n3285;
wire n3287;
wire n3288;
wire n3290;
wire n3291;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3298;
wire n3299;
wire n3301;
wire n3302;
wire n3304;
wire n3305;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3315;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3322;
wire n3324;
wire n3325;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3334;
wire n3335;
wire n3337;
wire n3339;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3357;
wire n3358;
wire n3360;
wire n3361;
wire n3363;
wire n3364;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3371;
wire n3372;
wire n3374;
wire n3375;
wire n3377;
wire n3378;
wire n3381;
wire n3382;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3390;
wire n3392;
wire n3394;
wire n3396;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3406;
wire n3408;
wire n3410;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3430;
wire n3431;
wire n3433;
wire n3434;
wire n3436;
wire n3437;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3444;
wire n3445;
wire n3447;
wire n3448;
wire n3450;
wire n3451;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3462;
wire n3464;
wire n3466;
wire n3468;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3478;
wire n3480;
wire n3482;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3497;
wire n3498;
wire n3500;
wire n3501;
wire n3503;
wire n3504;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3511;
wire n3512;
wire n3514;
wire n3515;
wire n3517;
wire n3518;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3535;
wire n3537;
wire n3539;
wire n3541;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3550;
wire n3552;
wire n3554;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3852;
wire n3854;
wire n3855;
wire n3856;
wire n3858;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3865;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3885;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3893;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3910;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3978;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3992;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4012;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4094;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4521;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5456;
wire n5457;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5468;
wire n5469;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5551;
wire n5552;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5584;
wire n5585;
wire n5586;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5621;
wire n5622;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5663;
wire n5664;
wire n5665;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5711;
wire n5712;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5747;
wire n5748;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5790;
wire n5791;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5826;
wire n5827;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5868;
wire n5869;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5929;
wire n5930;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n6001;
wire n6002;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6164;
wire n6165;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6183;
wire n6184;
wire n6185;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6208;
wire n6209;
wire n6210;
wire n6212;
wire n6213;
wire n6214;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6238;
wire n6239;
wire n6241;
wire n6243;
wire n6244;
wire n6245;
wire n6247;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6263;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6287;
wire n6288;
wire n6290;
wire n6292;
wire n6293;
wire n6294;
wire n6296;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6312;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6336;
wire n6337;
wire n6339;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6357;
wire n6359;
wire n6360;
wire n6362;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6390;
wire n6391;
wire n6393;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6416;
wire n6418;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6442;
wire n6443;
wire n6445;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6463;
wire n6465;
wire n6466;
wire n6468;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6495;
wire n6496;
wire n6498;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6521;
wire n6523;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6542;
wire n6544;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6577;
wire n6579;
wire n6580;
wire n6582;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6762;
wire n6763;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6878;
wire n6879;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6972;
wire n6973;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7100;
wire n7101;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7358;
wire n7359;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7377;
wire n7378;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7511;
wire n7512;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7620;
wire n7621;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7744;
wire n7745;
wire n7747;
wire n7749;
wire n7751;
wire n7752;
wire n7753;
wire n7755;
wire n7756;
wire n7758;
wire n7760;
wire n7762;
wire n7763;
wire n7764;
wire n7766;
wire n7767;
wire n7769;
wire n7771;
wire n7773;
wire n7774;
wire n7775;
wire n7777;
wire n7778;
wire n7780;
wire n7782;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7792;
wire n7793;
wire n7795;
wire n7797;
wire n7799;
wire n7800;
wire n7801;
wire n7803;
wire n7804;
wire n7806;
wire n7808;
wire n7810;
wire n7811;
wire n7812;
wire n7814;
wire n7815;
wire n7817;
wire n7819;
wire n7821;
wire n7822;
wire n7823;
wire n7825;
wire n7826;
wire n7828;
wire n7830;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10449;
wire n10450;
wire n10451;
wire n10452;
wire n10453;
wire n10454;
wire n10455;
xor (out,n0,n9707);
nand (n0,n1,n7724);
not (n1,n2);
nand (n2,n3,n7714);
or (n3,n4,n7711);
nor (n4,n5,n7705);
and (n5,n6,n7485);
nand (n6,n7,n7477);
or (n7,n8,n6963);
nand (n8,n9,n6851);
nand (n9,n10,n6757);
not (n10,n11);
or (n11,1'b0,n13,n4652,n4654,n4656);
and (n13,n14,n912);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n4648);
and (s0n14,notn14,1'b0);
and (s1n14,n4648,n15);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n4628);
and (s0n15,notn15,n16);
and (s1n15,n4628,1'b0);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n4502);
and (s0n16,notn16,n17);
and (s1n16,n4502,1'b1);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n28);
and (s0n17,notn17,n18);
and (s1n17,n28,n3841);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n28);
and (s0n18,notn18,n19);
and (s1n18,n28,n3840);
xor (n19,n20,n3823);
xor (n20,n21,n3778);
xor (n21,n22,n3723);
xor (n22,n23,n3713);
xor (n23,n24,n1992);
xor (n24,n25,n921);
xor (n25,n26,n919);
wire s0n26,s1n26,notn26;
or (n26,s0n26,s1n26);
not(notn26,n28);
and (s0n26,notn26,1'b0);
and (s1n26,n28,n27);
or (n28,n29,n916);
or (n29,n30,n911);
and (n30,n31,n897);
and (n31,n32,n677,n750,n824);
not (n32,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n676);
and (s0n33,notn33,1'b0);
and (s1n33,n676,n34);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n676);
and (s0n34,notn34,n35);
and (s1n34,n676,n628);
wire s0n35,s1n35,notn35;
or (n35,s0n35,s1n35);
not(notn35,n626);
and (s0n35,notn35,1'b0);
and (s1n35,n626,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n625);
and (s0n36,notn36,n37);
and (s1n36,n625,n616);
or (n37,n38,n592,n603,n614);
and (n38,n39,n62);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n56);
and (s0n39,notn39,n40);
and (s1n39,n56,n41);
or (n41,n42,n47,n51,n54);
and (n42,n43,n44);
nor (n44,n45,n46);
and (n47,n48,n49);
and (n49,n45,n50);
not (n50,n46);
and (n51,n52,n53);
nor (n53,n45,n50);
and (n54,n40,n55);
and (n55,n45,n46);
nor (n56,n57,n90);
nor (n57,n58,n77);
and (n58,n59,n76);
or (n59,n60,n65,n70,n73);
and (n60,n61,n62);
and (n62,n63,n64);
and (n65,n66,n67);
not (n67,n68);
nand (n68,n69,n64);
not (n69,n63);
and (n70,n71,n72);
nor (n72,n69,n64);
and (n73,n74,n75);
nor (n75,n63,n64);
nor (n77,n78,n86,n76);
and (n78,n79,n84);
nand (n79,n80,n82);
or (n80,n81,n74);
or (n82,n83,n66);
not (n83,n81);
not (n84,n85);
and (n86,n87,n85);
nand (n87,n88,n89);
or (n88,n81,n71);
or (n89,n83,n61);
nand (n90,n91,n100);
or (n91,n92,n94);
not (n92,n93);
not (n94,n95);
nand (n95,n96,n99);
nor (n96,n97,n98);
nand (n100,n101,n556);
nand (n101,n102,n548);
or (n102,n103,n472);
not (n103,n104);
or (n104,1'b0,n105,n392,n470);
and (n105,n106,n391);
wire s0n106,s1n106,notn106;
or (n106,s0n106,s1n106);
not(notn106,n382);
and (s0n106,notn106,n107);
and (s1n106,n382,1'b0);
wire s0n107,s1n107,notn107;
or (n107,s0n107,s1n107);
not(notn107,n318);
and (s0n107,notn107,1'b0);
and (s1n107,n318,n108);
or (n108,n109,n292,n298,n304,n309,1'b0,1'b0,1'b0);
and (n109,n110,n118);
xnor (n110,n111,n112);
not (n112,n113);
nor (n113,n114,n117);
or (n114,n115,n116);
and (n118,n119,n261,n280,n288);
wire s0n119,s1n119,notn119;
or (n119,s0n119,s1n119);
not(notn119,n152);
and (s0n119,notn119,n120);
and (s1n119,n152,1'b0);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n150);
and (s0n120,notn120,n121);
and (s1n120,n150,n148);
wire s0n121,s1n121,notn121;
or (n121,s0n121,s1n121);
not(notn121,n143);
and (s0n121,notn121,n122);
and (s1n121,n143,n137);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n136);
and (s0n122,notn122,n123);
and (s1n122,n136,1'b0);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n135);
and (s0n123,notn123,n124);
and (s1n123,n135,1'b1);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n134);
and (s0n124,notn124,n125);
and (s1n124,n134,1'b0);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n133);
and (s0n125,notn125,n126);
and (s1n125,n133,1'b1);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n132);
and (s0n126,notn126,n127);
and (s1n126,n132,1'b0);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n111);
and (s0n127,notn127,n128);
and (s1n127,n111,1'b1);
wire s0n128,s1n128,notn128;
or (n128,s0n128,s1n128);
not(notn128,n117);
and (s0n128,notn128,n129);
and (s1n128,n117,1'b0);
wire s0n129,s1n129,notn129;
or (n129,s0n129,s1n129);
not(notn129,n115);
and (s0n129,notn129,n130);
and (s1n129,n115,1'b1);
not (n130,n116);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n142);
and (s0n137,notn137,n138);
and (s1n137,n142,1'b0);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n141);
and (s0n138,notn138,n139);
and (s1n138,n141,1'b1);
not (n139,n140);
or (n143,n144,n147);
or (n144,n142,n145);
not (n145,n146);
nor (n146,n141,n140);
not (n148,n149);
or (n150,n149,n151);
not (n152,n153);
or (n153,n154,n259);
or (n154,n155,n257);
or (n155,n156,n251);
or (n156,n157,n250);
or (n157,n158,n246);
or (n158,n159,n245);
or (n159,n160,n240);
or (n160,n161,n239);
or (n161,n162,n238);
or (n162,n163,n236);
or (n163,n164,n233);
or (n164,n165,n232);
or (n165,n166,n231);
or (n166,n167,n230);
or (n167,n168,n229);
or (n168,n169,n227);
or (n169,n170,n225);
or (n170,n171,n224);
or (n171,n172,n222);
or (n172,n173,n216);
or (n173,n174,n215);
or (n174,n175,n214);
or (n175,n176,n213);
or (n176,n177,n212);
or (n177,n178,n211);
or (n178,n179,n209);
or (n179,n180,n207);
or (n180,n181,n201);
or (n181,n182,n200);
or (n182,n183,n199);
or (n183,n184,n198);
or (n184,n185,n197);
or (n185,n186,n195);
or (n186,n187,n193);
nor (n187,n188,n189,n191,n192);
not (n189,n190);
nor (n193,n188,n189,n194,n192);
not (n194,n191);
and (n195,n188,n190,n191,n196);
not (n196,n192);
and (n197,n188,n189,n191,n196);
nor (n198,n188,n190,n194,n192);
and (n199,n188,n189,n191,n192);
and (n200,n188,n190,n191,n192);
nor (n201,n202,n204,n205,n206);
not (n202,n203);
nor (n207,n202,n208,n205,n206);
not (n208,n204);
and (n209,n202,n204,n205,n210);
not (n210,n206);
and (n211,n203,n204,n205,n210);
and (n212,n203,n208,n205,n210);
and (n213,n202,n208,n205,n206);
and (n214,n203,n208,n205,n206);
and (n215,n203,n204,n205,n206);
nor (n216,n217,n219,n220,n221);
not (n217,n218);
nor (n222,n217,n223,n220,n221);
not (n223,n219);
nor (n224,n218,n223,n220,n221);
nor (n225,n217,n223,n226,n221);
not (n226,n220);
nor (n227,n218,n219,n226,n228);
not (n228,n221);
and (n229,n217,n219,n220,n221);
and (n230,n217,n219,n226,n221);
and (n231,n218,n219,n226,n221);
and (n232,n218,n223,n226,n221);
nor (n233,n234,n99,n97,n98);
not (n234,n235);
nor (n236,n235,n237,n97,n98);
not (n237,n99);
and (n238,n234,n237,n97,n98);
and (n239,n235,n237,n97,n98);
nor (n240,n241,n242,n244);
not (n242,n243);
and (n245,n241,n243,n244);
nor (n246,n247,n249);
not (n247,n248);
and (n250,n247,n249);
nor (n251,n252,n253,n255,n256);
not (n253,n254);
and (n257,n252,n254,n255,n258);
not (n258,n256);
and (n259,n260,n253,n255,n258);
not (n260,n252);
not (n261,n262);
or (n262,n152,n263);
nand (n263,n264,n279);
or (n264,n265,n278);
nor (n265,n266,n276);
nor (n266,n267,n273);
and (n267,n268,n272);
nand (n268,n269,n270);
or (n269,n115,n117);
wire s0n270,s1n270,notn270;
or (n270,s0n270,s1n270);
not(notn270,n132);
and (s0n270,notn270,n271);
and (s1n270,n132,1'b0);
not (n271,n111);
nor (n272,n133,n134);
not (n273,n274);
wire s0n274,s1n274,notn274;
or (n274,s0n274,s1n274);
not(notn274,n136);
and (s0n274,notn274,n275);
and (s1n274,n136,1'b0);
not (n275,n135);
nand (n276,n277,n139);
not (n277,n147);
or (n278,n142,n141);
not (n279,n150);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n152);
and (s0n280,notn280,n281);
and (s1n280,n152,1'b0);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n150);
and (s0n281,notn281,n282);
and (s1n281,n150,1'b0);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n143);
and (s0n282,notn282,n283);
and (s1n282,n143,n287);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n136);
and (s0n283,notn283,n284);
and (s1n283,n136,1'b1);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n135);
and (s0n284,notn284,n285);
and (s1n284,n135,1'b1);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n134);
and (s0n285,notn285,n286);
and (s1n285,n134,1'b0);
wire s0n286,s1n286,notn286;
or (n286,s0n286,s1n286);
not(notn286,n133);
and (s0n286,notn286,n270);
and (s1n286,n133,1'b0);
not (n287,n278);
not (n288,n289);
wire s0n289,s1n289,notn289;
or (n289,s0n289,s1n289);
not(notn289,n152);
and (s0n289,notn289,n290);
and (s1n289,n152,1'b0);
wire s0n290,s1n290,notn290;
or (n290,s0n290,s1n290);
not(notn290,n150);
and (s0n290,notn290,n291);
and (s1n290,n150,1'b0);
wire s0n291,s1n291,notn291;
or (n291,s0n291,s1n291);
not(notn291,n143);
and (s0n291,notn291,n274);
and (s1n291,n143,1'b0);
and (n292,n293,n296);
xnor (n293,n133,n294);
or (n294,n132,n295);
or (n295,n111,n117);
and (n296,n297,n261,n280,n288);
not (n297,n119);
and (n298,n299,n303);
xnor (n299,n135,n300);
not (n300,n301);
nor (n301,n302,n134);
or (n302,n133,n132);
and (n303,n119,n262,n280,n288);
and (n304,n305,n308);
xnor (n305,n147,n306);
or (n306,n136,n307);
or (n307,n135,n134);
and (n308,n297,n262,n280,n288);
and (n309,n310,n313);
not (n310,n311);
nand (n311,n312,n288,n119,n261);
not (n312,n280);
not (n313,n314);
nand (n314,n315,n141);
or (n315,n140,n316);
not (n316,n317);
nor (n317,n136,n147);
or (n318,n319,n365);
or (n319,n320,n341,n349,n355);
nand (n320,n321,n332);
or (n321,n322,n241);
nand (n322,n323,n330,n243);
nor (n323,n324,n98);
not (n324,n325);
and (n325,n326,n327,n228);
nor (n326,n220,n219);
nor (n327,n328,n218);
not (n328,n329);
nor (n330,n331,n235);
nand (n331,n237,n97);
nor (n332,n333,n335);
and (n333,n323,n334,n248);
nor (n334,n234,n331);
nand (n335,n336,n340);
or (n336,n337,n339);
nor (n337,n338,n326);
and (n338,n219,n228);
nand (n339,n218,n329);
nand (n340,n226,n327,n219);
nor (n341,n342,n347,n206);
nand (n342,n323,n343);
and (n343,n344,n346,n237);
not (n344,n345);
or (n345,n188,n190,n191,n192);
nor (n346,n97,n235);
nor (n347,n348,n203);
and (n348,n205,n204);
nor (n349,n350,n351,n352,n344);
not (n350,n346);
not (n351,n323);
nor (n352,n353,n354);
and (n353,n191,n188);
nor (n354,n188,n192);
nor (n355,n356,n363);
nor (n356,n357,n330);
and (n357,n358,n362);
not (n358,n359);
nor (n359,n360,n361);
and (n360,n346,n99);
and (n361,n235,n237);
not (n362,n98);
nand (n363,n364,n325);
or (n364,n331,n98);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n328);
and (s0n365,notn365,n366);
and (s1n365,n328,1'b0);
wire s0n366,s1n366,notn366;
or (n366,s0n366,s1n366);
not(notn366,n381);
and (s0n366,notn366,n367);
and (s1n366,n381,n380);
wire s0n367,s1n367,notn367;
or (n367,s0n367,s1n367);
not(notn367,n379);
and (s0n367,notn367,n368);
and (s1n367,n379,n371);
wire s0n368,s1n368,notn368;
or (n368,s0n368,s1n368);
not(notn368,n345);
and (s0n368,notn368,n369);
and (s1n368,n345,1'b0);
or (n369,n370,n215);
or (n370,n213,n214);
or (n371,1'b0,n239,n372,n377,1'b0);
and (n372,n373,n376);
or (n373,1'b0,n245,n374,1'b0);
and (n374,n375,n243,n244);
not (n375,n241);
and (n376,n234,n237,n97,n362);
and (n377,n249,n378);
and (n378,n235,n237,n97,n362);
or (n379,n235,n99,n97,n98);
or (n380,n229,n231);
or (n381,n218,n219,n220,n221);
nor (n382,n383,n385,n388);
not (n383,n384);
not (n385,n386);
xor (n386,n387,n384);
xor (n388,n389,n390);
and (n390,n387,n384);
and (n391,n319,n365);
and (n392,n393,n468);
wire s0n393,s1n393,notn393;
or (n393,s0n393,s1n393);
not(notn393,n453);
and (s0n393,notn393,n394);
and (s1n393,n453,n449);
xor (n394,n395,n411);
not (n395,n396);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n318);
and (s0n396,notn396,1'b0);
and (s1n396,n318,n397);
or (n397,n398,n401,n404,n408,1'b0,1'b0,1'b0,1'b0);
and (n398,n399,n118);
xnor (n399,n132,n400);
or (n400,n114,n295);
and (n401,n402,n296);
xnor (n402,n134,n403);
or (n403,n133,n294);
and (n404,n405,n303);
xnor (n405,n136,n406);
not (n406,n407);
and (n407,n301,n275);
and (n408,n409,n308);
xnor (n409,n140,n410);
or (n410,n147,n306);
and (n411,n412,n413);
not (n412,n107);
and (n413,n414,n431);
not (n414,n415);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n318);
and (s0n415,notn415,1'b0);
and (s1n415,n318,n416);
or (n416,n417,n419,n421,n423,n425,n428,1'b0,1'b0);
and (n417,n418,n118);
xnor (n418,n117,n114);
and (n419,n420,n296);
xnor (n420,n132,n295);
and (n421,n422,n303);
xnor (n422,n134,n302);
and (n423,n424,n308);
xnor (n424,n136,n307);
nor (n425,n426,n311);
not (n426,n427);
xnor (n427,n140,n316);
and (n428,n429,n430);
xnor (n429,n142,n145);
nor (n430,n119,n262,n280,n289);
not (n431,n432);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n318);
and (s0n432,notn432,1'b0);
and (s1n432,n318,n433);
or (n433,n434,n436,n438,n440,n442,n444,n446,1'b0);
and (n434,n435,n118);
xnor (n435,n115,n116);
and (n436,n437,n296);
xnor (n437,n111,n117);
and (n438,n439,n303);
xnor (n439,n133,n132);
and (n440,n441,n308);
xnor (n441,n135,n134);
and (n442,n443,n310);
xnor (n443,n147,n136);
and (n444,n445,n430);
xnor (n445,n141,n140);
and (n446,n447,n448);
xnor (n447,n151,n142);
nor (n448,n297,n261,n280,n289);
xor (n449,n396,n450);
and (n450,n107,n451);
and (n451,n415,n452);
and (n452,n432,n453);
wire s0n453,s1n453,notn453;
or (n453,s0n453,s1n453);
not(notn453,n318);
and (s0n453,notn453,1'b0);
and (s1n453,n318,n454);
or (n454,n455,n456,n458,n460,n462,n465,n466,1'b0);
and (n455,n130,n118);
and (n456,n457,n296);
not (n457,n117);
and (n458,n459,n303);
not (n459,n132);
and (n460,n461,n308);
not (n461,n134);
not (n462,n463);
nand (n463,n310,n464);
not (n464,n136);
and (n465,n139,n430);
and (n466,n467,n448);
not (n467,n142);
nor (n468,n469,n319);
not (n469,n365);
and (n470,n107,n471);
and (n471,n319,n469);
not (n472,n473);
nand (n473,n474,n498);
or (n474,n475,n482);
or (n475,n476,n481);
nor (n476,n477,n478,n480);
not (n478,n479);
and (n481,n477,n479,n480);
not (n482,n483);
nand (n483,n484,n492);
or (n484,1'b0,n485,n487,n491);
and (n485,n486,n391);
wire s0n486,s1n486,notn486;
or (n486,s0n486,s1n486);
not(notn486,n382);
and (s0n486,notn486,n415);
and (s1n486,n382,1'b0);
and (n487,n488,n468);
wire s0n488,s1n488,notn488;
or (n488,s0n488,s1n488);
not(notn488,n453);
and (s0n488,notn488,n489);
and (s1n488,n453,n490);
xor (n489,n412,n413);
xor (n490,n107,n451);
and (n491,n415,n471);
or (n492,1'b0,n493,n495,n497);
and (n493,n494,n391);
wire s0n494,s1n494,notn494;
or (n494,s0n494,s1n494);
not(notn494,n382);
and (s0n494,notn494,n432);
and (s1n494,n382,1'b0);
and (n495,n496,n468);
xor (n496,n414,n431);
and (n497,n432,n471);
nor (n498,n499,n522);
not (n499,n500);
or (n500,1'b0,n501,n503,n521);
and (n501,n502,n391);
wire s0n502,s1n502,notn502;
or (n502,s0n502,s1n502);
not(notn502,n382);
and (s0n502,notn502,n396);
and (s1n502,n382,1'b0);
and (n503,n504,n468);
wire s0n504,s1n504,notn504;
or (n504,s0n504,s1n504);
not(notn504,n453);
and (s0n504,notn504,n505);
and (s1n504,n453,n519);
xor (n505,n506,n518);
not (n506,n507);
wire s0n507,s1n507,notn507;
or (n507,s0n507,s1n507);
not(notn507,n318);
and (s0n507,notn507,1'b0);
and (s1n507,n318,n508);
or (n508,n509,n512,n515,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n509,n510,n118);
xnor (n510,n133,n511);
or (n511,n400,n132);
and (n512,n513,n296);
xnor (n513,n135,n514);
or (n514,n134,n403);
and (n515,n516,n303);
xnor (n516,n147,n517);
or (n517,n136,n406);
and (n518,n395,n411);
xor (n519,n507,n520);
and (n520,n396,n450);
and (n521,n396,n471);
nor (n522,n523,n526);
nand (n523,n524,n525);
not (n524,n484);
not (n525,n492);
or (n526,1'b0,n527,n545,n547);
and (n527,n528,n391);
wire s0n528,s1n528,notn528;
or (n528,s0n528,s1n528);
not(notn528,n382);
and (s0n528,notn528,n453);
and (s1n528,n382,n529);
not (n529,n530);
nor (n530,n453,n432,n415,n107,n396,n507,n531,n542);
wire s0n531,s1n531,notn531;
or (n531,s0n531,s1n531);
not(notn531,n318);
and (s0n531,notn531,1'b0);
and (s1n531,n318,n532);
or (n532,n533,n539,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n533,n534,n118);
nand (n534,n535,n537);
or (n535,n536,n461);
nor (n536,n400,n302);
nand (n537,n538,n301);
not (n538,n400);
and (n539,n540,n296);
xnor (n540,n136,n541);
or (n541,n135,n514);
wire s0n542,s1n542,notn542;
or (n542,s0n542,s1n542);
not(notn542,n318);
and (s0n542,notn542,1'b0);
and (s1n542,n318,n543);
and (n543,n544,n118);
xnor (n544,n135,n537);
and (n545,n546,n468);
xor (n546,n432,n453);
and (n547,n453,n471);
nand (n548,n549,n103);
or (n549,n550,n552);
not (n550,n551);
nor (n551,n500,n475);
not (n552,n553);
nand (n553,n554,n484);
nand (n554,n555,n525);
not (n555,n526);
nor (n556,n557,n591);
nand (n557,n558,n573,n582);
not (n558,n559);
or (n559,1'b0,n560,n562,n572);
and (n560,n561,n391);
wire s0n561,s1n561,notn561;
or (n561,s0n561,s1n561);
not(notn561,n382);
and (s0n561,notn561,n531);
and (s1n561,n382,1'b0);
and (n562,n563,n468);
wire s0n563,s1n563,notn563;
or (n563,s0n563,s1n563);
not(notn563,n453);
and (s0n563,notn563,n564);
and (s1n563,n453,n569);
xor (n564,n565,n566);
not (n565,n542);
and (n566,n567,n568);
not (n567,n531);
and (n568,n506,n518);
xor (n569,n542,n570);
and (n570,n531,n571);
and (n571,n507,n520);
and (n572,n531,n471);
not (n573,n574);
or (n574,1'b0,n575,n577,n581);
and (n575,n576,n391);
wire s0n576,s1n576,notn576;
or (n576,s0n576,s1n576);
not(notn576,n382);
and (s0n576,notn576,n507);
and (s1n576,n382,1'b0);
and (n577,n578,n468);
wire s0n578,s1n578,notn578;
or (n578,s0n578,s1n578);
not(notn578,n453);
and (s0n578,notn578,n579);
and (s1n578,n453,n580);
xor (n579,n567,n568);
xor (n580,n531,n571);
and (n581,n507,n471);
not (n582,n583);
or (n583,1'b0,n584,n586,n590);
and (n584,n585,n391);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n382);
and (s0n585,notn585,n542);
and (s1n585,n382,1'b0);
and (n586,n587,n468);
wire s0n587,s1n587,notn587;
or (n587,s0n587,s1n587);
not(notn587,n453);
and (s0n587,notn587,n588);
and (s1n587,n453,1'b0);
not (n588,n589);
and (n589,n565,n566);
and (n590,n542,n471);
not (n591,n236);
and (n592,n593,n67);
wire s0n593,s1n593,notn593;
or (n593,s0n593,s1n593);
not(notn593,n56);
and (s0n593,notn593,n594);
and (s1n593,n56,n595);
or (n595,n596,n598,n600,n602);
and (n596,n597,n44);
and (n598,n599,n49);
and (n600,n601,n53);
and (n602,n594,n55);
and (n603,n604,n72);
wire s0n604,s1n604,notn604;
or (n604,s0n604,s1n604);
not(notn604,n56);
and (s0n604,notn604,n605);
and (s1n604,n56,n606);
or (n606,n607,n609,n611,n613);
and (n607,n608,n44);
and (n609,n610,n49);
and (n611,n612,n53);
and (n613,n605,n55);
and (n614,n615,n75);
wire s0n615,s1n615,notn615;
or (n615,s0n615,s1n615);
not(notn615,n56);
and (s0n615,notn615,n616);
and (s1n615,n56,n617);
or (n617,n618,n620,n622,n624);
and (n618,n619,n44);
and (n620,n621,n49);
and (n622,n623,n53);
and (n624,n616,n55);
and (n626,n627,n76);
not (n627,n90);
wire s0n628,s1n628,notn628;
or (n628,s0n628,s1n628);
not(notn628,n625);
and (s0n628,notn628,n629);
and (s1n628,n625,n616);
wire s0n629,s1n629,notn629;
or (n629,s0n629,s1n629);
not(notn629,n56);
and (s0n629,notn629,n630);
and (s1n629,n56,n641);
or (n630,n631,n633,n635,n638);
and (n631,n40,n632);
and (n632,n85,n81);
and (n633,n594,n634);
and (n634,n84,n81);
and (n635,n605,n636);
not (n636,n637);
or (n637,n81,n84);
and (n638,n616,n639);
not (n639,n640);
or (n640,n85,n81);
or (n641,1'b0,n642,n645,n647,n650,n652,n654,n656,n658,n660,n662,n664,n666,n668,n670,n672,n674);
and (n642,n43,n643);
and (n643,n63,n64,n85,n81,n644);
not (n644,n76);
and (n645,n48,n646);
and (n646,n69,n64,n85,n81,n644);
and (n647,n52,n648);
and (n648,n63,n649,n85,n81,n644);
not (n649,n64);
and (n650,n40,n651);
and (n651,n69,n649,n85,n81,n644);
and (n652,n597,n653);
and (n653,n63,n64,n84,n81,n644);
and (n654,n599,n655);
and (n655,n69,n64,n84,n81,n644);
and (n656,n601,n657);
and (n657,n63,n649,n84,n81,n644);
and (n658,n594,n659);
and (n659,n69,n649,n84,n81,n644);
and (n660,n608,n661);
nor (n661,n69,n649,n84,n81,n76);
and (n662,n610,n663);
nor (n663,n63,n649,n84,n81,n76);
and (n664,n612,n665);
nor (n665,n69,n64,n84,n81,n76);
and (n666,n605,n667);
nor (n667,n63,n64,n84,n81,n76);
and (n668,n619,n669);
nor (n669,n69,n649,n85,n81,n76);
and (n670,n621,n671);
nor (n671,n63,n649,n85,n81,n76);
and (n672,n623,n673);
nor (n673,n69,n64,n85,n81,n76);
and (n674,n616,n675);
nor (n675,n63,n64,n85,n81,n76);
and (n676,n627,n644);
wire s0n677,s1n677,notn677;
or (n677,s0n677,s1n677);
not(notn677,n676);
and (s0n677,notn677,1'b0);
and (s1n677,n676,n678);
wire s0n678,s1n678,notn678;
or (n678,s0n678,s1n678);
not(notn678,n676);
and (s0n678,notn678,n679);
and (s1n678,n676,n726);
wire s0n679,s1n679,notn679;
or (n679,s0n679,s1n679);
not(notn679,n626);
and (s0n679,notn679,1'b0);
and (s1n679,n626,n680);
wire s0n680,s1n680,notn680;
or (n680,s0n680,s1n680);
not(notn680,n625);
and (s0n680,notn680,n681);
and (s1n680,n625,n717);
or (n681,n682,n693,n704,n715);
and (n682,n683,n62);
wire s0n683,s1n683,notn683;
or (n683,s0n683,s1n683);
not(notn683,n56);
and (s0n683,notn683,n684);
and (s1n683,n56,n685);
or (n685,n686,n688,n690,n692);
and (n686,n687,n44);
and (n688,n689,n49);
and (n690,n691,n53);
and (n692,n684,n55);
and (n693,n694,n67);
wire s0n694,s1n694,notn694;
or (n694,s0n694,s1n694);
not(notn694,n56);
and (s0n694,notn694,n695);
and (s1n694,n56,n696);
or (n696,n697,n699,n701,n703);
and (n697,n698,n44);
and (n699,n700,n49);
and (n701,n702,n53);
and (n703,n695,n55);
and (n704,n705,n72);
wire s0n705,s1n705,notn705;
or (n705,s0n705,s1n705);
not(notn705,n56);
and (s0n705,notn705,n706);
and (s1n705,n56,n707);
or (n707,n708,n710,n712,n714);
and (n708,n709,n44);
and (n710,n711,n49);
and (n712,n713,n53);
and (n714,n706,n55);
and (n715,n716,n75);
wire s0n716,s1n716,notn716;
or (n716,s0n716,s1n716);
not(notn716,n56);
and (s0n716,notn716,n717);
and (s1n716,n56,n718);
or (n718,n719,n721,n723,n725);
and (n719,n720,n44);
and (n721,n722,n49);
and (n723,n724,n53);
and (n725,n717,n55);
wire s0n726,s1n726,notn726;
or (n726,s0n726,s1n726);
not(notn726,n625);
and (s0n726,notn726,n727);
and (s1n726,n625,n717);
wire s0n727,s1n727,notn727;
or (n727,s0n727,s1n727);
not(notn727,n56);
and (s0n727,notn727,n728);
and (s1n727,n56,n733);
or (n728,n729,n730,n731,n732);
and (n729,n684,n632);
and (n730,n695,n634);
and (n731,n706,n636);
and (n732,n717,n639);
or (n733,1'b0,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749);
and (n734,n687,n643);
and (n735,n689,n646);
and (n736,n691,n648);
and (n737,n684,n651);
and (n738,n698,n653);
and (n739,n700,n655);
and (n740,n702,n657);
and (n741,n695,n659);
and (n742,n709,n661);
and (n743,n711,n663);
and (n744,n713,n665);
and (n745,n706,n667);
and (n746,n720,n669);
and (n747,n722,n671);
and (n748,n724,n673);
and (n749,n717,n675);
not (n750,n751);
wire s0n751,s1n751,notn751;
or (n751,s0n751,s1n751);
not(notn751,n676);
and (s0n751,notn751,1'b0);
and (s1n751,n676,n752);
wire s0n752,s1n752,notn752;
or (n752,s0n752,s1n752);
not(notn752,n676);
and (s0n752,notn752,n753);
and (s1n752,n676,n800);
wire s0n753,s1n753,notn753;
or (n753,s0n753,s1n753);
not(notn753,n626);
and (s0n753,notn753,1'b0);
and (s1n753,n626,n754);
wire s0n754,s1n754,notn754;
or (n754,s0n754,s1n754);
not(notn754,n625);
and (s0n754,notn754,n755);
and (s1n754,n625,n791);
or (n755,n756,n767,n778,n789);
and (n756,n757,n62);
wire s0n757,s1n757,notn757;
or (n757,s0n757,s1n757);
not(notn757,n56);
and (s0n757,notn757,n758);
and (s1n757,n56,n759);
or (n759,n760,n762,n764,n766);
and (n760,n761,n44);
and (n762,n763,n49);
and (n764,n765,n53);
and (n766,n758,n55);
and (n767,n768,n67);
wire s0n768,s1n768,notn768;
or (n768,s0n768,s1n768);
not(notn768,n56);
and (s0n768,notn768,n769);
and (s1n768,n56,n770);
or (n770,n771,n773,n775,n777);
and (n771,n772,n44);
and (n773,n774,n49);
and (n775,n776,n53);
and (n777,n769,n55);
and (n778,n779,n72);
wire s0n779,s1n779,notn779;
or (n779,s0n779,s1n779);
not(notn779,n56);
and (s0n779,notn779,n780);
and (s1n779,n56,n781);
or (n781,n782,n784,n786,n788);
and (n782,n783,n44);
and (n784,n785,n49);
and (n786,n787,n53);
and (n788,n780,n55);
and (n789,n790,n75);
wire s0n790,s1n790,notn790;
or (n790,s0n790,s1n790);
not(notn790,n56);
and (s0n790,notn790,n791);
and (s1n790,n56,n792);
or (n792,n793,n795,n797,n799);
and (n793,n794,n44);
and (n795,n796,n49);
and (n797,n798,n53);
and (n799,n791,n55);
wire s0n800,s1n800,notn800;
or (n800,s0n800,s1n800);
not(notn800,n625);
and (s0n800,notn800,n801);
and (s1n800,n625,n791);
wire s0n801,s1n801,notn801;
or (n801,s0n801,s1n801);
not(notn801,n56);
and (s0n801,notn801,n802);
and (s1n801,n56,n807);
or (n802,n803,n804,n805,n806);
and (n803,n758,n632);
and (n804,n769,n634);
and (n805,n780,n636);
and (n806,n791,n639);
or (n807,1'b0,n808,n809,n810,n811,n812,n813,n814,n815,n816,n817,n818,n819,n820,n821,n822,n823);
and (n808,n761,n643);
and (n809,n763,n646);
and (n810,n765,n648);
and (n811,n758,n651);
and (n812,n772,n653);
and (n813,n774,n655);
and (n814,n776,n657);
and (n815,n769,n659);
and (n816,n783,n661);
and (n817,n785,n663);
and (n818,n787,n665);
and (n819,n780,n667);
and (n820,n794,n669);
and (n821,n796,n671);
and (n822,n798,n673);
and (n823,n791,n675);
wire s0n824,s1n824,notn824;
or (n824,s0n824,s1n824);
not(notn824,n676);
and (s0n824,notn824,1'b0);
and (s1n824,n676,n825);
wire s0n825,s1n825,notn825;
or (n825,s0n825,s1n825);
not(notn825,n676);
and (s0n825,notn825,n826);
and (s1n825,n676,n873);
wire s0n826,s1n826,notn826;
or (n826,s0n826,s1n826);
not(notn826,n626);
and (s0n826,notn826,1'b0);
and (s1n826,n626,n827);
wire s0n827,s1n827,notn827;
or (n827,s0n827,s1n827);
not(notn827,n625);
and (s0n827,notn827,n828);
and (s1n827,n625,n864);
or (n828,n829,n840,n851,n862);
and (n829,n830,n62);
wire s0n830,s1n830,notn830;
or (n830,s0n830,s1n830);
not(notn830,n56);
and (s0n830,notn830,n831);
and (s1n830,n56,n832);
or (n832,n833,n835,n837,n839);
and (n833,n834,n44);
and (n835,n836,n49);
and (n837,n838,n53);
and (n839,n831,n55);
and (n840,n841,n67);
wire s0n841,s1n841,notn841;
or (n841,s0n841,s1n841);
not(notn841,n56);
and (s0n841,notn841,n842);
and (s1n841,n56,n843);
or (n843,n844,n846,n848,n850);
and (n844,n845,n44);
and (n846,n847,n49);
and (n848,n849,n53);
and (n850,n842,n55);
and (n851,n852,n72);
wire s0n852,s1n852,notn852;
or (n852,s0n852,s1n852);
not(notn852,n56);
and (s0n852,notn852,n853);
and (s1n852,n56,n854);
or (n854,n855,n857,n859,n861);
and (n855,n856,n44);
and (n857,n858,n49);
and (n859,n860,n53);
and (n861,n853,n55);
and (n862,n863,n75);
wire s0n863,s1n863,notn863;
or (n863,s0n863,s1n863);
not(notn863,n56);
and (s0n863,notn863,n864);
and (s1n863,n56,n865);
or (n865,n866,n868,n870,n872);
and (n866,n867,n44);
and (n868,n869,n49);
and (n870,n871,n53);
and (n872,n864,n55);
wire s0n873,s1n873,notn873;
or (n873,s0n873,s1n873);
not(notn873,n625);
and (s0n873,notn873,n874);
and (s1n873,n625,n864);
wire s0n874,s1n874,notn874;
or (n874,s0n874,s1n874);
not(notn874,n56);
and (s0n874,notn874,n875);
and (s1n874,n56,n880);
or (n875,n876,n877,n878,n879);
and (n876,n831,n632);
and (n877,n842,n634);
and (n878,n853,n636);
and (n879,n864,n639);
or (n880,1'b0,n881,n882,n883,n884,n885,n886,n887,n888,n889,n890,n891,n892,n893,n894,n895,n896);
and (n881,n834,n643);
and (n882,n836,n646);
and (n883,n838,n648);
and (n884,n831,n651);
and (n885,n845,n653);
and (n886,n847,n655);
and (n887,n849,n657);
and (n888,n842,n659);
and (n889,n856,n661);
and (n890,n858,n663);
and (n891,n860,n665);
and (n892,n853,n667);
and (n893,n867,n669);
and (n894,n869,n671);
and (n895,n871,n673);
and (n896,n864,n675);
or (n897,n898,n910);
or (n898,n899,n909);
or (n899,n900,n906);
nor (n900,n901,n902,n903,n905);
not (n903,n904);
nor (n906,n907,n908,n904,n905);
not (n907,n901);
not (n908,n902);
nor (n909,n901,n908,n904,n905);
nor (n910,n907,n902,n904,n905);
and (n911,n912,n897);
or (n912,n913,n915);
nor (n913,n32,n677,n751,n914);
not (n914,n824);
and (n915,n33,n677,n750,n824);
and (n916,n917,n676,n918);
and (n917,n751,n32,n677);
nor (n918,n907,n905);
wire s0n919,s1n919,notn919;
or (n919,s0n919,s1n919);
not(notn919,n28);
and (s0n919,notn919,1'b0);
and (s1n919,n28,n920);
or (n921,n922,n927,n1991);
and (n922,n923,n925);
wire s0n923,s1n923,notn923;
or (n923,s0n923,s1n923);
not(notn923,n28);
and (s0n923,notn923,1'b0);
and (s1n923,n28,n924);
wire s0n925,s1n925,notn925;
or (n925,s0n925,s1n925);
not(notn925,n28);
and (s0n925,notn925,1'b0);
and (s1n925,n28,n926);
and (n927,n925,n928);
or (n928,n929,n934,n1990);
and (n929,n930,n932);
wire s0n930,s1n930,notn930;
or (n930,s0n930,s1n930);
not(notn930,n28);
and (s0n930,notn930,1'b0);
and (s1n930,n28,n931);
wire s0n932,s1n932,notn932;
or (n932,s0n932,s1n932);
not(notn932,n28);
and (s0n932,notn932,1'b0);
and (s1n932,n28,n933);
and (n934,n932,n935);
or (n935,n936,n1129,n1989);
and (n936,n937,n1058);
wire s0n937,s1n937,notn937;
or (n937,s0n937,s1n937);
not(notn937,n28);
and (s0n937,notn937,n938);
and (s1n937,n28,n1057);
nand (n938,n939,n1003,n1015,n1027);
nor (n939,n940,n998);
nand (n940,n941,n988,n993);
nor (n941,n942,n976);
and (n942,n943,n975);
and (n943,n944,n970);
or (n944,n945,n962);
not (n945,n946);
nand (n946,n947,n957,n914);
nand (n947,n948,n955);
or (n948,n949,n950);
not (n949,n910);
not (n950,n951);
nand (n951,n952,n953);
nand (n952,n750,n914,n677);
nand (n953,n954,n33);
or (n954,n914,n751);
not (n955,n956);
and (n956,n751,n32,n677,n909);
not (n957,n958);
nand (n958,n959,n961);
or (n959,n960,n950);
not (n960,n909);
nand (n961,n751,n32,n677,n900);
not (n962,n963);
nand (n963,n964,n958,n966,n824);
and (n964,n965,n948);
nand (n965,n951,n906);
and (n966,n955,n967);
nand (n967,n32,n751,n677,n968);
and (n968,n907,n902,n904,n969);
not (n969,n905);
not (n970,n971);
nand (n971,n972,n973,n676);
or (n972,n56,n649);
not (n973,n974);
nor (n974,n69,n56);
and (n976,n977,n987);
not (n977,n978);
nand (n978,n979,n970);
not (n979,n980);
nand (n980,n981,n914);
nand (n981,n982,n984);
or (n982,n983,n950);
not (n983,n900);
not (n984,n985);
and (n985,n917,n986);
nor (n986,n901,n902,n904,n969);
nand (n988,n989,n992);
and (n989,n944,n990);
and (n990,n974,n991);
and (n991,n676,n649);
nand (n993,n994,n997);
and (n994,n995,n990);
and (n995,n996,n947,n957,n824);
and (n996,n965,n967);
and (n998,n999,n1002);
nand (n999,n1000,n1001);
nand (n1000,n995,n970);
nand (n1001,n979,n990);
nor (n1003,n1004,n1011);
and (n1004,n1005,n1010);
not (n1005,n1006);
nand (n1006,n1007,n990);
nand (n1007,n1008,n1009);
or (n1008,n914,n996);
nand (n1009,n964,n958,n966,n914);
nor (n1011,n1012,n1014);
not (n1012,n1013);
nand (n1014,n1007,n970);
nor (n1015,n1016,n1023);
and (n1016,n1017,n1022);
not (n1017,n1018);
nand (n1018,n1019,n990);
nand (n1019,n1020,n1021);
or (n1020,n824,n996);
nand (n1021,n981,n824);
and (n1023,n1024,n1026);
not (n1024,n1025);
nand (n1025,n1019,n970);
nor (n1027,n1028,n1044);
and (n1028,n1029,n1041);
nand (n1029,n1030,n1035,n1037,n1039);
nor (n1030,n1031,n1033);
and (n1031,n995,n1032);
and (n1033,n979,n1034);
nand (n1035,n944,n1036);
nand (n1037,n1007,n1038);
nand (n1039,n1019,n1040);
and (n1041,n1042,n1043);
and (n1042,n676,n64);
nor (n1043,n56,n63);
and (n1044,n1045,n1056);
nand (n1045,n1046,n1050,n1052,n1054);
nor (n1046,n1047,n1049);
and (n1047,n995,n1048);
and (n1049,n979,n1032);
nand (n1050,n944,n1051);
nand (n1052,n1007,n1053);
nand (n1054,n1019,n1055);
and (n1056,n1042,n974);
wire s0n1058,s1n1058,notn1058;
or (n1058,s0n1058,s1n1058);
not(notn1058,n28);
and (s0n1058,notn1058,n1059);
and (s1n1058,n28,n1128);
or (n1059,1'b0,n1060,n1083,n1097,n1110);
and (n1060,n1061,n1056);
or (n1061,1'b0,n1062,n1073,n1076,n1080);
and (n1062,n1063,n947);
wire s0n1063,s1n1063,notn1063;
or (n1063,s0n1063,s1n1063);
not(notn1063,n1066);
and (s0n1063,notn1063,n1064);
and (s1n1063,n1066,n1065);
or (n1066,n1067,n1071);
or (n1067,n1068,n1070);
and (n1068,n33,n1069,n751,n824);
not (n1069,n677);
and (n1070,n33,n677,n751,n824);
not (n1071,n1072);
nand (n1072,n32,n677,n751,n824);
and (n1073,n1074,n958);
wire s0n1074,s1n1074,notn1074;
or (n1074,s0n1074,s1n1074);
not(notn1074,n1066);
and (s0n1074,notn1074,n1075);
and (s1n1074,n1066,n1064);
and (n1076,n1077,n1079);
wire s0n1077,s1n1077,notn1077;
or (n1077,s0n1077,s1n1077);
not(notn1077,n1066);
and (s0n1077,notn1077,n1078);
and (s1n1077,n1066,n1075);
not (n1079,n996);
and (n1080,n1081,n981);
wire s0n1081,s1n1081,notn1081;
or (n1081,s0n1081,s1n1081);
not(notn1081,n1066);
and (s0n1081,notn1081,n1082);
and (s1n1081,n1066,n1078);
and (n1083,n1084,n1041);
or (n1084,1'b0,n1085,n1088,n1091,n1094);
and (n1085,n1086,n947);
wire s0n1086,s1n1086,notn1086;
or (n1086,s0n1086,s1n1086);
not(notn1086,n1066);
and (s0n1086,notn1086,n1087);
and (s1n1086,n1066,n1082);
and (n1088,n1089,n958);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n1066);
and (s0n1089,notn1089,n1090);
and (s1n1089,n1066,n1087);
and (n1091,n1092,n1079);
wire s0n1092,s1n1092,notn1092;
or (n1092,s0n1092,s1n1092);
not(notn1092,n1066);
and (s0n1092,notn1092,n1093);
and (s1n1092,n1066,n1090);
and (n1094,n1095,n981);
wire s0n1095,s1n1095,notn1095;
or (n1095,s0n1095,s1n1095);
not(notn1095,n1066);
and (s0n1095,notn1095,n1096);
and (s1n1095,n1066,n1093);
and (n1097,n1098,n990);
nand (n1098,n1099,n1104,n1106,n1108);
nor (n1099,n1100,n1102);
and (n1100,n995,n1101);
and (n1102,n979,n1103);
nand (n1104,n944,n1105);
nand (n1106,n1007,n1107);
nand (n1108,n1019,n1109);
and (n1110,n1111,n970);
nand (n1111,n1112,n1117);
nor (n1112,n1113,n1115);
and (n1113,n1007,n1114);
and (n1115,n1019,n1116);
nor (n1117,n1118,n1124);
nand (n1118,n1119,n1122);
or (n1119,n1120,n1121);
not (n1120,n1103);
not (n1121,n995);
nand (n1122,n979,n1123);
nor (n1124,n1125,n1127);
not (n1125,n1126);
not (n1127,n944);
and (n1129,n1058,n1130);
or (n1130,n1131,n1254,n1988);
and (n1131,n1132,n1185);
wire s0n1132,s1n1132,notn1132;
or (n1132,s0n1132,s1n1132);
not(notn1132,n28);
and (s0n1132,notn1132,n1133);
and (s1n1132,n28,n1184);
nand (n1133,n1134,n1147,n1173,n1179);
nor (n1134,n1135,n1145);
nand (n1135,n1136,n1141,n1143);
nor (n1136,n1137,n1139);
and (n1137,n943,n1138);
and (n1139,n977,n1140);
nand (n1141,n989,n1142);
nand (n1143,n994,n1144);
and (n1145,n999,n1146);
nor (n1147,n1148,n1161);
and (n1148,n1149,n1041);
nand (n1149,n1150,n1152,n1154,n1159);
nand (n1150,n1007,n1151);
nand (n1152,n1019,n1153);
nor (n1154,n1155,n1157);
and (n1155,n995,n1156);
and (n1157,n979,n1158);
nand (n1159,n944,n1160);
and (n1161,n1162,n1056);
nand (n1162,n1163,n1165,n1167,n1171);
nand (n1163,n1007,n1164);
nand (n1165,n1019,n1166);
nor (n1167,n1168,n1170);
and (n1168,n995,n1169);
and (n1170,n979,n1156);
nand (n1171,n944,n1172);
nor (n1173,n1174,n1177);
and (n1174,n1175,n1176);
not (n1175,n1014);
and (n1177,n1005,n1178);
nor (n1179,n1180,n1182);
and (n1180,n1024,n1181);
and (n1182,n1017,n1183);
wire s0n1185,s1n1185,notn1185;
or (n1185,s0n1185,s1n1185);
not(notn1185,n28);
and (s0n1185,notn1185,n1186);
and (s1n1185,n28,n1253);
nand (n1186,n1187,n1210,n1236,n1244);
nor (n1187,n1188,n1193);
and (n1188,n1189,n1192);
nand (n1189,n1190,n1191);
nand (n1190,n995,n1041);
nand (n1191,n979,n1056);
nand (n1193,n1194,n1202,n1206);
nor (n1194,n1195,n1198);
and (n1195,n1196,n1197);
and (n1196,n944,n1041);
and (n1198,n1199,n1201);
not (n1199,n1200);
nand (n1200,n979,n1041);
nand (n1202,n1203,n1205);
not (n1203,n1204);
nand (n1204,n944,n1056);
nand (n1206,n1207,n1209);
not (n1207,n1208);
nand (n1208,n995,n1056);
nor (n1210,n1211,n1224);
and (n1211,n1212,n970);
nand (n1212,n1213,n1215,n1217,n1222);
nand (n1213,n1007,n1214);
nand (n1215,n1019,n1216);
nor (n1217,n1218,n1220);
and (n1218,n995,n1219);
and (n1220,n979,n1221);
nand (n1222,n944,n1223);
and (n1224,n1225,n990);
nand (n1225,n1226,n1228,n1230,n1234);
nand (n1226,n1007,n1227);
nand (n1228,n1019,n1229);
nor (n1230,n1231,n1233);
and (n1231,n995,n1232);
and (n1233,n979,n1219);
nand (n1234,n944,n1235);
nor (n1236,n1237,n1240);
and (n1237,n1238,n1239);
and (n1238,n1007,n1041);
and (n1240,n1241,n1243);
not (n1241,n1242);
nand (n1242,n1007,n1056);
nor (n1244,n1245,n1249);
and (n1245,n1246,n1248);
not (n1246,n1247);
nand (n1247,n1019,n1041);
and (n1249,n1250,n1252);
not (n1250,n1251);
nand (n1251,n1019,n1056);
and (n1254,n1185,n1255);
or (n1255,n1256,n1378,n1987);
and (n1256,n1257,n1314);
wire s0n1257,s1n1257,notn1257;
or (n1257,s0n1257,s1n1257);
not(notn1257,n28);
and (s0n1257,notn1257,n1258);
and (s1n1257,n28,n1313);
or (n1258,1'b0,n1259,n1272,n1284,n1299);
and (n1259,n1260,n1056);
nand (n1260,n1261,n1266,n1268,n1270);
nor (n1261,n1262,n1264);
and (n1262,n995,n1263);
and (n1264,n979,n1265);
nand (n1266,n944,n1267);
nand (n1268,n1007,n1269);
nand (n1270,n1019,n1271);
and (n1272,n1273,n1041);
nand (n1273,n1274,n1278,n1280,n1282);
nor (n1274,n1275,n1276);
and (n1275,n995,n1265);
and (n1276,n979,n1277);
nand (n1278,n944,n1279);
nand (n1280,n1007,n1281);
nand (n1282,n1019,n1283);
and (n1284,n1285,n990);
or (n1285,1'b0,n1286,n1290,n1293,n1296);
and (n1286,n1287,n947);
wire s0n1287,s1n1287,notn1287;
or (n1287,s0n1287,s1n1287);
not(notn1287,n1066);
and (s0n1287,notn1287,n1288);
and (s1n1287,n1066,n1289);
and (n1290,n1291,n958);
wire s0n1291,s1n1291,notn1291;
or (n1291,s0n1291,s1n1291);
not(notn1291,n1066);
and (s0n1291,notn1291,n1292);
and (s1n1291,n1066,n1288);
and (n1293,n1294,n1079);
wire s0n1294,s1n1294,notn1294;
or (n1294,s0n1294,s1n1294);
not(notn1294,n1066);
and (s0n1294,notn1294,n1295);
and (s1n1294,n1066,n1292);
and (n1296,n1297,n981);
wire s0n1297,s1n1297,notn1297;
or (n1297,s0n1297,s1n1297);
not(notn1297,n1066);
and (s0n1297,notn1297,n1298);
and (s1n1297,n1066,n1295);
and (n1299,n1300,n970);
or (n1300,1'b0,n1301,n1304,n1307,n1310);
and (n1301,n1302,n947);
wire s0n1302,s1n1302,notn1302;
or (n1302,s0n1302,s1n1302);
not(notn1302,n1066);
and (s0n1302,notn1302,n1303);
and (s1n1302,n1066,n1298);
and (n1304,n1305,n958);
wire s0n1305,s1n1305,notn1305;
or (n1305,s0n1305,s1n1305);
not(notn1305,n1066);
and (s0n1305,notn1305,n1306);
and (s1n1305,n1066,n1303);
and (n1307,n1308,n1079);
wire s0n1308,s1n1308,notn1308;
or (n1308,s0n1308,s1n1308);
not(notn1308,n1066);
and (s0n1308,notn1308,n1309);
and (s1n1308,n1066,n1306);
and (n1310,n1311,n981);
wire s0n1311,s1n1311,notn1311;
or (n1311,s0n1311,s1n1311);
not(notn1311,n1066);
and (s0n1311,notn1311,n1312);
and (s1n1311,n1066,n1309);
wire s0n1314,s1n1314,notn1314;
or (n1314,s0n1314,s1n1314);
not(notn1314,n28);
and (s0n1314,notn1314,n1315);
and (s1n1314,n28,n1377);
or (n1315,1'b0,n1316,n1331,n1345,n1361);
and (n1316,n1317,n1056);
or (n1317,1'b0,n1318,n1322,n1325,n1328);
and (n1318,n1319,n947);
wire s0n1319,s1n1319,notn1319;
or (n1319,s0n1319,s1n1319);
not(notn1319,n1066);
and (s0n1319,notn1319,n1320);
and (s1n1319,n1066,n1321);
and (n1322,n1323,n958);
wire s0n1323,s1n1323,notn1323;
or (n1323,s0n1323,s1n1323);
not(notn1323,n1066);
and (s0n1323,notn1323,n1324);
and (s1n1323,n1066,n1320);
and (n1325,n1326,n1079);
wire s0n1326,s1n1326,notn1326;
or (n1326,s0n1326,s1n1326);
not(notn1326,n1066);
and (s0n1326,notn1326,n1327);
and (s1n1326,n1066,n1324);
and (n1328,n1329,n981);
wire s0n1329,s1n1329,notn1329;
or (n1329,s0n1329,s1n1329);
not(notn1329,n1066);
and (s0n1329,notn1329,n1330);
and (s1n1329,n1066,n1327);
and (n1331,n1332,n1041);
or (n1332,1'b0,n1333,n1336,n1339,n1342);
and (n1333,n1334,n947);
wire s0n1334,s1n1334,notn1334;
or (n1334,s0n1334,s1n1334);
not(notn1334,n1066);
and (s0n1334,notn1334,n1335);
and (s1n1334,n1066,n1330);
and (n1336,n1337,n958);
wire s0n1337,s1n1337,notn1337;
or (n1337,s0n1337,s1n1337);
not(notn1337,n1066);
and (s0n1337,notn1337,n1338);
and (s1n1337,n1066,n1335);
and (n1339,n1340,n1079);
wire s0n1340,s1n1340,notn1340;
or (n1340,s0n1340,s1n1340);
not(notn1340,n1066);
and (s0n1340,notn1340,n1341);
and (s1n1340,n1066,n1338);
and (n1342,n1343,n981);
wire s0n1343,s1n1343,notn1343;
or (n1343,s0n1343,s1n1343);
not(notn1343,n1066);
and (s0n1343,notn1343,n1344);
and (s1n1343,n1066,n1341);
and (n1345,n1346,n990);
nand (n1346,n1347,n1352);
nor (n1347,n1348,n1350);
and (n1348,n1007,n1349);
and (n1350,n1019,n1351);
nor (n1352,n1353,n1355);
and (n1353,n944,n1354);
nand (n1355,n1356,n1359);
or (n1356,n1357,n1121);
not (n1357,n1358);
nand (n1359,n979,n1360);
and (n1361,n1362,n970);
nand (n1362,n1363,n1368);
nor (n1363,n1364,n1366);
and (n1364,n1007,n1365);
and (n1366,n1019,n1367);
nor (n1368,n1369,n1374);
nand (n1369,n1370,n1372);
or (n1370,n1371,n1121);
not (n1371,n1360);
nand (n1372,n979,n1373);
nor (n1374,n1375,n1127);
not (n1375,n1376);
and (n1378,n1314,n1379);
or (n1379,n1380,n1493,n1986);
and (n1380,n1381,n1433);
wire s0n1381,s1n1381,notn1381;
or (n1381,s0n1381,s1n1381);
not(notn1381,n28);
and (s0n1381,notn1381,n1382);
and (s1n1381,n28,n1432);
nand (n1382,n1383,n1396,n1401,n1427);
nor (n1383,n1384,n1394);
nand (n1384,n1385,n1390,n1392);
nor (n1385,n1386,n1388);
and (n1386,n943,n1387);
and (n1388,n977,n1389);
nand (n1390,n989,n1391);
nand (n1392,n994,n1393);
and (n1394,n999,n1395);
nor (n1396,n1397,n1399);
and (n1397,n1175,n1398);
and (n1399,n1005,n1400);
nor (n1401,n1402,n1415);
and (n1402,n1403,n1041);
nand (n1403,n1404,n1409,n1411,n1413);
nor (n1404,n1405,n1407);
and (n1405,n995,n1406);
and (n1407,n979,n1408);
nand (n1409,n944,n1410);
nand (n1411,n1007,n1412);
nand (n1413,n1019,n1414);
and (n1415,n1416,n1056);
nand (n1416,n1417,n1421,n1423,n1425);
nor (n1417,n1418,n1420);
and (n1418,n995,n1419);
and (n1420,n979,n1406);
nand (n1421,n944,n1422);
nand (n1423,n1007,n1424);
nand (n1425,n1019,n1426);
nor (n1427,n1428,n1430);
and (n1428,n1024,n1429);
and (n1430,n1017,n1431);
wire s0n1433,s1n1433,notn1433;
or (n1433,s0n1433,s1n1433);
not(notn1433,n28);
and (s0n1433,notn1433,n1434);
and (s1n1433,n28,n1492);
or (n1434,1'b0,n1435,n1450,n1464,n1477);
and (n1435,n1436,n1056);
or (n1436,1'b0,n1437,n1441,n1444,n1447);
and (n1437,n1438,n947);
wire s0n1438,s1n1438,notn1438;
or (n1438,s0n1438,s1n1438);
not(notn1438,n1066);
and (s0n1438,notn1438,n1439);
and (s1n1438,n1066,n1440);
and (n1441,n1442,n958);
wire s0n1442,s1n1442,notn1442;
or (n1442,s0n1442,s1n1442);
not(notn1442,n1066);
and (s0n1442,notn1442,n1443);
and (s1n1442,n1066,n1439);
and (n1444,n1445,n1079);
wire s0n1445,s1n1445,notn1445;
or (n1445,s0n1445,s1n1445);
not(notn1445,n1066);
and (s0n1445,notn1445,n1446);
and (s1n1445,n1066,n1443);
and (n1447,n1448,n981);
wire s0n1448,s1n1448,notn1448;
or (n1448,s0n1448,s1n1448);
not(notn1448,n1066);
and (s0n1448,notn1448,n1449);
and (s1n1448,n1066,n1446);
and (n1450,n1451,n1041);
or (n1451,1'b0,n1452,n1455,n1458,n1461);
and (n1452,n1453,n947);
wire s0n1453,s1n1453,notn1453;
or (n1453,s0n1453,s1n1453);
not(notn1453,n1066);
and (s0n1453,notn1453,n1454);
and (s1n1453,n1066,n1449);
and (n1455,n1456,n958);
wire s0n1456,s1n1456,notn1456;
or (n1456,s0n1456,s1n1456);
not(notn1456,n1066);
and (s0n1456,notn1456,n1457);
and (s1n1456,n1066,n1454);
and (n1458,n1459,n1079);
wire s0n1459,s1n1459,notn1459;
or (n1459,s0n1459,s1n1459);
not(notn1459,n1066);
and (s0n1459,notn1459,n1460);
and (s1n1459,n1066,n1457);
and (n1461,n1462,n981);
wire s0n1462,s1n1462,notn1462;
or (n1462,s0n1462,s1n1462);
not(notn1462,n1066);
and (s0n1462,notn1462,n1463);
and (s1n1462,n1066,n1460);
and (n1464,n1465,n990);
nand (n1465,n1466,n1471,n1473,n1475);
nor (n1466,n1467,n1469);
and (n1467,n979,n1468);
and (n1469,n995,n1470);
nand (n1471,n944,n1472);
nand (n1473,n1007,n1474);
nand (n1475,n1019,n1476);
and (n1477,n1478,n970);
nand (n1478,n1479,n1484);
nor (n1479,n1480,n1482);
and (n1480,n1007,n1481);
and (n1482,n1019,n1483);
nor (n1484,n1485,n1490);
nand (n1485,n1486,n1488);
or (n1486,n1487,n1121);
not (n1487,n1468);
nand (n1488,n979,n1489);
and (n1490,n944,n1491);
and (n1493,n1433,n1494);
or (n1494,n1495,n1617,n1985);
and (n1495,n1496,n1553);
wire s0n1496,s1n1496,notn1496;
or (n1496,s0n1496,s1n1496);
not(notn1496,n28);
and (s0n1496,notn1496,n1497);
and (s1n1496,n28,n1552);
or (n1497,1'b0,n1498,n1511,n1523,n1538);
and (n1498,n1499,n1056);
nand (n1499,n1500,n1505,n1507,n1509);
nor (n1500,n1501,n1503);
and (n1501,n995,n1502);
and (n1503,n979,n1504);
nand (n1505,n944,n1506);
nand (n1507,n1007,n1508);
nand (n1509,n1019,n1510);
and (n1511,n1512,n1041);
nand (n1512,n1513,n1517,n1519,n1521);
nor (n1513,n1514,n1515);
and (n1514,n995,n1504);
and (n1515,n979,n1516);
nand (n1517,n944,n1518);
nand (n1519,n1007,n1520);
nand (n1521,n1019,n1522);
and (n1523,n1524,n990);
or (n1524,1'b0,n1525,n1529,n1532,n1535);
and (n1525,n1526,n947);
wire s0n1526,s1n1526,notn1526;
or (n1526,s0n1526,s1n1526);
not(notn1526,n1066);
and (s0n1526,notn1526,n1527);
and (s1n1526,n1066,n1528);
and (n1529,n1530,n958);
wire s0n1530,s1n1530,notn1530;
or (n1530,s0n1530,s1n1530);
not(notn1530,n1066);
and (s0n1530,notn1530,n1531);
and (s1n1530,n1066,n1527);
and (n1532,n1533,n1079);
wire s0n1533,s1n1533,notn1533;
or (n1533,s0n1533,s1n1533);
not(notn1533,n1066);
and (s0n1533,notn1533,n1534);
and (s1n1533,n1066,n1531);
and (n1535,n1536,n981);
wire s0n1536,s1n1536,notn1536;
or (n1536,s0n1536,s1n1536);
not(notn1536,n1066);
and (s0n1536,notn1536,n1537);
and (s1n1536,n1066,n1534);
and (n1538,n1539,n970);
or (n1539,1'b0,n1540,n1543,n1546,n1549);
and (n1540,n1541,n947);
wire s0n1541,s1n1541,notn1541;
or (n1541,s0n1541,s1n1541);
not(notn1541,n1066);
and (s0n1541,notn1541,n1542);
and (s1n1541,n1066,n1537);
and (n1543,n1544,n958);
wire s0n1544,s1n1544,notn1544;
or (n1544,s0n1544,s1n1544);
not(notn1544,n1066);
and (s0n1544,notn1544,n1545);
and (s1n1544,n1066,n1542);
and (n1546,n1547,n1079);
wire s0n1547,s1n1547,notn1547;
or (n1547,s0n1547,s1n1547);
not(notn1547,n1066);
and (s0n1547,notn1547,n1548);
and (s1n1547,n1066,n1545);
and (n1549,n1550,n981);
wire s0n1550,s1n1550,notn1550;
or (n1550,s0n1550,s1n1550);
not(notn1550,n1066);
and (s0n1550,notn1550,n1551);
and (s1n1550,n1066,n1548);
wire s0n1553,s1n1553,notn1553;
or (n1553,s0n1553,s1n1553);
not(notn1553,n28);
and (s0n1553,notn1553,n1554);
and (s1n1553,n28,n1616);
or (n1554,1'b0,n1555,n1570,n1584,n1600);
and (n1555,n1556,n1056);
or (n1556,1'b0,n1557,n1561,n1564,n1567);
and (n1557,n1558,n947);
wire s0n1558,s1n1558,notn1558;
or (n1558,s0n1558,s1n1558);
not(notn1558,n1066);
and (s0n1558,notn1558,n1559);
and (s1n1558,n1066,n1560);
and (n1561,n1562,n958);
wire s0n1562,s1n1562,notn1562;
or (n1562,s0n1562,s1n1562);
not(notn1562,n1066);
and (s0n1562,notn1562,n1563);
and (s1n1562,n1066,n1559);
and (n1564,n1565,n1079);
wire s0n1565,s1n1565,notn1565;
or (n1565,s0n1565,s1n1565);
not(notn1565,n1066);
and (s0n1565,notn1565,n1566);
and (s1n1565,n1066,n1563);
and (n1567,n1568,n981);
wire s0n1568,s1n1568,notn1568;
or (n1568,s0n1568,s1n1568);
not(notn1568,n1066);
and (s0n1568,notn1568,n1569);
and (s1n1568,n1066,n1566);
and (n1570,n1571,n1041);
or (n1571,1'b0,n1572,n1575,n1578,n1581);
and (n1572,n1573,n947);
wire s0n1573,s1n1573,notn1573;
or (n1573,s0n1573,s1n1573);
not(notn1573,n1066);
and (s0n1573,notn1573,n1574);
and (s1n1573,n1066,n1569);
and (n1575,n1576,n958);
wire s0n1576,s1n1576,notn1576;
or (n1576,s0n1576,s1n1576);
not(notn1576,n1066);
and (s0n1576,notn1576,n1577);
and (s1n1576,n1066,n1574);
and (n1578,n1579,n1079);
wire s0n1579,s1n1579,notn1579;
or (n1579,s0n1579,s1n1579);
not(notn1579,n1066);
and (s0n1579,notn1579,n1580);
and (s1n1579,n1066,n1577);
and (n1581,n1582,n981);
wire s0n1582,s1n1582,notn1582;
or (n1582,s0n1582,s1n1582);
not(notn1582,n1066);
and (s0n1582,notn1582,n1583);
and (s1n1582,n1066,n1580);
and (n1584,n1585,n990);
nand (n1585,n1586,n1591);
nor (n1586,n1587,n1589);
and (n1587,n1007,n1588);
and (n1589,n1019,n1590);
nor (n1591,n1592,n1594);
and (n1592,n944,n1593);
nand (n1594,n1595,n1598);
or (n1595,n1596,n1121);
not (n1596,n1597);
nand (n1598,n979,n1599);
and (n1600,n1601,n970);
nand (n1601,n1602,n1607);
nor (n1602,n1603,n1605);
and (n1603,n1007,n1604);
and (n1605,n1019,n1606);
nor (n1607,n1608,n1613);
nand (n1608,n1609,n1611);
or (n1609,n1610,n1121);
not (n1610,n1599);
nand (n1611,n979,n1612);
nor (n1613,n1614,n1127);
not (n1614,n1615);
and (n1617,n1553,n1618);
or (n1618,n1619,n1740,n1984);
and (n1619,n1620,n1677);
wire s0n1620,s1n1620,notn1620;
or (n1620,s0n1620,s1n1620);
not(notn1620,n28);
and (s0n1620,notn1620,n1621);
and (s1n1620,n28,n1676);
or (n1621,1'b0,n1622,n1635,n1647,n1662);
and (n1622,n1623,n1056);
nand (n1623,n1624,n1629,n1631,n1633);
nor (n1624,n1625,n1627);
and (n1625,n995,n1626);
and (n1627,n979,n1628);
nand (n1629,n944,n1630);
nand (n1631,n1007,n1632);
nand (n1633,n1019,n1634);
and (n1635,n1636,n1041);
nand (n1636,n1637,n1641,n1643,n1645);
nor (n1637,n1638,n1639);
and (n1638,n995,n1628);
and (n1639,n979,n1640);
nand (n1641,n944,n1642);
nand (n1643,n1007,n1644);
nand (n1645,n1019,n1646);
and (n1647,n1648,n990);
or (n1648,1'b0,n1649,n1653,n1656,n1659);
and (n1649,n1650,n947);
wire s0n1650,s1n1650,notn1650;
or (n1650,s0n1650,s1n1650);
not(notn1650,n1066);
and (s0n1650,notn1650,n1651);
and (s1n1650,n1066,n1652);
and (n1653,n1654,n958);
wire s0n1654,s1n1654,notn1654;
or (n1654,s0n1654,s1n1654);
not(notn1654,n1066);
and (s0n1654,notn1654,n1655);
and (s1n1654,n1066,n1651);
and (n1656,n1657,n1079);
wire s0n1657,s1n1657,notn1657;
or (n1657,s0n1657,s1n1657);
not(notn1657,n1066);
and (s0n1657,notn1657,n1658);
and (s1n1657,n1066,n1655);
and (n1659,n1660,n981);
wire s0n1660,s1n1660,notn1660;
or (n1660,s0n1660,s1n1660);
not(notn1660,n1066);
and (s0n1660,notn1660,n1661);
and (s1n1660,n1066,n1658);
and (n1662,n1663,n970);
or (n1663,1'b0,n1664,n1667,n1670,n1673);
and (n1664,n1665,n947);
wire s0n1665,s1n1665,notn1665;
or (n1665,s0n1665,s1n1665);
not(notn1665,n1066);
and (s0n1665,notn1665,n1666);
and (s1n1665,n1066,n1661);
and (n1667,n1668,n958);
wire s0n1668,s1n1668,notn1668;
or (n1668,s0n1668,s1n1668);
not(notn1668,n1066);
and (s0n1668,notn1668,n1669);
and (s1n1668,n1066,n1666);
and (n1670,n1671,n1079);
wire s0n1671,s1n1671,notn1671;
or (n1671,s0n1671,s1n1671);
not(notn1671,n1066);
and (s0n1671,notn1671,n1672);
and (s1n1671,n1066,n1669);
and (n1673,n1674,n981);
wire s0n1674,s1n1674,notn1674;
or (n1674,s0n1674,s1n1674);
not(notn1674,n1066);
and (s0n1674,notn1674,n1675);
and (s1n1674,n1066,n1672);
wire s0n1677,s1n1677,notn1677;
or (n1677,s0n1677,s1n1677);
not(notn1677,n28);
and (s0n1677,notn1677,n1678);
and (s1n1677,n28,n1739);
or (n1678,1'b0,n1679,n1694,n1708,n1724);
and (n1679,n1680,n1056);
or (n1680,1'b0,n1681,n1685,n1688,n1691);
and (n1681,n1682,n947);
wire s0n1682,s1n1682,notn1682;
or (n1682,s0n1682,s1n1682);
not(notn1682,n1066);
and (s0n1682,notn1682,n1683);
and (s1n1682,n1066,n1684);
and (n1685,n1686,n958);
wire s0n1686,s1n1686,notn1686;
or (n1686,s0n1686,s1n1686);
not(notn1686,n1066);
and (s0n1686,notn1686,n1687);
and (s1n1686,n1066,n1683);
and (n1688,n1689,n1079);
wire s0n1689,s1n1689,notn1689;
or (n1689,s0n1689,s1n1689);
not(notn1689,n1066);
and (s0n1689,notn1689,n1690);
and (s1n1689,n1066,n1687);
and (n1691,n1692,n981);
wire s0n1692,s1n1692,notn1692;
or (n1692,s0n1692,s1n1692);
not(notn1692,n1066);
and (s0n1692,notn1692,n1693);
and (s1n1692,n1066,n1690);
and (n1694,n1695,n1041);
or (n1695,1'b0,n1696,n1699,n1702,n1705);
and (n1696,n1697,n947);
wire s0n1697,s1n1697,notn1697;
or (n1697,s0n1697,s1n1697);
not(notn1697,n1066);
and (s0n1697,notn1697,n1698);
and (s1n1697,n1066,n1693);
and (n1699,n1700,n958);
wire s0n1700,s1n1700,notn1700;
or (n1700,s0n1700,s1n1700);
not(notn1700,n1066);
and (s0n1700,notn1700,n1701);
and (s1n1700,n1066,n1698);
and (n1702,n1703,n1079);
wire s0n1703,s1n1703,notn1703;
or (n1703,s0n1703,s1n1703);
not(notn1703,n1066);
and (s0n1703,notn1703,n1704);
and (s1n1703,n1066,n1701);
and (n1705,n1706,n981);
wire s0n1706,s1n1706,notn1706;
or (n1706,s0n1706,s1n1706);
not(notn1706,n1066);
and (s0n1706,notn1706,n1707);
and (s1n1706,n1066,n1704);
and (n1708,n1709,n990);
nand (n1709,n1710,n1715);
nor (n1710,n1711,n1713);
and (n1711,n1007,n1712);
and (n1713,n1019,n1714);
nor (n1715,n1716,n1718);
and (n1716,n944,n1717);
nand (n1718,n1719,n1722);
or (n1719,n1720,n1121);
not (n1720,n1721);
nand (n1722,n979,n1723);
and (n1724,n1725,n970);
nand (n1725,n1726,n1731);
nor (n1726,n1727,n1729);
and (n1727,n1007,n1728);
and (n1729,n1019,n1730);
nor (n1731,n1732,n1734);
and (n1732,n944,n1733);
nand (n1734,n1735,n1737);
or (n1735,n1736,n1121);
not (n1736,n1723);
nand (n1737,n979,n1738);
and (n1740,n1677,n1741);
or (n1741,n1742,n1861,n1983);
and (n1742,n1743,n1800);
wire s0n1743,s1n1743,notn1743;
or (n1743,s0n1743,s1n1743);
not(notn1743,n28);
and (s0n1743,notn1743,n1744);
and (s1n1743,n28,n1799);
or (n1744,1'b0,n1745,n1758,n1770,n1785);
and (n1745,n1746,n1056);
nand (n1746,n1747,n1749,n1751,n1756);
nand (n1747,n1007,n1748);
nand (n1749,n1019,n1750);
nor (n1751,n1752,n1754);
and (n1752,n995,n1753);
and (n1754,n979,n1755);
nand (n1756,n944,n1757);
and (n1758,n1759,n1041);
nand (n1759,n1760,n1762,n1764,n1768);
nand (n1760,n1007,n1761);
nand (n1762,n1019,n1763);
nor (n1764,n1765,n1766);
and (n1765,n995,n1755);
and (n1766,n979,n1767);
nand (n1768,n944,n1769);
and (n1770,n1771,n990);
or (n1771,1'b0,n1772,n1776,n1779,n1782);
and (n1772,n1773,n947);
wire s0n1773,s1n1773,notn1773;
or (n1773,s0n1773,s1n1773);
not(notn1773,n1066);
and (s0n1773,notn1773,n1774);
and (s1n1773,n1066,n1775);
and (n1776,n1777,n958);
wire s0n1777,s1n1777,notn1777;
or (n1777,s0n1777,s1n1777);
not(notn1777,n1066);
and (s0n1777,notn1777,n1778);
and (s1n1777,n1066,n1774);
and (n1779,n1780,n1079);
wire s0n1780,s1n1780,notn1780;
or (n1780,s0n1780,s1n1780);
not(notn1780,n1066);
and (s0n1780,notn1780,n1781);
and (s1n1780,n1066,n1778);
and (n1782,n1783,n981);
wire s0n1783,s1n1783,notn1783;
or (n1783,s0n1783,s1n1783);
not(notn1783,n1066);
and (s0n1783,notn1783,n1784);
and (s1n1783,n1066,n1781);
and (n1785,n1786,n970);
or (n1786,1'b0,n1787,n1790,n1793,n1796);
and (n1787,n1788,n947);
wire s0n1788,s1n1788,notn1788;
or (n1788,s0n1788,s1n1788);
not(notn1788,n1066);
and (s0n1788,notn1788,n1789);
and (s1n1788,n1066,n1784);
and (n1790,n1791,n958);
wire s0n1791,s1n1791,notn1791;
or (n1791,s0n1791,s1n1791);
not(notn1791,n1066);
and (s0n1791,notn1791,n1792);
and (s1n1791,n1066,n1789);
and (n1793,n1794,n1079);
wire s0n1794,s1n1794,notn1794;
or (n1794,s0n1794,s1n1794);
not(notn1794,n1066);
and (s0n1794,notn1794,n1795);
and (s1n1794,n1066,n1792);
and (n1796,n1797,n981);
wire s0n1797,s1n1797,notn1797;
or (n1797,s0n1797,s1n1797);
not(notn1797,n1066);
and (s0n1797,notn1797,n1798);
and (s1n1797,n1066,n1795);
wire s0n1800,s1n1800,notn1800;
or (n1800,s0n1800,s1n1800);
not(notn1800,n28);
and (s0n1800,notn1800,n1801);
and (s1n1800,n28,n1860);
or (n1801,1'b0,n1802,n1817,n1831,n1845);
and (n1802,n1803,n1056);
or (n1803,1'b0,n1804,n1808,n1811,n1814);
and (n1804,n1805,n947);
wire s0n1805,s1n1805,notn1805;
or (n1805,s0n1805,s1n1805);
not(notn1805,n1066);
and (s0n1805,notn1805,n1806);
and (s1n1805,n1066,n1807);
and (n1808,n1809,n958);
wire s0n1809,s1n1809,notn1809;
or (n1809,s0n1809,s1n1809);
not(notn1809,n1066);
and (s0n1809,notn1809,n1810);
and (s1n1809,n1066,n1806);
and (n1811,n1812,n1079);
wire s0n1812,s1n1812,notn1812;
or (n1812,s0n1812,s1n1812);
not(notn1812,n1066);
and (s0n1812,notn1812,n1813);
and (s1n1812,n1066,n1810);
and (n1814,n1815,n981);
wire s0n1815,s1n1815,notn1815;
or (n1815,s0n1815,s1n1815);
not(notn1815,n1066);
and (s0n1815,notn1815,n1816);
and (s1n1815,n1066,n1813);
and (n1817,n1818,n1041);
or (n1818,1'b0,n1819,n1822,n1825,n1828);
and (n1819,n1820,n947);
wire s0n1820,s1n1820,notn1820;
or (n1820,s0n1820,s1n1820);
not(notn1820,n1066);
and (s0n1820,notn1820,n1821);
and (s1n1820,n1066,n1816);
and (n1822,n1823,n958);
wire s0n1823,s1n1823,notn1823;
or (n1823,s0n1823,s1n1823);
not(notn1823,n1066);
and (s0n1823,notn1823,n1824);
and (s1n1823,n1066,n1821);
and (n1825,n1826,n1079);
wire s0n1826,s1n1826,notn1826;
or (n1826,s0n1826,s1n1826);
not(notn1826,n1066);
and (s0n1826,notn1826,n1827);
and (s1n1826,n1066,n1824);
and (n1828,n1829,n981);
wire s0n1829,s1n1829,notn1829;
or (n1829,s0n1829,s1n1829);
not(notn1829,n1066);
and (s0n1829,notn1829,n1830);
and (s1n1829,n1066,n1827);
not (n1831,n1832);
nand (n1832,n1833,n990);
nand (n1833,n1834,n1839,n1841,n1843);
nor (n1834,n1835,n1837);
and (n1835,n995,n1836);
and (n1837,n979,n1838);
nand (n1839,n1007,n1840);
nand (n1841,n1019,n1842);
nand (n1843,n944,n1844);
not (n1845,n1846);
or (n1846,n971,n1847);
not (n1847,n1848);
nand (n1848,n1849,n1854,n1856,n1858);
nor (n1849,n1850,n1851);
and (n1850,n995,n1838);
nor (n1851,n1852,n980);
not (n1852,n1853);
nand (n1854,n1007,n1855);
nand (n1856,n1019,n1857);
nand (n1858,n944,n1859);
and (n1861,n1800,n1862);
and (n1862,n1863,n1920);
wire s0n1863,s1n1863,notn1863;
or (n1863,s0n1863,s1n1863);
not(notn1863,n28);
and (s0n1863,notn1863,n1864);
and (s1n1863,n28,n1919);
or (n1864,1'b0,n1865,n1878,n1890,n1905);
and (n1865,n1866,n1056);
nand (n1866,n1867,n1872,n1874,n1876);
nor (n1867,n1868,n1870);
and (n1868,n979,n1869);
and (n1870,n995,n1871);
nand (n1872,n944,n1873);
nand (n1874,n1007,n1875);
nand (n1876,n1019,n1877);
and (n1878,n1879,n1041);
nand (n1879,n1880,n1884,n1886,n1888);
nor (n1880,n1881,n1883);
and (n1881,n979,n1882);
and (n1883,n995,n1869);
nand (n1884,n944,n1885);
nand (n1886,n1007,n1887);
nand (n1888,n1019,n1889);
and (n1890,n1891,n990);
or (n1891,1'b0,n1892,n1896,n1899,n1902);
and (n1892,n1893,n947);
wire s0n1893,s1n1893,notn1893;
or (n1893,s0n1893,s1n1893);
not(notn1893,n1066);
and (s0n1893,notn1893,n1894);
and (s1n1893,n1066,n1895);
and (n1896,n1897,n958);
wire s0n1897,s1n1897,notn1897;
or (n1897,s0n1897,s1n1897);
not(notn1897,n1066);
and (s0n1897,notn1897,n1898);
and (s1n1897,n1066,n1894);
and (n1899,n1900,n1079);
wire s0n1900,s1n1900,notn1900;
or (n1900,s0n1900,s1n1900);
not(notn1900,n1066);
and (s0n1900,notn1900,n1901);
and (s1n1900,n1066,n1898);
and (n1902,n1903,n981);
wire s0n1903,s1n1903,notn1903;
or (n1903,s0n1903,s1n1903);
not(notn1903,n1066);
and (s0n1903,notn1903,n1904);
and (s1n1903,n1066,n1901);
and (n1905,n1906,n970);
or (n1906,1'b0,n1907,n1910,n1913,n1916);
and (n1907,n1908,n947);
wire s0n1908,s1n1908,notn1908;
or (n1908,s0n1908,s1n1908);
not(notn1908,n1066);
and (s0n1908,notn1908,n1909);
and (s1n1908,n1066,n1904);
and (n1910,n1911,n958);
wire s0n1911,s1n1911,notn1911;
or (n1911,s0n1911,s1n1911);
not(notn1911,n1066);
and (s0n1911,notn1911,n1912);
and (s1n1911,n1066,n1909);
and (n1913,n1914,n1079);
wire s0n1914,s1n1914,notn1914;
or (n1914,s0n1914,s1n1914);
not(notn1914,n1066);
and (s0n1914,notn1914,n1915);
and (s1n1914,n1066,n1912);
and (n1916,n1917,n981);
wire s0n1917,s1n1917,notn1917;
or (n1917,s0n1917,s1n1917);
not(notn1917,n1066);
and (s0n1917,notn1917,n1918);
and (s1n1917,n1066,n1915);
wire s0n1920,s1n1920,notn1920;
or (n1920,s0n1920,s1n1920);
not(notn1920,n28);
and (s0n1920,notn1920,n1921);
and (s1n1920,n28,n1982);
or (n1921,1'b0,n1922,n1937,n1951,n1967);
and (n1922,n1923,n1056);
or (n1923,1'b0,n1924,n1928,n1931,n1934);
and (n1924,n1925,n947);
wire s0n1925,s1n1925,notn1925;
or (n1925,s0n1925,s1n1925);
not(notn1925,n1066);
and (s0n1925,notn1925,n1926);
and (s1n1925,n1066,n1927);
and (n1928,n1929,n958);
wire s0n1929,s1n1929,notn1929;
or (n1929,s0n1929,s1n1929);
not(notn1929,n1066);
and (s0n1929,notn1929,n1930);
and (s1n1929,n1066,n1926);
and (n1931,n1932,n1079);
wire s0n1932,s1n1932,notn1932;
or (n1932,s0n1932,s1n1932);
not(notn1932,n1066);
and (s0n1932,notn1932,n1933);
and (s1n1932,n1066,n1930);
and (n1934,n1935,n981);
wire s0n1935,s1n1935,notn1935;
or (n1935,s0n1935,s1n1935);
not(notn1935,n1066);
and (s0n1935,notn1935,n1936);
and (s1n1935,n1066,n1933);
and (n1937,n1938,n1041);
or (n1938,1'b0,n1939,n1942,n1945,n1948);
and (n1939,n1940,n947);
wire s0n1940,s1n1940,notn1940;
or (n1940,s0n1940,s1n1940);
not(notn1940,n1066);
and (s0n1940,notn1940,n1941);
and (s1n1940,n1066,n1936);
and (n1942,n1943,n958);
wire s0n1943,s1n1943,notn1943;
or (n1943,s0n1943,s1n1943);
not(notn1943,n1066);
and (s0n1943,notn1943,n1944);
and (s1n1943,n1066,n1941);
and (n1945,n1946,n1079);
wire s0n1946,s1n1946,notn1946;
or (n1946,s0n1946,s1n1946);
not(notn1946,n1066);
and (s0n1946,notn1946,n1947);
and (s1n1946,n1066,n1944);
and (n1948,n1949,n981);
wire s0n1949,s1n1949,notn1949;
or (n1949,s0n1949,s1n1949);
not(notn1949,n1066);
and (s0n1949,notn1949,n1950);
and (s1n1949,n1066,n1947);
and (n1951,n1952,n990);
nand (n1952,n1953,n1958);
nor (n1953,n1954,n1956);
and (n1954,n1019,n1955);
and (n1956,n1007,n1957);
nor (n1958,n1959,n1961);
and (n1959,n944,n1960);
nand (n1961,n1962,n1965);
or (n1962,n1963,n1121);
not (n1963,n1964);
nand (n1965,n979,n1966);
and (n1967,n1968,n970);
nand (n1968,n1969,n1974);
nor (n1969,n1970,n1972);
and (n1970,n1019,n1971);
and (n1972,n1007,n1973);
nor (n1974,n1975,n1977);
and (n1975,n944,n1976);
nand (n1977,n1978,n1980);
or (n1978,n1979,n1121);
not (n1979,n1966);
nand (n1980,n979,n1981);
and (n1983,n1743,n1862);
and (n1984,n1620,n1741);
and (n1985,n1496,n1618);
and (n1986,n1381,n1494);
and (n1987,n1257,n1379);
and (n1988,n1132,n1255);
and (n1989,n937,n1130);
and (n1990,n930,n935);
and (n1991,n923,n928);
xor (n1992,n1993,n3684);
xor (n1993,n1994,n3573);
xor (n1994,n1995,n2960);
xor (n1995,n1996,n2001);
xor (n1996,n1997,n1999);
wire s0n1997,s1n1997,notn1997;
or (n1997,s0n1997,s1n1997);
not(notn1997,n28);
and (s0n1997,notn1997,1'b0);
and (s1n1997,n28,n1998);
wire s0n1999,s1n1999,notn1999;
or (n1999,s0n1999,s1n1999);
not(notn1999,n28);
and (s0n1999,notn1999,1'b0);
and (s1n1999,n28,n2000);
or (n2001,n2002,n2106,n2959);
and (n2002,n2003,n2054);
wire s0n2003,s1n2003,notn2003;
or (n2003,s0n2003,s1n2003);
not(notn2003,n28);
and (s0n2003,notn2003,n2004);
and (s1n2003,n28,n2053);
nand (n2004,n2005,n2031,n2043,n2048);
nor (n2005,n2006,n2019);
and (n2006,n2007,n1041);
nand (n2007,n2008,n2013,n2015,n2017);
nor (n2008,n2009,n2011);
and (n2009,n995,n2010);
and (n2011,n979,n2012);
nand (n2013,n944,n2014);
nand (n2015,n1007,n2016);
nand (n2017,n1019,n2018);
and (n2019,n2020,n1056);
nand (n2020,n2021,n2025,n2027,n2029);
nor (n2021,n2022,n2024);
and (n2022,n995,n2023);
and (n2024,n979,n2010);
nand (n2025,n944,n2026);
nand (n2027,n1007,n2028);
nand (n2029,n1019,n2030);
nor (n2031,n2032,n2034);
and (n2032,n999,n2033);
nand (n2034,n2035,n2037,n2039,n2041);
nand (n2035,n989,n2036);
nand (n2037,n943,n2038);
nand (n2039,n994,n2040);
nand (n2041,n977,n2042);
nor (n2043,n2044,n2046);
and (n2044,n1005,n2045);
and (n2046,n1017,n2047);
nor (n2048,n2049,n2051);
and (n2049,n1175,n2050);
and (n2051,n1024,n2052);
wire s0n2054,s1n2054,notn2054;
or (n2054,s0n2054,s1n2054);
not(notn2054,n28);
and (s0n2054,notn2054,n2055);
and (s1n2054,n28,n2105);
nand (n2055,n2056,n2069,n2095,n2100);
nor (n2056,n2057,n2067);
nand (n2057,n2058,n2063,n2065);
nor (n2058,n2059,n2061);
and (n2059,n943,n2060);
and (n2061,n977,n2062);
nand (n2063,n989,n2064);
nand (n2065,n994,n2066);
and (n2067,n999,n2068);
nor (n2069,n2070,n2083);
and (n2070,n2071,n1041);
nand (n2071,n2072,n2077,n2079,n2081);
nor (n2072,n2073,n2075);
and (n2073,n995,n2074);
and (n2075,n979,n2076);
nand (n2077,n944,n2078);
nand (n2079,n1007,n2080);
nand (n2081,n1019,n2082);
and (n2083,n2084,n1056);
nand (n2084,n2085,n2089,n2091,n2093);
nor (n2085,n2086,n2088);
and (n2086,n995,n2087);
and (n2088,n979,n2074);
nand (n2089,n944,n2090);
nand (n2091,n1007,n2092);
nand (n2093,n1019,n2094);
nor (n2095,n2096,n2098);
and (n2096,n1175,n2097);
and (n2098,n1005,n2099);
nor (n2100,n2101,n2103);
and (n2101,n1024,n2102);
and (n2103,n1017,n2104);
and (n2106,n2054,n2107);
or (n2107,n2108,n2226,n2958);
and (n2108,n2109,n2161);
wire s0n2109,s1n2109,notn2109;
or (n2109,s0n2109,s1n2109);
not(notn2109,n28);
and (s0n2109,notn2109,n2110);
and (s1n2109,n28,n2160);
nand (n2110,n2111,n2137,n2150,n2155);
nor (n2111,n2112,n2125);
and (n2112,n2113,n1041);
nand (n2113,n2114,n2119,n2121,n2123);
nor (n2114,n2115,n2117);
and (n2115,n995,n2116);
and (n2117,n979,n2118);
nand (n2119,n944,n2120);
nand (n2121,n1007,n2122);
nand (n2123,n1019,n2124);
and (n2125,n2126,n1056);
nand (n2126,n2127,n2131,n2133,n2135);
nor (n2127,n2128,n2130);
and (n2128,n995,n2129);
and (n2130,n979,n2116);
nand (n2131,n944,n2132);
nand (n2133,n1007,n2134);
nand (n2135,n1019,n2136);
nor (n2137,n2138,n2140);
and (n2138,n999,n2139);
nand (n2140,n2141,n2146,n2148);
nor (n2141,n2142,n2144);
and (n2142,n977,n2143);
and (n2144,n943,n2145);
nand (n2146,n994,n2147);
nand (n2148,n989,n2149);
nor (n2150,n2151,n2153);
and (n2151,n1175,n2152);
and (n2153,n1005,n2154);
nor (n2155,n2156,n2158);
and (n2156,n1024,n2157);
and (n2158,n1017,n2159);
wire s0n2161,s1n2161,notn2161;
or (n2161,s0n2161,s1n2161);
not(notn2161,n28);
and (s0n2161,notn2161,n2162);
and (s1n2161,n28,n2225);
or (n2162,1'b0,n2163,n2180,n2196,n2211);
and (n2163,n2164,n1056);
nand (n2164,n2165,n2170);
nor (n2165,n2166,n2168);
and (n2166,n1007,n2167);
and (n2168,n1019,n2169);
nor (n2170,n2171,n2177);
nand (n2171,n2172,n2175);
or (n2172,n2173,n1121);
not (n2173,n2174);
nand (n2175,n979,n2176);
nor (n2177,n2178,n1127);
not (n2178,n2179);
and (n2180,n2181,n1041);
nand (n2181,n2182,n2187);
nor (n2182,n2183,n2185);
and (n2183,n1007,n2184);
and (n2185,n1019,n2186);
nor (n2187,n2188,n2193);
nand (n2188,n2189,n2191);
or (n2189,n2190,n1121);
not (n2190,n2176);
nand (n2191,n979,n2192);
nor (n2193,n2194,n1127);
not (n2194,n2195);
and (n2196,n2197,n990);
or (n2197,1'b0,n2198,n2202,n2205,n2208);
and (n2198,n2199,n947);
wire s0n2199,s1n2199,notn2199;
or (n2199,s0n2199,s1n2199);
not(notn2199,n1066);
and (s0n2199,notn2199,n2200);
and (s1n2199,n1066,n2201);
and (n2202,n2203,n958);
wire s0n2203,s1n2203,notn2203;
or (n2203,s0n2203,s1n2203);
not(notn2203,n1066);
and (s0n2203,notn2203,n2204);
and (s1n2203,n1066,n2200);
and (n2205,n2206,n1079);
wire s0n2206,s1n2206,notn2206;
or (n2206,s0n2206,s1n2206);
not(notn2206,n1066);
and (s0n2206,notn2206,n2207);
and (s1n2206,n1066,n2204);
and (n2208,n2209,n981);
wire s0n2209,s1n2209,notn2209;
or (n2209,s0n2209,s1n2209);
not(notn2209,n1066);
and (s0n2209,notn2209,n2210);
and (s1n2209,n1066,n2207);
and (n2211,n2212,n970);
or (n2212,1'b0,n2213,n2216,n2219,n2222);
and (n2213,n2214,n947);
wire s0n2214,s1n2214,notn2214;
or (n2214,s0n2214,s1n2214);
not(notn2214,n1066);
and (s0n2214,notn2214,n2215);
and (s1n2214,n1066,n2210);
and (n2216,n2217,n958);
wire s0n2217,s1n2217,notn2217;
or (n2217,s0n2217,s1n2217);
not(notn2217,n1066);
and (s0n2217,notn2217,n2218);
and (s1n2217,n1066,n2215);
and (n2219,n2220,n1079);
wire s0n2220,s1n2220,notn2220;
or (n2220,s0n2220,s1n2220);
not(notn2220,n1066);
and (s0n2220,notn2220,n2221);
and (s1n2220,n1066,n2218);
and (n2222,n2223,n981);
wire s0n2223,s1n2223,notn2223;
or (n2223,s0n2223,s1n2223);
not(notn2223,n1066);
and (s0n2223,notn2223,n2224);
and (s1n2223,n1066,n2221);
and (n2226,n2161,n2227);
or (n2227,n2228,n2334,n2957);
and (n2228,n2229,n2282);
wire s0n2229,s1n2229,notn2229;
or (n2229,s0n2229,s1n2229);
not(notn2229,n28);
and (s0n2229,notn2229,n2230);
and (s1n2229,n28,n2281);
nand (n2230,n2231,n2245,n2271,n2276);
nor (n2231,n2232,n2234);
and (n2232,n999,n2233);
nand (n2234,n2235,n2241,n2243);
nor (n2235,n2236,n2238);
and (n2236,n943,n2237);
nor (n2238,n2239,n978);
not (n2239,n2240);
nand (n2241,n994,n2242);
nand (n2243,n989,n2244);
nor (n2245,n2246,n2259);
and (n2246,n2247,n1041);
nand (n2247,n2248,n2250,n2252,n2257);
nand (n2248,n1007,n2249);
nand (n2250,n1019,n2251);
nor (n2252,n2253,n2255);
and (n2253,n995,n2254);
and (n2255,n979,n2256);
nand (n2257,n944,n2258);
and (n2259,n2260,n1056);
nand (n2260,n2261,n2263,n2265,n2269);
nand (n2261,n1007,n2262);
nand (n2263,n1019,n2264);
nor (n2265,n2266,n2268);
and (n2266,n995,n2267);
and (n2268,n979,n2254);
nand (n2269,n944,n2270);
nor (n2271,n2272,n2274);
and (n2272,n1175,n2273);
and (n2274,n1005,n2275);
nor (n2276,n2277,n2279);
and (n2277,n1024,n2278);
and (n2279,n1017,n2280);
wire s0n2282,s1n2282,notn2282;
or (n2282,s0n2282,s1n2282);
not(notn2282,n28);
and (s0n2282,notn2282,n2283);
and (s1n2282,n28,n2333);
nand (n2283,n2284,n2297,n2313,n2328);
nor (n2284,n2285,n2287);
and (n2285,n999,n2286);
nand (n2287,n2288,n2290,n2295);
nand (n2288,n943,n2289);
nor (n2290,n2291,n2293);
and (n2291,n989,n2292);
and (n2293,n977,n2294);
nand (n2295,n994,n2296);
nor (n2297,n2298,n2311);
and (n2298,n2299,n1056);
nand (n2299,n2300,n2305,n2307,n2309);
nor (n2300,n2301,n2303);
and (n2301,n995,n2302);
and (n2303,n979,n2304);
nand (n2305,n944,n2306);
nand (n2307,n1007,n2308);
nand (n2309,n1019,n2310);
and (n2311,n1175,n2312);
nor (n2313,n2314,n2326);
and (n2314,n2315,n1041);
nand (n2315,n2316,n2320,n2322,n2324);
nor (n2316,n2317,n2318);
and (n2317,n995,n2304);
and (n2318,n979,n2319);
nand (n2320,n944,n2321);
nand (n2322,n1007,n2323);
nand (n2324,n1019,n2325);
and (n2326,n1017,n2327);
nor (n2328,n2329,n2331);
and (n2329,n1005,n2330);
and (n2331,n1024,n2332);
and (n2334,n2282,n2335);
or (n2335,n2336,n2462,n2956);
and (n2336,n2337,n2402);
wire s0n2337,s1n2337,notn2337;
or (n2337,s0n2337,s1n2337);
not(notn2337,n28);
and (s0n2337,notn2337,n2338);
and (s1n2337,n28,n2401);
or (n2338,1'b0,n2339,n2356,n2372,n2387);
and (n2339,n2340,n1056);
nand (n2340,n2341,n2346);
nor (n2341,n2342,n2344);
and (n2342,n1019,n2343);
and (n2344,n1007,n2345);
nor (n2346,n2347,n2353);
nand (n2347,n2348,n2351);
or (n2348,n2349,n1121);
not (n2349,n2350);
nand (n2351,n979,n2352);
nor (n2353,n2354,n1127);
not (n2354,n2355);
and (n2356,n2357,n1041);
nand (n2357,n2358,n2363);
nor (n2358,n2359,n2361);
and (n2359,n1019,n2360);
and (n2361,n1007,n2362);
nor (n2363,n2364,n2369);
nand (n2364,n2365,n2367);
or (n2365,n2366,n1121);
not (n2366,n2352);
nand (n2367,n979,n2368);
nor (n2369,n1127,n2370);
not (n2370,n2371);
and (n2372,n2373,n990);
or (n2373,1'b0,n2374,n2378,n2381,n2384);
and (n2374,n2375,n947);
wire s0n2375,s1n2375,notn2375;
or (n2375,s0n2375,s1n2375);
not(notn2375,n1066);
and (s0n2375,notn2375,n2376);
and (s1n2375,n1066,n2377);
and (n2378,n2379,n958);
wire s0n2379,s1n2379,notn2379;
or (n2379,s0n2379,s1n2379);
not(notn2379,n1066);
and (s0n2379,notn2379,n2380);
and (s1n2379,n1066,n2376);
and (n2381,n2382,n1079);
wire s0n2382,s1n2382,notn2382;
or (n2382,s0n2382,s1n2382);
not(notn2382,n1066);
and (s0n2382,notn2382,n2383);
and (s1n2382,n1066,n2380);
and (n2384,n2385,n981);
wire s0n2385,s1n2385,notn2385;
or (n2385,s0n2385,s1n2385);
not(notn2385,n1066);
and (s0n2385,notn2385,n2386);
and (s1n2385,n1066,n2383);
and (n2387,n2388,n970);
or (n2388,1'b0,n2389,n2392,n2395,n2398);
and (n2389,n2390,n947);
wire s0n2390,s1n2390,notn2390;
or (n2390,s0n2390,s1n2390);
not(notn2390,n1066);
and (s0n2390,notn2390,n2391);
and (s1n2390,n1066,n2386);
and (n2392,n2393,n958);
wire s0n2393,s1n2393,notn2393;
or (n2393,s0n2393,s1n2393);
not(notn2393,n1066);
and (s0n2393,notn2393,n2394);
and (s1n2393,n1066,n2391);
and (n2395,n2396,n1079);
wire s0n2396,s1n2396,notn2396;
or (n2396,s0n2396,s1n2396);
not(notn2396,n1066);
and (s0n2396,notn2396,n2397);
and (s1n2396,n1066,n2394);
and (n2398,n2399,n981);
wire s0n2399,s1n2399,notn2399;
or (n2399,s0n2399,s1n2399);
not(notn2399,n1066);
and (s0n2399,notn2399,n2400);
and (s1n2399,n1066,n2397);
wire s0n2402,s1n2402,notn2402;
or (n2402,s0n2402,s1n2402);
not(notn2402,n28);
and (s0n2402,notn2402,n2403);
and (s1n2402,n28,n2461);
or (n2403,1'b0,n2404,n2417,n2432,n2447);
and (n2404,n2405,n1056);
nand (n2405,n2406,n2411,n2413,n2415);
nor (n2406,n2407,n2409);
and (n2407,n995,n2408);
and (n2409,n979,n2410);
nand (n2411,n944,n2412);
nand (n2413,n1007,n2414);
nand (n2415,n1019,n2416);
and (n2417,n2418,n1041);
nand (n2418,n2419,n2424);
nor (n2419,n2420,n2422);
and (n2420,n1007,n2421);
and (n2422,n1019,n2423);
nor (n2424,n2425,n2430);
nand (n2425,n2426,n2428);
or (n2426,n2427,n1121);
not (n2427,n2410);
nand (n2428,n979,n2429);
and (n2430,n944,n2431);
and (n2432,n2433,n990);
or (n2433,1'b0,n2434,n2438,n2441,n2444);
and (n2434,n2435,n947);
wire s0n2435,s1n2435,notn2435;
or (n2435,s0n2435,s1n2435);
not(notn2435,n1066);
and (s0n2435,notn2435,n2436);
and (s1n2435,n1066,n2437);
and (n2438,n2439,n958);
wire s0n2439,s1n2439,notn2439;
or (n2439,s0n2439,s1n2439);
not(notn2439,n1066);
and (s0n2439,notn2439,n2440);
and (s1n2439,n1066,n2436);
and (n2441,n2442,n1079);
wire s0n2442,s1n2442,notn2442;
or (n2442,s0n2442,s1n2442);
not(notn2442,n1066);
and (s0n2442,notn2442,n2443);
and (s1n2442,n1066,n2440);
and (n2444,n2445,n981);
wire s0n2445,s1n2445,notn2445;
or (n2445,s0n2445,s1n2445);
not(notn2445,n1066);
and (s0n2445,notn2445,n2446);
and (s1n2445,n1066,n2443);
and (n2447,n2448,n970);
or (n2448,1'b0,n2449,n2452,n2455,n2458);
and (n2449,n2450,n947);
wire s0n2450,s1n2450,notn2450;
or (n2450,s0n2450,s1n2450);
not(notn2450,n1066);
and (s0n2450,notn2450,n2451);
and (s1n2450,n1066,n2446);
and (n2452,n2453,n958);
wire s0n2453,s1n2453,notn2453;
or (n2453,s0n2453,s1n2453);
not(notn2453,n1066);
and (s0n2453,notn2453,n2454);
and (s1n2453,n1066,n2451);
and (n2455,n2456,n1079);
wire s0n2456,s1n2456,notn2456;
or (n2456,s0n2456,s1n2456);
not(notn2456,n1066);
and (s0n2456,notn2456,n2457);
and (s1n2456,n1066,n2454);
and (n2458,n2459,n981);
wire s0n2459,s1n2459,notn2459;
or (n2459,s0n2459,s1n2459);
not(notn2459,n1066);
and (s0n2459,notn2459,n2460);
and (s1n2459,n1066,n2457);
and (n2462,n2402,n2463);
or (n2463,n2464,n2587,n2955);
and (n2464,n2465,n2530);
wire s0n2465,s1n2465,notn2465;
or (n2465,s0n2465,s1n2465);
not(notn2465,n28);
and (s0n2465,notn2465,n2466);
and (s1n2465,n28,n2529);
or (n2466,1'b0,n2467,n2484,n2500,n2515);
and (n2467,n2468,n1056);
nand (n2468,n2469,n2474);
nor (n2469,n2470,n2472);
and (n2470,n1007,n2471);
and (n2472,n1019,n2473);
nor (n2474,n2475,n2481);
nand (n2475,n2476,n2479);
or (n2476,n2477,n1121);
not (n2477,n2478);
nand (n2479,n979,n2480);
nor (n2481,n2482,n1127);
not (n2482,n2483);
and (n2484,n2485,n1041);
nand (n2485,n2486,n2491);
nor (n2486,n2487,n2489);
and (n2487,n1007,n2488);
and (n2489,n1019,n2490);
nor (n2491,n2492,n2497);
nand (n2492,n2493,n2495);
or (n2493,n2494,n1121);
not (n2494,n2480);
nand (n2495,n979,n2496);
nor (n2497,n2498,n1127);
not (n2498,n2499);
and (n2500,n2501,n990);
or (n2501,1'b0,n2502,n2506,n2509,n2512);
and (n2502,n2503,n947);
wire s0n2503,s1n2503,notn2503;
or (n2503,s0n2503,s1n2503);
not(notn2503,n1066);
and (s0n2503,notn2503,n2504);
and (s1n2503,n1066,n2505);
and (n2506,n2507,n958);
wire s0n2507,s1n2507,notn2507;
or (n2507,s0n2507,s1n2507);
not(notn2507,n1066);
and (s0n2507,notn2507,n2508);
and (s1n2507,n1066,n2504);
and (n2509,n2510,n1079);
wire s0n2510,s1n2510,notn2510;
or (n2510,s0n2510,s1n2510);
not(notn2510,n1066);
and (s0n2510,notn2510,n2511);
and (s1n2510,n1066,n2508);
and (n2512,n2513,n981);
wire s0n2513,s1n2513,notn2513;
or (n2513,s0n2513,s1n2513);
not(notn2513,n1066);
and (s0n2513,notn2513,n2514);
and (s1n2513,n1066,n2511);
and (n2515,n2516,n970);
or (n2516,1'b0,n2517,n2520,n2523,n2526);
and (n2517,n2518,n947);
wire s0n2518,s1n2518,notn2518;
or (n2518,s0n2518,s1n2518);
not(notn2518,n1066);
and (s0n2518,notn2518,n2519);
and (s1n2518,n1066,n2514);
and (n2520,n2521,n958);
wire s0n2521,s1n2521,notn2521;
or (n2521,s0n2521,s1n2521);
not(notn2521,n1066);
and (s0n2521,notn2521,n2522);
and (s1n2521,n1066,n2519);
and (n2523,n2524,n1079);
wire s0n2524,s1n2524,notn2524;
or (n2524,s0n2524,s1n2524);
not(notn2524,n1066);
and (s0n2524,notn2524,n2525);
and (s1n2524,n1066,n2522);
and (n2526,n2527,n981);
wire s0n2527,s1n2527,notn2527;
or (n2527,s0n2527,s1n2527);
not(notn2527,n1066);
and (s0n2527,notn2527,n2528);
and (s1n2527,n1066,n2525);
wire s0n2530,s1n2530,notn2530;
or (n2530,s0n2530,s1n2530);
not(notn2530,n28);
and (s0n2530,notn2530,n2531);
and (s1n2530,n28,n2586);
or (n2531,1'b0,n2532,n2545,n2557,n2572);
and (n2532,n2533,n1056);
nand (n2533,n2534,n2536,n2538,n2543);
nand (n2534,n1007,n2535);
nand (n2536,n1019,n2537);
nor (n2538,n2539,n2541);
and (n2539,n995,n2540);
and (n2541,n979,n2542);
nand (n2543,n944,n2544);
and (n2545,n2546,n1041);
nand (n2546,n2547,n2549,n2551,n2555);
nand (n2547,n1007,n2548);
nand (n2549,n1019,n2550);
nor (n2551,n2552,n2553);
and (n2552,n995,n2542);
and (n2553,n979,n2554);
nand (n2555,n944,n2556);
and (n2557,n2558,n990);
or (n2558,1'b0,n2559,n2563,n2566,n2569);
and (n2559,n2560,n947);
wire s0n2560,s1n2560,notn2560;
or (n2560,s0n2560,s1n2560);
not(notn2560,n1066);
and (s0n2560,notn2560,n2561);
and (s1n2560,n1066,n2562);
and (n2563,n2564,n958);
wire s0n2564,s1n2564,notn2564;
or (n2564,s0n2564,s1n2564);
not(notn2564,n1066);
and (s0n2564,notn2564,n2565);
and (s1n2564,n1066,n2561);
and (n2566,n2567,n1079);
wire s0n2567,s1n2567,notn2567;
or (n2567,s0n2567,s1n2567);
not(notn2567,n1066);
and (s0n2567,notn2567,n2568);
and (s1n2567,n1066,n2565);
and (n2569,n2570,n981);
wire s0n2570,s1n2570,notn2570;
or (n2570,s0n2570,s1n2570);
not(notn2570,n1066);
and (s0n2570,notn2570,n2571);
and (s1n2570,n1066,n2568);
and (n2572,n2573,n970);
or (n2573,1'b0,n2574,n2577,n2580,n2583);
and (n2574,n2575,n947);
wire s0n2575,s1n2575,notn2575;
or (n2575,s0n2575,s1n2575);
not(notn2575,n1066);
and (s0n2575,notn2575,n2576);
and (s1n2575,n1066,n2571);
and (n2577,n2578,n958);
wire s0n2578,s1n2578,notn2578;
or (n2578,s0n2578,s1n2578);
not(notn2578,n1066);
and (s0n2578,notn2578,n2579);
and (s1n2578,n1066,n2576);
and (n2580,n2581,n1079);
wire s0n2581,s1n2581,notn2581;
or (n2581,s0n2581,s1n2581);
not(notn2581,n1066);
and (s0n2581,notn2581,n2582);
and (s1n2581,n1066,n2579);
and (n2583,n2584,n981);
wire s0n2584,s1n2584,notn2584;
or (n2584,s0n2584,s1n2584);
not(notn2584,n1066);
and (s0n2584,notn2584,n2585);
and (s1n2584,n1066,n2582);
and (n2587,n2530,n2588);
or (n2588,n2589,n2704,n2954);
and (n2589,n2590,n2647);
wire s0n2590,s1n2590,notn2590;
or (n2590,s0n2590,s1n2590);
not(notn2590,n28);
and (s0n2590,notn2590,n2591);
and (s1n2590,n28,n2646);
or (n2591,1'b0,n2592,n2605,n2617,n2632);
and (n2592,n2593,n1056);
nand (n2593,n2594,n2599,n2601,n2603);
nor (n2594,n2595,n2597);
and (n2595,n995,n2596);
and (n2597,n979,n2598);
nand (n2599,n944,n2600);
nand (n2601,n1007,n2602);
nand (n2603,n1019,n2604);
and (n2605,n2606,n1041);
nand (n2606,n2607,n2611,n2613,n2615);
nor (n2607,n2608,n2609);
and (n2608,n995,n2598);
and (n2609,n979,n2610);
nand (n2611,n944,n2612);
nand (n2613,n1007,n2614);
nand (n2615,n1019,n2616);
and (n2617,n2618,n990);
or (n2618,1'b0,n2619,n2623,n2626,n2629);
and (n2619,n2620,n947);
wire s0n2620,s1n2620,notn2620;
or (n2620,s0n2620,s1n2620);
not(notn2620,n1066);
and (s0n2620,notn2620,n2621);
and (s1n2620,n1066,n2622);
and (n2623,n2624,n958);
wire s0n2624,s1n2624,notn2624;
or (n2624,s0n2624,s1n2624);
not(notn2624,n1066);
and (s0n2624,notn2624,n2625);
and (s1n2624,n1066,n2621);
and (n2626,n2627,n1079);
wire s0n2627,s1n2627,notn2627;
or (n2627,s0n2627,s1n2627);
not(notn2627,n1066);
and (s0n2627,notn2627,n2628);
and (s1n2627,n1066,n2625);
and (n2629,n2630,n981);
wire s0n2630,s1n2630,notn2630;
or (n2630,s0n2630,s1n2630);
not(notn2630,n1066);
and (s0n2630,notn2630,n2631);
and (s1n2630,n1066,n2628);
and (n2632,n2633,n970);
or (n2633,1'b0,n2634,n2637,n2640,n2643);
and (n2634,n2635,n947);
wire s0n2635,s1n2635,notn2635;
or (n2635,s0n2635,s1n2635);
not(notn2635,n1066);
and (s0n2635,notn2635,n2636);
and (s1n2635,n1066,n2631);
and (n2637,n2638,n958);
wire s0n2638,s1n2638,notn2638;
or (n2638,s0n2638,s1n2638);
not(notn2638,n1066);
and (s0n2638,notn2638,n2639);
and (s1n2638,n1066,n2636);
and (n2640,n2641,n1079);
wire s0n2641,s1n2641,notn2641;
or (n2641,s0n2641,s1n2641);
not(notn2641,n1066);
and (s0n2641,notn2641,n2642);
and (s1n2641,n1066,n2639);
and (n2643,n2644,n981);
wire s0n2644,s1n2644,notn2644;
or (n2644,s0n2644,s1n2644);
not(notn2644,n1066);
and (s0n2644,notn2644,n2645);
and (s1n2644,n1066,n2642);
wire s0n2647,s1n2647,notn2647;
or (n2647,s0n2647,s1n2647);
not(notn2647,n28);
and (s0n2647,notn2647,n2648);
and (s1n2647,n28,n2703);
or (n2648,1'b0,n2649,n2662,n2674,n2689);
and (n2649,n2650,n1056);
nand (n2650,n2651,n2656,n2658,n2660);
nor (n2651,n2652,n2654);
and (n2652,n995,n2653);
and (n2654,n979,n2655);
nand (n2656,n944,n2657);
nand (n2658,n1007,n2659);
nand (n2660,n1019,n2661);
and (n2662,n2663,n1041);
nand (n2663,n2664,n2668,n2670,n2672);
nor (n2664,n2665,n2667);
and (n2665,n979,n2666);
and (n2667,n995,n2655);
nand (n2668,n944,n2669);
nand (n2670,n1007,n2671);
nand (n2672,n1019,n2673);
and (n2674,n2675,n990);
or (n2675,1'b0,n2676,n2680,n2683,n2686);
and (n2676,n2677,n947);
wire s0n2677,s1n2677,notn2677;
or (n2677,s0n2677,s1n2677);
not(notn2677,n1066);
and (s0n2677,notn2677,n2678);
and (s1n2677,n1066,n2679);
and (n2680,n2681,n958);
wire s0n2681,s1n2681,notn2681;
or (n2681,s0n2681,s1n2681);
not(notn2681,n1066);
and (s0n2681,notn2681,n2682);
and (s1n2681,n1066,n2678);
and (n2683,n2684,n1079);
wire s0n2684,s1n2684,notn2684;
or (n2684,s0n2684,s1n2684);
not(notn2684,n1066);
and (s0n2684,notn2684,n2685);
and (s1n2684,n1066,n2682);
and (n2686,n2687,n981);
wire s0n2687,s1n2687,notn2687;
or (n2687,s0n2687,s1n2687);
not(notn2687,n1066);
and (s0n2687,notn2687,n2688);
and (s1n2687,n1066,n2685);
and (n2689,n2690,n970);
or (n2690,1'b0,n2691,n2694,n2697,n2700);
and (n2691,n2692,n947);
wire s0n2692,s1n2692,notn2692;
or (n2692,s0n2692,s1n2692);
not(notn2692,n1066);
and (s0n2692,notn2692,n2693);
and (s1n2692,n1066,n2688);
and (n2694,n2695,n958);
wire s0n2695,s1n2695,notn2695;
or (n2695,s0n2695,s1n2695);
not(notn2695,n1066);
and (s0n2695,notn2695,n2696);
and (s1n2695,n1066,n2693);
and (n2697,n2698,n1079);
wire s0n2698,s1n2698,notn2698;
or (n2698,s0n2698,s1n2698);
not(notn2698,n1066);
and (s0n2698,notn2698,n2699);
and (s1n2698,n1066,n2696);
and (n2700,n2701,n981);
wire s0n2701,s1n2701,notn2701;
or (n2701,s0n2701,s1n2701);
not(notn2701,n1066);
and (s0n2701,notn2701,n2702);
and (s1n2701,n1066,n2699);
and (n2704,n2647,n2705);
or (n2705,n2706,n2828,n2953);
and (n2706,n2707,n2767);
wire s0n2707,s1n2707,notn2707;
or (n2707,s0n2707,s1n2707);
not(notn2707,n28);
and (s0n2707,notn2707,n2708);
and (s1n2707,n28,n2766);
or (n2708,1'b0,n2709,n2724,n2737,n2752);
and (n2709,n2710,n1056);
or (n2710,1'b0,n2711,n2715,n2718,n2721);
and (n2711,n2712,n947);
wire s0n2712,s1n2712,notn2712;
or (n2712,s0n2712,s1n2712);
not(notn2712,n1066);
and (s0n2712,notn2712,n2713);
and (s1n2712,n1066,n2714);
and (n2715,n2716,n958);
wire s0n2716,s1n2716,notn2716;
or (n2716,s0n2716,s1n2716);
not(notn2716,n1066);
and (s0n2716,notn2716,n2717);
and (s1n2716,n1066,n2713);
and (n2718,n2719,n1079);
wire s0n2719,s1n2719,notn2719;
or (n2719,s0n2719,s1n2719);
not(notn2719,n1066);
and (s0n2719,notn2719,n2720);
and (s1n2719,n1066,n2717);
and (n2721,n2722,n981);
wire s0n2722,s1n2722,notn2722;
or (n2722,s0n2722,s1n2722);
not(notn2722,n1066);
and (s0n2722,notn2722,n2723);
and (s1n2722,n1066,n2720);
and (n2724,n2725,n1041);
nand (n2725,n2726,n2731);
nor (n2726,n2727,n2729);
and (n2727,n1019,n2728);
and (n2729,n1007,n2730);
and (n2731,n2732,n2733,n2735);
nand (n2732,n995,n2723);
nand (n2733,n944,n2734);
nand (n2735,n979,n2736);
and (n2737,n2738,n990);
or (n2738,1'b0,n2739,n2743,n2746,n2749);
and (n2739,n2740,n947);
wire s0n2740,s1n2740,notn2740;
or (n2740,s0n2740,s1n2740);
not(notn2740,n1066);
and (s0n2740,notn2740,n2741);
and (s1n2740,n1066,n2742);
and (n2743,n2744,n958);
wire s0n2744,s1n2744,notn2744;
or (n2744,s0n2744,s1n2744);
not(notn2744,n1066);
and (s0n2744,notn2744,n2745);
and (s1n2744,n1066,n2741);
and (n2746,n2747,n1079);
wire s0n2747,s1n2747,notn2747;
or (n2747,s0n2747,s1n2747);
not(notn2747,n1066);
and (s0n2747,notn2747,n2748);
and (s1n2747,n1066,n2745);
and (n2749,n2750,n981);
wire s0n2750,s1n2750,notn2750;
or (n2750,s0n2750,s1n2750);
not(notn2750,n1066);
and (s0n2750,notn2750,n2751);
and (s1n2750,n1066,n2748);
and (n2752,n2753,n970);
or (n2753,1'b0,n2754,n2757,n2760,n2763);
and (n2754,n2755,n947);
wire s0n2755,s1n2755,notn2755;
or (n2755,s0n2755,s1n2755);
not(notn2755,n1066);
and (s0n2755,notn2755,n2756);
and (s1n2755,n1066,n2751);
and (n2757,n2758,n958);
wire s0n2758,s1n2758,notn2758;
or (n2758,s0n2758,s1n2758);
not(notn2758,n1066);
and (s0n2758,notn2758,n2759);
and (s1n2758,n1066,n2756);
and (n2760,n2761,n1079);
wire s0n2761,s1n2761,notn2761;
or (n2761,s0n2761,s1n2761);
not(notn2761,n1066);
and (s0n2761,notn2761,n2762);
and (s1n2761,n1066,n2759);
and (n2763,n2764,n981);
wire s0n2764,s1n2764,notn2764;
or (n2764,s0n2764,s1n2764);
not(notn2764,n1066);
and (s0n2764,notn2764,n2765);
and (s1n2764,n1066,n2762);
wire s0n2767,s1n2767,notn2767;
or (n2767,s0n2767,s1n2767);
not(notn2767,n28);
and (s0n2767,notn2767,n2768);
and (s1n2767,n28,n2827);
or (n2768,1'b0,n2769,n2785,n2798,n2813);
not (n2769,n2770);
or (n2770,n2771,n2772);
not (n2771,n1056);
not (n2772,n2773);
nand (n2773,n2774,n2779,n2781,n2783);
nor (n2774,n2775,n2777);
and (n2775,n995,n2776);
and (n2777,n979,n2778);
nand (n2779,n944,n2780);
nand (n2781,n1007,n2782);
nand (n2783,n1019,n2784);
not (n2785,n2786);
nand (n2786,n2787,n1041);
nand (n2787,n2788,n2792,n2794,n2796);
nor (n2788,n2789,n2790);
and (n2789,n995,n2778);
and (n2790,n979,n2791);
nand (n2792,n944,n2793);
nand (n2794,n1007,n2795);
nand (n2796,n1019,n2797);
and (n2798,n2799,n990);
or (n2799,1'b0,n2800,n2804,n2807,n2810);
and (n2800,n2801,n947);
wire s0n2801,s1n2801,notn2801;
or (n2801,s0n2801,s1n2801);
not(notn2801,n1066);
and (s0n2801,notn2801,n2802);
and (s1n2801,n1066,n2803);
and (n2804,n2805,n958);
wire s0n2805,s1n2805,notn2805;
or (n2805,s0n2805,s1n2805);
not(notn2805,n1066);
and (s0n2805,notn2805,n2806);
and (s1n2805,n1066,n2802);
and (n2807,n2808,n1079);
wire s0n2808,s1n2808,notn2808;
or (n2808,s0n2808,s1n2808);
not(notn2808,n1066);
and (s0n2808,notn2808,n2809);
and (s1n2808,n1066,n2806);
and (n2810,n2811,n981);
wire s0n2811,s1n2811,notn2811;
or (n2811,s0n2811,s1n2811);
not(notn2811,n1066);
and (s0n2811,notn2811,n2812);
and (s1n2811,n1066,n2809);
and (n2813,n2814,n970);
or (n2814,1'b0,n2815,n2818,n2821,n2824);
and (n2815,n2816,n947);
wire s0n2816,s1n2816,notn2816;
or (n2816,s0n2816,s1n2816);
not(notn2816,n1066);
and (s0n2816,notn2816,n2817);
and (s1n2816,n1066,n2812);
and (n2818,n2819,n958);
wire s0n2819,s1n2819,notn2819;
or (n2819,s0n2819,s1n2819);
not(notn2819,n1066);
and (s0n2819,notn2819,n2820);
and (s1n2819,n1066,n2817);
and (n2821,n2822,n1079);
wire s0n2822,s1n2822,notn2822;
or (n2822,s0n2822,s1n2822);
not(notn2822,n1066);
and (s0n2822,notn2822,n2823);
and (s1n2822,n1066,n2820);
and (n2824,n2825,n981);
wire s0n2825,s1n2825,notn2825;
or (n2825,s0n2825,s1n2825);
not(notn2825,n1066);
and (s0n2825,notn2825,n2826);
and (s1n2825,n1066,n2823);
and (n2828,n2767,n2829);
and (n2829,n2830,n2890);
wire s0n2830,s1n2830,notn2830;
or (n2830,s0n2830,s1n2830);
not(notn2830,n28);
and (s0n2830,notn2830,n2831);
and (s1n2830,n28,n2889);
or (n2831,1'b0,n2832,n2847,n2860,n2875);
not (n2832,n2833);
nand (n2833,n2834,n1056);
nand (n2834,n2835,n2840);
nor (n2835,n2836,n2838);
and (n2836,n1019,n2837);
and (n2838,n1007,n2839);
and (n2840,n2841,n2843,n2845);
nand (n2841,n995,n2842);
nand (n2843,n944,n2844);
nand (n2845,n979,n2846);
and (n2847,n2848,n1041);
nand (n2848,n2849,n2854);
nor (n2849,n2850,n2852);
and (n2850,n1007,n2851);
and (n2852,n1019,n2853);
and (n2854,n2855,n2856,n2858);
nand (n2855,n995,n2846);
nand (n2856,n944,n2857);
nand (n2858,n979,n2859);
and (n2860,n2861,n990);
or (n2861,1'b0,n2862,n2866,n2869,n2872);
and (n2862,n2863,n947);
wire s0n2863,s1n2863,notn2863;
or (n2863,s0n2863,s1n2863);
not(notn2863,n1066);
and (s0n2863,notn2863,n2864);
and (s1n2863,n1066,n2865);
and (n2866,n2867,n958);
wire s0n2867,s1n2867,notn2867;
or (n2867,s0n2867,s1n2867);
not(notn2867,n1066);
and (s0n2867,notn2867,n2868);
and (s1n2867,n1066,n2864);
and (n2869,n2870,n1079);
wire s0n2870,s1n2870,notn2870;
or (n2870,s0n2870,s1n2870);
not(notn2870,n1066);
and (s0n2870,notn2870,n2871);
and (s1n2870,n1066,n2868);
and (n2872,n2873,n981);
wire s0n2873,s1n2873,notn2873;
or (n2873,s0n2873,s1n2873);
not(notn2873,n1066);
and (s0n2873,notn2873,n2874);
and (s1n2873,n1066,n2871);
and (n2875,n2876,n970);
or (n2876,1'b0,n2877,n2880,n2883,n2886);
and (n2877,n2878,n947);
wire s0n2878,s1n2878,notn2878;
or (n2878,s0n2878,s1n2878);
not(notn2878,n1066);
and (s0n2878,notn2878,n2879);
and (s1n2878,n1066,n2874);
and (n2880,n2881,n958);
wire s0n2881,s1n2881,notn2881;
or (n2881,s0n2881,s1n2881);
not(notn2881,n1066);
and (s0n2881,notn2881,n2882);
and (s1n2881,n1066,n2879);
and (n2883,n2884,n1079);
wire s0n2884,s1n2884,notn2884;
or (n2884,s0n2884,s1n2884);
not(notn2884,n1066);
and (s0n2884,notn2884,n2885);
and (s1n2884,n1066,n2882);
and (n2886,n2887,n981);
wire s0n2887,s1n2887,notn2887;
or (n2887,s0n2887,s1n2887);
not(notn2887,n1066);
and (s0n2887,notn2887,n2888);
and (s1n2887,n1066,n2885);
wire s0n2890,s1n2890,notn2890;
or (n2890,s0n2890,s1n2890);
not(notn2890,n28);
and (s0n2890,notn2890,n2891);
and (s1n2890,n28,n2952);
or (n2891,1'b0,n2892,n2908,n2923,n2938);
and (n2892,n2893,n1056);
nand (n2893,n2894,n2899);
nor (n2894,n2895,n2897);
and (n2895,n1007,n2896);
and (n2897,n1019,n2898);
nor (n2899,n2900,n2902);
and (n2900,n944,n2901);
nand (n2902,n2903,n2906);
or (n2903,n2904,n1121);
not (n2904,n2905);
nand (n2906,n979,n2907);
and (n2908,n2909,n1041);
nand (n2909,n2910,n2915);
nor (n2910,n2911,n2913);
and (n2911,n1007,n2912);
and (n2913,n1019,n2914);
nor (n2915,n2916,n2918);
and (n2916,n944,n2917);
nand (n2918,n2919,n2921);
or (n2919,n2920,n1121);
not (n2920,n2907);
nand (n2921,n979,n2922);
and (n2923,n2924,n990);
or (n2924,1'b0,n2925,n2929,n2932,n2935);
and (n2925,n2926,n947);
wire s0n2926,s1n2926,notn2926;
or (n2926,s0n2926,s1n2926);
not(notn2926,n1066);
and (s0n2926,notn2926,n2927);
and (s1n2926,n1066,n2928);
and (n2929,n2930,n958);
wire s0n2930,s1n2930,notn2930;
or (n2930,s0n2930,s1n2930);
not(notn2930,n1066);
and (s0n2930,notn2930,n2931);
and (s1n2930,n1066,n2927);
and (n2932,n2933,n1079);
wire s0n2933,s1n2933,notn2933;
or (n2933,s0n2933,s1n2933);
not(notn2933,n1066);
and (s0n2933,notn2933,n2934);
and (s1n2933,n1066,n2931);
and (n2935,n2936,n981);
wire s0n2936,s1n2936,notn2936;
or (n2936,s0n2936,s1n2936);
not(notn2936,n1066);
and (s0n2936,notn2936,n2937);
and (s1n2936,n1066,n2934);
and (n2938,n2939,n970);
or (n2939,1'b0,n2940,n2943,n2946,n2949);
and (n2940,n2941,n947);
wire s0n2941,s1n2941,notn2941;
or (n2941,s0n2941,s1n2941);
not(notn2941,n1066);
and (s0n2941,notn2941,n2942);
and (s1n2941,n1066,n2937);
and (n2943,n2944,n958);
wire s0n2944,s1n2944,notn2944;
or (n2944,s0n2944,s1n2944);
not(notn2944,n1066);
and (s0n2944,notn2944,n2945);
and (s1n2944,n1066,n2942);
and (n2946,n2947,n1079);
wire s0n2947,s1n2947,notn2947;
or (n2947,s0n2947,s1n2947);
not(notn2947,n1066);
and (s0n2947,notn2947,n2948);
and (s1n2947,n1066,n2945);
and (n2949,n2950,n981);
wire s0n2950,s1n2950,notn2950;
or (n2950,s0n2950,s1n2950);
not(notn2950,n1066);
and (s0n2950,notn2950,n2951);
and (s1n2950,n1066,n2948);
and (n2953,n2707,n2829);
and (n2954,n2590,n2705);
and (n2955,n2465,n2588);
and (n2956,n2337,n2463);
and (n2957,n2229,n2335);
and (n2958,n2109,n2227);
and (n2959,n2003,n2107);
not (n2960,n2961);
nor (n2961,n2962,n3572);
and (n2962,n2963,n2969);
not (n2963,n2964);
xor (n2964,n2965,n2967);
wire s0n2965,s1n2965,notn2965;
or (n2965,s0n2965,s1n2965);
not(notn2965,n28);
and (s0n2965,notn2965,1'b0);
and (s1n2965,n28,n2966);
wire s0n2967,s1n2967,notn2967;
or (n2967,s0n2967,s1n2967);
not(notn2967,n28);
and (s0n2967,notn2967,1'b0);
and (s1n2967,n28,n2968);
not (n2969,n2970);
nand (n2970,n2971,n3564);
or (n2971,n2972,n3130);
not (n2972,n2973);
and (n2973,n2974,n3119);
nand (n2974,n2975,n3115);
not (n2975,n2976);
nand (n2976,n2977,n3113);
or (n2977,n2978,n3045);
not (n2978,n2979);
and (n2979,n2980,n3014);
wire s0n2980,s1n2980,notn2980;
or (n2980,s0n2980,s1n2980);
not(notn2980,n28);
and (s0n2980,notn2980,n2981);
and (s1n2980,n28,n3013);
or (n2981,1'b0,n2982,n2983,n2984,n2999);
and (n2982,n1225,n1056);
and (n2983,n1212,n1041);
and (n2984,n2985,n990);
or (n2985,1'b0,n2986,n2990,n2993,n2996);
and (n2986,n2987,n947);
wire s0n2987,s1n2987,notn2987;
or (n2987,s0n2987,s1n2987);
not(notn2987,n1066);
and (s0n2987,notn2987,n2988);
and (s1n2987,n1066,n2989);
and (n2990,n2991,n958);
wire s0n2991,s1n2991,notn2991;
or (n2991,s0n2991,s1n2991);
not(notn2991,n1066);
and (s0n2991,notn2991,n2992);
and (s1n2991,n1066,n2988);
and (n2993,n2994,n1079);
wire s0n2994,s1n2994,notn2994;
or (n2994,s0n2994,s1n2994);
not(notn2994,n1066);
and (s0n2994,notn2994,n2995);
and (s1n2994,n1066,n2992);
and (n2996,n2997,n981);
wire s0n2997,s1n2997,notn2997;
or (n2997,s0n2997,s1n2997);
not(notn2997,n1066);
and (s0n2997,notn2997,n2998);
and (s1n2997,n1066,n2995);
and (n2999,n3000,n970);
or (n3000,1'b0,n3001,n3004,n3007,n3010);
and (n3001,n3002,n947);
wire s0n3002,s1n3002,notn3002;
or (n3002,s0n3002,s1n3002);
not(notn3002,n1066);
and (s0n3002,notn3002,n3003);
and (s1n3002,n1066,n2998);
and (n3004,n3005,n958);
wire s0n3005,s1n3005,notn3005;
or (n3005,s0n3005,s1n3005);
not(notn3005,n1066);
and (s0n3005,notn3005,n3006);
and (s1n3005,n1066,n3003);
and (n3007,n3008,n1079);
wire s0n3008,s1n3008,notn3008;
or (n3008,s0n3008,s1n3008);
not(notn3008,n1066);
and (s0n3008,notn3008,n3009);
and (s1n3008,n1066,n3006);
and (n3010,n3011,n981);
wire s0n3011,s1n3011,notn3011;
or (n3011,s0n3011,s1n3011);
not(notn3011,n1066);
and (s0n3011,notn3011,n3012);
and (s1n3011,n1066,n3009);
or (n3014,n3015,n3017);
and (n3015,n28,n3016);
nand (n3017,n3018,n3031,n3032,n3033);
nand (n3018,n3019,n1056);
nand (n3019,n3020,n3022,n3024,n3029);
nand (n3020,n1007,n3021);
nand (n3022,n1019,n3023);
nor (n3024,n3025,n3027);
and (n3025,n995,n3026);
and (n3027,n979,n3028);
nand (n3029,n944,n3030);
nand (n3031,n1149,n970);
nand (n3032,n1162,n990);
nand (n3033,n3034,n1041);
nand (n3034,n3035,n3037,n3039,n3043);
nand (n3035,n1007,n3036);
nand (n3037,n1019,n3038);
nor (n3039,n3040,n3041);
and (n3040,n995,n3028);
and (n3041,n979,n3042);
nand (n3043,n944,n3044);
not (n3045,n3046);
nand (n3046,n3047,n3082);
not (n3047,n3048);
wire s0n3048,s1n3048,notn3048;
or (n3048,s0n3048,s1n3048);
not(notn3048,n28);
and (s0n3048,notn3048,n3049);
and (s1n3048,n28,n3081);
or (n3049,1'b0,n3050,n3051,n3052,n3067);
and (n3050,n1098,n1056);
and (n3051,n1111,n1041);
and (n3052,n3053,n990);
or (n3053,1'b0,n3054,n3058,n3061,n3064);
and (n3054,n3055,n947);
wire s0n3055,s1n3055,notn3055;
or (n3055,s0n3055,s1n3055);
not(notn3055,n1066);
and (s0n3055,notn3055,n3056);
and (s1n3055,n1066,n3057);
and (n3058,n3059,n958);
wire s0n3059,s1n3059,notn3059;
or (n3059,s0n3059,s1n3059);
not(notn3059,n1066);
and (s0n3059,notn3059,n3060);
and (s1n3059,n1066,n3056);
and (n3061,n3062,n1079);
wire s0n3062,s1n3062,notn3062;
or (n3062,s0n3062,s1n3062);
not(notn3062,n1066);
and (s0n3062,notn3062,n3063);
and (s1n3062,n1066,n3060);
and (n3064,n3065,n981);
wire s0n3065,s1n3065,notn3065;
or (n3065,s0n3065,s1n3065);
not(notn3065,n1066);
and (s0n3065,notn3065,n3066);
and (s1n3065,n1066,n3063);
and (n3067,n3068,n970);
or (n3068,1'b0,n3069,n3072,n3075,n3078);
and (n3069,n3070,n947);
wire s0n3070,s1n3070,notn3070;
or (n3070,s0n3070,s1n3070);
not(notn3070,n1066);
and (s0n3070,notn3070,n3071);
and (s1n3070,n1066,n3066);
and (n3072,n3073,n958);
wire s0n3073,s1n3073,notn3073;
or (n3073,s0n3073,s1n3073);
not(notn3073,n1066);
and (s0n3073,notn3073,n3074);
and (s1n3073,n1066,n3071);
and (n3075,n3076,n1079);
wire s0n3076,s1n3076,notn3076;
or (n3076,s0n3076,s1n3076);
not(notn3076,n1066);
and (s0n3076,notn3076,n3077);
and (s1n3076,n1066,n3074);
and (n3078,n3079,n981);
wire s0n3079,s1n3079,notn3079;
or (n3079,s0n3079,s1n3079);
not(notn3079,n1066);
and (s0n3079,notn3079,n3080);
and (s1n3079,n1066,n3077);
not (n3082,n3083);
wire s0n3083,s1n3083,notn3083;
or (n3083,s0n3083,s1n3083);
not(notn3083,n28);
and (s0n3083,notn3083,n3084);
and (s1n3083,n28,n3112);
nand (n3084,n3085,n3086,n3087,n3100);
nand (n3085,n1029,n970);
nand (n3086,n1045,n990);
nand (n3087,n3088,n1056);
nand (n3088,n3089,n3094,n3096,n3098);
nor (n3089,n3090,n3092);
and (n3090,n995,n3091);
and (n3092,n979,n3093);
nand (n3094,n944,n3095);
nand (n3096,n1007,n3097);
nand (n3098,n1019,n3099);
nand (n3100,n3101,n1041);
nand (n3101,n3102,n3106,n3108,n3110);
nor (n3102,n3103,n3104);
and (n3103,n995,n3093);
and (n3104,n979,n3105);
nand (n3106,n944,n3107);
nand (n3108,n1007,n3109);
nand (n3110,n1019,n3111);
not (n3113,n3114);
and (n3114,n3048,n3083);
nand (n3115,n3116,n3046);
nand (n3116,n3117,n3118);
not (n3117,n2980);
not (n3118,n3014);
and (n3119,n3120,n3125);
or (n3120,n3121,n3123);
wire s0n3121,s1n3121,notn3121;
or (n3121,s0n3121,s1n3121);
not(notn3121,n28);
and (s0n3121,notn3121,1'b0);
and (s1n3121,n28,n3122);
wire s0n3123,s1n3123,notn3123;
or (n3123,s0n3123,s1n3123);
not(notn3123,n28);
and (s0n3123,notn3123,1'b0);
and (s1n3123,n28,n3124);
or (n3125,n3126,n3128);
wire s0n3126,s1n3126,notn3126;
or (n3126,s0n3126,s1n3126);
not(notn3126,n28);
and (s0n3126,notn3126,1'b0);
and (s1n3126,n28,n3127);
wire s0n3128,s1n3128,notn3128;
or (n3128,s0n3128,s1n3128);
not(notn3128,n28);
and (s0n3128,notn3128,1'b0);
and (s1n3128,n28,n3129);
not (n3130,n3131);
nand (n3131,n3132,n3556);
or (n3132,n3133,n3414);
not (n3133,n3134);
nand (n3134,n3135,n3344);
nand (n3135,n3136,n3204,n3271);
nand (n3136,n3137,n3172);
not (n3137,n3138);
wire s0n3138,s1n3138,notn3138;
or (n3138,s0n3138,s1n3138);
not(notn3138,n28);
and (s0n3138,notn3138,n3139);
and (s1n3138,n28,n3171);
or (n3139,1'b0,n3140,n3141,n3142,n3157);
and (n3140,n1709,n1056);
and (n3141,n1725,n1041);
and (n3142,n3143,n990);
or (n3143,1'b0,n3144,n3148,n3151,n3154);
and (n3144,n3145,n947);
wire s0n3145,s1n3145,notn3145;
or (n3145,s0n3145,s1n3145);
not(notn3145,n1066);
and (s0n3145,notn3145,n3146);
and (s1n3145,n1066,n3147);
and (n3148,n3149,n958);
wire s0n3149,s1n3149,notn3149;
or (n3149,s0n3149,s1n3149);
not(notn3149,n1066);
and (s0n3149,notn3149,n3150);
and (s1n3149,n1066,n3146);
and (n3151,n3152,n1079);
wire s0n3152,s1n3152,notn3152;
or (n3152,s0n3152,s1n3152);
not(notn3152,n1066);
and (s0n3152,notn3152,n3153);
and (s1n3152,n1066,n3150);
and (n3154,n3155,n981);
wire s0n3155,s1n3155,notn3155;
or (n3155,s0n3155,s1n3155);
not(notn3155,n1066);
and (s0n3155,notn3155,n3156);
and (s1n3155,n1066,n3153);
and (n3157,n3158,n970);
or (n3158,1'b0,n3159,n3162,n3165,n3168);
and (n3159,n3160,n947);
wire s0n3160,s1n3160,notn3160;
or (n3160,s0n3160,s1n3160);
not(notn3160,n1066);
and (s0n3160,notn3160,n3161);
and (s1n3160,n1066,n3156);
and (n3162,n3163,n958);
wire s0n3163,s1n3163,notn3163;
or (n3163,s0n3163,s1n3163);
not(notn3163,n1066);
and (s0n3163,notn3163,n3164);
and (s1n3163,n1066,n3161);
and (n3165,n3166,n1079);
wire s0n3166,s1n3166,notn3166;
or (n3166,s0n3166,s1n3166);
not(notn3166,n1066);
and (s0n3166,notn3166,n3167);
and (s1n3166,n1066,n3164);
and (n3168,n3169,n981);
wire s0n3169,s1n3169,notn3169;
or (n3169,s0n3169,s1n3169);
not(notn3169,n1066);
and (s0n3169,notn3169,n3170);
and (s1n3169,n1066,n3167);
not (n3172,n3173);
or (n3173,n3174,n3176);
and (n3174,n28,n3175);
nand (n3176,n3177,n3178,n3191,n3192);
nand (n3177,n1623,n990);
nand (n3178,n3179,n1041);
nand (n3179,n3180,n3185,n3187,n3189);
nor (n3180,n3181,n3183);
and (n3181,n995,n3182);
and (n3183,n979,n3184);
nand (n3185,n944,n3186);
nand (n3187,n1007,n3188);
nand (n3189,n1019,n3190);
nand (n3191,n1636,n970);
nand (n3192,n3193,n1056);
nand (n3193,n3194,n3198,n3200,n3202);
nor (n3194,n3195,n3197);
and (n3195,n995,n3196);
and (n3197,n979,n3182);
nand (n3198,n944,n3199);
nand (n3200,n1007,n3201);
nand (n3202,n1019,n3203);
or (n3204,n3205,n3239);
wire s0n3205,s1n3205,notn3205;
or (n3205,s0n3205,s1n3205);
not(notn3205,n28);
and (s0n3205,notn3205,n3206);
and (s1n3205,n28,n3238);
or (n3206,1'b0,n3207,n3208,n3209,n3224);
and (n3207,n1833,n1056);
and (n3208,n1848,n1041);
and (n3209,n3210,n990);
or (n3210,1'b0,n3211,n3215,n3218,n3221);
and (n3211,n3212,n947);
wire s0n3212,s1n3212,notn3212;
or (n3212,s0n3212,s1n3212);
not(notn3212,n1066);
and (s0n3212,notn3212,n3213);
and (s1n3212,n1066,n3214);
and (n3215,n3216,n958);
wire s0n3216,s1n3216,notn3216;
or (n3216,s0n3216,s1n3216);
not(notn3216,n1066);
and (s0n3216,notn3216,n3217);
and (s1n3216,n1066,n3213);
and (n3218,n3219,n1079);
wire s0n3219,s1n3219,notn3219;
or (n3219,s0n3219,s1n3219);
not(notn3219,n1066);
and (s0n3219,notn3219,n3220);
and (s1n3219,n1066,n3217);
and (n3221,n3222,n981);
wire s0n3222,s1n3222,notn3222;
or (n3222,s0n3222,s1n3222);
not(notn3222,n1066);
and (s0n3222,notn3222,n3223);
and (s1n3222,n1066,n3220);
and (n3224,n3225,n970);
or (n3225,1'b0,n3226,n3229,n3232,n3235);
and (n3226,n3227,n947);
wire s0n3227,s1n3227,notn3227;
or (n3227,s0n3227,s1n3227);
not(notn3227,n1066);
and (s0n3227,notn3227,n3228);
and (s1n3227,n1066,n3223);
and (n3229,n3230,n958);
wire s0n3230,s1n3230,notn3230;
or (n3230,s0n3230,s1n3230);
not(notn3230,n1066);
and (s0n3230,notn3230,n3231);
and (s1n3230,n1066,n3228);
and (n3232,n3233,n1079);
wire s0n3233,s1n3233,notn3233;
or (n3233,s0n3233,s1n3233);
not(notn3233,n1066);
and (s0n3233,notn3233,n3234);
and (s1n3233,n1066,n3231);
and (n3235,n3236,n981);
wire s0n3236,s1n3236,notn3236;
or (n3236,s0n3236,s1n3236);
not(notn3236,n1066);
and (s0n3236,notn3236,n3237);
and (s1n3236,n1066,n3234);
not (n3239,n3240);
nor (n3240,n3241,n3269);
nand (n3241,n3242,n3255,n3256,n3257);
nand (n3242,n3243,n1056);
nand (n3243,n3244,n3246,n3248,n3253);
nand (n3244,n1007,n3245);
nand (n3246,n1019,n3247);
nor (n3248,n3249,n3251);
and (n3249,n995,n3250);
and (n3251,n979,n3252);
nand (n3253,n944,n3254);
nand (n3255,n1759,n970);
nand (n3256,n1746,n990);
nand (n3257,n3258,n1041);
nand (n3258,n3259,n3261,n3263,n3267);
nand (n3259,n1007,n3260);
nand (n3261,n1019,n3262);
nor (n3263,n3264,n3265);
and (n3264,n995,n3252);
and (n3265,n979,n3266);
nand (n3267,n944,n3268);
and (n3269,n28,n3270);
nand (n3271,n3272,n3342);
not (n3272,n3273);
and (n3273,n3274,n3308);
wire s0n3274,s1n3274,notn3274;
or (n3274,s0n3274,s1n3274);
not(notn3274,n28);
and (s0n3274,notn3274,n3275);
and (s1n3274,n28,n3307);
or (n3275,1'b0,n3276,n3277,n3278,n3293);
and (n3276,n1952,n1056);
and (n3277,n1968,n1041);
and (n3278,n3279,n990);
or (n3279,1'b0,n3280,n3284,n3287,n3290);
and (n3280,n3281,n947);
wire s0n3281,s1n3281,notn3281;
or (n3281,s0n3281,s1n3281);
not(notn3281,n1066);
and (s0n3281,notn3281,n3282);
and (s1n3281,n1066,n3283);
and (n3284,n3285,n958);
wire s0n3285,s1n3285,notn3285;
or (n3285,s0n3285,s1n3285);
not(notn3285,n1066);
and (s0n3285,notn3285,n3286);
and (s1n3285,n1066,n3282);
and (n3287,n3288,n1079);
wire s0n3288,s1n3288,notn3288;
or (n3288,s0n3288,s1n3288);
not(notn3288,n1066);
and (s0n3288,notn3288,n3289);
and (s1n3288,n1066,n3286);
and (n3290,n3291,n981);
wire s0n3291,s1n3291,notn3291;
or (n3291,s0n3291,s1n3291);
not(notn3291,n1066);
and (s0n3291,notn3291,n3292);
and (s1n3291,n1066,n3289);
and (n3293,n3294,n970);
or (n3294,1'b0,n3295,n3298,n3301,n3304);
and (n3295,n3296,n947);
wire s0n3296,s1n3296,notn3296;
or (n3296,s0n3296,s1n3296);
not(notn3296,n1066);
and (s0n3296,notn3296,n3297);
and (s1n3296,n1066,n3292);
and (n3298,n3299,n958);
wire s0n3299,s1n3299,notn3299;
or (n3299,s0n3299,s1n3299);
not(notn3299,n1066);
and (s0n3299,notn3299,n3300);
and (s1n3299,n1066,n3297);
and (n3301,n3302,n1079);
wire s0n3302,s1n3302,notn3302;
or (n3302,s0n3302,s1n3302);
not(notn3302,n1066);
and (s0n3302,notn3302,n3303);
and (s1n3302,n1066,n3300);
and (n3304,n3305,n981);
wire s0n3305,s1n3305,notn3305;
or (n3305,s0n3305,s1n3305);
not(notn3305,n1066);
and (s0n3305,notn3305,n3306);
and (s1n3305,n1066,n3303);
wire s0n3308,s1n3308,notn3308;
or (n3308,s0n3308,s1n3308);
not(notn3308,n28);
and (s0n3308,notn3308,n3309);
and (s1n3308,n28,n3341);
nand (n3309,n3310,n3327,n3328,n3329);
nand (n3310,n3311,n1056);
nand (n3311,n3312,n3317);
nor (n3312,n3313,n3315);
and (n3313,n1007,n3314);
and (n3315,n1019,n3316);
nor (n3317,n3318,n3324);
nand (n3318,n3319,n3322);
or (n3319,n3320,n1121);
not (n3320,n3321);
nand (n3322,n979,n3323);
nor (n3324,n3325,n1127);
not (n3325,n3326);
nand (n3327,n1866,n990);
nand (n3328,n1879,n970);
nand (n3329,n3330,n1041);
nand (n3330,n3331,n3335,n3337,n3339);
nor (n3331,n3332,n3334);
and (n3332,n979,n3333);
and (n3334,n995,n3323);
nand (n3335,n944,n3336);
nand (n3337,n1007,n3338);
nand (n3339,n1019,n3340);
not (n3342,n3343);
and (n3343,n3205,n3239);
and (n3344,n3345,n3412);
not (n3345,n3346);
and (n3346,n3347,n3381);
wire s0n3347,s1n3347,notn3347;
or (n3347,s0n3347,s1n3347);
not(notn3347,n28);
and (s0n3347,notn3347,n3348);
and (s1n3347,n28,n3380);
or (n3348,1'b0,n3349,n3350,n3351,n3366);
and (n3349,n1585,n1056);
and (n3350,n1601,n1041);
and (n3351,n3352,n990);
or (n3352,1'b0,n3353,n3357,n3360,n3363);
and (n3353,n3354,n947);
wire s0n3354,s1n3354,notn3354;
or (n3354,s0n3354,s1n3354);
not(notn3354,n1066);
and (s0n3354,notn3354,n3355);
and (s1n3354,n1066,n3356);
and (n3357,n3358,n958);
wire s0n3358,s1n3358,notn3358;
or (n3358,s0n3358,s1n3358);
not(notn3358,n1066);
and (s0n3358,notn3358,n3359);
and (s1n3358,n1066,n3355);
and (n3360,n3361,n1079);
wire s0n3361,s1n3361,notn3361;
or (n3361,s0n3361,s1n3361);
not(notn3361,n1066);
and (s0n3361,notn3361,n3362);
and (s1n3361,n1066,n3359);
and (n3363,n3364,n981);
wire s0n3364,s1n3364,notn3364;
or (n3364,s0n3364,s1n3364);
not(notn3364,n1066);
and (s0n3364,notn3364,n3365);
and (s1n3364,n1066,n3362);
and (n3366,n3367,n970);
or (n3367,1'b0,n3368,n3371,n3374,n3377);
and (n3368,n3369,n947);
wire s0n3369,s1n3369,notn3369;
or (n3369,s0n3369,s1n3369);
not(notn3369,n1066);
and (s0n3369,notn3369,n3370);
and (s1n3369,n1066,n3365);
and (n3371,n3372,n958);
wire s0n3372,s1n3372,notn3372;
or (n3372,s0n3372,s1n3372);
not(notn3372,n1066);
and (s0n3372,notn3372,n3373);
and (s1n3372,n1066,n3370);
and (n3374,n3375,n1079);
wire s0n3375,s1n3375,notn3375;
or (n3375,s0n3375,s1n3375);
not(notn3375,n1066);
and (s0n3375,notn3375,n3376);
and (s1n3375,n1066,n3373);
and (n3377,n3378,n981);
wire s0n3378,s1n3378,notn3378;
or (n3378,s0n3378,s1n3378);
not(notn3378,n1066);
and (s0n3378,notn3378,n3379);
and (s1n3378,n1066,n3376);
or (n3381,n3382,n3384);
and (n3382,n28,n3383);
nand (n3384,n3385,n3398,n3399,n3400);
nand (n3385,n3386,n1056);
nand (n3386,n3387,n3392,n3394,n3396);
nor (n3387,n3388,n3390);
and (n3388,n995,n3389);
and (n3390,n979,n3391);
nand (n3392,n944,n3393);
nand (n3394,n1007,n3395);
nand (n3396,n1019,n3397);
nand (n3398,n1499,n990);
nand (n3399,n1512,n970);
nand (n3400,n3401,n1041);
nand (n3401,n3402,n3406,n3408,n3410);
nor (n3402,n3403,n3404);
and (n3403,n995,n3391);
and (n3404,n979,n3405);
nand (n3406,n944,n3407);
nand (n3408,n1007,n3409);
nand (n3410,n1019,n3411);
not (n3412,n3413);
and (n3413,n3138,n3173);
not (n3414,n3415);
nor (n3415,n3416,n3417);
nor (n3416,n3347,n3381);
nand (n3417,n3418,n3485);
nand (n3418,n3419,n3454);
not (n3419,n3420);
wire s0n3420,s1n3420,notn3420;
or (n3420,s0n3420,s1n3420);
not(notn3420,n28);
and (s0n3420,notn3420,n3421);
and (s1n3420,n28,n3453);
or (n3421,1'b0,n3422,n3423,n3424,n3439);
and (n3422,n1346,n1056);
and (n3423,n1362,n1041);
and (n3424,n3425,n990);
or (n3425,1'b0,n3426,n3430,n3433,n3436);
and (n3426,n3427,n947);
wire s0n3427,s1n3427,notn3427;
or (n3427,s0n3427,s1n3427);
not(notn3427,n1066);
and (s0n3427,notn3427,n3428);
and (s1n3427,n1066,n3429);
and (n3430,n3431,n958);
wire s0n3431,s1n3431,notn3431;
or (n3431,s0n3431,s1n3431);
not(notn3431,n1066);
and (s0n3431,notn3431,n3432);
and (s1n3431,n1066,n3428);
and (n3433,n3434,n1079);
wire s0n3434,s1n3434,notn3434;
or (n3434,s0n3434,s1n3434);
not(notn3434,n1066);
and (s0n3434,notn3434,n3435);
and (s1n3434,n1066,n3432);
and (n3436,n3437,n981);
wire s0n3437,s1n3437,notn3437;
or (n3437,s0n3437,s1n3437);
not(notn3437,n1066);
and (s0n3437,notn3437,n3438);
and (s1n3437,n1066,n3435);
and (n3439,n3440,n970);
or (n3440,1'b0,n3441,n3444,n3447,n3450);
and (n3441,n3442,n947);
wire s0n3442,s1n3442,notn3442;
or (n3442,s0n3442,s1n3442);
not(notn3442,n1066);
and (s0n3442,notn3442,n3443);
and (s1n3442,n1066,n3438);
and (n3444,n3445,n958);
wire s0n3445,s1n3445,notn3445;
or (n3445,s0n3445,s1n3445);
not(notn3445,n1066);
and (s0n3445,notn3445,n3446);
and (s1n3445,n1066,n3443);
and (n3447,n3448,n1079);
wire s0n3448,s1n3448,notn3448;
or (n3448,s0n3448,s1n3448);
not(notn3448,n1066);
and (s0n3448,notn3448,n3449);
and (s1n3448,n1066,n3446);
and (n3450,n3451,n981);
wire s0n3451,s1n3451,notn3451;
or (n3451,s0n3451,s1n3451);
not(notn3451,n1066);
and (s0n3451,notn3451,n3452);
and (s1n3451,n1066,n3449);
not (n3454,n3455);
wire s0n3455,s1n3455,notn3455;
or (n3455,s0n3455,s1n3455);
not(notn3455,n28);
and (s0n3455,notn3455,n3456);
and (s1n3455,n28,n3484);
nand (n3456,n3457,n3470,n3471,n3472);
nand (n3457,n3458,n1056);
nand (n3458,n3459,n3464,n3466,n3468);
nor (n3459,n3460,n3462);
and (n3460,n995,n3461);
and (n3462,n979,n3463);
nand (n3464,n944,n3465);
nand (n3466,n1007,n3467);
nand (n3468,n1019,n3469);
nand (n3470,n1260,n990);
nand (n3471,n1273,n970);
nand (n3472,n3473,n1041);
nand (n3473,n3474,n3478,n3480,n3482);
nor (n3474,n3475,n3476);
and (n3475,n995,n3463);
and (n3476,n979,n3477);
nand (n3478,n944,n3479);
nand (n3480,n1007,n3481);
nand (n3482,n1019,n3483);
nand (n3485,n3486,n3521);
not (n3486,n3487);
wire s0n3487,s1n3487,notn3487;
or (n3487,s0n3487,s1n3487);
not(notn3487,n28);
and (s0n3487,notn3487,n3488);
and (s1n3487,n28,n3520);
or (n3488,1'b0,n3489,n3490,n3491,n3506);
and (n3489,n1465,n1056);
and (n3490,n1478,n1041);
and (n3491,n3492,n990);
or (n3492,1'b0,n3493,n3497,n3500,n3503);
and (n3493,n3494,n947);
wire s0n3494,s1n3494,notn3494;
or (n3494,s0n3494,s1n3494);
not(notn3494,n1066);
and (s0n3494,notn3494,n3495);
and (s1n3494,n1066,n3496);
and (n3497,n3498,n958);
wire s0n3498,s1n3498,notn3498;
or (n3498,s0n3498,s1n3498);
not(notn3498,n1066);
and (s0n3498,notn3498,n3499);
and (s1n3498,n1066,n3495);
and (n3500,n3501,n1079);
wire s0n3501,s1n3501,notn3501;
or (n3501,s0n3501,s1n3501);
not(notn3501,n1066);
and (s0n3501,notn3501,n3502);
and (s1n3501,n1066,n3499);
and (n3503,n3504,n981);
wire s0n3504,s1n3504,notn3504;
or (n3504,s0n3504,s1n3504);
not(notn3504,n1066);
and (s0n3504,notn3504,n3505);
and (s1n3504,n1066,n3502);
and (n3506,n3507,n970);
or (n3507,1'b0,n3508,n3511,n3514,n3517);
and (n3508,n3509,n947);
wire s0n3509,s1n3509,notn3509;
or (n3509,s0n3509,s1n3509);
not(notn3509,n1066);
and (s0n3509,notn3509,n3510);
and (s1n3509,n1066,n3505);
and (n3511,n3512,n958);
wire s0n3512,s1n3512,notn3512;
or (n3512,s0n3512,s1n3512);
not(notn3512,n1066);
and (s0n3512,notn3512,n3513);
and (s1n3512,n1066,n3510);
and (n3514,n3515,n1079);
wire s0n3515,s1n3515,notn3515;
or (n3515,s0n3515,s1n3515);
not(notn3515,n1066);
and (s0n3515,notn3515,n3516);
and (s1n3515,n1066,n3513);
and (n3517,n3518,n981);
wire s0n3518,s1n3518,notn3518;
or (n3518,s0n3518,s1n3518);
not(notn3518,n1066);
and (s0n3518,notn3518,n3519);
and (s1n3518,n1066,n3516);
not (n3521,n3522);
nand (n3522,n3523,n3527);
or (n3523,n3524,n3526);
not (n3524,n3525);
not (n3526,n28);
not (n3527,n3528);
nand (n3528,n3529,n3530,n3543,n3544);
nand (n3529,n1403,n970);
nand (n3530,n3531,n1056);
nand (n3531,n3532,n3537,n3539,n3541);
nor (n3532,n3533,n3535);
and (n3533,n995,n3534);
and (n3535,n979,n3536);
nand (n3537,n944,n3538);
nand (n3539,n1007,n3540);
nand (n3541,n1019,n3542);
nand (n3543,n1416,n990);
nand (n3544,n3545,n1041);
nand (n3545,n3546,n3550,n3552,n3554);
nor (n3546,n3547,n3548);
and (n3547,n995,n3536);
and (n3548,n979,n3549);
nand (n3550,n944,n3551);
nand (n3552,n1007,n3553);
nand (n3554,n1019,n3555);
nor (n3556,n2976,n3557);
nand (n3557,n3558,n3562);
or (n3558,n3559,n3561);
not (n3559,n3560);
and (n3560,n3487,n3522);
not (n3561,n3418);
not (n3562,n3563);
and (n3563,n3420,n3455);
not (n3564,n3565);
nand (n3565,n3566,n3570);
or (n3566,n3567,n3568);
not (n3567,n3125);
not (n3568,n3569);
and (n3569,n3123,n3121);
not (n3570,n3571);
and (n3571,n3128,n3126);
and (n3572,n2964,n2970);
or (n3573,n3574,n3593,n3683);
and (n3574,n3575,n3577);
xor (n3575,n3576,n2107);
xor (n3576,n2003,n2054);
not (n3577,n3578);
nor (n3578,n3579,n3590);
and (n3579,n3580,n3581);
xor (n3580,n3128,n3126);
nand (n3581,n3582,n3587,n3589);
nand (n3582,n3134,n3583,n3585,n3586);
and (n3583,n3584,n3120);
not (n3584,n3416);
not (n3585,n3115);
not (n3586,n3417);
nor (n3587,n3588,n3569);
and (n3588,n2976,n3120);
nand (n3589,n3557,n3585,n3120);
and (n3590,n3591,n3592);
not (n3591,n3580);
not (n3592,n3581);
and (n3593,n3577,n3594);
or (n3594,n3595,n3608,n3682);
and (n3595,n3596,n3598);
xor (n3596,n3597,n2227);
xor (n3597,n2109,n2161);
not (n3598,n3599);
nand (n3599,n3600,n3607);
or (n3600,n3601,n3602);
xor (n3601,n3123,n3121);
not (n3602,n3603);
nand (n3603,n3604,n3606);
nor (n3604,n3605,n2976);
and (n3605,n3557,n3585);
nand (n3606,n3134,n3415,n3585);
nand (n3607,n3602,n3601);
and (n3608,n3598,n3609);
or (n3609,n3610,n3633,n3681);
and (n3610,n3611,n3613);
xor (n3611,n3612,n2335);
xor (n3612,n2229,n2282);
not (n3613,n3614);
xor (n3614,n3615,n3616);
xor (n3615,n3048,n3083);
nand (n3616,n3617,n3631);
or (n3617,n3618,n3621);
not (n3618,n3619);
nor (n3619,n3620,n3417);
not (n3620,n3116);
not (n3621,n3622);
or (n3622,n3346,n3623,n3630);
and (n3623,n3381,n3624);
or (n3624,n3413,n3625,n3629);
and (n3625,n3173,n3626);
or (n3626,n3343,n3627,n3628);
and (n3627,n3239,n3273);
and (n3628,n3205,n3273);
and (n3629,n3138,n3626);
and (n3630,n3347,n3624);
nor (n3631,n3632,n2979);
and (n3632,n3557,n3116);
and (n3633,n3613,n3634);
or (n3634,n3635,n3647,n3680);
and (n3635,n3636,n3638);
xor (n3636,n3637,n2463);
xor (n3637,n2337,n2402);
not (n3638,n3639);
xor (n3639,n3640,n3641);
xor (n3640,n2980,n3014);
or (n3641,n3563,n3642,n3646);
and (n3642,n3455,n3643);
or (n3643,n3560,n3644,n3645);
and (n3644,n3522,n3622);
and (n3645,n3487,n3622);
and (n3646,n3420,n3643);
and (n3647,n3638,n3648);
or (n3648,n3649,n3655,n3679);
and (n3649,n3650,n3652);
xor (n3650,n3651,n2588);
xor (n3651,n2465,n2530);
not (n3652,n3653);
xor (n3653,n3654,n3643);
xor (n3654,n3420,n3455);
and (n3655,n3652,n3656);
or (n3656,n3657,n3663,n3678);
and (n3657,n3658,n3660);
xor (n3658,n3659,n2705);
xor (n3659,n2590,n2647);
not (n3660,n3661);
xor (n3661,n3662,n3622);
xor (n3662,n3487,n3522);
and (n3663,n3660,n3664);
or (n3664,n3665,n3671,n3677);
and (n3665,n3666,n3668);
xor (n3666,n3667,n2829);
xor (n3667,n2707,n2767);
not (n3668,n3669);
xor (n3669,n3670,n3624);
xor (n3670,n3347,n3381);
and (n3671,n3668,n3672);
and (n3672,n3673,n3674);
xor (n3673,n2830,n2890);
not (n3674,n3675);
xor (n3675,n3676,n3626);
xor (n3676,n3138,n3173);
and (n3677,n3666,n3672);
and (n3678,n3658,n3664);
and (n3679,n3650,n3656);
and (n3680,n3636,n3648);
and (n3681,n3611,n3634);
and (n3682,n3596,n3609);
and (n3683,n3575,n3594);
and (n3684,n3685,n3687);
xor (n3685,n3686,n3594);
xor (n3686,n3575,n3577);
and (n3687,n3688,n3690);
xor (n3688,n3689,n3609);
xor (n3689,n3596,n3598);
and (n3690,n3691,n3693);
xor (n3691,n3692,n3634);
xor (n3692,n3611,n3613);
and (n3693,n3694,n3696);
xor (n3694,n3695,n3648);
xor (n3695,n3636,n3638);
and (n3696,n3697,n3699);
xor (n3697,n3698,n3656);
xor (n3698,n3650,n3652);
and (n3699,n3700,n3702);
xor (n3700,n3701,n3664);
xor (n3701,n3658,n3660);
and (n3702,n3703,n3705);
xor (n3703,n3704,n3672);
xor (n3704,n3666,n3668);
and (n3705,n3706,n3707);
xor (n3706,n3673,n3674);
and (n3707,n3708,n3711);
not (n3708,n3709);
xor (n3709,n3710,n3273);
xor (n3710,n3205,n3239);
not (n3711,n3712);
xor (n3712,n3274,n3308);
or (n3713,n3714,n3718,n3777);
and (n3714,n3715,n3717);
xor (n3715,n3716,n928);
xor (n3716,n923,n925);
xor (n3717,n3685,n3687);
and (n3718,n3717,n3719);
or (n3719,n3720,n3724,n3776);
and (n3720,n3721,n3723);
xor (n3721,n3722,n935);
xor (n3722,n930,n932);
xor (n3723,n3688,n3690);
and (n3724,n3723,n3725);
or (n3725,n3726,n3730,n3775);
and (n3726,n3727,n3729);
xor (n3727,n3728,n1130);
xor (n3728,n937,n1058);
xor (n3729,n3691,n3693);
and (n3730,n3729,n3731);
or (n3731,n3732,n3736,n3774);
and (n3732,n3733,n3735);
xor (n3733,n3734,n1255);
xor (n3734,n1132,n1185);
xor (n3735,n3694,n3696);
and (n3736,n3735,n3737);
or (n3737,n3738,n3742,n3773);
and (n3738,n3739,n3741);
xor (n3739,n3740,n1379);
xor (n3740,n1257,n1314);
xor (n3741,n3697,n3699);
and (n3742,n3741,n3743);
or (n3743,n3744,n3748,n3772);
and (n3744,n3745,n3747);
xor (n3745,n3746,n1494);
xor (n3746,n1381,n1433);
xor (n3747,n3700,n3702);
and (n3748,n3747,n3749);
or (n3749,n3750,n3754,n3771);
and (n3750,n3751,n3753);
xor (n3751,n3752,n1618);
xor (n3752,n1496,n1553);
xor (n3753,n3703,n3705);
and (n3754,n3753,n3755);
or (n3755,n3756,n3760,n3770);
and (n3756,n3757,n3759);
xor (n3757,n3758,n1741);
xor (n3758,n1620,n1677);
xor (n3759,n3706,n3707);
and (n3760,n3759,n3761);
or (n3761,n3762,n3766,n3769);
and (n3762,n3763,n3765);
xor (n3763,n3764,n1862);
xor (n3764,n1743,n1800);
xor (n3765,n3708,n3711);
and (n3766,n3765,n3767);
and (n3767,n3768,n3712);
xor (n3768,n1863,n1920);
and (n3769,n3763,n3767);
and (n3770,n3757,n3761);
and (n3771,n3751,n3755);
and (n3772,n3745,n3749);
and (n3773,n3739,n3743);
and (n3774,n3733,n3737);
and (n3775,n3727,n3731);
and (n3776,n3721,n3725);
and (n3777,n3715,n3719);
or (n3778,n3779,n3782,n3822);
and (n3779,n3780,n3729);
xor (n3780,n3781,n3719);
xor (n3781,n3715,n3717);
and (n3782,n3729,n3783);
or (n3783,n3784,n3787,n3821);
and (n3784,n3785,n3735);
xor (n3785,n3786,n3725);
xor (n3786,n3721,n3723);
and (n3787,n3735,n3788);
or (n3788,n3789,n3792,n3820);
and (n3789,n3790,n3741);
xor (n3790,n3791,n3731);
xor (n3791,n3727,n3729);
and (n3792,n3741,n3793);
or (n3793,n3794,n3797,n3819);
and (n3794,n3795,n3747);
xor (n3795,n3796,n3737);
xor (n3796,n3733,n3735);
and (n3797,n3747,n3798);
or (n3798,n3799,n3802,n3818);
and (n3799,n3800,n3753);
xor (n3800,n3801,n3743);
xor (n3801,n3739,n3741);
and (n3802,n3753,n3803);
or (n3803,n3804,n3807,n3817);
and (n3804,n3805,n3759);
xor (n3805,n3806,n3749);
xor (n3806,n3745,n3747);
and (n3807,n3759,n3808);
or (n3808,n3809,n3812,n3816);
and (n3809,n3810,n3765);
xor (n3810,n3811,n3755);
xor (n3811,n3751,n3753);
and (n3812,n3765,n3813);
and (n3813,n3814,n3712);
xor (n3814,n3815,n3761);
xor (n3815,n3757,n3759);
and (n3816,n3810,n3813);
and (n3817,n3805,n3808);
and (n3818,n3800,n3803);
and (n3819,n3795,n3798);
and (n3820,n3790,n3793);
and (n3821,n3785,n3788);
and (n3822,n3780,n3783);
and (n3823,n3824,n3826);
xor (n3824,n3825,n3783);
xor (n3825,n3780,n3729);
and (n3826,n3827,n3829);
xor (n3827,n3828,n3788);
xor (n3828,n3785,n3735);
and (n3829,n3830,n3832);
xor (n3830,n3831,n3793);
xor (n3831,n3790,n3741);
and (n3832,n3833,n3835);
xor (n3833,n3834,n3798);
xor (n3834,n3795,n3747);
and (n3835,n3836,n3838);
xor (n3836,n3837,n3803);
xor (n3837,n3800,n3753);
xor (n3838,n3839,n3808);
xor (n3839,n3805,n3759);
xor (n3840,n20,n3824);
wire s0n3841,s1n3841,notn3841;
or (n3841,s0n3841,s1n3841);
not(notn3841,n28);
and (s0n3841,notn3841,n3842);
and (s1n3841,n28,n4496);
xor (n3842,n3843,n4483);
xor (n3843,n3844,n4334);
xor (n3844,n3845,n3966);
xor (n3845,n3846,n3959);
xor (n3846,n3847,n3915);
xor (n3847,n3848,n3874);
xor (n3848,n3849,n3854);
xor (n3849,n3850,n3852);
wire s0n3850,s1n3850,notn3850;
or (n3850,s0n3850,s1n3850);
not(notn3850,n28);
and (s0n3850,notn3850,1'b0);
and (s1n3850,n28,n3851);
wire s0n3852,s1n3852,notn3852;
or (n3852,s0n3852,s1n3852);
not(notn3852,n28);
and (s0n3852,notn3852,1'b0);
and (s1n3852,n28,n3853);
or (n3854,n3855,n3860,n3873);
and (n3855,n3856,n3858);
wire s0n3856,s1n3856,notn3856;
or (n3856,s0n3856,s1n3856);
not(notn3856,n28);
and (s0n3856,notn3856,1'b0);
and (s1n3856,n28,n3857);
wire s0n3858,s1n3858,notn3858;
or (n3858,s0n3858,s1n3858);
not(notn3858,n28);
and (s0n3858,notn3858,1'b0);
and (s1n3858,n28,n3859);
and (n3860,n3858,n3861);
or (n3861,n3862,n3867,n3872);
and (n3862,n3863,n3865);
wire s0n3863,s1n3863,notn3863;
or (n3863,s0n3863,s1n3863);
not(notn3863,n28);
and (s0n3863,notn3863,1'b0);
and (s1n3863,n28,n3864);
wire s0n3865,s1n3865,notn3865;
or (n3865,s0n3865,s1n3865);
not(notn3865,n28);
and (s0n3865,notn3865,1'b0);
and (s1n3865,n28,n3866);
and (n3867,n3865,n3868);
or (n3868,n3869,n3870,n3871);
and (n3869,n1997,n1999);
and (n3870,n1999,n2001);
and (n3871,n1997,n2001);
and (n3872,n3863,n3868);
and (n3873,n3856,n3861);
not (n3874,n3875);
nor (n3875,n3876,n3912);
and (n3876,n3877,n3907);
nand (n3877,n3878,n3896);
or (n3878,n3879,n3602);
not (n3879,n3880);
nor (n3880,n3881,n3887);
not (n3881,n3882);
or (n3882,n3883,n3885);
wire s0n3883,s1n3883,notn3883;
or (n3883,s0n3883,s1n3883);
not(notn3883,n28);
and (s0n3883,notn3883,1'b0);
and (s1n3883,n28,n3884);
wire s0n3885,s1n3885,notn3885;
or (n3885,s0n3885,s1n3885);
not(notn3885,n28);
and (s0n3885,notn3885,1'b0);
and (s1n3885,n28,n3886);
not (n3887,n3888);
and (n3888,n3119,n3889);
nor (n3889,n3890,n3895);
nor (n3890,n3891,n3893);
wire s0n3891,s1n3891,notn3891;
or (n3891,s0n3891,s1n3891);
not(notn3891,n28);
and (s0n3891,notn3891,1'b0);
and (s1n3891,n28,n3892);
wire s0n3893,s1n3893,notn3893;
or (n3893,s0n3893,s1n3893);
not(notn3893,n28);
and (s0n3893,notn3893,1'b0);
and (s1n3893,n28,n3894);
nor (n3895,n2967,n2965);
nor (n3896,n3897,n3906);
and (n3897,n3898,n3882);
nand (n3898,n3899,n3901);
or (n3899,n3900,n3564);
not (n3900,n3889);
nor (n3901,n3902,n3905);
and (n3902,n3903,n3904);
not (n3903,n3890);
and (n3904,n2965,n2967);
and (n3905,n3893,n3891);
and (n3906,n3885,n3883);
xor (n3907,n3908,n3910);
wire s0n3908,s1n3908,notn3908;
or (n3908,s0n3908,s1n3908);
not(notn3908,n28);
and (s0n3908,notn3908,1'b0);
and (s1n3908,n28,n3909);
wire s0n3910,s1n3910,notn3910;
or (n3910,s0n3910,s1n3910);
not(notn3910,n28);
and (s0n3910,notn3910,1'b0);
and (s1n3910,n28,n3911);
and (n3912,n3913,n3914);
not (n3913,n3877);
not (n3914,n3907);
or (n3915,n3916,n3931,n3958);
and (n3916,n3917,n3919);
xor (n3917,n3918,n3861);
xor (n3918,n3856,n3858);
not (n3919,n3920);
nor (n3920,n3921,n3930);
and (n3921,n3922,n3924);
not (n3922,n3923);
xor (n3923,n3885,n3883);
not (n3924,n3925);
nand (n3925,n3926,n3929);
or (n3926,n3927,n3130);
not (n3927,n3928);
and (n3928,n2974,n3888);
not (n3929,n3898);
and (n3930,n3923,n3925);
and (n3931,n3919,n3932);
or (n3932,n3933,n3952,n3957);
and (n3933,n3934,n3936);
xor (n3934,n3935,n3868);
xor (n3935,n3863,n3865);
not (n3936,n3937);
nor (n3937,n3938,n3949);
and (n3938,n3939,n3940);
xor (n3939,n3893,n3891);
nand (n3940,n3941,n3946);
or (n3941,n3942,n3130);
not (n3942,n3943);
and (n3943,n2974,n3944);
nor (n3944,n3945,n3895);
not (n3945,n3119);
nor (n3946,n3947,n3904);
and (n3947,n3565,n3948);
not (n3948,n3895);
and (n3949,n3950,n3951);
not (n3950,n3939);
not (n3951,n3940);
and (n3952,n3936,n3953);
or (n3953,n3954,n3955,n3956);
and (n3954,n1995,n2960);
and (n3955,n2960,n3573);
and (n3956,n1995,n3573);
and (n3957,n3934,n3953);
and (n3958,n3917,n3932);
and (n3959,n3960,n3962);
xor (n3960,n3961,n3932);
xor (n3961,n3917,n3919);
and (n3962,n3963,n3965);
xor (n3963,n3964,n3953);
xor (n3964,n3934,n3936);
and (n3965,n1993,n3684);
nand (n3966,n3967,n4333);
or (n3967,n3968,n4067);
not (n3968,n3969);
nor (n3969,n3970,n4063);
not (n3970,n3971);
nand (n3971,n3972,n4040);
xor (n3972,n3973,n4027);
xor (n3973,n3974,n4006);
xor (n3974,n3975,n3980);
xor (n3975,n3976,n3978);
wire s0n3976,s1n3976,notn3976;
or (n3976,s0n3976,s1n3976);
not(notn3976,n28);
and (s0n3976,notn3976,1'b0);
and (s1n3976,n28,n3977);
wire s0n3978,s1n3978,notn3978;
or (n3978,s0n3978,s1n3978);
not(notn3978,n28);
and (s0n3978,notn3978,1'b0);
and (s1n3978,n28,n3979);
not (n3980,n3981);
nor (n3981,n3982,n3994);
and (n3982,n3603,n3983);
nor (n3983,n3887,n3984);
nand (n3984,n3985,n3988);
not (n3985,n3986);
nand (n3986,n3987,n3882);
or (n3987,n3910,n3908);
not (n3988,n3989);
and (n3989,n3990,n3992);
wire s0n3990,s1n3990,notn3990;
or (n3990,s0n3990,s1n3990);
not(notn3990,n28);
and (s0n3990,notn3990,1'b0);
and (s1n3990,n28,n3991);
wire s0n3992,s1n3992,notn3992;
or (n3992,s0n3992,s1n3992);
not(notn3992,n28);
and (s0n3992,notn3992,1'b0);
and (s1n3992,n28,n3993);
nand (n3994,n3995,n3996);
or (n3995,n3929,n3984);
nor (n3996,n3997,n4004);
and (n3997,n3998,n3988);
nand (n3998,n3999,n4002);
or (n3999,n4000,n4001);
not (n4000,n3906);
not (n4001,n3987);
not (n4002,n4003);
and (n4003,n3908,n3910);
not (n4004,n4005);
or (n4005,n3992,n3990);
not (n4006,n4007);
or (n4007,n4008,n4026);
and (n4008,n4009,n4014);
xor (n4009,n4010,n4012);
wire s0n4010,s1n4010,notn4010;
or (n4010,s0n4010,s1n4010);
not(notn4010,n28);
and (s0n4010,notn4010,1'b0);
and (s1n4010,n28,n4011);
wire s0n4012,s1n4012,notn4012;
or (n4012,s0n4012,s1n4012);
not(notn4012,n28);
and (s0n4012,notn4012,1'b0);
and (s1n4012,n28,n4013);
not (n4014,n4015);
nand (n4015,n4016,n4025);
or (n4016,n4017,n4019);
not (n4017,n4018);
xor (n4018,n3990,n3992);
nand (n4019,n4020,n4023);
or (n4020,n4021,n3602);
not (n4021,n4022);
nor (n4022,n3887,n3986);
nor (n4023,n4024,n3998);
and (n4024,n3898,n3985);
nand (n4025,n4019,n4017);
and (n4026,n4010,n4012);
nand (n4027,n4028,n4039);
nand (n4028,n4029,n4036);
or (n4029,n4030,n4033);
not (n4030,n4031);
wire s0n4031,s1n4031,notn4031;
or (n4031,s0n4031,s1n4031);
not(notn4031,n28);
and (s0n4031,notn4031,1'b0);
and (s1n4031,n28,n4032);
or (n4033,n4034,n4035);
and (n4034,n3849,n3874);
and (n4035,n3850,n3852);
not (n4036,n4037);
wire s0n4037,s1n4037,notn4037;
or (n4037,s0n4037,s1n4037);
not(notn4037,n28);
and (s0n4037,notn4037,1'b0);
and (s1n4037,n28,n4038);
nand (n4039,n4030,n4033);
or (n4040,n4041,n4062);
and (n4041,n4042,n4050);
xor (n4042,n4043,n4044);
xor (n4043,n4009,n4014);
nor (n4044,n4045,n4049);
and (n4045,n4046,n4048);
not (n4046,n4047);
xor (n4047,n4031,n4037);
not (n4048,n4033);
and (n4049,n4047,n4033);
nand (n4050,n4051,n4058);
or (n4051,n4052,n4055);
not (n4052,n4053);
wire s0n4053,s1n4053,notn4053;
or (n4053,s0n4053,s1n4053);
not(notn4053,n28);
and (s0n4053,notn4053,1'b0);
and (s1n4053,n28,n4054);
not (n4055,n4056);
or (n4056,n4057,n3855);
and (n4057,n3918,n3919);
nand (n4058,n4059,n4060);
or (n4059,n4053,n4056);
wire s0n4060,s1n4060,notn4060;
or (n4060,s0n4060,s1n4060);
not(notn4060,n28);
and (s0n4060,notn4060,1'b0);
and (s1n4060,n28,n4061);
and (n4062,n4043,n4044);
not (n4063,n4064);
nand (n4064,n4065,n4066);
not (n4065,n3972);
not (n4066,n4040);
nand (n4067,n4068,n4309,n4323);
nand (n4068,n4069,n4140,n4258);
and (n4069,n4070,n4133);
and (n4070,n4071,n4115);
nand (n4071,n4072,n4099);
not (n4072,n4073);
xor (n4073,n4074,n4088);
xor (n4074,n4075,n4076);
xor (n4075,n3918,n3919);
nand (n4076,n4077,n4084);
or (n4077,n4078,n4081);
not (n4078,n4079);
wire s0n4079,s1n4079,notn4079;
or (n4079,s0n4079,s1n4079);
not(notn4079,n28);
and (s0n4079,notn4079,1'b0);
and (s1n4079,n28,n4080);
not (n4081,n4082);
or (n4082,n4083,n3869);
and (n4083,n1996,n2960);
nand (n4084,n4085,n4086);
or (n4085,n4079,n4082);
wire s0n4086,s1n4086,notn4086;
or (n4086,s0n4086,s1n4086);
not(notn4086,n28);
and (s0n4086,notn4086,1'b0);
and (s1n4086,n28,n4087);
nand (n4088,n4089,n4098);
or (n4089,n4090,n4096);
not (n4090,n4091);
xor (n4091,n4092,n4094);
wire s0n4092,s1n4092,notn4092;
or (n4092,s0n4092,s1n4092);
not(notn4092,n28);
and (s0n4092,notn4092,1'b0);
and (s1n4092,n28,n4093);
wire s0n4094,s1n4094,notn4094;
or (n4094,s0n4094,s1n4094);
not(notn4094,n28);
and (s0n4094,notn4094,1'b0);
and (s1n4094,n28,n4095);
or (n4096,n4097,n3862);
and (n4097,n3935,n3936);
nand (n4098,n4090,n4096);
not (n4099,n4100);
or (n4100,n4101,n4114);
and (n4101,n4102,n4109);
xor (n4102,n4103,n4104);
xor (n4103,n3935,n3936);
or (n4104,n4105,n4108);
and (n4105,n25,n4106);
or (n4106,n4107,n2002);
and (n4107,n3576,n3577);
and (n4108,n26,n919);
nand (n4109,n4110,n4113);
or (n4110,n4111,n4082);
not (n4111,n4112);
xor (n4112,n4079,n4086);
nand (n4113,n4111,n4082);
and (n4114,n4103,n4104);
nand (n4115,n4116,n4129);
not (n4116,n4117);
xor (n4117,n4118,n4125);
xor (n4118,n4119,n4120);
xor (n4119,n3849,n3874);
nand (n4120,n4121,n4124);
or (n4121,n4122,n4056);
not (n4122,n4123);
xor (n4123,n4053,n4060);
nand (n4124,n4122,n4056);
nand (n4125,n4126,n4128);
nand (n4126,n4127,n4094);
or (n4127,n4092,n4096);
nand (n4128,n4096,n4092);
not (n4129,n4130);
or (n4130,n4131,n4132);
and (n4131,n4074,n4088);
and (n4132,n4075,n4076);
nand (n4133,n4134,n4136);
not (n4134,n4135);
xor (n4135,n4042,n4050);
not (n4136,n4137);
or (n4137,n4138,n4139);
and (n4138,n4118,n4125);
and (n4139,n4119,n4120);
nand (n4140,n4141,n4251);
or (n4141,n4142,n4186);
not (n4142,n4143);
and (n4143,n4144,n4172);
nand (n4144,n4145,n4158);
not (n4145,n4146);
xor (n4146,n4147,n4155);
xor (n4147,n4148,n4149);
xor (n4148,n3637,n3638);
nand (n4149,n4150,n4154);
nand (n4150,n4151,n1314);
or (n4151,n1257,n4152);
or (n4152,n4153,n2589);
and (n4153,n3659,n3660);
nand (n4154,n4152,n1257);
xor (n4155,n3734,n4156);
or (n4156,n4157,n2464);
and (n4157,n3651,n3652);
not (n4158,n4159);
or (n4159,n4160,n4171);
and (n4160,n4161,n4167);
xor (n4161,n4162,n4163);
xor (n4162,n3651,n3652);
or (n4163,n4164,n1380);
and (n4164,n3746,n4165);
or (n4165,n4166,n2706);
and (n4166,n3667,n3668);
nand (n4167,n4168,n4170);
or (n4168,n4169,n4152);
not (n4169,n3740);
nand (n4170,n4169,n4152);
and (n4171,n4162,n4163);
nand (n4172,n4173,n4182);
not (n4173,n4174);
xor (n4174,n4175,n4179);
xor (n4175,n4176,n4177);
xor (n4176,n3612,n3613);
or (n4177,n4178,n1131);
and (n4178,n3734,n4156);
xor (n4179,n3728,n4180);
or (n4180,n4181,n2336);
and (n4181,n3637,n3638);
not (n4182,n4183);
or (n4183,n4184,n4185);
and (n4184,n4147,n4155);
and (n4185,n4148,n4149);
not (n4186,n4187);
nand (n4187,n4188,n4245);
or (n4188,n4189,n4228);
not (n4189,n4190);
or (n4190,n4191,n4227);
and (n4191,n4192,n4208);
xor (n4192,n4193,n4202);
or (n4193,n4194,n4201);
and (n4194,n4195,n4197);
xor (n4195,n4196,n1620);
xor (n4196,n1677,n2830);
nand (n4197,n4198,n4200);
or (n4198,n4199,n3674);
not (n4199,n2890);
nand (n4200,n4199,n3674);
and (n4201,n4196,n1620);
xor (n4202,n4203,n4206);
xor (n4203,n4204,n4205);
and (n4204,n1677,n2830);
xor (n4205,n3667,n3668);
xor (n4206,n3752,n4207);
and (n4207,n3674,n2890);
or (n4208,n4209,n4226);
and (n4209,n4210,n4225);
xor (n4210,n4211,n4213);
or (n4211,n4212,n1742);
and (n4212,n3764,n3708);
nand (n4213,n4214,n4224);
or (n4214,n4215,n4217);
nor (n4215,n4216,n3711);
xor (n4216,n3764,n3708);
nor (n4217,n4218,n4222);
nand (n4218,n4219,n4221);
or (n4219,n4220,n3711);
not (n4220,n1863);
not (n4221,n1862);
nor (n4222,n4223,n3711);
not (n4223,n1920);
nand (n4224,n4216,n3711);
xor (n4225,n4195,n4197);
and (n4226,n4211,n4213);
and (n4227,n4193,n4202);
not (n4228,n4229);
nor (n4229,n4230,n4240);
nor (n4230,n4231,n4232);
xor (n4231,n4161,n4167);
or (n4232,n4233,n4239);
and (n4233,n4234,n4238);
xor (n4234,n4235,n4236);
xor (n4235,n3659,n3660);
or (n4236,n4237,n1495);
and (n4237,n3752,n4207);
xor (n4238,n3746,n4165);
and (n4239,n4235,n4236);
nor (n4240,n4241,n4242);
xor (n4241,n4234,n4238);
or (n4242,n4243,n4244);
and (n4243,n4203,n4206);
and (n4244,n4204,n4205);
nor (n4245,n4246,n4250);
and (n4246,n4247,n4248);
not (n4247,n4230);
not (n4248,n4249);
nand (n4249,n4241,n4242);
and (n4250,n4231,n4232);
not (n4251,n4252);
nand (n4252,n4253,n4257);
or (n4253,n4254,n4256);
not (n4254,n4255);
and (n4255,n4146,n4159);
not (n4256,n4172);
nand (n4257,n4183,n4174);
and (n4258,n4259,n4290);
and (n4259,n4260,n4274);
nand (n4260,n4261,n4263);
not (n4261,n4262);
xor (n4262,n4102,n4109);
not (n4263,n4264);
or (n4264,n4265,n4273);
and (n4265,n4266,n4269);
xor (n4266,n4267,n4268);
xor (n4267,n1996,n2960);
xor (n4268,n25,n4106);
or (n4269,n4270,n922);
and (n4270,n3716,n4271);
or (n4271,n4272,n2108);
and (n4272,n3597,n3598);
and (n4273,n4267,n4268);
nand (n4274,n4275,n4277);
not (n4275,n4276);
xor (n4276,n4266,n4269);
not (n4277,n4278);
or (n4278,n4279,n4289);
and (n4279,n4280,n4283);
xor (n4280,n4281,n4282);
xor (n4281,n3576,n3577);
xor (n4282,n3716,n4271);
nand (n4283,n4284,n4288);
nand (n4284,n4285,n932);
or (n4285,n930,n4286);
or (n4286,n4287,n2228);
and (n4287,n3612,n3613);
nand (n4288,n4286,n930);
and (n4289,n4281,n4282);
nor (n4290,n4291,n4304);
nor (n4291,n4292,n4293);
xor (n4292,n4280,n4283);
or (n4293,n4294,n4303);
and (n4294,n4295,n4301);
xor (n4295,n4296,n4297);
xor (n4296,n3597,n3598);
nand (n4297,n4298,n4300);
or (n4298,n4299,n4286);
not (n4299,n3722);
nand (n4300,n4286,n4299);
or (n4301,n4302,n936);
and (n4302,n3728,n4180);
and (n4303,n4296,n4297);
nor (n4304,n4305,n4306);
xor (n4305,n4295,n4301);
or (n4306,n4307,n4308);
and (n4307,n4175,n4179);
and (n4308,n4176,n4177);
nand (n4309,n4069,n4310);
not (n4310,n4311);
nor (n4311,n4312,n4317);
and (n4312,n4259,n4313);
nand (n4313,n4314,n4316);
or (n4314,n4291,n4315);
nand (n4315,n4305,n4306);
nand (n4316,n4292,n4293);
nand (n4317,n4318,n4322);
or (n4318,n4319,n4321);
not (n4319,n4320);
nor (n4320,n4275,n4277);
not (n4321,n4260);
nand (n4322,n4262,n4264);
nor (n4323,n4324,n4332);
and (n4324,n4325,n4133);
not (n4325,n4326);
or (n4326,n4327,n4328);
not (n4327,n4115);
not (n4328,n4329);
nand (n4329,n4330,n4331);
nand (n4330,n4117,n4130);
nand (n4331,n4073,n4100);
and (n4332,n4135,n4137);
nand (n4333,n3968,n4067);
or (n4334,n4335,n4459,n4482);
and (n4335,n4336,n4445);
xor (n4336,n4337,n4438);
xor (n4337,n4338,n4354);
xor (n4338,n4047,n4339);
or (n4339,n4340,n4341,n4353);
and (n4340,n4053,n4060);
and (n4341,n4060,n4342);
or (n4342,n4343,n4344,n4352);
and (n4343,n4092,n4094);
and (n4344,n4094,n4345);
or (n4345,n4346,n4347,n4351);
and (n4346,n4079,n4086);
and (n4347,n4086,n4348);
or (n4348,n4108,n4349,n4350);
and (n4349,n919,n921);
and (n4350,n26,n921);
and (n4351,n4079,n4348);
and (n4352,n4092,n4345);
and (n4353,n4053,n4342);
nand (n4354,n4355,n4437);
or (n4355,n4356,n4362);
not (n4356,n4357);
nor (n4357,n4358,n4361);
not (n4358,n4359);
nand (n4359,n4360,n4048);
not (n4360,n4043);
nor (n4361,n4048,n4360);
nand (n4362,n4363,n4371,n4398);
not (n4363,n4364);
nand (n4364,n4365,n4370);
or (n4365,n4366,n4368);
not (n4366,n4367);
and (n4367,n4096,n4075);
not (n4368,n4369);
or (n4369,n4119,n4056);
nand (n4370,n4119,n4056);
nand (n4371,n4372,n4396);
not (n4372,n4373);
nor (n4373,n4374,n4390);
and (n4374,n4375,n4380);
and (n4375,n4376,n4377);
or (n4376,n4103,n4082);
nand (n4377,n4378,n4379);
not (n4378,n4267);
not (n4379,n4106);
not (n4380,n4381);
nor (n4381,n4382,n4389);
and (n4382,n4383,n4386);
nand (n4383,n4384,n4385);
not (n4384,n4271);
not (n4385,n4281);
nor (n4386,n4387,n4388);
not (n4387,n4286);
not (n4388,n4296);
nor (n4389,n4384,n4385);
nand (n4390,n4391,n4395);
or (n4391,n4392,n4394);
not (n4392,n4393);
nor (n4393,n4378,n4379);
not (n4394,n4376);
nand (n4395,n4103,n4082);
and (n4396,n4369,n4397);
or (n4397,n4075,n4096);
nand (n4398,n4399,n4403,n4396);
and (n4399,n4375,n4400);
nor (n4400,n4401,n4402);
not (n4401,n4383);
and (n4402,n4387,n4388);
nand (n4403,n4404,n4423);
nor (n4404,n4405,n4417);
and (n4405,n4406,n4411);
and (n4406,n4407,n4408);
or (n4407,n4176,n4180);
nand (n4408,n4409,n4410);
not (n4409,n4156);
not (n4410,n4148);
nor (n4411,n4412,n4415);
and (n4412,n4413,n4414);
nand (n4413,n4152,n4162);
nand (n4414,n4165,n4235);
not (n4415,n4416);
or (n4416,n4162,n4152);
nand (n4417,n4418,n4422);
or (n4418,n4419,n4421);
not (n4419,n4420);
nor (n4420,n4409,n4410);
not (n4421,n4407);
nand (n4422,n4176,n4180);
nand (n4423,n4406,n4424,n4426);
and (n4424,n4416,n4425);
or (n4425,n4165,n4235);
nand (n4426,n4427,n4433);
or (n4427,n4428,n4431);
not (n4428,n4429);
and (n4429,n4430,n3707);
or (n4430,n4197,n2830);
not (n4431,n4432);
or (n4432,n4205,n4207);
nor (n4433,n4434,n4436);
and (n4434,n4432,n4435);
and (n4435,n4197,n2830);
and (n4436,n4205,n4207);
nand (n4437,n4356,n4362);
or (n4438,n4439,n4441,n4458);
and (n4439,n4440,n3845);
xor (n4440,n4123,n4342);
and (n4441,n3845,n4442);
or (n4442,n4443,n4446,n4457);
and (n4443,n4444,n4445);
xor (n4444,n4091,n4345);
xor (n4445,n3960,n3962);
and (n4446,n4445,n4447);
or (n4447,n4448,n4451,n4456);
and (n4448,n4449,n4450);
xor (n4449,n4112,n4348);
xor (n4450,n3963,n3965);
and (n4451,n4450,n4452);
or (n4452,n4453,n4454,n4455);
and (n4453,n24,n1992);
and (n4454,n1992,n3713);
and (n4455,n24,n3713);
and (n4456,n4449,n4452);
and (n4457,n4444,n4447);
and (n4458,n4440,n4442);
and (n4459,n4445,n4460);
or (n4460,n4461,n4464,n4481);
and (n4461,n4462,n4450);
xor (n4462,n4463,n4442);
xor (n4463,n4440,n3845);
and (n4464,n4450,n4465);
or (n4465,n4466,n4469,n4480);
and (n4466,n4467,n1992);
xor (n4467,n4468,n4447);
xor (n4468,n4444,n4445);
and (n4469,n1992,n4470);
or (n4470,n4471,n4474,n4479);
and (n4471,n4472,n3717);
xor (n4472,n4473,n4452);
xor (n4473,n4449,n4450);
and (n4474,n3717,n4475);
or (n4475,n4476,n4477,n4478);
and (n4476,n22,n3723);
and (n4477,n3723,n3778);
and (n4478,n22,n3778);
and (n4479,n4472,n4475);
and (n4480,n4467,n4470);
and (n4481,n4462,n4465);
and (n4482,n4336,n4460);
and (n4483,n4484,n4486);
xor (n4484,n4485,n4460);
xor (n4485,n4336,n4445);
and (n4486,n4487,n4489);
xor (n4487,n4488,n4465);
xor (n4488,n4462,n4450);
and (n4489,n4490,n4492);
xor (n4490,n4491,n4470);
xor (n4491,n4467,n1992);
and (n4492,n4493,n4495);
xor (n4493,n4494,n4475);
xor (n4494,n4472,n3717);
and (n4495,n20,n3823);
xor (n4496,n3843,n4497);
and (n4497,n4484,n4498);
and (n4498,n4487,n4499);
and (n4499,n4490,n4500);
and (n4500,n4493,n4501);
and (n4501,n20,n3824);
wire s0n4502,s1n4502,notn4502;
or (n4502,s0n4502,s1n4502);
not(notn4502,n28);
and (s0n4502,notn4502,n4503);
and (s1n4502,n28,n4506);
wire s0n4503,s1n4503,notn4503;
or (n4503,s0n4503,s1n4503);
not(notn4503,n28);
and (s0n4503,notn4503,n4504);
and (s1n4503,n28,n4505);
xor (n4504,n4487,n4489);
xor (n4505,n4487,n4499);
wire s0n4506,s1n4506,notn4506;
or (n4506,s0n4506,s1n4506);
not(notn4506,n28);
and (s0n4506,notn4506,n4507);
and (s1n4506,n28,n4624);
xor (n4507,n4508,n4614);
xor (n4508,n4509,n4577);
nand (n4509,n4510,n4576);
or (n4510,n4511,n4536);
not (n4511,n4512);
xor (n4512,n4513,n4523);
xor (n4513,n4514,n4517);
or (n4514,n4515,n4516);
and (n4515,n3975,n3980);
and (n4516,n3976,n3978);
xor (n4517,n4518,n3980);
xor (n4518,n4519,n4521);
wire s0n4519,s1n4519,notn4519;
or (n4519,s0n4519,s1n4519);
not(notn4519,n28);
and (s0n4519,notn4519,1'b0);
and (s1n4519,n28,n4520);
wire s0n4521,s1n4521,notn4521;
or (n4521,s0n4521,s1n4521);
not(notn4521,n28);
and (s0n4521,notn4521,1'b0);
and (s1n4521,n28,n4522);
nand (n4523,n4524,n4528,n4529);
nand (n4524,n4372,n4525);
and (n4525,n4396,n4526);
and (n4526,n4527,n4359);
or (n4527,n4007,n3974);
nand (n4528,n4525,n4399,n4403);
nor (n4529,n4530,n4531);
and (n4530,n4364,n4526);
nand (n4531,n4532,n4535);
or (n4532,n4533,n4534);
not (n4533,n4527);
not (n4534,n4361);
nand (n4535,n4007,n3974);
nand (n4536,n4537,n4575);
or (n4537,n4538,n4557);
not (n4538,n4539);
xnor (n4539,n4540,n4545);
or (n4540,n4541,n4543);
and (n4541,n4542,n4007);
not (n4542,n4513);
and (n4543,n4517,n4544);
not (n4544,n4514);
nand (n4545,n4546,n4556);
or (n4546,n4544,n4547);
nand (n4547,n4548,n4555);
or (n4548,n3980,n4549);
not (n4549,n4550);
or (n4550,n4551,n4552);
and (n4551,n4518,n3980);
and (n4552,n4553,n4554);
not (n4553,n4519);
not (n4554,n4521);
or (n4555,n4550,n3981);
nand (n4556,n4547,n4544);
nand (n4557,n4558,n4572,n4574);
nand (n4558,n4559,n4560,n4311);
nand (n4559,n4140,n4258);
nand (n4560,n4561,n4570);
or (n4561,n4562,n4568);
nand (n4562,n3971,n4563);
nand (n4563,n4564,n4567);
or (n4564,n4565,n4566);
and (n4565,n3973,n4027);
and (n4566,n3974,n4006);
xor (n4567,n4542,n4007);
not (n4568,n4569);
nand (n4569,n4133,n4064);
nand (n4570,n4326,n4571);
nor (n4571,n4562,n4332);
nand (n4572,n4560,n4573);
nand (n4573,n4070,n4568);
or (n4574,n4564,n4567);
nand (n4575,n4538,n4557);
nand (n4576,n4536,n4511);
or (n4577,n4578,n4590,n4613);
and (n4578,n4536,n4579);
nand (n4579,n4580,n4589);
or (n4580,n4581,n4583);
not (n4581,n4582);
not (n4582,n3973);
nand (n4583,n4584,n4586,n4587);
nand (n4584,n4372,n4585);
and (n4585,n4396,n4359);
nand (n4586,n4585,n4399,n4403);
nor (n4587,n4588,n4361);
and (n4588,n4364,n4359);
nand (n4589,n4581,n4583);
and (n4590,n4579,n4591);
or (n4591,n4592,n4607,n4612);
and (n4592,n4354,n4593);
nand (n4593,n4594,n4606);
or (n4594,n4595,n4597);
not (n4595,n4596);
and (n4596,n4563,n4574);
nand (n4597,n4598,n4600,n4601);
nand (n4598,n4599,n4140,n4258);
not (n4599,n4573);
nand (n4600,n4599,n4310);
nor (n4601,n4602,n4603);
and (n4602,n4325,n4568);
nand (n4603,n4604,n3971);
or (n4604,n4605,n4063);
not (n4605,n4332);
nand (n4606,n4595,n4597);
and (n4607,n4354,n4608);
or (n4608,n4609,n4610,n4611);
and (n4609,n3845,n3966);
and (n4610,n3845,n4334);
and (n4611,n3966,n4334);
and (n4612,n4593,n4608);
and (n4613,n4536,n4591);
and (n4614,n4615,n4620);
xor (n4615,n4616,n4591);
nor (n4616,n4578,n4617);
and (n4617,n4618,n4619);
not (n4618,n4579);
not (n4619,n4536);
and (n4620,n4621,n4623);
xor (n4621,n4622,n4608);
xor (n4622,n4593,n4354);
and (n4623,n3843,n4483);
xor (n4624,n4508,n4625);
and (n4625,n4615,n4626);
and (n4626,n4621,n4627);
and (n4627,n3843,n4497);
wire s0n4628,s1n4628,notn4628;
or (n4628,s0n4628,s1n4628);
not(notn4628,n28);
and (s0n4628,notn4628,n4629);
and (s1n4628,n28,n4646);
xor (n4629,n4630,n4645);
xor (n4630,n4631,n4641);
nand (n4631,n4632,n4640);
or (n4632,n4633,n4536);
not (n4633,n4634);
nand (n4634,n4635,n4639);
or (n4635,n4636,n4547);
or (n4636,n4637,n4638);
and (n4637,n4513,n4523);
and (n4638,n4514,n4517);
nand (n4639,n4636,n4547);
nand (n4640,n4536,n4633);
or (n4641,n4642,n4643,n4644);
and (n4642,n4536,n4512);
and (n4643,n4512,n4577);
and (n4644,n4536,n4577);
and (n4645,n4508,n4614);
xor (n4646,n4630,n4647);
and (n4647,n4508,n4625);
and (n4648,n4649,n4651);
not (n4649,n4650);
nor (n4650,n907,n902,n903,n905);
or (n4651,n901,n902,n904,n905);
and (n4652,n4653,n917);
wire s0n4653,s1n4653,notn4653;
or (n4653,s0n4653,s1n4653);
not(notn4653,n918);
and (s0n4653,notn4653,1'b0);
and (s1n4653,n918,n15);
and (n4654,n15,n4655);
not (n4655,n953);
and (n4656,n4657,n6755);
wire s0n4657,s1n4657,notn4657;
or (n4657,s0n4657,s1n4657);
not(notn4657,n6750);
and (s0n4657,notn4657,n4658);
and (s1n4657,n6750,1'b0);
wire s0n4658,s1n4658,notn4658;
or (n4658,s0n4658,s1n4658);
not(notn4658,n6724);
and (s0n4658,notn4658,n4659);
and (s1n4658,n6724,1'b1);
wire s0n4659,s1n4659,notn4659;
or (n4659,s0n4659,s1n4659);
not(notn4659,n6717);
and (s0n4659,notn4659,1'b0);
and (s1n4659,n6717,n4660);
xor (n4660,n4661,n6700);
xor (n4661,n4662,n6656);
xor (n4662,n4663,n6591);
xor (n4663,n4664,n6152);
xor (n4664,n4665,n6120);
xnor (n4665,n4666,n5409);
or (n4666,n4667,n4822,n5408);
not (n4667,n4668);
or (n4668,n4669,n4779);
not (n4669,n4670);
nand (n4670,n4671,n4736);
nor (n4671,n4672,n4719);
nand (n4672,n4673,n4706,n4710,n4714);
nand (n4673,n4674,n4703);
not (n4674,n4675);
nand (n4675,n4676,n1056);
not (n4676,n4677);
nand (n4677,n4678,n4698);
nand (n4678,n4679,n4693);
not (n4679,n4680);
nand (n4680,n4681,n4687);
nand (n4681,n4682,n906);
nand (n4682,n4683,n4684,n4686);
nand (n4683,n32,n1069,n824);
not (n4684,n4685);
nor (n4685,n33,n677,n750,n824);
nand (n4686,n751,n33);
nor (n4687,n4688,n4692);
nor (n4688,n4689,n960);
nand (n4689,n4690,n4691);
or (n4690,n677,n33);
not (n4691,n954);
not (n4692,n967);
and (n4693,n4694,n4695,n955);
nand (n4694,n4682,n910);
not (n4695,n4696);
and (n4696,n4697,n900);
not (n4697,n4689);
nand (n4698,n4699,n4681,n4700,n4701);
nand (n4699,n909,n4682);
and (n4700,n4695,n961);
nor (n4701,n4702,n4692);
and (n4702,n4697,n906);
wire s0n4703,s1n4703,notn4703;
or (n4703,s0n4703,s1n4703);
not(notn4703,n4704);
and (s0n4703,notn4703,n2028);
and (s1n4703,n4704,n2092);
not (n4704,n4705);
nand (n4705,n751,n33,n677);
nand (n4706,n4707,n4709);
not (n4707,n4708);
nand (n4708,n4676,n1041);
wire s0n4709,s1n4709,notn4709;
or (n4709,s0n4709,s1n4709);
not(notn4709,n4704);
and (s0n4709,notn4709,n2016);
and (s1n4709,n4704,n2080);
nand (n4710,n4711,n4713);
not (n4711,n4712);
nand (n4712,n4676,n990);
wire s0n4713,s1n4713,notn4713;
or (n4713,s0n4713,s1n4713);
not(notn4713,n4704);
and (s0n4713,notn4713,n2045);
and (s1n4713,n4704,n2099);
nand (n4714,n4715,n4718);
and (n4715,n4716,n970);
and (n4716,n4678,n4717);
not (n4717,n4698);
wire s0n4718,s1n4718,notn4718;
or (n4718,s0n4718,s1n4718);
not(notn4718,n4704);
and (s0n4718,notn4718,n2033);
and (s1n4718,n4704,n2068);
nand (n4719,n4720,n4723,n4726,n4733);
nand (n4720,n4721,n4722);
and (n4721,n4716,n1041);
wire s0n4722,s1n4722,notn4722;
or (n4722,s0n4722,s1n4722);
not(notn4722,n4704);
and (s0n4722,notn4722,n2010);
and (s1n4722,n4704,n2074);
nand (n4723,n4724,n4725);
and (n4724,n4716,n990);
wire s0n4725,s1n4725,notn4725;
or (n4725,s0n4725,s1n4725);
not(notn4725,n4704);
and (s0n4725,notn4725,n2040);
and (s1n4725,n4704,n2066);
nand (n4726,n4727,n4732);
not (n4727,n4728);
nand (n4728,n4729,n970);
not (n4729,n4730);
nand (n4730,n4679,n4693,n4731);
nand (n4731,n4699,n4701,n961);
wire s0n4732,s1n4732,notn4732;
or (n4732,s0n4732,s1n4732);
not(notn4732,n4704);
and (s0n4732,notn4732,n2038);
and (s1n4732,n4704,n2060);
nand (n4733,n4734,n4735);
and (n4734,n4716,n1056);
wire s0n4735,s1n4735,notn4735;
or (n4735,s0n4735,s1n4735);
not(notn4735,n4704);
and (s0n4735,notn4735,n2023);
and (s1n4735,n4704,n2087);
nor (n4736,n4737,n4748);
nand (n4737,n4738,n4741,n4744);
nand (n4738,n4739,n4740);
and (n4739,n4729,n990);
wire s0n4740,s1n4740,notn4740;
or (n4740,s0n4740,s1n4740);
not(notn4740,n4704);
and (s0n4740,notn4740,n2036);
and (s1n4740,n4704,n2064);
nand (n4741,n4742,n4743);
and (n4742,n4729,n1056);
wire s0n4743,s1n4743,notn4743;
or (n4743,s0n4743,s1n4743);
not(notn4743,n4704);
and (s0n4743,notn4743,n2026);
and (s1n4743,n4704,n2090);
nand (n4744,n4745,n4747);
not (n4745,n4746);
nand (n4746,n4729,n1041);
wire s0n4747,s1n4747,notn4747;
or (n4747,s0n4747,s1n4747);
not(notn4747,n4704);
and (s0n4747,notn4747,n2014);
and (s1n4747,n4704,n2078);
nand (n4748,n4749,n4753);
or (n4749,n4750,n4752);
not (n4750,n4751);
wire s0n4751,s1n4751,notn4751;
or (n4751,s0n4751,s1n4751);
not(notn4751,n4704);
and (s0n4751,notn4751,n2050);
and (s1n4751,n4704,n2097);
nand (n4752,n4676,n970);
nor (n4753,n4754,n4769);
nand (n4754,n4755,n4764);
or (n4755,n4756,n4762);
not (n4756,n4757);
and (n4757,n4758,n1041);
nand (n4758,n984,n4759,n4761);
not (n4759,n4760);
and (n4760,n4697,n4650);
nand (n4761,n4682,n900);
not (n4762,n4763);
wire s0n4763,s1n4763,notn4763;
or (n4763,s0n4763,s1n4763);
not(notn4763,n4704);
and (s0n4763,notn4763,n2018);
and (s1n4763,n4704,n2082);
or (n4764,n4765,n4767);
not (n4765,n4766);
and (n4766,n4758,n970);
not (n4767,n4768);
wire s0n4768,s1n4768,notn4768;
or (n4768,s0n4768,s1n4768);
not(notn4768,n4704);
and (s0n4768,notn4768,n2052);
and (s1n4768,n4704,n2102);
nand (n4769,n4770,n4774);
or (n4770,n4771,n4772);
nand (n4771,n4758,n1056);
not (n4772,n4773);
wire s0n4773,s1n4773,notn4773;
or (n4773,s0n4773,s1n4773);
not(notn4773,n4704);
and (s0n4773,notn4773,n2030);
and (s1n4773,n4704,n2094);
or (n4774,n4775,n4777);
not (n4775,n4776);
and (n4776,n4758,n990);
not (n4777,n4778);
wire s0n4778,s1n4778,notn4778;
or (n4778,s0n4778,s1n4778);
not(notn4778,n4704);
and (s0n4778,notn4778,n2047);
and (s1n4778,n4704,n2104);
not (n4779,n4780);
nand (n4780,n4781,n4804,n4813);
nor (n4781,n4782,n4799);
nand (n4782,n4783,n4785,n4786);
nand (n4783,n4784,n4768);
not (n4784,n4752);
nand (n4785,n4745,n4709);
nor (n4786,n4787,n4792);
nand (n4787,n4788,n4790);
or (n4788,n4771,n4789);
not (n4789,n4722);
or (n4790,n4775,n4791);
not (n4791,n4718);
nand (n4792,n4793,n4796);
or (n4793,n4756,n4794);
not (n4794,n4795);
wire s0n4795,s1n4795,notn4795;
or (n4795,s0n4795,s1n4795);
not(notn4795,n4704);
and (s0n4795,notn4795,n2012);
and (s1n4795,n4704,n2076);
or (n4796,n4765,n4797);
not (n4797,n4798);
wire s0n4798,s1n4798,notn4798;
or (n4798,s0n4798,s1n4798);
not(notn4798,n4704);
and (s0n4798,notn4798,n2042);
and (s1n4798,n4704,n2062);
nand (n4799,n4800,n4803);
or (n4800,n4801,n4802);
not (n4801,n4713);
not (n4802,n4739);
nand (n4803,n4742,n4703);
nor (n4804,n4805,n4808);
nand (n4805,n4806,n4807);
or (n4806,n4777,n4712);
nand (n4807,n4674,n4773);
nand (n4808,n4809,n4812);
or (n4809,n4810,n4811);
not (n4810,n4743);
not (n4811,n4734);
nand (n4812,n4715,n4732);
nor (n4813,n4814,n4819);
nand (n4814,n4815,n4818);
or (n4815,n4816,n4817);
not (n4816,n4740);
not (n4817,n4724);
nand (n4818,n4721,n4747);
nand (n4819,n4820,n4821);
or (n4820,n4750,n4728);
nand (n4821,n4707,n4763);
and (n4822,n4670,n4823);
or (n4823,n4824,n4908,n5407);
and (n4824,n4825,n4879);
nand (n4825,n4826,n4852,n4865);
nor (n4826,n4827,n4846);
nand (n4827,n4828,n4830,n4832);
nand (n4828,n4784,n4829);
wire s0n4829,s1n4829,notn4829;
or (n4829,s0n4829,s1n4829);
not(notn4829,n4704);
and (s0n4829,notn4829,n2152);
and (s1n4829,n4704,n2218);
nand (n4830,n4742,n4831);
wire s0n4831,s1n4831,notn4831;
or (n4831,s0n4831,s1n4831);
not(notn4831,n4704);
and (s0n4831,notn4831,n2132);
and (s1n4831,n4704,n2179);
nor (n4832,n4833,n4840);
nand (n4833,n4834,n4837);
or (n4834,n4835,n4775);
not (n4835,n4836);
wire s0n4836,s1n4836,notn4836;
or (n4836,s0n4836,s1n4836);
not(notn4836,n4704);
and (s0n4836,notn4836,n2159);
and (s1n4836,n4704,n2207);
nand (n4837,n4838,n4839);
not (n4838,n4771);
wire s0n4839,s1n4839,notn4839;
or (n4839,s0n4839,s1n4839);
not(notn4839,n4704);
and (s0n4839,notn4839,n2136);
and (s1n4839,n4704,n2169);
nand (n4840,n4841,n4844);
or (n4841,n4842,n4765);
not (n4842,n4843);
wire s0n4843,s1n4843,notn4843;
or (n4843,s0n4843,s1n4843);
not(notn4843,n4704);
and (s0n4843,notn4843,n2157);
and (s1n4843,n4704,n2221);
nand (n4844,n4757,n4845);
wire s0n4845,s1n4845,notn4845;
or (n4845,s0n4845,s1n4845);
not(notn4845,n4704);
and (s0n4845,notn4845,n2124);
and (s1n4845,n4704,n2186);
nand (n4846,n4847,n4850);
or (n4847,n4848,n4802);
not (n4848,n4849);
wire s0n4849,s1n4849,notn4849;
or (n4849,s0n4849,s1n4849);
not(notn4849,n4704);
and (s0n4849,notn4849,n2149);
and (s1n4849,n4704,n2200);
nand (n4850,n4745,n4851);
wire s0n4851,s1n4851,notn4851;
or (n4851,s0n4851,s1n4851);
not(notn4851,n4704);
and (s0n4851,notn4851,n2120);
and (s1n4851,n4704,n2195);
nor (n4852,n4853,n4859);
nand (n4853,n4854,n4857);
or (n4854,n4855,n4712);
not (n4855,n4856);
wire s0n4856,s1n4856,notn4856;
or (n4856,s0n4856,s1n4856);
not(notn4856,n4704);
and (s0n4856,notn4856,n2154);
and (s1n4856,n4704,n2204);
nand (n4857,n4707,n4858);
wire s0n4858,s1n4858,notn4858;
or (n4858,s0n4858,s1n4858);
not(notn4858,n4704);
and (s0n4858,notn4858,n2122);
and (s1n4858,n4704,n2184);
nand (n4859,n4860,n4863);
or (n4860,n4861,n4675);
not (n4861,n4862);
wire s0n4862,s1n4862,notn4862;
or (n4862,s0n4862,s1n4862);
not(notn4862,n4704);
and (s0n4862,notn4862,n2134);
and (s1n4862,n4704,n2167);
nand (n4863,n4721,n4864);
wire s0n4864,s1n4864,notn4864;
or (n4864,s0n4864,s1n4864);
not(notn4864,n4704);
and (s0n4864,notn4864,n2116);
and (s1n4864,n4704,n2176);
nor (n4865,n4866,n4873);
nand (n4866,n4867,n4871);
or (n4867,n4868,n4870);
not (n4868,n4869);
wire s0n4869,s1n4869,notn4869;
or (n4869,s0n4869,s1n4869);
not(notn4869,n4704);
and (s0n4869,notn4869,n2139);
and (s1n4869,n4704,n2210);
not (n4870,n4715);
nand (n4871,n4724,n4872);
wire s0n4872,s1n4872,notn4872;
or (n4872,s0n4872,s1n4872);
not(notn4872,n4704);
and (s0n4872,notn4872,n2147);
and (s1n4872,n4704,n2201);
nand (n4873,n4874,n4877);
or (n4874,n4875,n4728);
not (n4875,n4876);
wire s0n4876,s1n4876,notn4876;
or (n4876,s0n4876,s1n4876);
not(notn4876,n4704);
and (s0n4876,notn4876,n2145);
and (s1n4876,n4704,n2215);
nand (n4877,n4734,n4878);
wire s0n4878,s1n4878,notn4878;
or (n4878,s0n4878,s1n4878);
not(notn4878,n4704);
and (s0n4878,notn4878,n2129);
and (s1n4878,n4704,n2174);
nand (n4879,n4880,n4891);
nor (n4880,n4881,n4886);
nand (n4881,n4882,n4883,n4884,n4885);
nand (n4882,n4674,n4839);
nand (n4883,n4707,n4845);
nand (n4884,n4711,n4836);
nand (n4885,n4715,n4876);
nand (n4886,n4887,n4888,n4889,n4890);
nand (n4887,n4721,n4851);
nand (n4888,n4727,n4829);
nand (n4889,n4734,n4831);
nand (n4890,n4724,n4849);
nor (n4891,n4892,n4905);
nand (n4892,n4893,n4894,n4895);
nand (n4893,n4784,n4843);
nand (n4894,n4742,n4862);
nor (n4895,n4896,n4899);
nand (n4896,n4897,n4898);
or (n4897,n4868,n4775);
nand (n4898,n4838,n4864);
nand (n4899,n4900,n4903);
or (n4900,n4901,n4756);
not (n4901,n4902);
wire s0n4902,s1n4902,notn4902;
or (n4902,s0n4902,s1n4902);
not(notn4902,n4704);
and (s0n4902,notn4902,n2118);
and (s1n4902,n4704,n2192);
nand (n4903,n4904,n4766);
wire s0n4904,s1n4904,notn4904;
or (n4904,s0n4904,s1n4904);
not(notn4904,n4704);
and (s0n4904,notn4904,n2143);
and (s1n4904,n4704,n2224);
nand (n4905,n4906,n4907);
or (n4906,n4855,n4802);
nand (n4907,n4745,n4858);
and (n4908,n4825,n4909);
or (n4909,n4910,n4987,n5406);
and (n4910,n4911,n4956);
nand (n4911,n4912,n4931);
nor (n4912,n4913,n4922);
nand (n4913,n4914,n4916,n4918,n4920);
nand (n4914,n4711,n4915);
wire s0n4915,s1n4915,notn4915;
or (n4915,s0n4915,s1n4915);
not(notn4915,n4704);
and (s0n4915,notn4915,n2275);
and (s1n4915,n4704,n2330);
nand (n4916,n4674,n4917);
wire s0n4917,s1n4917,notn4917;
or (n4917,s0n4917,s1n4917);
not(notn4917,n4704);
and (s0n4917,notn4917,n2262);
and (s1n4917,n4704,n2308);
nand (n4918,n4715,n4919);
wire s0n4919,s1n4919,notn4919;
or (n4919,s0n4919,s1n4919);
not(notn4919,n4704);
and (s0n4919,notn4919,n2233);
and (s1n4919,n4704,n2286);
nand (n4920,n4707,n4921);
wire s0n4921,s1n4921,notn4921;
or (n4921,s0n4921,s1n4921);
not(notn4921,n4704);
and (s0n4921,notn4921,n2249);
and (s1n4921,n4704,n2323);
nand (n4922,n4923,n4925,n4927,n4929);
nand (n4923,n4721,n4924);
wire s0n4924,s1n4924,notn4924;
or (n4924,s0n4924,s1n4924);
not(notn4924,n4704);
and (s0n4924,notn4924,n2254);
and (s1n4924,n4704,n2304);
nand (n4925,n4727,n4926);
wire s0n4926,s1n4926,notn4926;
or (n4926,s0n4926,s1n4926);
not(notn4926,n4704);
and (s0n4926,notn4926,n2237);
and (s1n4926,n4704,n2289);
nand (n4927,n4724,n4928);
wire s0n4928,s1n4928,notn4928;
or (n4928,s0n4928,s1n4928);
not(notn4928,n4704);
and (s0n4928,notn4928,n2242);
and (s1n4928,n4704,n2296);
nand (n4929,n4734,n4930);
wire s0n4930,s1n4930,notn4930;
or (n4930,s0n4930,s1n4930);
not(notn4930,n4704);
and (s0n4930,notn4930,n2267);
and (s1n4930,n4704,n2302);
nor (n4931,n4932,n4950);
nand (n4932,n4933,n4935,n4937);
nand (n4933,n4784,n4934);
wire s0n4934,s1n4934,notn4934;
or (n4934,s0n4934,s1n4934);
not(notn4934,n4704);
and (s0n4934,notn4934,n2273);
and (s1n4934,n4704,n2312);
nand (n4935,n4742,n4936);
wire s0n4936,s1n4936,notn4936;
or (n4936,s0n4936,s1n4936);
not(notn4936,n4704);
and (s0n4936,notn4936,n2270);
and (s1n4936,n4704,n2306);
nor (n4937,n4938,n4944);
nand (n4938,n4939,n4942);
or (n4939,n4940,n4771);
not (n4940,n4941);
wire s0n4941,s1n4941,notn4941;
or (n4941,s0n4941,s1n4941);
not(notn4941,n4704);
and (s0n4941,notn4941,n2264);
and (s1n4941,n4704,n2310);
nand (n4942,n4776,n4943);
wire s0n4943,s1n4943,notn4943;
or (n4943,s0n4943,s1n4943);
not(notn4943,n4704);
and (s0n4943,notn4943,n2280);
and (s1n4943,n4704,n2327);
nand (n4944,n4945,n4948);
or (n4945,n4946,n4765);
not (n4946,n4947);
wire s0n4947,s1n4947,notn4947;
or (n4947,s0n4947,s1n4947);
not(notn4947,n4704);
and (s0n4947,notn4947,n2278);
and (s1n4947,n4704,n2332);
nand (n4948,n4757,n4949);
wire s0n4949,s1n4949,notn4949;
or (n4949,s0n4949,s1n4949);
not(notn4949,n4704);
and (s0n4949,notn4949,n2251);
and (s1n4949,n4704,n2325);
nand (n4950,n4951,n4954);
or (n4951,n4952,n4802);
not (n4952,n4953);
wire s0n4953,s1n4953,notn4953;
or (n4953,s0n4953,s1n4953);
not(notn4953,n4704);
and (s0n4953,notn4953,n2244);
and (s1n4953,n4704,n2292);
nand (n4954,n4745,n4955);
wire s0n4955,s1n4955,notn4955;
or (n4955,s0n4955,s1n4955);
not(notn4955,n4704);
and (s0n4955,notn4955,n2258);
and (s1n4955,n4704,n2321);
nand (n4956,n4957,n4968);
nor (n4957,n4958,n4963);
nand (n4958,n4959,n4960,n4961,n4962);
nand (n4959,n4721,n4955);
nand (n4960,n4707,n4949);
nand (n4961,n4711,n4943);
nand (n4962,n4674,n4941);
nand (n4963,n4964,n4965,n4966,n4967);
nand (n4964,n4727,n4934);
nand (n4965,n4715,n4926);
nand (n4966,n4724,n4953);
nand (n4967,n4734,n4936);
nor (n4968,n4969,n4983);
nand (n4969,n4970,n4971,n4972);
nand (n4970,n4784,n4947);
nand (n4971,n4742,n4917);
nor (n4972,n4973,n4977);
nand (n4973,n4974,n4976);
or (n4974,n4975,n4775);
not (n4975,n4919);
nand (n4976,n4838,n4924);
nand (n4977,n4978,n4981);
or (n4978,n4979,n4756);
not (n4979,n4980);
wire s0n4980,s1n4980,notn4980;
or (n4980,s0n4980,s1n4980);
not(notn4980,n4704);
and (s0n4980,notn4980,n2256);
and (s1n4980,n4704,n2319);
nand (n4981,n4766,n4982);
wire s0n4982,s1n4982,notn4982;
or (n4982,s0n4982,s1n4982);
not(notn4982,n4704);
and (s0n4982,notn4982,n2240);
and (s1n4982,n4704,n2294);
nand (n4983,n4984,n4986);
or (n4984,n4985,n4746);
not (n4985,n4921);
nand (n4986,n4739,n4915);
and (n4987,n4911,n4988);
or (n4988,n4989,n5064,n5405);
and (n4989,n4990,n5034);
nand (n4990,n4991,n5010);
nor (n4991,n4992,n5001);
nand (n4992,n4993,n4995,n4997,n4999);
nand (n4993,n4721,n4994);
wire s0n4994,s1n4994,notn4994;
or (n4994,s0n4994,s1n4994);
not(notn4994,n4704);
and (s0n4994,notn4994,n2371);
and (s1n4994,n4704,n2431);
nand (n4995,n4711,n4996);
wire s0n4996,s1n4996,notn4996;
or (n4996,s0n4996,s1n4996);
not(notn4996,n4704);
and (s0n4996,notn4996,n2383);
and (s1n4996,n4704,n2443);
nand (n4997,n4674,n4998);
wire s0n4998,s1n4998,notn4998;
or (n4998,s0n4998,s1n4998);
not(notn4998,n4704);
and (s0n4998,notn4998,n2343);
and (s1n4998,n4704,n2416);
nand (n4999,n4707,n5000);
wire s0n5000,s1n5000,notn5000;
or (n5000,s0n5000,s1n5000);
not(notn5000,n4704);
and (s0n5000,notn5000,n2360);
and (s1n5000,n4704,n2423);
nand (n5001,n5002,n5004,n5006,n5008);
nand (n5002,n4727,n5003);
wire s0n5003,s1n5003,notn5003;
or (n5003,s0n5003,s1n5003);
not(notn5003,n4704);
and (s0n5003,notn5003,n2394);
and (s1n5003,n4704,n2454);
nand (n5004,n4715,n5005);
wire s0n5005,s1n5005,notn5005;
or (n5005,s0n5005,s1n5005);
not(notn5005,n4704);
and (s0n5005,notn5005,n2391);
and (s1n5005,n4704,n2451);
nand (n5006,n4724,n5007);
wire s0n5007,s1n5007,notn5007;
or (n5007,s0n5007,s1n5007);
not(notn5007,n4704);
and (s0n5007,notn5007,n2376);
and (s1n5007,n4704,n2436);
nand (n5008,n4734,n5009);
wire s0n5009,s1n5009,notn5009;
or (n5009,s0n5009,s1n5009);
not(notn5009,n4704);
and (s0n5009,notn5009,n2355);
and (s1n5009,n4704,n2412);
nor (n5010,n5011,n5018);
nand (n5011,n5012,n5014,n5016);
nand (n5012,n4745,n5013);
wire s0n5013,s1n5013,notn5013;
or (n5013,s0n5013,s1n5013);
not(notn5013,n4704);
and (s0n5013,notn5013,n2362);
and (s1n5013,n4704,n2421);
nand (n5014,n4739,n5015);
wire s0n5015,s1n5015,notn5015;
or (n5015,s0n5015,s1n5015);
not(notn5015,n4704);
and (s0n5015,notn5015,n2380);
and (s1n5015,n4704,n2440);
nand (n5016,n4742,n5017);
wire s0n5017,s1n5017,notn5017;
or (n5017,s0n5017,s1n5017);
not(notn5017,n4704);
and (s0n5017,notn5017,n2345);
and (s1n5017,n4704,n2414);
nand (n5018,n5019,n5022);
or (n5019,n5020,n4752);
not (n5020,n5021);
wire s0n5021,s1n5021,notn5021;
or (n5021,s0n5021,s1n5021);
not(notn5021,n4704);
and (s0n5021,notn5021,n2397);
and (s1n5021,n4704,n2457);
nor (n5022,n5023,n5029);
nand (n5023,n5024,n5027);
or (n5024,n5025,n4775);
not (n5025,n5026);
wire s0n5026,s1n5026,notn5026;
or (n5026,s0n5026,s1n5026);
not(notn5026,n4704);
and (s0n5026,notn5026,n2386);
and (s1n5026,n4704,n2446);
nand (n5027,n4838,n5028);
wire s0n5028,s1n5028,notn5028;
or (n5028,s0n5028,s1n5028);
not(notn5028,n4704);
and (s0n5028,notn5028,n2352);
and (s1n5028,n4704,n2410);
nand (n5029,n5030,n5032);
nand (n5030,n4757,n5031);
wire s0n5031,s1n5031,notn5031;
or (n5031,s0n5031,s1n5031);
not(notn5031,n4704);
and (s0n5031,notn5031,n2368);
and (s1n5031,n4704,n2429);
nand (n5032,n4766,n5033);
wire s0n5033,s1n5033,notn5033;
or (n5033,s0n5033,s1n5033);
not(notn5033,n4704);
and (s0n5033,notn5033,n2400);
and (s1n5033,n4704,n2460);
nand (n5034,n5035,n5048);
nor (n5035,n5036,n5041);
nand (n5036,n5037,n5038,n5039,n5040);
nand (n5037,n4711,n5015);
nand (n5038,n4674,n5017);
nand (n5039,n4721,n5028);
nand (n5040,n4707,n5013);
nand (n5041,n5042,n5043,n5044,n5046);
nand (n5042,n4715,n5026);
nand (n5043,n4727,n5005);
nand (n5044,n4734,n5045);
wire s0n5045,s1n5045,notn5045;
or (n5045,s0n5045,s1n5045);
not(notn5045,n4704);
and (s0n5045,notn5045,n2350);
and (s1n5045,n4704,n2408);
nand (n5046,n4724,n5047);
wire s0n5047,s1n5047,notn5047;
or (n5047,s0n5047,s1n5047);
not(notn5047,n4704);
and (s0n5047,notn5047,n2377);
and (s1n5047,n4704,n2437);
nor (n5048,n5049,n5060);
nand (n5049,n5050,n5051,n5052);
nand (n5050,n4784,n5003);
nand (n5051,n4742,n5009);
nor (n5052,n5053,n5057);
nand (n5053,n5054,n5056);
or (n5054,n5055,n4775);
not (n5055,n4996);
nand (n5056,n4838,n4998);
nand (n5057,n5058,n5059);
or (n5058,n5020,n4765);
nand (n5059,n4757,n5000);
nand (n5060,n5061,n5063);
or (n5061,n5062,n4802);
not (n5062,n5007);
nand (n5063,n4745,n4994);
and (n5064,n5034,n5065);
or (n5065,n5066,n5149,n5404);
and (n5066,n5067,n5112);
nand (n5067,n5068,n5087);
nor (n5068,n5069,n5078);
nand (n5069,n5070,n5072,n5074,n5076);
nand (n5070,n4715,n5071);
wire s0n5071,s1n5071,notn5071;
or (n5071,s0n5071,s1n5071);
not(notn5071,n4704);
and (s0n5071,notn5071,n2519);
and (s1n5071,n4704,n2576);
nand (n5072,n4711,n5073);
wire s0n5073,s1n5073,notn5073;
or (n5073,s0n5073,s1n5073);
not(notn5073,n4704);
and (s0n5073,notn5073,n2511);
and (s1n5073,n4704,n2568);
nand (n5074,n4674,n5075);
wire s0n5075,s1n5075,notn5075;
or (n5075,s0n5075,s1n5075);
not(notn5075,n4704);
and (s0n5075,notn5075,n2473);
and (s1n5075,n4704,n2537);
nand (n5076,n4707,n5077);
wire s0n5077,s1n5077,notn5077;
or (n5077,s0n5077,s1n5077);
not(notn5077,n4704);
and (s0n5077,notn5077,n2490);
and (s1n5077,n4704,n2550);
nand (n5078,n5079,n5081,n5083,n5085);
nand (n5079,n4721,n5080);
wire s0n5080,s1n5080,notn5080;
or (n5080,s0n5080,s1n5080);
not(notn5080,n4704);
and (s0n5080,notn5080,n2499);
and (s1n5080,n4704,n2556);
nand (n5081,n4724,n5082);
wire s0n5082,s1n5082,notn5082;
or (n5082,s0n5082,s1n5082);
not(notn5082,n4704);
and (s0n5082,notn5082,n2504);
and (s1n5082,n4704,n2561);
nand (n5083,n4727,n5084);
wire s0n5084,s1n5084,notn5084;
or (n5084,s0n5084,s1n5084);
not(notn5084,n4704);
and (s0n5084,notn5084,n2522);
and (s1n5084,n4704,n2579);
nand (n5085,n4734,n5086);
wire s0n5086,s1n5086,notn5086;
or (n5086,s0n5086,s1n5086);
not(notn5086,n4704);
and (s0n5086,notn5086,n2483);
and (s1n5086,n4704,n2544);
nor (n5087,n5088,n5106);
nand (n5088,n5089,n5091,n5093);
nand (n5089,n5090,n4742);
wire s0n5090,s1n5090,notn5090;
or (n5090,s0n5090,s1n5090);
not(notn5090,n4704);
and (s0n5090,notn5090,n2471);
and (s1n5090,n4704,n2535);
nand (n5091,n4784,n5092);
wire s0n5092,s1n5092,notn5092;
or (n5092,s0n5092,s1n5092);
not(notn5092,n4704);
and (s0n5092,notn5092,n2525);
and (s1n5092,n4704,n2582);
nor (n5093,n5094,n5100);
nand (n5094,n5095,n5098);
or (n5095,n5096,n4775);
not (n5096,n5097);
wire s0n5097,s1n5097,notn5097;
or (n5097,s0n5097,s1n5097);
not(notn5097,n4704);
and (s0n5097,notn5097,n2514);
and (s1n5097,n4704,n2571);
nand (n5098,n4838,n5099);
wire s0n5099,s1n5099,notn5099;
or (n5099,s0n5099,s1n5099);
not(notn5099,n4704);
and (s0n5099,notn5099,n2480);
and (s1n5099,n4704,n2542);
nand (n5100,n5101,n5104);
or (n5101,n5102,n4756);
not (n5102,n5103);
wire s0n5103,s1n5103,notn5103;
or (n5103,s0n5103,s1n5103);
not(notn5103,n4704);
and (s0n5103,notn5103,n2496);
and (s1n5103,n4704,n2554);
nand (n5104,n4766,n5105);
wire s0n5105,s1n5105,notn5105;
or (n5105,s0n5105,s1n5105);
not(notn5105,n4704);
and (s0n5105,notn5105,n2528);
and (s1n5105,n4704,n2585);
nand (n5106,n5107,n5110);
or (n5107,n5108,n4802);
not (n5108,n5109);
wire s0n5109,s1n5109,notn5109;
or (n5109,s0n5109,s1n5109);
not(notn5109,n4704);
and (s0n5109,notn5109,n2508);
and (s1n5109,n4704,n2565);
nand (n5110,n4745,n5111);
wire s0n5111,s1n5111,notn5111;
or (n5111,s0n5111,s1n5111);
not(notn5111,n4704);
and (s0n5111,notn5111,n2488);
and (s1n5111,n4704,n2548);
nand (n5112,n5113,n5130,n5139);
nor (n5113,n5114,n5118);
nand (n5114,n5115,n5116,n5117);
nand (n5115,n4742,n5086);
nand (n5116,n4745,n5080);
nand (n5117,n4739,n5082);
nand (n5118,n5119,n5121);
or (n5119,n5120,n4752);
not (n5120,n5084);
nor (n5121,n5122,n5126);
nand (n5122,n5123,n5125);
or (n5123,n5124,n4775);
not (n5124,n5073);
nand (n5125,n4838,n5075);
nand (n5126,n5127,n5129);
or (n5127,n5128,n4765);
not (n5128,n5092);
nand (n5129,n4757,n5077);
nor (n5130,n5131,n5136);
nand (n5131,n5132,n5135);
or (n5132,n5133,n5134);
not (n5133,n5099);
not (n5134,n4721);
nand (n5135,n4674,n5090);
nand (n5136,n5137,n5138);
or (n5137,n5108,n4712);
nand (n5138,n4707,n5111);
nor (n5139,n5140,n5144);
nand (n5140,n5141,n5142);
or (n5141,n5096,n4870);
nand (n5142,n4724,n5143);
wire s0n5143,s1n5143,notn5143;
or (n5143,s0n5143,s1n5143);
not(notn5143,n4704);
and (s0n5143,notn5143,n2505);
and (s1n5143,n4704,n2562);
nand (n5144,n5145,n5147);
or (n5145,n5146,n4728);
not (n5146,n5071);
nand (n5147,n4734,n5148);
wire s0n5148,s1n5148,notn5148;
or (n5148,s0n5148,s1n5148);
not(notn5148,n4704);
and (s0n5148,notn5148,n2478);
and (s1n5148,n4704,n2540);
and (n5149,n5112,n5150);
or (n5150,n5151,n5227,n5403);
and (n5151,n5152,n5197);
nand (n5152,n5153,n5172);
nor (n5153,n5154,n5163);
nand (n5154,n5155,n5157,n5159,n5161);
nand (n5155,n4674,n5156);
wire s0n5156,s1n5156,notn5156;
or (n5156,s0n5156,s1n5156);
not(notn5156,n4704);
and (s0n5156,notn5156,n2604);
and (s1n5156,n4704,n2661);
nand (n5157,n4707,n5158);
wire s0n5158,s1n5158,notn5158;
or (n5158,s0n5158,s1n5158);
not(notn5158,n4704);
and (s0n5158,notn5158,n2616);
and (s1n5158,n4704,n2673);
nand (n5159,n4711,n5160);
wire s0n5160,s1n5160,notn5160;
or (n5160,s0n5160,s1n5160);
not(notn5160,n4704);
and (s0n5160,notn5160,n2628);
and (s1n5160,n4704,n2685);
nand (n5161,n4715,n5162);
wire s0n5162,s1n5162,notn5162;
or (n5162,s0n5162,s1n5162);
not(notn5162,n4704);
and (s0n5162,notn5162,n2636);
and (s1n5162,n4704,n2693);
nand (n5163,n5164,n5166,n5168,n5170);
nand (n5164,n4721,n5165);
wire s0n5165,s1n5165,notn5165;
or (n5165,s0n5165,s1n5165);
not(notn5165,n4704);
and (s0n5165,notn5165,n2612);
and (s1n5165,n4704,n2669);
nand (n5166,n4734,n5167);
wire s0n5167,s1n5167,notn5167;
or (n5167,s0n5167,s1n5167);
not(notn5167,n4704);
and (s0n5167,notn5167,n2600);
and (s1n5167,n4704,n2657);
nand (n5168,n4724,n5169);
wire s0n5169,s1n5169,notn5169;
or (n5169,s0n5169,s1n5169);
not(notn5169,n4704);
and (s0n5169,notn5169,n2621);
and (s1n5169,n4704,n2678);
nand (n5170,n4727,n5171);
wire s0n5171,s1n5171,notn5171;
or (n5171,s0n5171,s1n5171);
not(notn5171,n4704);
and (s0n5171,notn5171,n2639);
and (s1n5171,n4704,n2696);
nor (n5172,n5173,n5180);
nand (n5173,n5174,n5176,n5178);
nand (n5174,n4745,n5175);
wire s0n5175,s1n5175,notn5175;
or (n5175,s0n5175,s1n5175);
not(notn5175,n4704);
and (s0n5175,notn5175,n2614);
and (s1n5175,n4704,n2671);
nand (n5176,n4739,n5177);
wire s0n5177,s1n5177,notn5177;
or (n5177,s0n5177,s1n5177);
not(notn5177,n4704);
and (s0n5177,notn5177,n2625);
and (s1n5177,n4704,n2682);
nand (n5178,n4742,n5179);
wire s0n5179,s1n5179,notn5179;
or (n5179,s0n5179,s1n5179);
not(notn5179,n4704);
and (s0n5179,notn5179,n2602);
and (s1n5179,n4704,n2659);
nand (n5180,n5181,n5184);
or (n5181,n5182,n4752);
not (n5182,n5183);
wire s0n5183,s1n5183,notn5183;
or (n5183,s0n5183,s1n5183);
not(notn5183,n4704);
and (s0n5183,notn5183,n2642);
and (s1n5183,n4704,n2699);
nor (n5184,n5185,n5191);
nand (n5185,n5186,n5189);
or (n5186,n5187,n4756);
not (n5187,n5188);
wire s0n5188,s1n5188,notn5188;
or (n5188,s0n5188,s1n5188);
not(notn5188,n4704);
and (s0n5188,notn5188,n2610);
and (s1n5188,n4704,n2666);
nand (n5189,n4766,n5190);
wire s0n5190,s1n5190,notn5190;
or (n5190,s0n5190,s1n5190);
not(notn5190,n4704);
and (s0n5190,notn5190,n2645);
and (s1n5190,n4704,n2702);
nand (n5191,n5192,n5195);
or (n5192,n5193,n4775);
not (n5193,n5194);
wire s0n5194,s1n5194,notn5194;
or (n5194,s0n5194,s1n5194);
not(notn5194,n4704);
and (s0n5194,notn5194,n2631);
and (s1n5194,n4704,n2688);
nand (n5195,n4838,n5196);
wire s0n5196,s1n5196,notn5196;
or (n5196,s0n5196,s1n5196);
not(notn5196,n4704);
and (s0n5196,notn5196,n2598);
and (s1n5196,n4704,n2655);
nand (n5197,n5198,n5211);
nor (n5198,n5199,n5204);
nand (n5199,n5200,n5201,n5202,n5203);
nand (n5200,n4721,n5196);
nand (n5201,n4707,n5175);
nand (n5202,n4674,n5179);
nand (n5203,n4711,n5177);
nand (n5204,n5205,n5207,n5208,n5209);
nand (n5205,n4724,n5206);
wire s0n5206,s1n5206,notn5206;
or (n5206,s0n5206,s1n5206);
not(notn5206,n4704);
and (s0n5206,notn5206,n2622);
and (s1n5206,n4704,n2679);
nand (n5207,n5194,n4715);
nand (n5208,n4727,n5162);
nand (n5209,n4734,n5210);
wire s0n5210,s1n5210,notn5210;
or (n5210,s0n5210,s1n5210);
not(notn5210,n4704);
and (s0n5210,notn5210,n2596);
and (s1n5210,n4704,n2653);
nor (n5211,n5212,n5223);
nand (n5212,n5213,n5214,n5215);
nand (n5213,n4742,n5167);
nand (n5214,n4784,n5171);
nor (n5215,n5216,n5219);
nand (n5216,n5217,n5218);
or (n5217,n5182,n4765);
nand (n5218,n4757,n5158);
nand (n5219,n5220,n5222);
or (n5220,n5221,n4775);
not (n5221,n5160);
nand (n5222,n4838,n5156);
nand (n5223,n5224,n5226);
or (n5224,n5225,n4802);
not (n5225,n5169);
nand (n5226,n4745,n5165);
and (n5227,n5197,n5228);
nand (n5228,n5229,n5318);
or (n5229,n5230,n5283);
not (n5230,n5231);
nand (n5231,n5232,n5257,n5270);
nor (n5232,n5233,n5240);
nand (n5233,n5234,n5236,n5238);
nand (n5234,n4742,n5235);
wire s0n5235,s1n5235,notn5235;
or (n5235,s0n5235,s1n5235);
not(notn5235,n4704);
and (s0n5235,notn5235,n2713);
and (s1n5235,n4704,n2780);
nand (n5236,n4745,n5237);
wire s0n5237,s1n5237,notn5237;
or (n5237,s0n5237,s1n5237);
not(notn5237,n4704);
and (s0n5237,notn5237,n2734);
and (s1n5237,n4704,n2793);
nand (n5238,n4739,n5239);
wire s0n5239,s1n5239,notn5239;
or (n5239,s0n5239,s1n5239);
not(notn5239,n4704);
and (s0n5239,notn5239,n2741);
and (s1n5239,n4704,n2802);
nand (n5240,n5241,n5244);
or (n5241,n5242,n4752);
not (n5242,n5243);
wire s0n5243,s1n5243,notn5243;
or (n5243,s0n5243,s1n5243);
not(notn5243,n4704);
and (s0n5243,notn5243,n2759);
and (s1n5243,n4704,n2820);
nor (n5244,n5245,n5251);
nand (n5245,n5246,n5249);
or (n5246,n5247,n4775);
not (n5247,n5248);
wire s0n5248,s1n5248,notn5248;
or (n5248,s0n5248,s1n5248);
not(notn5248,n4704);
and (s0n5248,notn5248,n2748);
and (s1n5248,n4704,n2809);
nand (n5249,n4838,n5250);
wire s0n5250,s1n5250,notn5250;
or (n5250,s0n5250,s1n5250);
not(notn5250,n4704);
and (s0n5250,notn5250,n2720);
and (s1n5250,n4704,n2784);
nand (n5251,n5252,n5255);
or (n5252,n5253,n4765);
not (n5253,n5254);
wire s0n5254,s1n5254,notn5254;
or (n5254,s0n5254,s1n5254);
not(notn5254,n4704);
and (s0n5254,notn5254,n2762);
and (s1n5254,n4704,n2823);
nand (n5255,n4757,n5256);
wire s0n5256,s1n5256,notn5256;
or (n5256,s0n5256,s1n5256);
not(notn5256,n4704);
and (s0n5256,notn5256,n2728);
and (s1n5256,n4704,n2797);
nor (n5257,n5258,n5264);
nand (n5258,n5259,n5262);
or (n5259,n5260,n4712);
not (n5260,n5261);
wire s0n5261,s1n5261,notn5261;
or (n5261,s0n5261,s1n5261);
not(notn5261,n4704);
and (s0n5261,notn5261,n2745);
and (s1n5261,n4704,n2806);
nand (n5262,n4707,n5263);
wire s0n5263,s1n5263,notn5263;
or (n5263,s0n5263,s1n5263);
not(notn5263,n4704);
and (s0n5263,notn5263,n2730);
and (s1n5263,n4704,n2795);
nand (n5264,n5265,n5268);
or (n5265,n5266,n4675);
not (n5266,n5267);
wire s0n5267,s1n5267,notn5267;
or (n5267,s0n5267,s1n5267);
not(notn5267,n4704);
and (s0n5267,notn5267,n2717);
and (s1n5267,n4704,n2782);
nand (n5268,n4721,n5269);
wire s0n5269,s1n5269,notn5269;
or (n5269,s0n5269,s1n5269);
not(notn5269,n4704);
and (s0n5269,notn5269,n2723);
and (s1n5269,n4704,n2778);
nor (n5270,n5271,n5277);
nand (n5271,n5272,n5275);
or (n5272,n5273,n4811);
not (n5273,n5274);
wire s0n5274,s1n5274,notn5274;
or (n5274,s0n5274,s1n5274);
not(notn5274,n4704);
and (s0n5274,notn5274,n2714);
and (s1n5274,n4704,n2776);
nand (n5275,n4724,n5276);
wire s0n5276,s1n5276,notn5276;
or (n5276,s0n5276,s1n5276);
not(notn5276,n4704);
and (s0n5276,notn5276,n2742);
and (s1n5276,n4704,n2803);
nand (n5277,n5278,n5281);
or (n5278,n5279,n4870);
not (n5279,n5280);
wire s0n5280,s1n5280,notn5280;
or (n5280,s0n5280,s1n5280);
not(notn5280,n4704);
and (s0n5280,notn5280,n2751);
and (s1n5280,n4704,n2812);
nand (n5281,n4727,n5282);
wire s0n5282,s1n5282,notn5282;
or (n5282,s0n5282,s1n5282);
not(notn5282,n4704);
and (s0n5282,notn5282,n2756);
and (s1n5282,n4704,n2817);
not (n5283,n5284);
nand (n5284,n5285,n5302,n5310);
nor (n5285,n5286,n5299);
nand (n5286,n5287,n5288,n5289);
nand (n5287,n4784,n5254);
nand (n5288,n4742,n5267);
nor (n5289,n5290,n5296);
nand (n5290,n5291,n5294);
or (n5291,n5292,n4756);
not (n5292,n5293);
wire s0n5293,s1n5293,notn5293;
or (n5293,s0n5293,s1n5293);
not(notn5293,n4704);
and (s0n5293,notn5293,n2736);
and (s1n5293,n4704,n2791);
nand (n5294,n4766,n5295);
wire s0n5295,s1n5295,notn5295;
or (n5295,s0n5295,s1n5295);
not(notn5295,n4704);
and (s0n5295,notn5295,n2765);
and (s1n5295,n4704,n2826);
nand (n5296,n5297,n5298);
or (n5297,n5279,n4775);
nand (n5298,n4838,n5269);
nand (n5299,n5300,n5301);
or (n5300,n5260,n4802);
nand (n5301,n4745,n5263);
nor (n5302,n5303,n5307);
nand (n5303,n5304,n5306);
or (n5304,n5305,n4675);
not (n5305,n5250);
nand (n5306,n4707,n5256);
nand (n5307,n5308,n5309);
or (n5308,n5247,n4712);
nand (n5309,n4715,n5282);
nor (n5310,n5311,n5315);
nand (n5311,n5312,n5314);
or (n5312,n5313,n4811);
not (n5313,n5235);
nand (n5314,n4721,n5237);
nand (n5315,n5316,n5317);
or (n5316,n5242,n4728);
nand (n5317,n4724,n5239);
or (n5318,n5319,n5402);
not (n5319,n5320);
and (n5320,n5321,n5372);
nand (n5321,n5322,n5346,n5359);
nor (n5322,n5323,n5330);
nand (n5323,n5324,n5326,n5328);
nand (n5324,n4742,n5325);
wire s0n5325,s1n5325,notn5325;
or (n5325,s0n5325,s1n5325);
not(notn5325,n4704);
and (s0n5325,notn5325,n2844);
and (s1n5325,n4704,n2901);
nand (n5326,n4739,n5327);
wire s0n5327,s1n5327,notn5327;
or (n5327,s0n5327,s1n5327);
not(notn5327,n4704);
and (s0n5327,notn5327,n2864);
and (s1n5327,n4704,n2927);
nand (n5328,n4745,n5329);
wire s0n5329,s1n5329,notn5329;
or (n5329,s0n5329,s1n5329);
not(notn5329,n4704);
and (s0n5329,notn5329,n2857);
and (s1n5329,n4704,n2917);
nand (n5330,n5331,n5334);
or (n5331,n5332,n4752);
not (n5332,n5333);
wire s0n5333,s1n5333,notn5333;
or (n5333,s0n5333,s1n5333);
not(notn5333,n4704);
and (s0n5333,notn5333,n2882);
and (s1n5333,n4704,n2945);
nor (n5334,n5335,n5340);
nand (n5335,n5336,n5338);
nand (n5336,n4776,n5337);
wire s0n5337,s1n5337,notn5337;
or (n5337,s0n5337,s1n5337);
not(notn5337,n4704);
and (s0n5337,notn5337,n2871);
and (s1n5337,n4704,n2934);
nand (n5338,n4838,n5339);
wire s0n5339,s1n5339,notn5339;
or (n5339,s0n5339,s1n5339);
not(notn5339,n4704);
and (s0n5339,notn5339,n2837);
and (s1n5339,n4704,n2898);
nand (n5340,n5341,n5344);
or (n5341,n5342,n4765);
not (n5342,n5343);
wire s0n5343,s1n5343,notn5343;
or (n5343,s0n5343,s1n5343);
not(notn5343,n4704);
and (s0n5343,notn5343,n2885);
and (s1n5343,n4704,n2948);
nand (n5344,n4757,n5345);
wire s0n5345,s1n5345,notn5345;
or (n5345,s0n5345,s1n5345);
not(notn5345,n4704);
and (s0n5345,notn5345,n2853);
and (s1n5345,n4704,n2914);
nor (n5346,n5347,n5353);
nand (n5347,n5348,n5351);
or (n5348,n5349,n4712);
not (n5349,n5350);
wire s0n5350,s1n5350,notn5350;
or (n5350,s0n5350,s1n5350);
not(notn5350,n4704);
and (s0n5350,notn5350,n2868);
and (s1n5350,n4704,n2931);
nand (n5351,n4707,n5352);
wire s0n5352,s1n5352,notn5352;
or (n5352,s0n5352,s1n5352);
not(notn5352,n4704);
and (s0n5352,notn5352,n2851);
and (s1n5352,n4704,n2912);
nand (n5353,n5354,n5357);
or (n5354,n5355,n5134);
not (n5355,n5356);
wire s0n5356,s1n5356,notn5356;
or (n5356,s0n5356,s1n5356);
not(notn5356,n4704);
and (s0n5356,notn5356,n2846);
and (s1n5356,n4704,n2907);
nand (n5357,n4674,n5358);
wire s0n5358,s1n5358,notn5358;
or (n5358,s0n5358,s1n5358);
not(notn5358,n4704);
and (s0n5358,notn5358,n2839);
and (s1n5358,n4704,n2896);
nor (n5359,n5360,n5366);
nand (n5360,n5361,n5364);
or (n5361,n5362,n4817);
not (n5362,n5363);
wire s0n5363,s1n5363,notn5363;
or (n5363,s0n5363,s1n5363);
not(notn5363,n4704);
and (s0n5363,notn5363,n2865);
and (s1n5363,n4704,n2928);
nand (n5364,n4715,n5365);
wire s0n5365,s1n5365,notn5365;
or (n5365,s0n5365,s1n5365);
not(notn5365,n4704);
and (s0n5365,notn5365,n2874);
and (s1n5365,n4704,n2937);
nand (n5366,n5367,n5370);
or (n5367,n5368,n4728);
not (n5368,n5369);
wire s0n5369,s1n5369,notn5369;
or (n5369,s0n5369,s1n5369);
not(notn5369,n4704);
and (s0n5369,notn5369,n2879);
and (s1n5369,n4704,n2942);
nand (n5370,n4734,n5371);
wire s0n5371,s1n5371,notn5371;
or (n5371,s0n5371,s1n5371);
not(notn5371,n4704);
and (s0n5371,notn5371,n2842);
and (s1n5371,n4704,n2905);
nand (n5372,n5373,n5384);
nor (n5373,n5374,n5379);
nand (n5374,n5375,n5376,n5377,n5378);
nand (n5375,n4707,n5345);
nand (n5376,n4711,n5337);
nand (n5377,n4674,n5339);
nand (n5378,n4734,n5325);
nand (n5379,n5380,n5381,n5382,n5383);
nand (n5380,n4715,n5369);
nand (n5381,n4727,n5333);
nand (n5382,n4721,n5329);
nand (n5383,n4724,n5327);
nor (n5384,n5385,n5389);
nand (n5385,n5386,n5387,n5388);
nand (n5386,n4739,n5350);
nand (n5387,n4742,n5358);
nand (n5388,n4745,n5352);
nand (n5389,n5390,n5391);
or (n5390,n5342,n4752);
nor (n5391,n5392,n5398);
nand (n5392,n5393,n5396);
or (n5393,n5394,n4756);
not (n5394,n5395);
wire s0n5395,s1n5395,notn5395;
or (n5395,s0n5395,s1n5395);
not(notn5395,n4704);
and (s0n5395,notn5395,n2859);
and (s1n5395,n4704,n2922);
nand (n5396,n4766,n5397);
wire s0n5397,s1n5397,notn5397;
or (n5397,s0n5397,s1n5397);
not(notn5397,n4704);
and (s0n5397,notn5397,n2888);
and (s1n5397,n4704,n2951);
nand (n5398,n5399,n5401);
or (n5399,n5400,n4775);
not (n5400,n5365);
nand (n5401,n4838,n5356);
and (n5402,n5230,n5283);
and (n5403,n5152,n5228);
and (n5404,n5067,n5150);
and (n5405,n4990,n5065);
and (n5406,n4956,n4988);
and (n5407,n4879,n4909);
and (n5408,n4780,n4823);
or (n5409,n5410,n5414);
xor (n5410,n5411,n4823);
not (n5411,n5412);
nand (n5412,n4668,n5413);
or (n5413,n4780,n4670);
or (n5414,n5415,n6036,n6119);
and (n5415,n5416,n5418);
xor (n5416,n5417,n4909);
xor (n5417,n4825,n4879);
nand (n5418,n5419,n6035);
or (n5419,n5420,n5496);
not (n5420,n5421);
nand (n5421,n5422,n5461);
nand (n5422,n5423,n5440,n5448);
nor (n5423,n5424,n5434);
and (n5424,n5425,n990);
not (n5425,n5426);
nor (n5426,n5427,n5431);
nand (n5427,n5428,n5430);
or (n5428,n4801,n5429);
not (n5429,n4716);
nand (n5430,n4676,n4718);
nand (n5431,n5432,n5433);
or (n5432,n4777,n4730);
nand (n5433,n4758,n4732);
and (n5434,n5435,n1056);
nand (n5435,n5436,n5437,n5438,n5439);
nand (n5436,n4729,n4773);
nand (n5437,n4716,n4703);
nand (n5438,n4676,n4722);
nand (n5439,n4758,n4747);
nor (n5440,n5441,n5445);
nand (n5441,n5442,n5444);
or (n5442,n5443,n5134);
not (n5443,n4709);
nand (n5444,n4745,n4763);
nand (n5445,n5446,n5447);
or (n5446,n4750,n4870);
nand (n5447,n4784,n4798);
nor (n5448,n5449,n5460);
nand (n5449,n5450,n5451);
or (n5450,n4794,n4708);
nor (n5451,n5452,n5456);
and (n5452,n4757,n5453);
wire s0n5453,s1n5453,notn5453;
or (n5453,s0n5453,s1n5453);
not(notn5453,n4704);
and (s0n5453,notn5453,n5454);
and (s1n5453,n4704,n5455);
and (n5456,n4766,n5457);
wire s0n5457,s1n5457,notn5457;
or (n5457,s0n5457,s1n5457);
not(notn5457,n4704);
and (s0n5457,notn5457,n5458);
and (s1n5457,n4704,n5459);
and (n5460,n4727,n4768);
nand (n5461,n5462,n5480);
nor (n5462,n5463,n5474);
nand (n5463,n5464,n5468,n5472,n5473);
nand (n5464,n4724,n5465);
wire s0n5465,s1n5465,notn5465;
or (n5465,s0n5465,s1n5465);
not(notn5465,n4704);
and (s0n5465,notn5465,n5466);
and (s1n5465,n4704,n5467);
nand (n5468,n4734,n5469);
wire s0n5469,s1n5469,notn5469;
or (n5469,s0n5469,s1n5469);
not(notn5469,n4704);
and (s0n5469,notn5469,n5470);
and (s1n5469,n4704,n5471);
nand (n5472,n4711,n4740);
nand (n5473,n4742,n4735);
nand (n5474,n5475,n5476,n5477);
nand (n5475,n4739,n4725);
nand (n5476,n4674,n4743);
nor (n5477,n5478,n5479);
and (n5478,n4838,n4703);
and (n5479,n4776,n4713);
nor (n5480,n5481,n5490);
and (n5481,n5482,n970);
nand (n5482,n5483,n5487);
not (n5483,n5484);
nand (n5484,n5485,n5486);
or (n5485,n4777,n5429);
nand (n5486,n4676,n4732);
nor (n5487,n5488,n5489);
and (n5488,n4758,n4751);
and (n5489,n4729,n4718);
and (n5490,n5491,n1041);
nand (n5491,n5492,n5493,n5494,n5495);
nand (n5492,n4716,n4773);
nand (n5493,n4729,n4722);
nand (n5494,n4676,n4747);
nand (n5495,n4758,n4709);
nand (n5496,n5497,n6034);
or (n5497,n5498,n5570);
not (n5498,n5499);
or (n5499,n5500,n5536);
nand (n5500,n5501,n5520);
nor (n5501,n5502,n5513);
nand (n5502,n5503,n5507,n5508,n5509);
nand (n5503,n4724,n5504);
wire s0n5504,s1n5504,notn5504;
or (n5504,s0n5504,s1n5504);
not(notn5504,n4704);
and (s0n5504,notn5504,n5505);
and (s1n5504,n4704,n5506);
nand (n5507,n4711,n4849);
nand (n5508,n4742,n4878);
nand (n5509,n4734,n5510);
wire s0n5510,s1n5510,notn5510;
or (n5510,s0n5510,s1n5510);
not(notn5510,n4704);
and (s0n5510,notn5510,n5511);
and (s1n5510,n4704,n5512);
nand (n5513,n5514,n5518,n5519);
not (n5514,n5515);
nand (n5515,n5516,n5517);
or (n5516,n4855,n4775);
nand (n5517,n4838,n4862);
nand (n5518,n4739,n4872);
nand (n5519,n4674,n4831);
nor (n5520,n5521,n5530);
and (n5521,n5522,n970);
nand (n5522,n5523,n5527);
not (n5523,n5524);
nand (n5524,n5525,n5526);
or (n5525,n4835,n5429);
nand (n5526,n4676,n4876);
nor (n5527,n5528,n5529);
and (n5528,n4758,n4829);
and (n5529,n4729,n4869);
and (n5530,n5531,n1041);
nand (n5531,n5532,n5533,n5534,n5535);
nand (n5532,n4729,n4864);
nand (n5533,n4716,n4839);
nand (n5534,n4676,n4851);
nand (n5535,n4758,n4858);
nand (n5536,n5537,n5557);
nor (n5537,n5538,n5543);
nand (n5538,n5539,n5540,n5541,n5542);
nand (n5539,n4784,n4904);
nand (n5540,n4715,n4829);
nand (n5541,n4721,n4858);
nand (n5542,n4745,n4845);
nand (n5543,n5544,n5555,n5556);
not (n5544,n5545);
nand (n5545,n5546,n5551);
or (n5546,n5547,n4756);
not (n5547,n5548);
wire s0n5548,s1n5548,notn5548;
or (n5548,s0n5548,s1n5548);
not(notn5548,n4704);
and (s0n5548,notn5548,n5549);
and (s1n5548,n4704,n5550);
nand (n5551,n4766,n5552);
wire s0n5552,s1n5552,notn5552;
or (n5552,s0n5552,s1n5552);
not(notn5552,n4704);
and (s0n5552,notn5552,n5553);
and (s1n5552,n4704,n5554);
nand (n5555,n4707,n4902);
nand (n5556,n4727,n4843);
nor (n5557,n5558,n5564);
and (n5558,n5559,n1056);
nand (n5559,n5560,n5561,n5562,n5563);
nand (n5560,n4729,n4839);
nand (n5561,n4716,n4862);
nand (n5562,n4676,n4864);
nand (n5563,n4758,n4851);
and (n5564,n5565,n990);
nand (n5565,n5566,n5567,n5568,n5569);
nand (n5566,n4729,n4836);
nand (n5567,n4716,n4856);
nand (n5568,n4676,n4869);
nand (n5569,n4758,n4876);
not (n5570,n5571);
nand (n5571,n5572,n6027);
or (n5572,n5573,n5719);
not (n5573,n5574);
nor (n5574,n5575,n5644);
nor (n5575,n5576,n5610);
nand (n5576,n5577,n5595);
nor (n5577,n5578,n5589);
nand (n5578,n5579,n5580,n5584,n5585);
nand (n5579,n4674,n4936);
nand (n5580,n4734,n5581);
wire s0n5581,s1n5581,notn5581;
or (n5581,s0n5581,s1n5581);
not(notn5581,n4704);
and (s0n5581,notn5581,n5582);
and (s1n5581,n4704,n5583);
nand (n5584,n4739,n4928);
nand (n5585,n4724,n5586);
wire s0n5586,s1n5586,notn5586;
or (n5586,s0n5586,s1n5586);
not(notn5586,n4704);
and (s0n5586,notn5586,n5587);
and (s1n5586,n4704,n5588);
nand (n5589,n5590,n5591,n5592);
nand (n5590,n4711,n4953);
nand (n5591,n4742,n4930);
nor (n5592,n5593,n5594);
and (n5593,n4776,n4915);
and (n5594,n4838,n4917);
nor (n5595,n5596,n5604);
and (n5596,n5597,n970);
nand (n5597,n5598,n5601);
nor (n5598,n5599,n5600);
and (n5599,n4716,n4943);
and (n5600,n4676,n4926);
nor (n5601,n5602,n5603);
and (n5602,n4758,n4934);
and (n5603,n4729,n4919);
and (n5604,n5605,n1041);
nand (n5605,n5606,n5607,n5608,n5609);
nand (n5606,n4729,n4924);
nand (n5607,n4716,n4941);
nand (n5608,n4676,n4955);
nand (n5609,n4758,n4921);
nand (n5610,n5611,n5629);
nor (n5611,n5612,n5625);
nand (n5612,n5613,n5614,n5615,n5616);
nand (n5613,n4707,n4980);
nand (n5614,n4727,n4947);
nand (n5615,n4745,n4949);
nor (n5616,n5617,n5621);
and (n5617,n4766,n5618);
wire s0n5618,s1n5618,notn5618;
or (n5618,s0n5618,s1n5618);
not(notn5618,n4704);
and (s0n5618,notn5618,n5619);
and (s1n5618,n4704,n5620);
and (n5621,n4757,n5622);
wire s0n5622,s1n5622,notn5622;
or (n5622,s0n5622,s1n5622);
not(notn5622,n4704);
and (s0n5622,notn5622,n5623);
and (s1n5622,n4704,n5624);
nand (n5625,n5626,n5627,n5628);
nand (n5626,n4721,n4921);
nand (n5627,n4715,n4934);
nand (n5628,n4784,n4982);
nor (n5629,n5630,n5638);
and (n5630,n5631,n1056);
nand (n5631,n5632,n5635);
nor (n5632,n5633,n5634);
and (n5633,n4716,n4917);
and (n5634,n4676,n4924);
nor (n5635,n5636,n5637);
and (n5636,n4758,n4955);
and (n5637,n4729,n4941);
and (n5638,n5639,n990);
nand (n5639,n5640,n5641,n5642,n5643);
nand (n5640,n4676,n4919);
nand (n5641,n4716,n4915);
nand (n5642,n4729,n4943);
nand (n5643,n4758,n4926);
nor (n5644,n5645,n5683);
nand (n5645,n5646,n5668);
nor (n5646,n5647,n5658);
nand (n5647,n5648,n5655);
not (n5648,n5649);
nand (n5649,n5650,n5652);
or (n5650,n5651,n4802);
not (n5651,n5047);
nor (n5652,n5653,n5654);
and (n5653,n4838,n5017);
and (n5654,n4776,n5015);
nor (n5655,n5656,n5657);
and (n5656,n4742,n5045);
and (n5657,n4674,n5009);
nand (n5658,n5659,n5663,n5664);
nand (n5659,n4724,n5660);
wire s0n5660,s1n5660,notn5660;
or (n5660,s0n5660,s1n5660);
not(notn5660,n4704);
and (s0n5660,notn5660,n5661);
and (s1n5660,n4704,n5662);
nand (n5663,n4711,n5007);
nand (n5664,n4734,n5665);
wire s0n5665,s1n5665,notn5665;
or (n5665,s0n5665,s1n5665);
not(notn5665,n4704);
and (s0n5665,notn5665,n5666);
and (s1n5665,n4704,n5667);
nor (n5668,n5669,n5677);
and (n5669,n5670,n970);
nand (n5670,n5671,n5674);
nor (n5671,n5672,n5673);
and (n5672,n4676,n5005);
and (n5673,n4716,n4996);
nor (n5674,n5675,n5676);
and (n5675,n4758,n5003);
and (n5676,n4729,n5026);
and (n5677,n5678,n1041);
nand (n5678,n5679,n5680,n5681,n5682);
nand (n5679,n4676,n4994);
nand (n5680,n4716,n4998);
nand (n5681,n4729,n5028);
nand (n5682,n4758,n5013);
nand (n5683,n5684,n5701);
nor (n5684,n5685,n5693);
and (n5685,n5686,n1056);
nand (n5686,n5687,n5690);
nor (n5687,n5688,n5689);
and (n5688,n4676,n5028);
and (n5689,n4716,n5017);
nor (n5690,n5691,n5692);
and (n5691,n4758,n4994);
and (n5692,n4729,n4998);
and (n5693,n5694,n990);
nand (n5694,n5695,n5698);
nor (n5695,n5696,n5697);
and (n5696,n4676,n5026);
and (n5697,n4716,n5015);
nor (n5698,n5699,n5700);
and (n5699,n4758,n5005);
and (n5700,n4729,n4996);
nor (n5701,n5702,n5715);
nand (n5702,n5703,n5704,n5705,n5706);
nand (n5703,n4727,n5021);
nand (n5704,n4745,n5000);
nand (n5705,n4784,n5033);
nor (n5706,n5707,n5711);
and (n5707,n4766,n5708);
wire s0n5708,s1n5708,notn5708;
or (n5708,s0n5708,s1n5708);
not(notn5708,n4704);
and (s0n5708,notn5708,n5709);
and (s1n5708,n4704,n5710);
and (n5711,n4757,n5712);
wire s0n5712,s1n5712,notn5712;
or (n5712,s0n5712,s1n5712);
not(notn5712,n4704);
and (s0n5712,notn5712,n5713);
and (s1n5712,n4704,n5714);
nand (n5715,n5716,n5717,n5718);
nand (n5716,n4715,n5003);
nand (n5717,n4721,n5013);
nand (n5718,n4707,n5031);
not (n5719,n5720);
nand (n5720,n5721,n6020);
or (n5721,n5722,n5872);
not (n5722,n5723);
nor (n5723,n5724,n5794);
nor (n5724,n5725,n5759);
nand (n5725,n5726,n5741);
nor (n5726,n5727,n5735);
and (n5727,n5728,n970);
nand (n5728,n5729,n5732);
nor (n5729,n5730,n5731);
and (n5730,n4716,n5073);
and (n5731,n4676,n5071);
nor (n5732,n5733,n5734);
and (n5733,n4758,n5084);
and (n5734,n4729,n5097);
and (n5735,n5736,n1041);
nand (n5736,n5737,n5738,n5739,n5740);
nand (n5737,n4729,n5099);
nand (n5738,n4716,n5075);
nand (n5739,n4676,n5080);
nand (n5740,n4758,n5111);
nor (n5741,n5742,n5752);
nand (n5742,n5743,n5747,n5751);
nand (n5743,n4724,n5744);
wire s0n5744,s1n5744,notn5744;
or (n5744,s0n5744,s1n5744);
not(notn5744,n4704);
and (s0n5744,notn5744,n5745);
and (s1n5744,n4704,n5746);
nand (n5747,n4734,n5748);
wire s0n5748,s1n5748,notn5748;
or (n5748,s0n5748,s1n5748);
not(notn5748,n4704);
and (s0n5748,notn5748,n5749);
and (s1n5748,n4704,n5750);
nand (n5751,n4711,n5082);
nand (n5752,n5753,n5754,n5755,n5756);
nand (n5753,n4674,n5086);
nand (n5754,n4742,n5148);
nand (n5755,n4739,n5143);
nor (n5756,n5757,n5758);
and (n5757,n4838,n5090);
and (n5758,n4776,n5109);
nand (n5759,n5760,n5776);
not (n5760,n5761);
nand (n5761,n5762,n5770);
or (n5762,n5763,n5764);
not (n5763,n990);
not (n5764,n5765);
nand (n5765,n5766,n5767,n5768,n5769);
nand (n5766,n4716,n5109);
nand (n5767,n4729,n5073);
nand (n5768,n4676,n5097);
nand (n5769,n4758,n5071);
nand (n5770,n5771,n1056);
nand (n5771,n5772,n5773,n5774,n5775);
nand (n5772,n4716,n5090);
nand (n5773,n4729,n5075);
nand (n5774,n4676,n5099);
nand (n5775,n4758,n5080);
nor (n5776,n5777,n5781);
nand (n5777,n5778,n5779,n5780);
nand (n5778,n4721,n5111);
nand (n5779,n4784,n5105);
nand (n5780,n4715,n5084);
nand (n5781,n5782,n5783,n5784,n5785);
nand (n5782,n4745,n5077);
nand (n5783,n4707,n5103);
nand (n5784,n4727,n5092);
nor (n5785,n5786,n5790);
and (n5786,n4766,n5787);
wire s0n5787,s1n5787,notn5787;
or (n5787,s0n5787,s1n5787);
not(notn5787,n4704);
and (s0n5787,notn5787,n5788);
and (s1n5787,n4704,n5789);
and (n5790,n4757,n5791);
wire s0n5791,s1n5791,notn5791;
or (n5791,s0n5791,s1n5791);
not(notn5791,n4704);
and (s0n5791,notn5791,n5792);
and (s1n5791,n4704,n5793);
nor (n5794,n5795,n5834);
nand (n5795,n5796,n5816);
nor (n5796,n5797,n5808);
and (n5797,n5798,n1056);
not (n5798,n5799);
nor (n5799,n5800,n5804);
nand (n5800,n5801,n5803);
or (n5801,n5802,n4677);
not (n5802,n5196);
nand (n5803,n4716,n5179);
nand (n5804,n5805,n5807);
or (n5805,n5806,n4730);
not (n5806,n5156);
nand (n5807,n4758,n5165);
and (n5808,n5809,n990);
nand (n5809,n5810,n5813);
nor (n5810,n5811,n5812);
and (n5811,n4676,n5194);
and (n5812,n4716,n5177);
nor (n5813,n5814,n5815);
and (n5814,n4758,n5162);
and (n5815,n4729,n5160);
nor (n5816,n5817,n5830);
nand (n5817,n5818,n5819,n5820,n5821);
nand (n5818,n4707,n5188);
nand (n5819,n4727,n5183);
nand (n5820,n4745,n5158);
nor (n5821,n5822,n5826);
and (n5822,n4757,n5823);
wire s0n5823,s1n5823,notn5823;
or (n5823,s0n5823,s1n5823);
not(notn5823,n4704);
and (s0n5823,notn5823,n5824);
and (s1n5823,n4704,n5825);
and (n5826,n4766,n5827);
wire s0n5827,s1n5827,notn5827;
or (n5827,s0n5827,s1n5827);
not(notn5827,n4704);
and (s0n5827,notn5827,n5828);
and (s1n5827,n4704,n5829);
nand (n5830,n5831,n5832,n5833);
nand (n5831,n4784,n5190);
nand (n5832,n4715,n5171);
nand (n5833,n4721,n5175);
nand (n5834,n5835,n5854);
nor (n5835,n5836,n5846);
and (n5836,n5837,n970);
not (n5837,n5838);
nor (n5838,n5839,n5843);
nand (n5839,n5840,n5842);
or (n5840,n5841,n4677);
not (n5841,n5162);
nand (n5842,n4716,n5160);
nand (n5843,n5844,n5845);
or (n5844,n5193,n4730);
nand (n5845,n4758,n5171);
and (n5846,n5847,n1041);
nand (n5847,n5848,n5851);
nor (n5848,n5849,n5850);
and (n5849,n4676,n5165);
and (n5850,n4716,n5156);
nor (n5851,n5852,n5853);
and (n5852,n4758,n5175);
and (n5853,n4729,n5196);
nor (n5854,n5855,n5862);
nand (n5855,n5856,n5857,n5858,n5859);
nand (n5856,n4711,n5169);
nand (n5857,n4739,n5206);
nand (n5858,n4742,n5210);
nor (n5859,n5860,n5861);
and (n5860,n4838,n5179);
and (n5861,n4776,n5177);
nand (n5862,n5863,n5864,n5868);
nand (n5863,n4674,n5167);
nand (n5864,n4734,n5865);
wire s0n5865,s1n5865,notn5865;
or (n5865,s0n5865,s1n5865);
not(notn5865,n4704);
and (s0n5865,notn5865,n5866);
and (s1n5865,n4704,n5867);
nand (n5868,n4724,n5869);
wire s0n5869,s1n5869,notn5869;
or (n5869,s0n5869,s1n5869);
not(notn5869,n4704);
and (s0n5869,notn5869,n5870);
and (s1n5869,n4704,n5871);
not (n5872,n5873);
nand (n5873,n5874,n6019);
or (n5874,n5875,n5947);
nor (n5875,n5876,n5912);
nand (n5876,n5877,n5885,n5900,n5906);
nor (n5877,n5878,n5883);
nand (n5878,n5879,n5880);
or (n5879,n5313,n4675);
nor (n5880,n5881,n5882);
and (n5881,n4838,n5267);
and (n5882,n4776,n5261);
nor (n5883,n5884,n5273);
not (n5884,n4742);
nor (n5885,n5886,n5893);
nand (n5886,n5887,n5889);
or (n5887,n5888,n4712);
not (n5888,n5239);
nand (n5889,n4724,n5890);
wire s0n5890,s1n5890,notn5890;
or (n5890,s0n5890,s1n5890);
not(notn5890,n4704);
and (s0n5890,notn5890,n5891);
and (s1n5890,n4704,n5892);
nand (n5893,n5894,n5899);
or (n5894,n5895,n4811);
not (n5895,n5896);
wire s0n5896,s1n5896,notn5896;
or (n5896,s0n5896,s1n5896);
not(notn5896,n4704);
and (s0n5896,notn5896,n5897);
and (s1n5896,n4704,n5898);
nand (n5899,n4739,n5276);
nand (n5900,n5901,n1041);
nand (n5901,n5902,n5903,n5904,n5905);
nand (n5902,n4729,n5269);
nand (n5903,n4716,n5250);
nand (n5904,n4676,n5237);
nand (n5905,n4758,n5263);
nand (n5906,n5907,n970);
nand (n5907,n5908,n5909,n5910,n5911);
nand (n5908,n4729,n5280);
nand (n5909,n4716,n5248);
nand (n5910,n4676,n5282);
nand (n5911,n4758,n5243);
nand (n5912,n5913,n5921,n5935,n5941);
nor (n5913,n5914,n5917);
nand (n5914,n5915,n5916);
or (n5915,n5242,n4870);
nand (n5916,n4784,n5295);
nand (n5917,n5918,n5920);
or (n5918,n5919,n5134);
not (n5919,n5263);
nand (n5920,n4727,n5254);
nor (n5921,n5922,n5933);
nand (n5922,n5923,n5924);
or (n5923,n5292,n4708);
nor (n5924,n5925,n5929);
and (n5925,n4766,n5926);
wire s0n5926,s1n5926,notn5926;
or (n5926,s0n5926,s1n5926);
not(notn5926,n4704);
and (s0n5926,notn5926,n5927);
and (s1n5926,n4704,n5928);
and (n5929,n4757,n5930);
wire s0n5930,s1n5930,notn5930;
or (n5930,s0n5930,s1n5930);
not(notn5930,n4704);
and (s0n5930,notn5930,n5931);
and (s1n5930,n4704,n5932);
nor (n5933,n5934,n4746);
not (n5934,n5256);
nand (n5935,n5936,n990);
nand (n5936,n5937,n5938,n5939,n5940);
nand (n5937,n4729,n5248);
nand (n5938,n4716,n5261);
nand (n5939,n4676,n5280);
nand (n5940,n4758,n5282);
nand (n5941,n5942,n1056);
nand (n5942,n5943,n5944,n5945,n5946);
nand (n5943,n4729,n5250);
nand (n5944,n4716,n5267);
nand (n5945,n4676,n5269);
nand (n5946,n4758,n5237);
nand (n5947,n5948,n5984);
nand (n5948,n5949,n5957,n5972,n5978);
nor (n5949,n5950,n5951);
and (n5950,n4742,n5371);
nand (n5951,n5952,n5954);
or (n5952,n5953,n4675);
not (n5953,n5325);
nor (n5954,n5955,n5956);
and (n5955,n4838,n5358);
and (n5956,n4776,n5350);
nor (n5957,n5958,n5965);
nand (n5958,n5959,n5961);
or (n5959,n5960,n4712);
not (n5960,n5327);
nand (n5961,n4724,n5962);
wire s0n5962,s1n5962,notn5962;
or (n5962,s0n5962,s1n5962);
not(notn5962,n4704);
and (s0n5962,notn5962,n5963);
and (s1n5962,n4704,n5964);
nand (n5965,n5966,n5971);
or (n5966,n5967,n4811);
not (n5967,n5968);
wire s0n5968,s1n5968,notn5968;
or (n5968,s0n5968,s1n5968);
not(notn5968,n4704);
and (s0n5968,notn5968,n5969);
and (s1n5968,n4704,n5970);
nand (n5971,n4739,n5363);
nand (n5972,n5973,n1041);
nand (n5973,n5974,n5975,n5976,n5977);
nand (n5974,n4729,n5356);
nand (n5975,n4716,n5339);
nand (n5976,n4676,n5329);
nand (n5977,n4758,n5352);
nand (n5978,n5979,n970);
nand (n5979,n5980,n5981,n5982,n5983);
nand (n5980,n4729,n5365);
nand (n5981,n4716,n5337);
nand (n5982,n4676,n5369);
nand (n5983,n4758,n5333);
nand (n5984,n5985,n5992,n6007,n6013);
nor (n5985,n5986,n5989);
nand (n5986,n5987,n5988);
or (n5987,n5394,n4708);
nand (n5988,n4721,n5352);
nand (n5989,n5990,n5991);
or (n5990,n5332,n4870);
nand (n5991,n4727,n5343);
nor (n5992,n5993,n6005);
nand (n5993,n5994,n5996);
or (n5994,n5995,n4752);
not (n5995,n5397);
nor (n5996,n5997,n6001);
and (n5997,n4766,n5998);
wire s0n5998,s1n5998,notn5998;
or (n5998,s0n5998,s1n5998);
not(notn5998,n4704);
and (s0n5998,notn5998,n5999);
and (s1n5998,n4704,n6000);
and (n6001,n4757,n6002);
wire s0n6002,s1n6002,notn6002;
or (n6002,s0n6002,s1n6002);
not(notn6002,n4704);
and (s0n6002,notn6002,n6003);
and (s1n6002,n4704,n6004);
nor (n6005,n4746,n6006);
not (n6006,n5345);
nand (n6007,n6008,n990);
nand (n6008,n6009,n6010,n6011,n6012);
nand (n6009,n4729,n5337);
nand (n6010,n4716,n5350);
nand (n6011,n4676,n5365);
nand (n6012,n4758,n5369);
nand (n6013,n6014,n1056);
nand (n6014,n6015,n6016,n6017,n6018);
nand (n6015,n4729,n5339);
nand (n6016,n4716,n5358);
nand (n6017,n4676,n5356);
nand (n6018,n4758,n5329);
nand (n6019,n5876,n5912);
nor (n6020,n6021,n6025);
and (n6021,n6022,n6023);
not (n6022,n5724);
not (n6023,n6024);
nand (n6024,n5795,n5834);
not (n6025,n6026);
nand (n6026,n5725,n5759);
nand (n6027,n6028,n6033);
or (n6028,n6029,n6031);
not (n6029,n6030);
nand (n6030,n5610,n5576);
not (n6031,n6032);
nand (n6032,n5683,n5645);
not (n6033,n5575);
nand (n6034,n5536,n5500);
or (n6035,n5422,n5461);
and (n6036,n5418,n6037);
or (n6037,n6038,n6047,n6118);
and (n6038,n6039,n6041);
xor (n6039,n6040,n4988);
xor (n6040,n4911,n4956);
nor (n6041,n6042,n6044);
and (n6042,n6043,n5496);
nand (n6043,n6035,n5421);
and (n6044,n6045,n6046);
not (n6045,n6043);
not (n6046,n5496);
and (n6047,n6041,n6048);
or (n6048,n6049,n6058,n6117);
and (n6049,n6050,n6053);
xor (n6050,n6051,n5065);
not (n6051,n6052);
xnor (n6052,n5034,n4990);
nor (n6053,n6054,n6056);
and (n6054,n5571,n6055);
nand (n6055,n5499,n6034);
and (n6056,n5570,n6057);
not (n6057,n6055);
and (n6058,n6053,n6059);
or (n6059,n6060,n6073,n6116);
and (n6060,n6061,n6065);
xor (n6061,n6062,n5150);
not (n6062,n6063);
xor (n6063,n5067,n6064);
not (n6064,n5112);
nor (n6065,n6066,n6070);
and (n6066,n6067,n6069);
nand (n6067,n6068,n6032);
or (n6068,n5644,n5719);
nand (n6069,n6033,n6030);
and (n6070,n6071,n6072);
not (n6071,n6067);
not (n6072,n6069);
and (n6073,n6065,n6074);
or (n6074,n6075,n6089,n6115);
and (n6075,n6076,n6083);
xor (n6076,n6077,n5228);
not (n6077,n6078);
nor (n6078,n6079,n6081);
and (n6079,n5197,n6080);
not (n6080,n5152);
and (n6081,n6082,n5152);
not (n6082,n5197);
nand (n6083,n6084,n6088);
or (n6084,n6085,n5720);
not (n6085,n6086);
nand (n6086,n6087,n6032);
not (n6087,n5644);
nand (n6088,n6085,n5720);
and (n6089,n6083,n6090);
or (n6090,n6091,n6105,n6114);
not (n6091,n6092);
nand (n6092,n6093,n6101);
nand (n6093,n6094,n6100);
or (n6094,n6095,n6097);
not (n6095,n6096);
nor (n6096,n5724,n6025);
not (n6097,n6098);
nand (n6098,n6099,n6024);
or (n6099,n5794,n5872);
or (n6100,n6098,n6096);
nand (n6101,n6102,n6104);
or (n6102,n6103,n5319);
xor (n6103,n5230,n5283);
nand (n6104,n5319,n6103);
and (n6105,n6093,n6106);
not (n6106,n6107);
nand (n6107,n6108,n6113);
nand (n6108,n6109,n6112);
or (n6109,n6110,n5872);
nand (n6110,n6111,n6024);
not (n6111,n5794);
nand (n6112,n5872,n6110);
xor (n6113,n5321,n5372);
and (n6114,n6101,n6106);
and (n6115,n6076,n6090);
and (n6116,n6061,n6074);
and (n6117,n6050,n6059);
and (n6118,n6039,n6048);
and (n6119,n5416,n6037);
and (n6120,n6121,n6122);
xnor (n6121,n5410,n5414);
and (n6122,n6123,n6125);
xor (n6123,n6124,n6037);
xor (n6124,n5416,n5418);
and (n6125,n6126,n6128);
xor (n6126,n6127,n6048);
xor (n6127,n6039,n6041);
and (n6128,n6129,n6131);
xor (n6129,n6130,n6059);
xor (n6130,n6050,n6053);
and (n6131,n6132,n6134);
xor (n6132,n6133,n6074);
xor (n6133,n6061,n6065);
and (n6134,n6135,n6137);
xor (n6135,n6136,n6090);
xor (n6136,n6076,n6083);
and (n6137,n6138,n6140);
xor (n6138,n6139,n6106);
xor (n6139,n6101,n6093);
and (n6140,n6141,n6142);
xor (n6141,n6113,n6108);
not (n6142,n6143);
nand (n6143,n6144,n6150);
not (n6144,n6145);
xor (n6145,n6146,n6149);
not (n6146,n6147);
nand (n6147,n6148,n6019);
not (n6148,n5875);
not (n6149,n5947);
not (n6150,n6151);
xor (n6151,n5948,n5984);
and (n6152,n6153,n6154);
xor (n6153,n6121,n6122);
or (n6154,n6155,n6592,n6655);
and (n6155,n6156,n6591);
or (n6156,n6157,n6216,n6590);
and (n6157,n6158,n6187);
nand (n6158,n6159,n6167,n6179,n6183);
nor (n6159,n6160,n6164);
and (n6160,n6161,n6163);
not (n6161,n6162);
nand (n6162,n4724,n4705);
and (n6164,n6165,n6166);
nor (n6165,n4817,n4705);
nor (n6167,n6168,n6175);
nand (n6168,n6169,n6170,n6171,n6172);
nand (n6169,n5435,n1041);
nand (n6170,n4674,n4735);
nand (n6171,n4742,n5469);
nor (n6172,n6173,n6174);
and (n6173,n4838,n4743);
and (n6174,n4776,n4740);
nand (n6175,n6176,n6177,n6178);
nand (n6176,n5425,n970);
nand (n6177,n4711,n4725);
nand (n6178,n4739,n5465);
nand (n6179,n6180,n6182);
not (n6180,n6181);
nand (n6181,n4734,n4705);
nand (n6183,n6184,n6186);
not (n6184,n6185);
nand (n6185,n4734,n4704);
nand (n6187,n6188,n6197,n6208);
nor (n6188,n6189,n6194);
nand (n6189,n6190,n6191,n6192,n6193);
nand (n6190,n4784,n5457);
nand (n6191,n4707,n5453);
nand (n6192,n4715,n4768);
nand (n6193,n4721,n4763);
and (n6194,n6195,n6196);
and (n6195,n4766,n4704);
nor (n6197,n6198,n6202);
nand (n6198,n6199,n6200,n6201);
nand (n6199,n5482,n990);
nand (n6200,n4727,n4798);
nand (n6201,n4745,n4795);
nand (n6202,n6203,n6205);
or (n6203,n2771,n6204);
not (n6204,n5491);
nand (n6205,n6206,n6207);
and (n6206,n4766,n4705);
nor (n6208,n6209,n6212);
and (n6209,n6210,n6211);
and (n6210,n4757,n4705);
and (n6212,n6213,n6215);
not (n6213,n6214);
nand (n6214,n4757,n4704);
and (n6216,n6158,n6217);
or (n6217,n6218,n6265,n6589);
and (n6218,n6219,n6243);
nand (n6219,n6220,n6228,n6238);
nor (n6220,n6221,n6226);
nand (n6221,n6222,n6223,n6224,n6225);
nand (n6222,n4784,n5552);
nand (n6223,n4707,n5548);
nand (n6224,n4715,n4843);
nand (n6225,n4721,n4845);
and (n6226,n6213,n6227);
nor (n6228,n6229,n6233);
nand (n6229,n6230,n6231,n6232);
nand (n6230,n5522,n990);
nand (n6231,n4727,n4904);
nand (n6232,n4745,n4902);
nand (n6233,n6234,n6236);
or (n6234,n2771,n6235);
not (n6235,n5531);
nand (n6236,n6206,n6237);
nor (n6238,n6239,n6241);
and (n6239,n6210,n6240);
and (n6241,n6195,n6242);
nand (n6243,n6244,n6249,n6261,n6263);
nor (n6244,n6245,n6247);
and (n6245,n6161,n6246);
and (n6247,n6165,n6248);
nor (n6249,n6250,n6257);
nand (n6250,n6251,n6252,n6253,n6254);
nand (n6251,n5559,n1041);
nand (n6252,n4674,n4878);
nand (n6253,n4742,n5510);
nor (n6254,n6255,n6256);
and (n6255,n4838,n4831);
and (n6256,n4776,n4849);
nand (n6257,n6258,n6259,n6260);
nand (n6258,n5565,n970);
nand (n6259,n4711,n4872);
nand (n6260,n4739,n5504);
nand (n6261,n6180,n6262);
nand (n6263,n6184,n6264);
and (n6265,n6243,n6266);
or (n6266,n6267,n6314,n6588);
and (n6267,n6268,n6292);
nand (n6268,n6269,n6277,n6287);
nor (n6269,n6270,n6275);
nand (n6270,n6271,n6272,n6273,n6274);
nand (n6271,n5618,n4784);
nand (n6272,n4707,n5622);
nand (n6273,n4715,n4947);
nand (n6274,n4721,n4949);
and (n6275,n6195,n6276);
nor (n6277,n6278,n6282);
nand (n6278,n6279,n6280,n6281);
nand (n6279,n5597,n990);
nand (n6280,n4727,n4982);
nand (n6281,n4745,n4980);
nand (n6282,n6283,n6285);
or (n6283,n2771,n6284);
not (n6284,n5605);
nand (n6285,n6206,n6286);
nor (n6287,n6288,n6290);
and (n6288,n6213,n6289);
and (n6290,n6210,n6291);
nand (n6292,n6293,n6298,n6310,n6312);
nor (n6293,n6294,n6296);
and (n6294,n6161,n6295);
and (n6296,n6165,n6297);
nor (n6298,n6299,n6306);
nand (n6299,n6300,n6301,n6302,n6303);
nand (n6300,n5631,n1041);
nand (n6301,n4674,n4930);
nand (n6302,n4742,n5581);
nor (n6303,n6304,n6305);
and (n6304,n4838,n4936);
and (n6305,n4776,n4953);
nand (n6306,n6307,n6308,n6309);
nand (n6307,n5639,n970);
nand (n6308,n4711,n4928);
nand (n6309,n4739,n5586);
nand (n6310,n6180,n6311);
nand (n6312,n6184,n6313);
and (n6314,n6292,n6315);
or (n6315,n6316,n6364,n6587);
and (n6316,n6317,n6341);
nand (n6317,n6318,n6328,n6336);
nor (n6318,n6319,n6323);
nand (n6319,n6320,n6321,n6322);
nand (n6320,n5670,n990);
nand (n6321,n4727,n5033);
nand (n6322,n4745,n5031);
nand (n6323,n6324,n6326);
or (n6324,n2771,n6325);
not (n6325,n5678);
nand (n6326,n6206,n6327);
nor (n6328,n6329,n6334);
nand (n6329,n6330,n6331,n6332,n6333);
nand (n6330,n4721,n5000);
nand (n6331,n5708,n4784);
nand (n6332,n4707,n5712);
nand (n6333,n4715,n5021);
and (n6334,n6195,n6335);
nor (n6336,n6337,n6339);
and (n6337,n6213,n6338);
and (n6339,n6210,n6340);
nand (n6341,n6342,n6359);
and (n6342,n6343,n6355,n6357);
nor (n6343,n6344,n6351);
nand (n6344,n6345,n6346,n6347,n6348);
nand (n6345,n5694,n970);
nand (n6346,n4674,n5045);
nand (n6347,n4742,n5665);
nor (n6348,n6349,n6350);
and (n6349,n4838,n5009);
and (n6350,n4776,n5007);
nand (n6351,n6352,n6353,n6354);
nand (n6352,n5686,n1041);
nand (n6353,n4711,n5047);
nand (n6354,n4739,n5660);
nand (n6355,n6180,n6356);
nand (n6357,n6161,n6358);
nor (n6359,n6360,n6362);
and (n6360,n6165,n6361);
and (n6362,n6184,n6363);
and (n6364,n6341,n6365);
or (n6365,n6366,n6420,n6586);
and (n6366,n6367,n6395);
nand (n6367,n6368,n6380,n6390);
nor (n6368,n6369,n6372,n6376);
nand (n6369,n6370,n6371);
or (n6370,n5128,n4870);
nand (n6371,n4721,n5077);
nand (n6372,n6373,n6375);
or (n6373,n6374,n4708);
not (n6374,n5791);
nand (n6375,n5787,n4784);
nor (n6376,n6377,n6379);
not (n6377,n6378);
not (n6379,n6195);
nor (n6380,n6381,n6385);
nand (n6381,n6382,n6383,n6384);
nand (n6382,n5728,n990);
nand (n6383,n4727,n5105);
nand (n6384,n4745,n5103);
nand (n6385,n6386,n6388);
or (n6386,n2771,n6387);
not (n6387,n5736);
nand (n6388,n6206,n6389);
nor (n6390,n6391,n6393);
and (n6391,n6213,n6392);
and (n6393,n6210,n6394);
nand (n6395,n6396,n6413,n6418);
not (n6396,n6397);
nand (n6397,n6398,n6401);
or (n6398,n6399,n6181);
not (n6399,n6400);
nor (n6401,n6402,n6409);
nand (n6402,n6403,n6404,n6405,n6406);
nand (n6403,n5771,n1041);
nand (n6404,n4674,n5148);
nand (n6405,n4742,n5748);
nor (n6406,n6407,n6408);
and (n6407,n4838,n5086);
and (n6408,n4776,n5082);
nand (n6409,n6410,n6411,n6412);
nand (n6410,n5765,n970);
nand (n6411,n4739,n5744);
nand (n6412,n4711,n5143);
nor (n6413,n6414,n6416);
and (n6414,n6161,n6415);
and (n6416,n6165,n6417);
nand (n6418,n6184,n6419);
and (n6420,n6395,n6421);
or (n6421,n6422,n6470,n6585);
and (n6422,n6423,n6447);
nand (n6423,n6424,n6432,n6442);
nor (n6424,n6425,n6430);
nand (n6425,n6426,n6427,n6428,n6429);
nand (n6426,n4721,n5158);
nand (n6427,n4784,n5827);
nand (n6428,n5823,n4707);
nand (n6429,n4715,n5183);
and (n6430,n6195,n6431);
nor (n6432,n6433,n6437);
nand (n6433,n6434,n6435,n6436);
nand (n6434,n4727,n5190);
nand (n6435,n5837,n990);
nand (n6436,n4745,n5188);
nand (n6437,n6438,n6440);
or (n6438,n2771,n6439);
not (n6439,n5847);
nand (n6440,n6206,n6441);
nor (n6442,n6443,n6445);
and (n6443,n6213,n6444);
and (n6445,n6210,n6446);
nand (n6447,n6448,n6465);
and (n6448,n6449,n6461,n6463);
nor (n6449,n6450,n6457);
nand (n6450,n6451,n6452,n6453,n6454);
nand (n6451,n5798,n1041);
nand (n6452,n4674,n5210);
nand (n6453,n4742,n5865);
nor (n6454,n6455,n6456);
and (n6455,n4838,n5167);
and (n6456,n4776,n5169);
nand (n6457,n6458,n6459,n6460);
nand (n6458,n5809,n970);
nand (n6459,n4739,n5869);
nand (n6460,n5206,n4711);
nand (n6461,n6180,n6462);
nand (n6463,n6184,n6464);
nor (n6465,n6466,n6468);
and (n6466,n6161,n6467);
and (n6468,n6165,n6469);
and (n6470,n6447,n6471);
or (n6471,n6472,n6525,n6584);
and (n6472,n6473,n6500);
nand (n6473,n6474,n6485,n6495);
nor (n6474,n6475,n6478,n6482);
nand (n6475,n6476,n6477);
or (n6476,n5253,n4870);
nand (n6477,n4721,n5256);
nand (n6478,n6479,n6481);
or (n6479,n6480,n4708);
not (n6480,n5930);
nand (n6481,n5926,n4784);
nor (n6482,n6483,n6379);
not (n6483,n6484);
nor (n6485,n6486,n6490);
nand (n6486,n6487,n6488,n6489);
nand (n6487,n5907,n990);
nand (n6488,n4727,n5295);
nand (n6489,n4745,n5293);
nand (n6490,n6491,n6493);
or (n6491,n2771,n6492);
not (n6492,n5901);
nand (n6493,n6206,n6494);
nor (n6495,n6496,n6498);
and (n6496,n6213,n6497);
and (n6498,n6210,n6499);
nand (n6500,n6501,n6518,n6523);
not (n6501,n6502);
nand (n6502,n6503,n6506);
or (n6503,n6504,n6181);
not (n6504,n6505);
nor (n6506,n6507,n6514);
nand (n6507,n6508,n6509,n6510,n6511);
nand (n6508,n5942,n1041);
nand (n6509,n4674,n5274);
nand (n6510,n4742,n5896);
nor (n6511,n6512,n6513);
and (n6512,n4838,n5235);
and (n6513,n4776,n5239);
nand (n6514,n6515,n6516,n6517);
nand (n6515,n5936,n970);
nand (n6516,n4739,n5890);
nand (n6517,n4711,n5276);
nor (n6518,n6519,n6521);
and (n6519,n6161,n6520);
and (n6521,n6165,n6522);
nand (n6523,n6184,n6524);
and (n6525,n6500,n6526);
and (n6526,n6527,n6559);
nand (n6527,n6528,n6546);
not (n6528,n6529);
nand (n6529,n6530,n6536,n6539,n6544);
not (n6530,n6531);
nand (n6531,n6532,n6534);
or (n6532,n4708,n6533);
not (n6533,n6002);
or (n6534,n4752,n6535);
not (n6535,n5998);
nor (n6536,n6537,n6538);
and (n6537,n4721,n5345);
and (n6538,n4715,n5343);
nor (n6539,n6540,n6542);
and (n6540,n6213,n6541);
and (n6542,n6210,n6543);
nand (n6544,n6195,n6545);
nor (n6546,n6547,n6552);
nand (n6547,n6548,n6550,n6551);
or (n6548,n6549,n5763);
not (n6549,n5979);
or (n6550,n4728,n5995);
or (n6551,n4746,n5394);
nand (n6552,n6553,n6557);
or (n6553,n6554,n6556);
not (n6554,n6555);
not (n6556,n6206);
or (n6557,n6558,n2771);
not (n6558,n5973);
nand (n6559,n6560,n6579);
and (n6560,n6561,n6575,n6577);
nor (n6561,n6562,n6569);
nand (n6562,n6563,n6564,n6565,n6566);
nand (n6563,n6014,n1041);
nand (n6564,n4739,n5962);
nand (n6565,n4711,n5363);
nor (n6566,n6567,n6568);
and (n6567,n4776,n5327);
and (n6568,n4838,n5325);
nand (n6569,n6570,n6572,n6574);
or (n6570,n6571,n971);
not (n6571,n6008);
or (n6572,n4675,n6573);
not (n6573,n5371);
nand (n6574,n4742,n5968);
nand (n6575,n6180,n6576);
nand (n6577,n6184,n6578);
nor (n6579,n6580,n6582);
and (n6580,n6161,n6581);
and (n6582,n6165,n6583);
and (n6584,n6473,n6526);
and (n6585,n6423,n6471);
and (n6586,n6367,n6421);
and (n6587,n6317,n6365);
and (n6588,n6268,n6315);
and (n6589,n6219,n6266);
and (n6590,n6187,n6217);
xor (n6591,n6123,n6125);
and (n6592,n6591,n6593);
or (n6593,n6594,n6598,n6654);
and (n6594,n6595,n6597);
xor (n6595,n6596,n6217);
xor (n6596,n6158,n6187);
xor (n6597,n6126,n6128);
and (n6598,n6597,n6599);
or (n6599,n6600,n6604,n6653);
and (n6600,n6601,n6603);
xor (n6601,n6602,n6266);
xor (n6602,n6219,n6243);
xor (n6603,n6129,n6131);
and (n6604,n6603,n6605);
or (n6605,n6606,n6610,n6652);
and (n6606,n6607,n6609);
xor (n6607,n6608,n6315);
xor (n6608,n6268,n6292);
xor (n6609,n6132,n6134);
and (n6610,n6609,n6611);
or (n6611,n6612,n6627,n6651);
and (n6612,n6613,n6615);
xor (n6613,n6614,n6365);
xor (n6614,n6317,n6341);
xor (n6615,n6616,n6624);
xor (n6616,n5228,n6617);
nand (n6617,n6618,n6092);
or (n6618,n6619,n6623);
not (n6619,n6620);
nand (n6620,n6621,n6107);
or (n6621,n6622,n6143);
nor (n6622,n6108,n6113);
nor (n6623,n6093,n6101);
nand (n6624,n6625,n6626);
or (n6625,n6078,n6083);
nand (n6626,n6083,n6078);
and (n6627,n6615,n6628);
or (n6628,n6629,n6633,n6650);
and (n6629,n6630,n6632);
xor (n6630,n6631,n6421);
xor (n6631,n6367,n6395);
xor (n6632,n6138,n6140);
and (n6633,n6632,n6634);
or (n6634,n6635,n6639,n6649);
and (n6635,n6636,n6638);
xor (n6636,n6637,n6471);
xor (n6637,n6423,n6447);
xor (n6638,n6141,n6142);
and (n6639,n6638,n6640);
or (n6640,n6641,n6645,n6648);
and (n6641,n6642,n6644);
xor (n6642,n6643,n6526);
xor (n6643,n6473,n6500);
xor (n6644,n6144,n6150);
and (n6645,n6644,n6646);
and (n6646,n6647,n6151);
xor (n6647,n6527,n6559);
and (n6648,n6642,n6646);
and (n6649,n6636,n6640);
and (n6650,n6630,n6634);
and (n6651,n6613,n6628);
and (n6652,n6607,n6611);
and (n6653,n6601,n6605);
and (n6654,n6595,n6599);
and (n6655,n6156,n6593);
or (n6656,n6657,n6659,n6699);
and (n6657,n6658,n6597);
xor (n6658,n6153,n6154);
and (n6659,n6597,n6660);
or (n6660,n6661,n6664,n6698);
and (n6661,n6662,n6603);
xor (n6662,n6663,n6593);
xor (n6663,n6156,n6591);
and (n6664,n6603,n6665);
or (n6665,n6666,n6669,n6697);
and (n6666,n6667,n6609);
xor (n6667,n6668,n6599);
xor (n6668,n6595,n6597);
and (n6669,n6609,n6670);
or (n6670,n6671,n6674,n6696);
and (n6671,n6672,n6615);
xor (n6672,n6673,n6605);
xor (n6673,n6601,n6603);
and (n6674,n6615,n6675);
or (n6675,n6676,n6679,n6695);
and (n6676,n6677,n6632);
xor (n6677,n6678,n6611);
xor (n6678,n6607,n6609);
and (n6679,n6632,n6680);
or (n6680,n6681,n6684,n6694);
and (n6681,n6682,n6638);
xor (n6682,n6683,n6628);
xor (n6683,n6613,n6615);
and (n6684,n6638,n6685);
or (n6685,n6686,n6689,n6693);
and (n6686,n6687,n6644);
xor (n6687,n6688,n6634);
xor (n6688,n6630,n6632);
and (n6689,n6644,n6690);
and (n6690,n6691,n6151);
xor (n6691,n6692,n6640);
xor (n6692,n6636,n6638);
and (n6693,n6687,n6690);
and (n6694,n6682,n6685);
and (n6695,n6677,n6680);
and (n6696,n6672,n6675);
and (n6697,n6667,n6670);
and (n6698,n6662,n6665);
and (n6699,n6658,n6660);
and (n6700,n6701,n6703);
xor (n6701,n6702,n6660);
xor (n6702,n6658,n6597);
and (n6703,n6704,n6706);
xor (n6704,n6705,n6665);
xor (n6705,n6662,n6603);
and (n6706,n6707,n6709);
xor (n6707,n6708,n6670);
xor (n6708,n6667,n6609);
and (n6709,n6710,n6712);
xor (n6710,n6711,n6675);
xor (n6711,n6672,n6615);
and (n6712,n6713,n6715);
xor (n6713,n6714,n6680);
xor (n6714,n6677,n6632);
xor (n6715,n6716,n6685);
xor (n6716,n6682,n6638);
nor (n6717,n6718,n31);
not (n6718,n6719);
nor (n6719,n6720,n917,n6723);
and (n6720,n6721,n6722);
nor (n6721,n751,n824);
nand (n6722,n32,n677);
not (n6723,n4651);
wire s0n6724,s1n6724,notn6724;
or (n6724,s0n6724,s1n6724);
not(notn6724,n6717);
and (s0n6724,notn6724,1'b0);
and (s1n6724,n6717,n6725);
xor (n6725,n6726,n6742);
xor (n6726,n6727,n6733);
and (n6727,n6728,n6732);
xor (n6728,n6729,n6731);
not (n6729,n6730);
or (n6730,n4666,n5409);
and (n6731,n4665,n6120);
and (n6732,n4664,n6152);
and (n6733,n4664,n6734);
or (n6734,n6735,n6736,n6741);
xor (n6735,n6728,n6732);
and (n6736,n6153,n6737);
or (n6737,n6738,n6739,n6740);
and (n6738,n4663,n6591);
and (n6739,n6591,n6656);
and (n6740,n4663,n6656);
and (n6741,n6735,n6737);
and (n6742,n6743,n6746);
xor (n6743,n6744,n6734);
xor (n6744,n6745,n4664);
xor (n6745,n6728,n6727);
and (n6746,n6747,n6749);
xor (n6747,n6748,n6737);
xor (n6748,n6735,n6153);
and (n6749,n4661,n6700);
wire s0n6750,s1n6750,notn6750;
or (n6750,s0n6750,s1n6750);
not(notn6750,n6717);
and (s0n6750,notn6750,1'b0);
and (s1n6750,n6717,n6751);
xor (n6751,n6752,n6754);
xor (n6752,n6727,n6753);
and (n6753,n6728,n6733);
and (n6754,n6726,n6742);
or (n6755,n4685,n6756);
and (n6756,n32,n1069,n751,n824);
not (n6757,n6758);
or (n6758,1'b0,n6759,n6762,n6765,n6767);
and (n6759,n6760,n912);
wire s0n6760,s1n6760,notn6760;
or (n6760,s0n6760,s1n6760);
not(notn6760,n4648);
and (s0n6760,notn6760,1'b0);
and (s1n6760,n4648,n6761);
and (n6762,n6763,n917);
wire s0n6763,s1n6763,notn6763;
or (n6763,s0n6763,s1n6763);
not(notn6763,n918);
and (s0n6763,notn6763,1'b0);
and (s1n6763,n918,n6764);
and (n6765,n4657,n6766);
not (n6766,n4686);
or (n6767,1'b0,n6768,n6791,n6811,n6831);
and (n6768,n6769,n1056);
or (n6769,1'b0,n6770,n6777,n6783);
and (n6770,n6771,n6776);
or (n6771,1'b0,n6772,n6773,n6774,n6775);
and (n6772,n2306,n910);
and (n6773,n2308,n909);
and (n6774,n2310,n906);
and (n6775,n2304,n900);
nor (n6776,n32,n1069,n751,n824);
and (n6777,n6778,n6756);
or (n6778,1'b0,n6779,n6780,n6781,n6782);
and (n6779,n2267,n910);
and (n6780,n2270,n909);
and (n6781,n2262,n906);
and (n6782,n2264,n900);
and (n6783,n6784,n6789);
or (n6784,1'b0,n6785,n6786,n6787,n6788);
and (n6785,n2270,n910);
and (n6786,n2262,n909);
and (n6787,n2264,n906);
and (n6788,n2254,n900);
or (n6789,n4685,n6790);
nor (n6790,n32,n677,n751,n824);
and (n6791,n6792,n1041);
or (n6792,1'b0,n6793,n6799,n6805);
and (n6793,n6794,n6776);
or (n6794,1'b0,n6795,n6796,n6797,n6798);
and (n6795,n2321,n910);
and (n6796,n2323,n909);
and (n6797,n2325,n906);
and (n6798,n2319,n900);
and (n6799,n6800,n6756);
or (n6800,1'b0,n6801,n6802,n6803,n6804);
and (n6801,n2254,n910);
and (n6802,n2258,n909);
and (n6803,n2249,n906);
and (n6804,n2251,n900);
and (n6805,n6806,n6789);
or (n6806,1'b0,n6807,n6808,n6809,n6810);
and (n6807,n2258,n910);
and (n6808,n2249,n909);
and (n6809,n2251,n906);
and (n6810,n2256,n900);
and (n6811,n6812,n990);
or (n6812,1'b0,n6813,n6819,n6825);
and (n6813,n6814,n6776);
or (n6814,1'b0,n6815,n6816,n6817,n6818);
and (n6815,n2292,n910);
and (n6816,n2330,n909);
and (n6817,n2327,n906);
and (n6818,n2286,n900);
and (n6819,n6820,n6756);
or (n6820,1'b0,n6821,n6822,n6823,n6824);
and (n6821,n2242,n910);
and (n6822,n2244,n909);
and (n6823,n2275,n906);
and (n6824,n2280,n900);
and (n6825,n6826,n6789);
or (n6826,1'b0,n6827,n6828,n6829,n6830);
and (n6827,n2244,n910);
and (n6828,n2275,n909);
and (n6829,n2280,n906);
and (n6830,n2233,n900);
and (n6831,n6832,n970);
or (n6832,1'b0,n6833,n6839,n6845);
and (n6833,n6834,n6776);
or (n6834,1'b0,n6835,n6836,n6837,n6838);
and (n6835,n2289,n910);
and (n6836,n2312,n909);
and (n6837,n2332,n906);
and (n6838,n2294,n900);
and (n6839,n6840,n6756);
or (n6840,1'b0,n6841,n6842,n6843,n6844);
and (n6841,n2233,n910);
and (n6842,n2237,n909);
and (n6843,n2273,n906);
and (n6844,n2278,n900);
and (n6845,n6846,n6789);
or (n6846,1'b0,n6847,n6848,n6849,n6850);
and (n6847,n2237,n910);
and (n6848,n2273,n909);
and (n6849,n2278,n906);
and (n6850,n2240,n900);
nand (n6851,n6852,n6873);
not (n6852,n6853);
or (n6853,1'b0,n6854,n6865,n6867,n6868);
and (n6854,n6855,n912);
wire s0n6855,s1n6855,notn6855;
or (n6855,s0n6855,s1n6855);
not(notn6855,n4648);
and (s0n6855,notn6855,1'b0);
and (s1n6855,n4648,n6856);
wire s0n6856,s1n6856,notn6856;
or (n6856,s0n6856,s1n6856);
not(notn6856,n4628);
and (s0n6856,notn6856,n6857);
and (s1n6856,n4628,1'b0);
wire s0n6857,s1n6857,notn6857;
or (n6857,s0n6857,s1n6857);
not(notn6857,n4502);
and (s0n6857,notn6857,n6858);
and (s1n6857,n4502,1'b1);
wire s0n6858,s1n6858,notn6858;
or (n6858,s0n6858,s1n6858);
not(notn6858,n28);
and (s0n6858,notn6858,n6859);
and (s1n6858,n28,n6862);
wire s0n6859,s1n6859,notn6859;
or (n6859,s0n6859,s1n6859);
not(notn6859,n28);
and (s0n6859,notn6859,n6860);
and (s1n6859,n28,n6861);
xor (n6860,n3824,n3826);
not (n6861,n3824);
wire s0n6862,s1n6862,notn6862;
or (n6862,s0n6862,s1n6862);
not(notn6862,n28);
and (s0n6862,notn6862,n6863);
and (s1n6862,n28,n6864);
xor (n6863,n4484,n4486);
xor (n6864,n4484,n4498);
and (n6865,n6866,n917);
wire s0n6866,s1n6866,notn6866;
or (n6866,s0n6866,s1n6866);
not(notn6866,n918);
and (s0n6866,notn6866,1'b0);
and (s1n6866,n918,n6856);
and (n6867,n6856,n4655);
and (n6868,n6869,n6755);
wire s0n6869,s1n6869,notn6869;
or (n6869,s0n6869,s1n6869);
not(notn6869,n6750);
and (s0n6869,notn6869,n6870);
and (s1n6869,n6750,1'b0);
wire s0n6870,s1n6870,notn6870;
or (n6870,s0n6870,s1n6870);
not(notn6870,n6724);
and (s0n6870,notn6870,n6871);
and (s1n6870,n6724,1'b1);
wire s0n6871,s1n6871,notn6871;
or (n6871,s0n6871,s1n6871);
not(notn6871,n6717);
and (s0n6871,notn6871,1'b0);
and (s1n6871,n6717,n6872);
xor (n6872,n6701,n6703);
not (n6873,n6874);
or (n6874,1'b0,n6875,n6878,n6881,n6882);
and (n6875,n6876,n912);
wire s0n6876,s1n6876,notn6876;
or (n6876,s0n6876,s1n6876);
not(notn6876,n4648);
and (s0n6876,notn6876,1'b0);
and (s1n6876,n4648,n6877);
and (n6878,n6879,n917);
wire s0n6879,s1n6879,notn6879;
or (n6879,s0n6879,s1n6879);
not(notn6879,n918);
and (s0n6879,notn6879,1'b0);
and (s1n6879,n918,n6880);
and (n6881,n6869,n6766);
or (n6882,1'b0,n6883,n6903,n6923,n6943);
and (n6883,n6884,n1056);
or (n6884,1'b0,n6885,n6891,n6897);
and (n6885,n6886,n6776);
or (n6886,1'b0,n6887,n6888,n6889,n6890);
and (n6887,n2412,n910);
and (n6888,n2414,n909);
and (n6889,n2416,n906);
and (n6890,n2410,n900);
and (n6891,n6892,n6756);
or (n6892,1'b0,n6893,n6894,n6895,n6896);
and (n6893,n2350,n910);
and (n6894,n2355,n909);
and (n6895,n2345,n906);
and (n6896,n2343,n900);
and (n6897,n6898,n6789);
or (n6898,1'b0,n6899,n6900,n6901,n6902);
and (n6899,n2355,n910);
and (n6900,n2345,n909);
and (n6901,n2343,n906);
and (n6902,n2352,n900);
and (n6903,n6904,n1041);
or (n6904,1'b0,n6905,n6911,n6917);
and (n6905,n6906,n6776);
or (n6906,1'b0,n6907,n6908,n6909,n6910);
and (n6907,n2431,n910);
and (n6908,n2421,n909);
and (n6909,n2423,n906);
and (n6910,n2429,n900);
and (n6911,n6912,n6756);
or (n6912,1'b0,n6913,n6914,n6915,n6916);
and (n6913,n2352,n910);
and (n6914,n2371,n909);
and (n6915,n2362,n906);
and (n6916,n2360,n900);
and (n6917,n6918,n6789);
or (n6918,1'b0,n6919,n6920,n6921,n6922);
and (n6919,n2371,n910);
and (n6920,n2362,n909);
and (n6921,n2360,n906);
and (n6922,n2368,n900);
and (n6923,n6924,n990);
or (n6924,1'b0,n6925,n6931,n6937);
and (n6925,n6926,n6776);
or (n6926,1'b0,n6927,n6928,n6929,n6930);
and (n6927,n2436,n910);
and (n6928,n2440,n909);
and (n6929,n2443,n906);
and (n6930,n2446,n900);
and (n6931,n6932,n6756);
or (n6932,1'b0,n6933,n6934,n6935,n6936);
and (n6933,n2377,n910);
and (n6934,n2376,n909);
and (n6935,n2380,n906);
and (n6936,n2383,n900);
and (n6937,n6938,n6789);
or (n6938,1'b0,n6939,n6940,n6941,n6942);
and (n6939,n2376,n910);
and (n6940,n2380,n909);
and (n6941,n2383,n906);
and (n6942,n2386,n900);
and (n6943,n6944,n970);
or (n6944,1'b0,n6945,n6951,n6957);
and (n6945,n6946,n6776);
or (n6946,1'b0,n6947,n6948,n6949,n6950);
and (n6947,n2451,n910);
and (n6948,n2454,n909);
and (n6949,n2457,n906);
and (n6950,n2460,n900);
and (n6951,n6952,n6756);
or (n6952,1'b0,n6953,n6954,n6955,n6956);
and (n6953,n2386,n910);
and (n6954,n2391,n909);
and (n6955,n2394,n906);
and (n6956,n2397,n900);
and (n6957,n6958,n6789);
or (n6958,1'b0,n6959,n6960,n6961,n6962);
and (n6959,n2391,n910);
and (n6960,n2394,n909);
and (n6961,n2397,n906);
and (n6962,n2400,n900);
nand (n6963,n6964,n7476);
or (n6964,n6965,n7073);
not (n6965,n6966);
not (n6966,n6967);
and (n6967,n6968,n7061);
or (n6968,1'b0,n6969,n6972,n6975,n6980);
and (n6969,n6970,n912);
wire s0n6970,s1n6970,notn6970;
or (n6970,s0n6970,s1n6970);
not(notn6970,n4648);
and (s0n6970,notn6970,1'b0);
and (s1n6970,n4648,n6971);
and (n6972,n6973,n917);
wire s0n6973,s1n6973,notn6973;
or (n6973,s0n6973,s1n6973);
not(notn6973,n918);
and (s0n6973,notn6973,1'b0);
and (s1n6973,n918,n6974);
and (n6975,n6976,n6766);
wire s0n6976,s1n6976,notn6976;
or (n6976,s0n6976,s1n6976);
not(notn6976,n6750);
and (s0n6976,notn6976,n6977);
and (s1n6976,n6750,1'b0);
wire s0n6977,s1n6977,notn6977;
or (n6977,s0n6977,s1n6977);
not(notn6977,n6724);
and (s0n6977,notn6977,n6978);
and (s1n6977,n6724,1'b1);
wire s0n6978,s1n6978,notn6978;
or (n6978,s0n6978,s1n6978);
not(notn6978,n6717);
and (s0n6978,notn6978,1'b0);
and (s1n6978,n6717,n6979);
xor (n6979,n6704,n6706);
or (n6980,1'b0,n6981,n7001,n7021,n7041);
and (n6981,n6982,n1056);
or (n6982,1'b0,n6983,n6989,n6995);
and (n6983,n6984,n6776);
or (n6984,1'b0,n6985,n6986,n6987,n6988);
and (n6985,n2544,n910);
and (n6986,n2535,n909);
and (n6987,n2537,n906);
and (n6988,n2542,n900);
and (n6989,n6990,n6756);
or (n6990,1'b0,n6991,n6992,n6993,n6994);
and (n6991,n2478,n910);
and (n6992,n2483,n909);
and (n6993,n2471,n906);
and (n6994,n2473,n900);
and (n6995,n6996,n6789);
or (n6996,1'b0,n6997,n6998,n6999,n7000);
and (n6997,n2483,n910);
and (n6998,n2471,n909);
and (n6999,n2473,n906);
and (n7000,n2480,n900);
and (n7001,n7002,n1041);
or (n7002,1'b0,n7003,n7009,n7015);
and (n7003,n7004,n6776);
or (n7004,1'b0,n7005,n7006,n7007,n7008);
and (n7005,n2556,n910);
and (n7006,n2548,n909);
and (n7007,n2550,n906);
and (n7008,n2554,n900);
and (n7009,n7010,n6756);
or (n7010,1'b0,n7011,n7012,n7013,n7014);
and (n7011,n2480,n910);
and (n7012,n2499,n909);
and (n7013,n2488,n906);
and (n7014,n2490,n900);
and (n7015,n7016,n6789);
or (n7016,1'b0,n7017,n7018,n7019,n7020);
and (n7017,n2499,n910);
and (n7018,n2488,n909);
and (n7019,n2490,n906);
and (n7020,n2496,n900);
and (n7021,n7022,n990);
or (n7022,1'b0,n7023,n7029,n7035);
and (n7023,n7024,n6776);
or (n7024,1'b0,n7025,n7026,n7027,n7028);
and (n7025,n2561,n910);
and (n7026,n2565,n909);
and (n7027,n2568,n906);
and (n7028,n2571,n900);
and (n7029,n7030,n6756);
or (n7030,1'b0,n7031,n7032,n7033,n7034);
and (n7031,n2505,n910);
and (n7032,n2504,n909);
and (n7033,n2508,n906);
and (n7034,n2511,n900);
and (n7035,n7036,n6789);
or (n7036,1'b0,n7037,n7038,n7039,n7040);
and (n7037,n2504,n910);
and (n7038,n2508,n909);
and (n7039,n2511,n906);
and (n7040,n2514,n900);
and (n7041,n7042,n970);
or (n7042,1'b0,n7043,n7049,n7055);
and (n7043,n7044,n6776);
or (n7044,1'b0,n7045,n7046,n7047,n7048);
and (n7045,n2576,n910);
and (n7046,n2579,n909);
and (n7047,n2582,n906);
and (n7048,n2585,n900);
and (n7049,n7050,n6756);
or (n7050,1'b0,n7051,n7052,n7053,n7054);
and (n7051,n2514,n910);
and (n7052,n2519,n909);
and (n7053,n2522,n906);
and (n7054,n2525,n900);
and (n7055,n7056,n6789);
or (n7056,1'b0,n7057,n7058,n7059,n7060);
and (n7057,n2519,n910);
and (n7058,n2522,n909);
and (n7059,n2525,n906);
and (n7060,n2528,n900);
or (n7061,1'b0,n7062,n7069,n7071,n7072);
and (n7062,n7063,n912);
wire s0n7063,s1n7063,notn7063;
or (n7063,s0n7063,s1n7063);
not(notn7063,n4648);
and (s0n7063,notn7063,1'b0);
and (s1n7063,n4648,n7064);
wire s0n7064,s1n7064,notn7064;
or (n7064,s0n7064,s1n7064);
not(notn7064,n4628);
and (s0n7064,notn7064,n7065);
and (s1n7064,n4628,1'b0);
wire s0n7065,s1n7065,notn7065;
or (n7065,s0n7065,s1n7065);
not(notn7065,n4502);
and (s0n7065,notn7065,n7066);
and (s1n7065,n4502,1'b1);
wire s0n7066,s1n7066,notn7066;
or (n7066,s0n7066,s1n7066);
not(notn7066,n28);
and (s0n7066,notn7066,n7067);
and (s1n7066,n28,n4503);
wire s0n7067,s1n7067,notn7067;
or (n7067,s0n7067,s1n7067);
not(notn7067,n28);
and (s0n7067,notn7067,n7068);
and (s1n7067,n28,n3827);
xor (n7068,n3827,n3829);
and (n7069,n7070,n917);
wire s0n7070,s1n7070,notn7070;
or (n7070,s0n7070,s1n7070);
not(notn7070,n918);
and (s0n7070,notn7070,1'b0);
and (s1n7070,n918,n7064);
and (n7071,n7064,n4655);
and (n7072,n6976,n6755);
not (n7073,n7074);
nor (n7074,n7075,n7475);
and (n7075,n7076,n7185);
or (n7076,n7077,n7096);
or (n7077,1'b0,n7078,n7088,n7090,n7091);
and (n7078,n7079,n912);
wire s0n7079,s1n7079,notn7079;
or (n7079,s0n7079,s1n7079);
not(notn7079,n4648);
and (s0n7079,notn7079,1'b0);
and (s1n7079,n4648,n7080);
wire s0n7080,s1n7080,notn7080;
or (n7080,s0n7080,s1n7080);
not(notn7080,n4628);
and (s0n7080,notn7080,n7081);
and (s1n7080,n4628,1'b0);
wire s0n7081,s1n7081,notn7081;
or (n7081,s0n7081,s1n7081);
not(notn7081,n4502);
and (s0n7081,notn7081,n7082);
and (s1n7081,n4502,1'b1);
wire s0n7082,s1n7082,notn7082;
or (n7082,s0n7082,s1n7082);
not(notn7082,n28);
and (s0n7082,notn7082,n7083);
and (s1n7082,n28,n7085);
wire s0n7083,s1n7083,notn7083;
or (n7083,s0n7083,s1n7083);
not(notn7083,n28);
and (s0n7083,notn7083,n7084);
and (s1n7083,n28,n3830);
xor (n7084,n3830,n3832);
wire s0n7085,s1n7085,notn7085;
or (n7085,s0n7085,s1n7085);
not(notn7085,n28);
and (s0n7085,notn7085,n7086);
and (s1n7085,n28,n7087);
xor (n7086,n4490,n4492);
xor (n7087,n4490,n4500);
and (n7088,n7089,n917);
wire s0n7089,s1n7089,notn7089;
or (n7089,s0n7089,s1n7089);
not(notn7089,n918);
and (s0n7089,notn7089,1'b0);
and (s1n7089,n918,n7080);
and (n7090,n7080,n4655);
and (n7091,n7092,n6755);
wire s0n7092,s1n7092,notn7092;
or (n7092,s0n7092,s1n7092);
not(notn7092,n6750);
and (s0n7092,notn7092,n7093);
and (s1n7092,n6750,1'b0);
wire s0n7093,s1n7093,notn7093;
or (n7093,s0n7093,s1n7093);
not(notn7093,n6724);
and (s0n7093,notn7093,n7094);
and (s1n7093,n6724,1'b1);
wire s0n7094,s1n7094,notn7094;
or (n7094,s0n7094,s1n7094);
not(notn7094,n6717);
and (s0n7094,notn7094,1'b0);
and (s1n7094,n6717,n7095);
xor (n7095,n6707,n6709);
or (n7096,1'b0,n7097,n7100,n7103,n7104);
and (n7097,n7098,n912);
wire s0n7098,s1n7098,notn7098;
or (n7098,s0n7098,s1n7098);
not(notn7098,n4648);
and (s0n7098,notn7098,1'b0);
and (s1n7098,n4648,n7099);
and (n7100,n7101,n917);
wire s0n7101,s1n7101,notn7101;
or (n7101,s0n7101,s1n7101);
not(notn7101,n918);
and (s0n7101,notn7101,1'b0);
and (s1n7101,n918,n7102);
and (n7103,n7092,n6766);
or (n7104,1'b0,n7105,n7125,n7145,n7165);
and (n7105,n7106,n1056);
or (n7106,1'b0,n7107,n7113,n7119);
and (n7107,n7108,n6776);
or (n7108,1'b0,n7109,n7110,n7111,n7112);
and (n7109,n2657,n910);
and (n7110,n2659,n909);
and (n7111,n2661,n906);
and (n7112,n2655,n900);
and (n7113,n7114,n6756);
or (n7114,1'b0,n7115,n7116,n7117,n7118);
and (n7115,n2596,n910);
and (n7116,n2600,n909);
and (n7117,n2602,n906);
and (n7118,n2604,n900);
and (n7119,n7120,n6789);
or (n7120,1'b0,n7121,n7122,n7123,n7124);
and (n7121,n2600,n910);
and (n7122,n2602,n909);
and (n7123,n2604,n906);
and (n7124,n2598,n900);
and (n7125,n7126,n1041);
or (n7126,1'b0,n7127,n7133,n7139);
and (n7127,n7128,n6776);
or (n7128,1'b0,n7129,n7130,n7131,n7132);
and (n7129,n2669,n910);
and (n7130,n2671,n909);
and (n7131,n2673,n906);
and (n7132,n2666,n900);
and (n7133,n7134,n6756);
or (n7134,1'b0,n7135,n7136,n7137,n7138);
and (n7135,n2598,n910);
and (n7136,n2612,n909);
and (n7137,n2614,n906);
and (n7138,n2616,n900);
and (n7139,n7140,n6789);
or (n7140,1'b0,n7141,n7142,n7143,n7144);
and (n7141,n2612,n910);
and (n7142,n2614,n909);
and (n7143,n2616,n906);
and (n7144,n2610,n900);
and (n7145,n7146,n990);
or (n7146,1'b0,n7147,n7153,n7159);
and (n7147,n7148,n6776);
or (n7148,1'b0,n7149,n7150,n7151,n7152);
and (n7149,n2678,n910);
and (n7150,n2682,n909);
and (n7151,n2685,n906);
and (n7152,n2688,n900);
and (n7153,n7154,n6756);
or (n7154,1'b0,n7155,n7156,n7157,n7158);
and (n7155,n2622,n910);
and (n7156,n2621,n909);
and (n7157,n2625,n906);
and (n7158,n2628,n900);
and (n7159,n7160,n6789);
or (n7160,1'b0,n7161,n7162,n7163,n7164);
and (n7161,n2621,n910);
and (n7162,n2625,n909);
and (n7163,n2628,n906);
and (n7164,n2631,n900);
and (n7165,n7166,n970);
or (n7166,1'b0,n7167,n7173,n7179);
and (n7167,n7168,n6776);
or (n7168,1'b0,n7169,n7170,n7171,n7172);
and (n7169,n2693,n910);
and (n7170,n2696,n909);
and (n7171,n2699,n906);
and (n7172,n2702,n900);
and (n7173,n7174,n6756);
or (n7174,1'b0,n7175,n7176,n7177,n7178);
and (n7175,n2631,n910);
and (n7176,n2636,n909);
and (n7177,n2639,n906);
and (n7178,n2642,n900);
and (n7179,n7180,n6789);
or (n7180,1'b0,n7181,n7182,n7183,n7184);
and (n7181,n2636,n910);
and (n7182,n2639,n909);
and (n7183,n2642,n906);
and (n7184,n2645,n900);
nand (n7185,n7186,n7467);
or (n7186,n7187,n7361);
not (n7187,n7188);
nand (n7188,n7189,n7203);
or (n7189,n7190,n7197);
not (n7190,n7191);
nand (n7191,n7192,n7193,n7194);
or (n7192,n953,n6723);
not (n7193,n916);
not (n7194,n7195);
and (n7195,n912,n7196,n4649);
and (n7196,n676,n4651);
not (n7197,n7198);
wire s0n7198,s1n7198,notn7198;
or (n7198,s0n7198,s1n7198);
not(notn7198,n4628);
and (s0n7198,notn7198,n7199);
and (s1n7198,n4628,1'b0);
wire s0n7199,s1n7199,notn7199;
or (n7199,s0n7199,s1n7199);
not(notn7199,n4502);
and (s0n7199,notn7199,n7200);
and (s1n7199,n4502,1'b1);
wire s0n7200,s1n7200,notn7200;
or (n7200,s0n7200,s1n7200);
not(notn7200,n28);
and (s0n7200,notn7200,n7201);
and (s1n7200,n28,n18);
wire s0n7201,s1n7201,notn7201;
or (n7201,s0n7201,s1n7201);
not(notn7201,n28);
and (s0n7201,notn7201,n7202);
and (s1n7201,n28,n3836);
xor (n7202,n3836,n3838);
nor (n7203,n7204,n7271);
and (n7204,n7205,n7263);
wire s0n7205,s1n7205,notn7205;
or (n7205,s0n7205,s1n7205);
not(notn7205,n6750);
and (s0n7205,notn7205,n7206);
and (s1n7205,n6750,1'b0);
wire s0n7206,s1n7206,notn7206;
or (n7206,s0n7206,s1n7206);
not(notn7206,n6724);
and (s0n7206,notn7206,n7207);
and (s1n7206,n6724,1'b1);
wire s0n7207,s1n7207,notn7207;
or (n7207,s0n7207,s1n7207);
not(notn7207,n6717);
and (s0n7207,notn7207,1'b0);
and (s1n7207,n6717,n7208);
xor (n7208,n7209,n7232);
xor (n7209,n7210,n7215);
xor (n7210,n7211,n6609);
xor (n7211,n7212,n7214);
or (n7212,n7213,n6316);
and (n7213,n6614,n6638);
xor (n7214,n6608,n6632);
nand (n7215,n7216,n7231);
or (n7216,n7217,n7223);
or (n7217,n7218,n7222);
and (n7218,n7219,n6632);
xor (n7219,n7220,n7221);
and (n7220,n6447,n6151);
xor (n7221,n6631,n6644);
and (n7222,n7220,n7221);
not (n7223,n7224);
or (n7224,n7225,n7230);
and (n7225,n7226,n6615);
xor (n7226,n7227,n7229);
or (n7227,n7228,n6366);
and (n7228,n6631,n6644);
xor (n7229,n6614,n6638);
and (n7230,n7227,n7229);
nand (n7231,n7223,n7217);
or (n7232,n7233,n7262);
and (n7233,n7234,n7237);
xor (n7234,n7235,n7236);
xor (n7235,n7226,n6615);
not (n7236,n7217);
or (n7237,n7238,n7261);
and (n7238,n7239,n7246);
xor (n7239,n7240,n7245);
or (n7240,n7241,n7244);
and (n7241,n7242,n6638);
xor (n7242,n6423,n7243);
xor (n7243,n6447,n6151);
and (n7244,n6423,n7243);
xor (n7245,n7219,n6632);
or (n7246,n7247,n7260);
and (n7247,n7248,n7252);
xor (n7248,n7249,n7251);
or (n7249,n7250,n6472);
and (n7250,n6643,n6644);
xor (n7251,n7242,n6638);
or (n7252,n7253,n7259);
and (n7253,n7254,n7257);
xor (n7254,n7255,n7256);
and (n7255,n6559,n6151);
xor (n7256,n6643,n6644);
and (n7257,n7258,n6527);
xor (n7258,n6559,n6151);
and (n7259,n7255,n7256);
and (n7260,n7249,n7251);
and (n7261,n7240,n7245);
and (n7262,n7235,n7236);
nand (n7263,n7264,n7266);
not (n7264,n7265);
and (n7265,n6766,n4651);
not (n7266,n7267);
and (n7267,n7268,n7269,n4651);
and (n7268,n1069,n751);
nor (n7269,n7270,n33);
not (n7270,n676);
nand (n7271,n7272,n7354);
not (n7272,n7273);
or (n7273,1'b0,n7274,n7294,n7314,n7334);
and (n7274,n7275,n1056);
or (n7275,1'b0,n7276,n7282,n7288);
and (n7276,n7277,n6776);
or (n7277,1'b0,n7278,n7279,n7280,n7281);
and (n7278,n2901,n910);
and (n7279,n2896,n909);
and (n7280,n2898,n906);
and (n7281,n2907,n900);
and (n7282,n7283,n6756);
or (n7283,1'b0,n7284,n7285,n7286,n7287);
and (n7284,n2842,n910);
and (n7285,n2844,n909);
and (n7286,n2839,n906);
and (n7287,n2837,n900);
and (n7288,n7289,n6789);
or (n7289,1'b0,n7290,n7291,n7292,n7293);
and (n7290,n2844,n910);
and (n7291,n2839,n909);
and (n7292,n2837,n906);
and (n7293,n2846,n900);
and (n7294,n7295,n1041);
or (n7295,1'b0,n7296,n7302,n7308);
and (n7296,n7297,n6776);
or (n7297,1'b0,n7298,n7299,n7300,n7301);
and (n7298,n2917,n910);
and (n7299,n2912,n909);
and (n7300,n2914,n906);
and (n7301,n2922,n900);
and (n7302,n7303,n6756);
or (n7303,1'b0,n7304,n7305,n7306,n7307);
and (n7304,n2846,n910);
and (n7305,n2857,n909);
and (n7306,n2851,n906);
and (n7307,n2853,n900);
and (n7308,n7309,n6789);
or (n7309,1'b0,n7310,n7311,n7312,n7313);
and (n7310,n2857,n910);
and (n7311,n2851,n909);
and (n7312,n2853,n906);
and (n7313,n2859,n900);
and (n7314,n7315,n990);
or (n7315,1'b0,n7316,n7322,n7328);
and (n7316,n7317,n6776);
or (n7317,1'b0,n7318,n7319,n7320,n7321);
and (n7318,n2927,n910);
and (n7319,n2931,n909);
and (n7320,n2934,n906);
and (n7321,n2937,n900);
and (n7322,n7323,n6756);
or (n7323,1'b0,n7324,n7325,n7326,n7327);
and (n7324,n2865,n910);
and (n7325,n2864,n909);
and (n7326,n2868,n906);
and (n7327,n2871,n900);
and (n7328,n7329,n6789);
or (n7329,1'b0,n7330,n7331,n7332,n7333);
and (n7330,n2864,n910);
and (n7331,n2868,n909);
and (n7332,n2871,n906);
and (n7333,n2874,n900);
and (n7334,n7335,n970);
or (n7335,1'b0,n7336,n7342,n7348);
and (n7336,n7337,n6776);
or (n7337,1'b0,n7338,n7339,n7340,n7341);
and (n7338,n2942,n910);
and (n7339,n2945,n909);
and (n7340,n2948,n906);
and (n7341,n2951,n900);
and (n7342,n7343,n6756);
or (n7343,1'b0,n7344,n7345,n7346,n7347);
and (n7344,n2874,n910);
and (n7345,n2879,n909);
and (n7346,n2882,n906);
and (n7347,n2885,n900);
and (n7348,n7349,n6789);
or (n7349,1'b0,n7350,n7351,n7352,n7353);
and (n7350,n2879,n910);
and (n7351,n2882,n909);
and (n7352,n2885,n906);
and (n7353,n2888,n900);
nor (n7354,n7355,n7358);
and (n7355,n7356,n912);
wire s0n7356,s1n7356,notn7356;
or (n7356,s0n7356,s1n7356);
not(notn7356,n4648);
and (s0n7356,notn7356,1'b0);
and (s1n7356,n4648,n7357);
and (n7358,n7359,n917);
wire s0n7359,s1n7359,notn7359;
or (n7359,s0n7359,s1n7359);
not(notn7359,n918);
and (s0n7359,notn7359,1'b0);
and (s1n7359,n918,n7360);
not (n7361,n7362);
nand (n7362,n7363,n7372);
nand (n7363,n7364,n7191);
wire s0n7364,s1n7364,notn7364;
or (n7364,s0n7364,s1n7364);
not(notn7364,n4628);
and (s0n7364,notn7364,n7365);
and (s1n7364,n4628,1'b0);
wire s0n7365,s1n7365,notn7365;
or (n7365,s0n7365,s1n7365);
not(notn7365,n4502);
and (s0n7365,notn7365,n7366);
and (s1n7365,n4502,1'b1);
wire s0n7366,s1n7366,notn7366;
or (n7366,s0n7366,s1n7366);
not(notn7366,n28);
and (s0n7366,notn7366,n7367);
and (s1n7366,n28,n7369);
wire s0n7367,s1n7367,notn7367;
or (n7367,s0n7367,s1n7367);
not(notn7367,n28);
and (s0n7367,notn7367,n7368);
and (s1n7367,n28,n3833);
xor (n7368,n3833,n3835);
wire s0n7369,s1n7369,notn7369;
or (n7369,s0n7369,s1n7369);
not(notn7369,n28);
and (s0n7369,notn7369,n7370);
and (s1n7369,n28,n7371);
xor (n7370,n4493,n4495);
xor (n7371,n4493,n4501);
nor (n7372,n7373,n7466);
or (n7373,1'b0,n7374,n7377,n7380,n7385);
and (n7374,n7375,n912);
wire s0n7375,s1n7375,notn7375;
or (n7375,s0n7375,s1n7375);
not(notn7375,n4648);
and (s0n7375,notn7375,1'b0);
and (s1n7375,n4648,n7376);
and (n7377,n7378,n917);
wire s0n7378,s1n7378,notn7378;
or (n7378,s0n7378,s1n7378);
not(notn7378,n918);
and (s0n7378,notn7378,1'b0);
and (s1n7378,n918,n7379);
and (n7380,n7381,n6766);
wire s0n7381,s1n7381,notn7381;
or (n7381,s0n7381,s1n7381);
not(notn7381,n6750);
and (s0n7381,notn7381,n7382);
and (s1n7381,n6750,1'b0);
wire s0n7382,s1n7382,notn7382;
or (n7382,s0n7382,s1n7382);
not(notn7382,n6724);
and (s0n7382,notn7382,n7383);
and (s1n7382,n6724,1'b1);
wire s0n7383,s1n7383,notn7383;
or (n7383,s0n7383,s1n7383);
not(notn7383,n6717);
and (s0n7383,notn7383,1'b0);
and (s1n7383,n6717,n7384);
xor (n7384,n6710,n6712);
or (n7385,1'b0,n7386,n7406,n7426,n7446);
and (n7386,n7387,n1056);
or (n7387,1'b0,n7388,n7394,n7400);
and (n7388,n7389,n6776);
or (n7389,1'b0,n7390,n7391,n7392,n7393);
and (n7390,n2780,n910);
and (n7391,n2782,n909);
and (n7392,n2784,n906);
and (n7393,n2778,n900);
and (n7394,n7395,n6756);
or (n7395,1'b0,n7396,n7397,n7398,n7399);
and (n7396,n2714,n910);
and (n7397,n2713,n909);
and (n7398,n2717,n906);
and (n7399,n2720,n900);
and (n7400,n7401,n6789);
or (n7401,1'b0,n7402,n7403,n7404,n7405);
and (n7402,n2713,n910);
and (n7403,n2717,n909);
and (n7404,n2720,n906);
and (n7405,n2723,n900);
and (n7406,n7407,n1041);
or (n7407,1'b0,n7408,n7414,n7420);
and (n7408,n7409,n6776);
or (n7409,1'b0,n7410,n7411,n7412,n7413);
and (n7410,n2793,n910);
and (n7411,n2795,n909);
and (n7412,n2797,n906);
and (n7413,n2791,n900);
and (n7414,n7415,n6756);
or (n7415,1'b0,n7416,n7417,n7418,n7419);
and (n7416,n2723,n910);
and (n7417,n2734,n909);
and (n7418,n2730,n906);
and (n7419,n2728,n900);
and (n7420,n7421,n6789);
or (n7421,1'b0,n7422,n7423,n7424,n7425);
and (n7422,n2734,n910);
and (n7423,n2730,n909);
and (n7424,n2728,n906);
and (n7425,n2736,n900);
and (n7426,n7427,n990);
or (n7427,1'b0,n7428,n7434,n7440);
and (n7428,n7429,n6776);
or (n7429,1'b0,n7430,n7431,n7432,n7433);
and (n7430,n2802,n910);
and (n7431,n2806,n909);
and (n7432,n2809,n906);
and (n7433,n2812,n900);
and (n7434,n7435,n6756);
or (n7435,1'b0,n7436,n7437,n7438,n7439);
and (n7436,n2742,n910);
and (n7437,n2741,n909);
and (n7438,n2745,n906);
and (n7439,n2748,n900);
and (n7440,n7441,n6789);
or (n7441,1'b0,n7442,n7443,n7444,n7445);
and (n7442,n2741,n910);
and (n7443,n2745,n909);
and (n7444,n2748,n906);
and (n7445,n2751,n900);
and (n7446,n7447,n970);
or (n7447,1'b0,n7448,n7454,n7460);
and (n7448,n7449,n6776);
or (n7449,1'b0,n7450,n7451,n7452,n7453);
and (n7450,n2817,n910);
and (n7451,n2820,n909);
and (n7452,n2823,n906);
and (n7453,n2826,n900);
and (n7454,n7455,n6756);
or (n7455,1'b0,n7456,n7457,n7458,n7459);
and (n7456,n2751,n910);
and (n7457,n2756,n909);
and (n7458,n2759,n906);
and (n7459,n2762,n900);
and (n7460,n7461,n6789);
or (n7461,1'b0,n7462,n7463,n7464,n7465);
and (n7462,n2756,n910);
and (n7463,n2759,n909);
and (n7464,n2762,n906);
and (n7465,n2765,n900);
and (n7466,n7381,n6755);
not (n7467,n7468);
and (n7468,n7373,n7469);
or (n7469,1'b0,n7470,n7472,n7474,n7466);
and (n7470,n7471,n912);
wire s0n7471,s1n7471,notn7471;
or (n7471,s0n7471,s1n7471);
not(notn7471,n4648);
and (s0n7471,notn7471,1'b0);
and (s1n7471,n4648,n7364);
and (n7472,n7473,n917);
wire s0n7473,s1n7473,notn7473;
or (n7473,s0n7473,s1n7473);
not(notn7473,n918);
and (s0n7473,notn7473,1'b0);
and (s1n7473,n918,n7364);
and (n7474,n7364,n4655);
and (n7475,n7096,n7077);
or (n7476,n7061,n6968);
not (n7477,n7478);
nand (n7478,n7479,n7483);
or (n7479,n7480,n7481);
not (n7480,n9);
not (n7481,n7482);
and (n7482,n6874,n6853);
not (n7483,n7484);
and (n7484,n6758,n11);
nor (n7485,n7486,n7596);
not (n7486,n7487);
nand (n7487,n7488,n7506);
not (n7488,n7489);
or (n7489,1'b0,n7490,n7498,n7500,n7501);
and (n7490,n7491,n912);
wire s0n7491,s1n7491,notn7491;
or (n7491,s0n7491,s1n7491);
not(notn7491,n4648);
and (s0n7491,notn7491,1'b0);
and (s1n7491,n4648,n7492);
wire s0n7492,s1n7492,notn7492;
or (n7492,s0n7492,s1n7492);
not(notn7492,n4628);
and (s0n7492,notn7492,n7493);
and (s1n7492,n4628,1'b0);
wire s0n7493,s1n7493,notn7493;
or (n7493,s0n7493,s1n7493);
not(notn7493,n4502);
and (s0n7493,notn7493,n7494);
and (s1n7493,n4502,1'b1);
wire s0n7494,s1n7494,notn7494;
or (n7494,s0n7494,s1n7494);
not(notn7494,n28);
and (s0n7494,notn7494,n7369);
and (s1n7494,n28,n7495);
wire s0n7495,s1n7495,notn7495;
or (n7495,s0n7495,s1n7495);
not(notn7495,n28);
and (s0n7495,notn7495,n7496);
and (s1n7495,n28,n7497);
xor (n7496,n4621,n4623);
xor (n7497,n4621,n4627);
and (n7498,n7499,n917);
wire s0n7499,s1n7499,notn7499;
or (n7499,s0n7499,s1n7499);
not(notn7499,n918);
and (s0n7499,notn7499,1'b0);
and (s1n7499,n918,n7492);
and (n7500,n7492,n4655);
and (n7501,n7502,n6755);
wire s0n7502,s1n7502,notn7502;
or (n7502,s0n7502,s1n7502);
not(notn7502,n6750);
and (s0n7502,notn7502,n7503);
and (s1n7502,n6750,1'b0);
wire s0n7503,s1n7503,notn7503;
or (n7503,s0n7503,s1n7503);
not(notn7503,n6724);
and (s0n7503,notn7503,n7504);
and (s1n7503,n6724,1'b1);
wire s0n7504,s1n7504,notn7504;
or (n7504,s0n7504,s1n7504);
not(notn7504,n6717);
and (s0n7504,notn7504,1'b0);
and (s1n7504,n6717,n7505);
xor (n7505,n6747,n6749);
not (n7506,n7507);
or (n7507,1'b0,n7508,n7511,n7514,n7515);
and (n7508,n7509,n912);
wire s0n7509,s1n7509,notn7509;
or (n7509,s0n7509,s1n7509);
not(notn7509,n4648);
and (s0n7509,notn7509,1'b0);
and (s1n7509,n4648,n7510);
and (n7511,n7512,n917);
wire s0n7512,s1n7512,notn7512;
or (n7512,s0n7512,s1n7512);
not(notn7512,n918);
and (s0n7512,notn7512,1'b0);
and (s1n7512,n918,n7513);
and (n7514,n7502,n6766);
or (n7515,1'b0,n7516,n7536,n7556,n7576);
and (n7516,n7517,n1056);
or (n7517,1'b0,n7518,n7524,n7530);
and (n7518,n7519,n6776);
or (n7519,1'b0,n7520,n7521,n7522,n7523);
and (n7520,n2179,n910);
and (n7521,n2167,n909);
and (n7522,n2169,n906);
and (n7523,n2176,n900);
and (n7524,n7525,n6756);
or (n7525,1'b0,n7526,n7527,n7528,n7529);
and (n7526,n2129,n910);
and (n7527,n2132,n909);
and (n7528,n2134,n906);
and (n7529,n2136,n900);
and (n7530,n7531,n6789);
or (n7531,1'b0,n7532,n7533,n7534,n7535);
and (n7532,n2132,n910);
and (n7533,n2134,n909);
and (n7534,n2136,n906);
and (n7535,n2116,n900);
and (n7536,n7537,n1041);
or (n7537,1'b0,n7538,n7544,n7550);
and (n7538,n7539,n6776);
or (n7539,1'b0,n7540,n7541,n7542,n7543);
and (n7540,n2195,n910);
and (n7541,n2184,n909);
and (n7542,n2186,n906);
and (n7543,n2192,n900);
and (n7544,n7545,n6756);
or (n7545,1'b0,n7546,n7547,n7548,n7549);
and (n7546,n2116,n910);
and (n7547,n2120,n909);
and (n7548,n2122,n906);
and (n7549,n2124,n900);
and (n7550,n7551,n6789);
or (n7551,1'b0,n7552,n7553,n7554,n7555);
and (n7552,n2120,n910);
and (n7553,n2122,n909);
and (n7554,n2124,n906);
and (n7555,n2118,n900);
and (n7556,n7557,n990);
or (n7557,1'b0,n7558,n7564,n7570);
and (n7558,n7559,n6776);
or (n7559,1'b0,n7560,n7561,n7562,n7563);
and (n7560,n2200,n910);
and (n7561,n2204,n909);
and (n7562,n2207,n906);
and (n7563,n2210,n900);
and (n7564,n7565,n6756);
or (n7565,1'b0,n7566,n7567,n7568,n7569);
and (n7566,n2147,n910);
and (n7567,n2149,n909);
and (n7568,n2154,n906);
and (n7569,n2159,n900);
and (n7570,n7571,n6789);
or (n7571,1'b0,n7572,n7573,n7574,n7575);
and (n7572,n2149,n910);
and (n7573,n2154,n909);
and (n7574,n2159,n906);
and (n7575,n2139,n900);
and (n7576,n7577,n970);
or (n7577,1'b0,n7578,n7584,n7590);
and (n7578,n7579,n6776);
or (n7579,1'b0,n7580,n7581,n7582,n7583);
and (n7580,n2215,n910);
and (n7581,n2218,n909);
and (n7582,n2221,n906);
and (n7583,n2224,n900);
and (n7584,n7585,n6756);
or (n7585,1'b0,n7586,n7587,n7588,n7589);
and (n7586,n2139,n910);
and (n7587,n2145,n909);
and (n7588,n2152,n906);
and (n7589,n2157,n900);
and (n7590,n7591,n6789);
or (n7591,1'b0,n7592,n7593,n7594,n7595);
and (n7592,n2145,n910);
and (n7593,n2152,n909);
and (n7594,n2157,n906);
and (n7595,n2143,n900);
and (n7596,n7597,n7615);
not (n7597,n7598);
or (n7598,1'b0,n7599,n7607,n7609,n7610);
and (n7599,n7600,n912);
wire s0n7600,s1n7600,notn7600;
or (n7600,s0n7600,s1n7600);
not(notn7600,n4648);
and (s0n7600,notn7600,1'b0);
and (s1n7600,n4648,n7601);
wire s0n7601,s1n7601,notn7601;
or (n7601,s0n7601,s1n7601);
not(notn7601,n4628);
and (s0n7601,notn7601,n7602);
and (s1n7601,n4628,1'b0);
wire s0n7602,s1n7602,notn7602;
or (n7602,s0n7602,s1n7602);
not(notn7602,n4502);
and (s0n7602,notn7602,n7603);
and (s1n7602,n4502,1'b1);
wire s0n7603,s1n7603,notn7603;
or (n7603,s0n7603,s1n7603);
not(notn7603,n28);
and (s0n7603,notn7603,n7085);
and (s1n7603,n28,n7604);
wire s0n7604,s1n7604,notn7604;
or (n7604,s0n7604,s1n7604);
not(notn7604,n28);
and (s0n7604,notn7604,n7605);
and (s1n7604,n28,n7606);
xor (n7605,n4615,n4620);
xor (n7606,n4615,n4626);
and (n7607,n7608,n917);
wire s0n7608,s1n7608,notn7608;
or (n7608,s0n7608,s1n7608);
not(notn7608,n918);
and (s0n7608,notn7608,1'b0);
and (s1n7608,n918,n7601);
and (n7609,n7601,n4655);
and (n7610,n7611,n6755);
wire s0n7611,s1n7611,notn7611;
or (n7611,s0n7611,s1n7611);
not(notn7611,n6750);
and (s0n7611,notn7611,n7612);
and (s1n7611,n6750,1'b0);
wire s0n7612,s1n7612,notn7612;
or (n7612,s0n7612,s1n7612);
not(notn7612,n6724);
and (s0n7612,notn7612,n7613);
and (s1n7612,n6724,1'b1);
wire s0n7613,s1n7613,notn7613;
or (n7613,s0n7613,s1n7613);
not(notn7613,n6717);
and (s0n7613,notn7613,1'b0);
and (s1n7613,n6717,n7614);
xor (n7614,n6743,n6746);
not (n7615,n7616);
or (n7616,1'b0,n7617,n7620,n7623,n7624);
and (n7617,n7618,n912);
wire s0n7618,s1n7618,notn7618;
or (n7618,s0n7618,s1n7618);
not(notn7618,n4648);
and (s0n7618,notn7618,1'b0);
and (s1n7618,n4648,n7619);
and (n7620,n7621,n917);
wire s0n7621,s1n7621,notn7621;
or (n7621,s0n7621,s1n7621);
not(notn7621,n918);
and (s0n7621,notn7621,1'b0);
and (s1n7621,n918,n7622);
and (n7623,n7611,n6766);
or (n7624,1'b0,n7625,n7645,n7665,n7685);
and (n7625,n7626,n1056);
or (n7626,1'b0,n7627,n7633,n7639);
and (n7627,n7628,n6776);
or (n7628,1'b0,n7629,n7630,n7631,n7632);
and (n7629,n2090,n910);
and (n7630,n2092,n909);
and (n7631,n2094,n906);
and (n7632,n2074,n900);
and (n7633,n7634,n6756);
or (n7634,1'b0,n7635,n7636,n7637,n7638);
and (n7635,n2023,n910);
and (n7636,n2026,n909);
and (n7637,n2028,n906);
and (n7638,n2030,n900);
and (n7639,n7640,n6789);
or (n7640,1'b0,n7641,n7642,n7643,n7644);
and (n7641,n2026,n910);
and (n7642,n2028,n909);
and (n7643,n2030,n906);
and (n7644,n2010,n900);
and (n7645,n7646,n1041);
or (n7646,1'b0,n7647,n7653,n7659);
and (n7647,n7648,n6776);
or (n7648,1'b0,n7649,n7650,n7651,n7652);
and (n7649,n2078,n910);
and (n7650,n2080,n909);
and (n7651,n2082,n906);
and (n7652,n2076,n900);
and (n7653,n7654,n6756);
or (n7654,1'b0,n7655,n7656,n7657,n7658);
and (n7655,n2010,n910);
and (n7656,n2014,n909);
and (n7657,n2016,n906);
and (n7658,n2018,n900);
and (n7659,n7660,n6789);
or (n7660,1'b0,n7661,n7662,n7663,n7664);
and (n7661,n2014,n910);
and (n7662,n2016,n909);
and (n7663,n2018,n906);
and (n7664,n2012,n900);
and (n7665,n7666,n990);
or (n7666,1'b0,n7667,n7673,n7679);
and (n7667,n7668,n6776);
or (n7668,1'b0,n7669,n7670,n7671,n7672);
and (n7669,n2064,n910);
and (n7670,n2099,n909);
and (n7671,n2104,n906);
and (n7672,n2068,n900);
and (n7673,n7674,n6756);
or (n7674,1'b0,n7675,n7676,n7677,n7678);
and (n7675,n2040,n910);
and (n7676,n2036,n909);
and (n7677,n2045,n906);
and (n7678,n2047,n900);
and (n7679,n7680,n6789);
or (n7680,1'b0,n7681,n7682,n7683,n7684);
and (n7681,n2036,n910);
and (n7682,n2045,n909);
and (n7683,n2047,n906);
and (n7684,n2033,n900);
and (n7685,n7686,n970);
or (n7686,1'b0,n7687,n7693,n7699);
and (n7687,n7688,n6776);
or (n7688,1'b0,n7689,n7690,n7691,n7692);
and (n7689,n2060,n910);
and (n7690,n2097,n909);
and (n7691,n2102,n906);
and (n7692,n2062,n900);
and (n7693,n7694,n6756);
or (n7694,1'b0,n7695,n7696,n7697,n7698);
and (n7695,n2033,n910);
and (n7696,n2038,n909);
and (n7697,n2050,n906);
and (n7698,n2052,n900);
and (n7699,n7700,n6789);
or (n7700,1'b0,n7701,n7702,n7703,n7704);
and (n7701,n2038,n910);
and (n7702,n2050,n909);
and (n7703,n2052,n906);
and (n7704,n2042,n900);
nand (n7705,n7706,n7709);
or (n7706,n7596,n7707);
not (n7707,n7708);
and (n7708,n7507,n7489);
not (n7709,n7710);
and (n7710,n7616,n7598);
and (n7711,n7193,n7712);
nand (n7712,n7713,n897);
or (n7713,n7268,n33);
nor (n7714,n7715,n7722);
and (n7715,n7601,n7716);
and (n7716,n7717,n7196);
nand (n7717,n7718,n7720);
or (n7718,n4650,n7719);
not (n7719,n31);
not (n7720,n7721);
nor (n7721,n33,n1069,n751,n824);
and (n7722,n7611,n7723);
nor (n7723,n33,n677,n751,n914);
nor (n7724,n7725,n7841);
wire s0n7725,s1n7725,notn7725;
or (n7725,s0n7725,s1n7725);
not(notn7725,n7838);
and (s0n7725,notn7725,n7726);
and (s1n7725,n7838,n7833);
wire s0n7726,s1n7726,notn7726;
or (n7726,s0n7726,s1n7726);
not(notn7726,n7735);
and (s0n7726,notn7726,1'b0);
and (s1n7726,n7735,n7727);
wire s0n7727,s1n7727,notn7727;
or (n7727,s0n7727,s1n7727);
not(notn7727,n56);
and (s0n7727,notn7727,n7728);
and (s1n7727,n56,n7734);
or (n7728,1'b0,n7729,n7730,n7731,n7732);
and (n7729,n2042,n910);
and (n7730,n6207,n909);
and (n7731,n987,n906);
and (n7732,n7733,n900);
wire s0n7734,s1n7734,notn7734;
or (n7734,s0n7734,s1n7734);
not(notn7734,n4651);
and (s0n7734,notn7734,1'b0);
and (s1n7734,n4651,n7733);
and (n7735,n7736,n7785);
and (n7736,n626,n7737);
nor (n7737,n753,n826,n7738);
wire s0n7738,s1n7738,notn7738;
or (n7738,s0n7738,s1n7738);
not(notn7738,n626);
and (s0n7738,notn7738,1'b0);
and (s1n7738,n626,n7739);
wire s0n7739,s1n7739,notn7739;
or (n7739,s0n7739,s1n7739);
not(notn7739,n625);
and (s0n7739,notn7739,n7740);
and (s1n7739,n625,n7776);
or (n7740,n7741,n7752,n7763,n7774);
and (n7741,n7742,n62);
wire s0n7742,s1n7742,notn7742;
or (n7742,s0n7742,s1n7742);
not(notn7742,n56);
and (s0n7742,notn7742,n7743);
and (s1n7742,n56,n7744);
or (n7744,n7745,n7747,n7749,n7751);
and (n7745,n7746,n44);
and (n7747,n7748,n49);
and (n7749,n7750,n53);
and (n7751,n7743,n55);
and (n7752,n7753,n67);
wire s0n7753,s1n7753,notn7753;
or (n7753,s0n7753,s1n7753);
not(notn7753,n56);
and (s0n7753,notn7753,n7754);
and (s1n7753,n56,n7755);
or (n7755,n7756,n7758,n7760,n7762);
and (n7756,n7757,n44);
and (n7758,n7759,n49);
and (n7760,n7761,n53);
and (n7762,n7754,n55);
and (n7763,n7764,n72);
wire s0n7764,s1n7764,notn7764;
or (n7764,s0n7764,s1n7764);
not(notn7764,n56);
and (s0n7764,notn7764,n7765);
and (s1n7764,n56,n7766);
or (n7766,n7767,n7769,n7771,n7773);
and (n7767,n7768,n44);
and (n7769,n7770,n49);
and (n7771,n7772,n53);
and (n7773,n7765,n55);
and (n7774,n7775,n75);
wire s0n7775,s1n7775,notn7775;
or (n7775,s0n7775,s1n7775);
not(notn7775,n56);
and (s0n7775,notn7775,n7776);
and (s1n7775,n56,n7777);
or (n7777,n7778,n7780,n7782,n7784);
and (n7778,n7779,n44);
and (n7780,n7781,n49);
and (n7782,n7783,n53);
and (n7784,n7776,n55);
nor (n7785,n35,n679,n7786);
wire s0n7786,s1n7786,notn7786;
or (n7786,s0n7786,s1n7786);
not(notn7786,n626);
and (s0n7786,notn7786,1'b0);
and (s1n7786,n626,n7787);
wire s0n7787,s1n7787,notn7787;
or (n7787,s0n7787,s1n7787);
not(notn7787,n625);
and (s0n7787,notn7787,n7788);
and (s1n7787,n625,n7824);
or (n7788,n7789,n7800,n7811,n7822);
and (n7789,n7790,n62);
wire s0n7790,s1n7790,notn7790;
or (n7790,s0n7790,s1n7790);
not(notn7790,n56);
and (s0n7790,notn7790,n7791);
and (s1n7790,n56,n7792);
or (n7792,n7793,n7795,n7797,n7799);
and (n7793,n7794,n44);
and (n7795,n7796,n49);
and (n7797,n7798,n53);
and (n7799,n7791,n55);
and (n7800,n7801,n67);
wire s0n7801,s1n7801,notn7801;
or (n7801,s0n7801,s1n7801);
not(notn7801,n56);
and (s0n7801,notn7801,n7802);
and (s1n7801,n56,n7803);
or (n7803,n7804,n7806,n7808,n7810);
and (n7804,n7805,n44);
and (n7806,n7807,n49);
and (n7808,n7809,n53);
and (n7810,n7802,n55);
and (n7811,n7812,n72);
wire s0n7812,s1n7812,notn7812;
or (n7812,s0n7812,s1n7812);
not(notn7812,n56);
and (s0n7812,notn7812,n7813);
and (s1n7812,n56,n7814);
or (n7814,n7815,n7817,n7819,n7821);
and (n7815,n7816,n44);
and (n7817,n7818,n49);
and (n7819,n7820,n53);
and (n7821,n7813,n55);
and (n7822,n7823,n75);
wire s0n7823,s1n7823,notn7823;
or (n7823,s0n7823,s1n7823);
not(notn7823,n56);
and (s0n7823,notn7823,n7824);
and (s1n7823,n56,n7825);
or (n7825,n7826,n7828,n7830,n7832);
and (n7826,n7827,n44);
and (n7828,n7829,n49);
and (n7830,n7831,n53);
and (n7832,n7824,n55);
or (n7833,1'b0,n7834,n7835,n7836,n7837);
and (n7834,n7640,n1056);
and (n7835,n7660,n1041);
and (n7836,n7680,n990);
and (n7837,n7700,n970);
and (n7838,n676,n7839);
not (n7839,n7840);
or (n7840,n33,n677,n751,n824);
and (n7841,n7842,n9704);
nand (n7842,n7843,n9675);
not (n7843,n7844);
or (n7844,n7845,n9674);
and (n7845,n7846,n9199);
xor (n7846,n7847,n9126);
xor (n7847,n7848,n9063);
xor (n7848,n7849,n9032);
or (n7849,n7850,n9031);
and (n7850,n7851,n8837);
xor (n7851,n7852,n8792);
xor (n7852,n7853,n8646);
xor (n7853,n7854,n8239);
xor (n7854,n7855,n8233);
xor (n7855,n7856,n8051);
wire s0n7856,s1n7856,notn7856;
or (n7856,s0n7856,s1n7856);
not(notn7856,n8048);
and (s0n7856,notn7856,1'b0);
and (s1n7856,n8048,n7857);
xor (n7857,n7858,n7868);
wire s0n7858,s1n7858,notn7858;
or (n7858,s0n7858,s1n7858);
not(notn7858,n7737);
and (s0n7858,notn7858,1'b0);
and (s1n7858,n7737,n7859);
nand (n7859,n7860,n7866);
or (n7860,n7861,n7862);
not (n7861,n7733);
not (n7862,n7863);
and (n7863,n7864,n626);
nor (n7864,n7865,n949);
not (n7865,n56);
nand (n7866,n7867,n7728);
and (n7867,n7865,n626);
or (n7868,n7869,n7989,n8047);
and (n7869,n7870,n7888);
xor (n7870,n7871,n7882);
wire s0n7871,s1n7871,notn7871;
or (n7871,s0n7871,s1n7871);
not(notn7871,n7737);
and (s0n7871,notn7871,1'b0);
and (s1n7871,n7737,n7872);
nand (n7872,n7873,n7876);
or (n7873,n7874,n7862);
not (n7874,n7875);
nand (n7876,n7867,n7877);
or (n7877,1'b0,n7878,n7879,n7880,n7881);
and (n7878,n2143,n910);
and (n7879,n6237,n909);
and (n7880,n1140,n906);
and (n7881,n7875,n900);
wire s0n7882,s1n7882,notn7882;
or (n7882,s0n7882,s1n7882);
not(notn7882,n7883);
and (s0n7882,notn7882,1'b0);
and (s1n7882,n7883,n7859);
xor (n7883,n7884,n7885);
not (n7884,n7738);
and (n7885,n7886,n7887);
not (n7886,n826);
not (n7887,n753);
and (n7888,n7889,n7891);
wire s0n7889,s1n7889,notn7889;
or (n7889,s0n7889,s1n7889);
not(notn7889,n7890);
and (s0n7889,notn7889,1'b0);
and (s1n7889,n7890,n7859);
xor (n7890,n7886,n7887);
or (n7891,n7892,n7895,n7988);
and (n7892,n7893,n7894);
wire s0n7893,s1n7893,notn7893;
or (n7893,s0n7893,s1n7893);
not(notn7893,n7890);
and (s0n7893,notn7893,1'b0);
and (s1n7893,n7890,n7872);
wire s0n7894,s1n7894,notn7894;
or (n7894,s0n7894,s1n7894);
not(notn7894,n753);
and (s0n7894,notn7894,1'b0);
and (s1n7894,n753,n7859);
and (n7895,n7894,n7896);
or (n7896,n7897,n7910,n7987);
and (n7897,n7898,n7909);
wire s0n7898,s1n7898,notn7898;
or (n7898,s0n7898,s1n7898);
not(notn7898,n7890);
and (s0n7898,notn7898,1'b0);
and (s1n7898,n7890,n7899);
nand (n7899,n7900,n7903);
or (n7900,n7901,n7862);
not (n7901,n7902);
nand (n7903,n7867,n7904);
or (n7904,1'b0,n7905,n7906,n7907,n7908);
and (n7905,n2240,n910);
and (n7906,n6286,n909);
and (n7907,n1312,n906);
and (n7908,n7902,n900);
wire s0n7909,s1n7909,notn7909;
or (n7909,s0n7909,s1n7909);
not(notn7909,n753);
and (s0n7909,notn7909,1'b0);
and (s1n7909,n753,n7872);
and (n7910,n7909,n7911);
or (n7911,n7912,n7925,n7986);
and (n7912,n7913,n7924);
wire s0n7913,s1n7913,notn7913;
or (n7913,s0n7913,s1n7913);
not(notn7913,n7890);
and (s0n7913,notn7913,1'b0);
and (s1n7913,n7890,n7914);
nand (n7914,n7915,n7918);
or (n7915,n7916,n7862);
not (n7916,n7917);
nand (n7918,n7867,n7919);
or (n7919,1'b0,n7920,n7921,n7922,n7923);
and (n7920,n2400,n910);
and (n7921,n6327,n909);
and (n7922,n1389,n906);
and (n7923,n7917,n900);
wire s0n7924,s1n7924,notn7924;
or (n7924,s0n7924,s1n7924);
not(notn7924,n753);
and (s0n7924,notn7924,1'b0);
and (s1n7924,n753,n7899);
and (n7925,n7924,n7926);
or (n7926,n7927,n7940,n7985);
and (n7927,n7928,n7939);
wire s0n7928,s1n7928,notn7928;
or (n7928,s0n7928,s1n7928);
not(notn7928,n7890);
and (s0n7928,notn7928,1'b0);
and (s1n7928,n7890,n7929);
nand (n7929,n7930,n7933);
or (n7930,n7931,n7862);
not (n7931,n7932);
nand (n7933,n7867,n7934);
or (n7934,1'b0,n7935,n7936,n7937,n7938);
and (n7935,n2528,n910);
and (n7936,n6389,n909);
and (n7937,n1551,n906);
and (n7938,n7932,n900);
wire s0n7939,s1n7939,notn7939;
or (n7939,s0n7939,s1n7939);
not(notn7939,n753);
and (s0n7939,notn7939,1'b0);
and (s1n7939,n753,n7914);
and (n7940,n7939,n7941);
or (n7941,n7942,n7955,n7957);
and (n7942,n7943,n7954);
wire s0n7943,s1n7943,notn7943;
or (n7943,s0n7943,s1n7943);
not(notn7943,n7890);
and (s0n7943,notn7943,1'b0);
and (s1n7943,n7890,n7944);
nand (n7944,n7945,n7948);
or (n7945,n7946,n7862);
not (n7946,n7947);
nand (n7948,n7867,n7949);
or (n7949,1'b0,n7950,n7951,n7952,n7953);
and (n7950,n2645,n910);
and (n7951,n6441,n909);
and (n7952,n1675,n906);
and (n7953,n7947,n900);
wire s0n7954,s1n7954,notn7954;
or (n7954,s0n7954,s1n7954);
not(notn7954,n753);
and (s0n7954,notn7954,1'b0);
and (s1n7954,n753,n7929);
and (n7955,n7954,n7956);
or (n7956,n7957,n7970,n7971);
and (n7957,n7958,n7969);
wire s0n7958,s1n7958,notn7958;
or (n7958,s0n7958,s1n7958);
not(notn7958,n7890);
and (s0n7958,notn7958,1'b0);
and (s1n7958,n7890,n7959);
nand (n7959,n7960,n7963);
or (n7960,n7961,n7862);
not (n7961,n7962);
nand (n7963,n7867,n7964);
or (n7964,1'b0,n7965,n7966,n7967,n7968);
and (n7965,n2765,n910);
and (n7966,n6494,n909);
and (n7967,n1798,n906);
and (n7968,n7962,n900);
wire s0n7969,s1n7969,notn7969;
or (n7969,s0n7969,s1n7969);
not(notn7969,n753);
and (s0n7969,notn7969,1'b0);
and (s1n7969,n753,n7944);
and (n7970,n7969,n7971);
and (n7971,n7972,n7984);
wire s0n7972,s1n7972,notn7972;
or (n7972,s0n7972,s1n7972);
not(notn7972,n7890);
and (s0n7972,notn7972,1'b0);
and (s1n7972,n7890,n7973);
nand (n7973,n7974,n7983);
or (n7974,n7975,n7982);
not (n7975,n7976);
or (n7976,1'b0,n7977,n7978,n7979,n7980);
and (n7977,n2888,n910);
and (n7978,n6555,n909);
and (n7979,n1918,n906);
and (n7980,n7981,n900);
not (n7982,n7867);
nand (n7983,n7863,n7981);
wire s0n7984,s1n7984,notn7984;
or (n7984,s0n7984,s1n7984);
not(notn7984,n753);
and (s0n7984,notn7984,1'b0);
and (s1n7984,n753,n7959);
and (n7985,n7928,n7941);
and (n7986,n7913,n7926);
and (n7987,n7898,n7911);
and (n7988,n7893,n7896);
and (n7989,n7888,n7990);
or (n7990,n7991,n7996,n8046);
and (n7991,n7992,n7995);
xor (n7992,n7993,n7994);
wire s0n7993,s1n7993,notn7993;
or (n7993,s0n7993,s1n7993);
not(notn7993,n7737);
and (s0n7993,notn7993,1'b0);
and (s1n7993,n7737,n7899);
wire s0n7994,s1n7994,notn7994;
or (n7994,s0n7994,s1n7994);
not(notn7994,n7883);
and (s0n7994,notn7994,1'b0);
and (s1n7994,n7883,n7872);
xor (n7995,n7889,n7891);
and (n7996,n7995,n7997);
or (n7997,n7998,n8004,n8045);
and (n7998,n7999,n8002);
xor (n7999,n8000,n8001);
wire s0n8000,s1n8000,notn8000;
or (n8000,s0n8000,s1n8000);
not(notn8000,n7737);
and (s0n8000,notn8000,1'b0);
and (s1n8000,n7737,n7914);
wire s0n8001,s1n8001,notn8001;
or (n8001,s0n8001,s1n8001);
not(notn8001,n7883);
and (s0n8001,notn8001,1'b0);
and (s1n8001,n7883,n7899);
xor (n8002,n8003,n7896);
xor (n8003,n7893,n7894);
and (n8004,n8002,n8005);
or (n8005,n8006,n8012,n8044);
and (n8006,n8007,n8010);
xor (n8007,n8008,n8009);
wire s0n8008,s1n8008,notn8008;
or (n8008,s0n8008,s1n8008);
not(notn8008,n7737);
and (s0n8008,notn8008,1'b0);
and (s1n8008,n7737,n7929);
wire s0n8009,s1n8009,notn8009;
or (n8009,s0n8009,s1n8009);
not(notn8009,n7883);
and (s0n8009,notn8009,1'b0);
and (s1n8009,n7883,n7914);
xor (n8010,n8011,n7911);
xor (n8011,n7898,n7909);
and (n8012,n8010,n8013);
or (n8013,n8014,n8020,n8043);
and (n8014,n8015,n8018);
xor (n8015,n8016,n8017);
wire s0n8016,s1n8016,notn8016;
or (n8016,s0n8016,s1n8016);
not(notn8016,n7737);
and (s0n8016,notn8016,1'b0);
and (s1n8016,n7737,n7944);
wire s0n8017,s1n8017,notn8017;
or (n8017,s0n8017,s1n8017);
not(notn8017,n7883);
and (s0n8017,notn8017,1'b0);
and (s1n8017,n7883,n7929);
xor (n8018,n8019,n7926);
xor (n8019,n7913,n7924);
and (n8020,n8018,n8021);
or (n8021,n8022,n8028,n8042);
and (n8022,n8023,n8026);
xor (n8023,n8024,n8025);
wire s0n8024,s1n8024,notn8024;
or (n8024,s0n8024,s1n8024);
not(notn8024,n7737);
and (s0n8024,notn8024,1'b0);
and (s1n8024,n7737,n7959);
wire s0n8025,s1n8025,notn8025;
or (n8025,s0n8025,s1n8025);
not(notn8025,n7883);
and (s0n8025,notn8025,1'b0);
and (s1n8025,n7883,n7944);
xor (n8026,n8027,n7941);
xor (n8027,n7928,n7939);
and (n8028,n8026,n8029);
or (n8029,n8030,n8036,n8041);
and (n8030,n8031,n8034);
xor (n8031,n8032,n8033);
wire s0n8032,s1n8032,notn8032;
or (n8032,s0n8032,s1n8032);
not(notn8032,n7737);
and (s0n8032,notn8032,1'b0);
and (s1n8032,n7737,n7973);
wire s0n8033,s1n8033,notn8033;
or (n8033,s0n8033,s1n8033);
not(notn8033,n7883);
and (s0n8033,notn8033,1'b0);
and (s1n8033,n7883,n7959);
xor (n8034,n8035,n7956);
xor (n8035,n7943,n7954);
and (n8036,n8034,n8037);
and (n8037,n8038,n8039);
wire s0n8038,s1n8038,notn8038;
or (n8038,s0n8038,s1n8038);
not(notn8038,n7883);
and (s0n8038,notn8038,1'b0);
and (s1n8038,n7883,n7973);
xor (n8039,n8040,n7971);
xor (n8040,n7958,n7969);
and (n8041,n8031,n8037);
and (n8042,n8023,n8029);
and (n8043,n8015,n8021);
and (n8044,n8007,n8013);
and (n8045,n7999,n8005);
and (n8046,n7992,n7997);
and (n8047,n7870,n7990);
xor (n8048,n8049,n8050);
not (n8049,n679);
not (n8050,n35);
wire s0n8051,s1n8051,notn8051;
or (n8051,s0n8051,s1n8051);
not(notn8051,n7786);
and (s0n8051,notn8051,1'b0);
and (s1n8051,n7786,n8052);
xor (n8052,n8053,n8176);
xor (n8053,n8054,n8077);
xor (n8054,n8055,n8066);
wire s0n8055,s1n8055,notn8055;
or (n8055,s0n8055,s1n8055);
not(notn8055,n7737);
and (s0n8055,notn8055,1'b0);
and (s1n8055,n7737,n8056);
nand (n8056,n8057,n8060);
or (n8057,n8058,n7862);
not (n8058,n8059);
nand (n8060,n7867,n8061);
or (n8061,1'b0,n8062,n8063,n8064,n8065);
and (n8062,n2224,n910);
and (n8063,n6242,n909);
and (n8064,n3012,n906);
and (n8065,n8059,n900);
wire s0n8066,s1n8066,notn8066;
or (n8066,s0n8066,s1n8066);
not(notn8066,n7883);
and (s0n8066,notn8066,1'b0);
and (s1n8066,n7883,n8067);
nand (n8067,n8068,n8071);
or (n8068,n8069,n7862);
not (n8069,n8070);
nand (n8071,n7867,n8072);
or (n8072,1'b0,n8073,n8074,n8075,n8076);
and (n8073,n2062,n910);
and (n8074,n6196,n909);
and (n8075,n3080,n906);
and (n8076,n8070,n900);
and (n8077,n8078,n8079);
wire s0n8078,s1n8078,notn8078;
or (n8078,s0n8078,s1n8078);
not(notn8078,n7890);
and (s0n8078,notn8078,1'b0);
and (s1n8078,n7890,n8067);
or (n8079,n8080,n8083,n8175);
and (n8080,n8081,n8082);
wire s0n8081,s1n8081,notn8081;
or (n8081,s0n8081,s1n8081);
not(notn8081,n7890);
and (s0n8081,notn8081,1'b0);
and (s1n8081,n7890,n8056);
wire s0n8082,s1n8082,notn8082;
or (n8082,s0n8082,s1n8082);
not(notn8082,n753);
and (s0n8082,notn8082,1'b0);
and (s1n8082,n753,n8067);
and (n8083,n8082,n8084);
or (n8084,n8085,n8098,n8174);
and (n8085,n8086,n8097);
wire s0n8086,s1n8086,notn8086;
or (n8086,s0n8086,s1n8086);
not(notn8086,n7890);
and (s0n8086,notn8086,1'b0);
and (s1n8086,n7890,n8087);
nand (n8087,n8088,n8091);
or (n8088,n8089,n7862);
not (n8089,n8090);
nand (n8091,n7867,n8092);
or (n8092,1'b0,n8093,n8094,n8095,n8096);
and (n8093,n2294,n910);
and (n8094,n6276,n909);
and (n8095,n3452,n906);
and (n8096,n8090,n900);
wire s0n8097,s1n8097,notn8097;
or (n8097,s0n8097,s1n8097);
not(notn8097,n753);
and (s0n8097,notn8097,1'b0);
and (s1n8097,n753,n8056);
and (n8098,n8097,n8099);
or (n8099,n8100,n8113,n8173);
and (n8100,n8101,n8112);
wire s0n8101,s1n8101,notn8101;
or (n8101,s0n8101,s1n8101);
not(notn8101,n7890);
and (s0n8101,notn8101,1'b0);
and (s1n8101,n7890,n8102);
nand (n8102,n8103,n8106);
or (n8103,n8104,n7862);
not (n8104,n8105);
nand (n8106,n7867,n8107);
or (n8107,1'b0,n8108,n8109,n8110,n8111);
and (n8108,n2460,n910);
and (n8109,n6335,n909);
and (n8110,n3519,n906);
and (n8111,n8105,n900);
wire s0n8112,s1n8112,notn8112;
or (n8112,s0n8112,s1n8112);
not(notn8112,n753);
and (s0n8112,notn8112,1'b0);
and (s1n8112,n753,n8087);
and (n8113,n8112,n8114);
or (n8114,n8115,n8128,n8172);
and (n8115,n8116,n8127);
wire s0n8116,s1n8116,notn8116;
or (n8116,s0n8116,s1n8116);
not(notn8116,n7890);
and (s0n8116,notn8116,1'b0);
and (s1n8116,n7890,n8117);
nand (n8117,n8118,n8121);
or (n8118,n8119,n7862);
not (n8119,n8120);
nand (n8121,n7867,n8122);
or (n8122,1'b0,n8123,n8124,n8125,n8126);
and (n8123,n2585,n910);
and (n8124,n6378,n909);
and (n8125,n3379,n906);
and (n8126,n8120,n900);
wire s0n8127,s1n8127,notn8127;
or (n8127,s0n8127,s1n8127);
not(notn8127,n753);
and (s0n8127,notn8127,1'b0);
and (s1n8127,n753,n8102);
and (n8128,n8127,n8129);
or (n8129,n8130,n8143,n8145);
and (n8130,n8131,n8142);
wire s0n8131,s1n8131,notn8131;
or (n8131,s0n8131,s1n8131);
not(notn8131,n7890);
and (s0n8131,notn8131,1'b0);
and (s1n8131,n7890,n8132);
nand (n8132,n8133,n8141);
or (n8133,n8134,n7982);
not (n8134,n8135);
or (n8135,1'b0,n8136,n8137,n8138,n8139);
and (n8136,n2702,n910);
and (n8137,n6431,n909);
and (n8138,n3170,n906);
and (n8139,n8140,n900);
nand (n8141,n7863,n8140);
wire s0n8142,s1n8142,notn8142;
or (n8142,s0n8142,s1n8142);
not(notn8142,n753);
and (s0n8142,notn8142,1'b0);
and (s1n8142,n753,n8117);
and (n8143,n8142,n8144);
or (n8144,n8145,n8158,n8159);
and (n8145,n8146,n8157);
wire s0n8146,s1n8146,notn8146;
or (n8146,s0n8146,s1n8146);
not(notn8146,n7890);
and (s0n8146,notn8146,1'b0);
and (s1n8146,n7890,n8147);
nand (n8147,n8148,n8156);
or (n8148,n8149,n7982);
not (n8149,n8150);
or (n8150,1'b0,n8151,n8152,n8153,n8154);
and (n8151,n2826,n910);
and (n8152,n6484,n909);
and (n8153,n3237,n906);
and (n8154,n8155,n900);
nand (n8156,n7863,n8155);
wire s0n8157,s1n8157,notn8157;
or (n8157,s0n8157,s1n8157);
not(notn8157,n753);
and (s0n8157,notn8157,1'b0);
and (s1n8157,n753,n8132);
and (n8158,n8157,n8159);
and (n8159,n8160,n8171);
wire s0n8160,s1n8160,notn8160;
or (n8160,s0n8160,s1n8160);
not(notn8160,n7890);
and (s0n8160,notn8160,1'b0);
and (s1n8160,n7890,n8161);
nand (n8161,n8162,n8165);
or (n8162,n8163,n7862);
not (n8163,n8164);
nand (n8165,n7867,n8166);
or (n8166,1'b0,n8167,n8168,n8169,n8170);
and (n8167,n2951,n910);
and (n8168,n6545,n909);
and (n8169,n3306,n906);
and (n8170,n8164,n900);
wire s0n8171,s1n8171,notn8171;
or (n8171,s0n8171,s1n8171);
not(notn8171,n753);
and (s0n8171,notn8171,1'b0);
and (s1n8171,n753,n8147);
and (n8172,n8116,n8129);
and (n8173,n8101,n8114);
and (n8174,n8086,n8099);
and (n8175,n8081,n8084);
or (n8176,n8177,n8182,n8232);
and (n8177,n8178,n8181);
xor (n8178,n8179,n8180);
wire s0n8179,s1n8179,notn8179;
or (n8179,s0n8179,s1n8179);
not(notn8179,n7737);
and (s0n8179,notn8179,1'b0);
and (s1n8179,n7737,n8087);
wire s0n8180,s1n8180,notn8180;
or (n8180,s0n8180,s1n8180);
not(notn8180,n7883);
and (s0n8180,notn8180,1'b0);
and (s1n8180,n7883,n8056);
xor (n8181,n8078,n8079);
and (n8182,n8181,n8183);
or (n8183,n8184,n8190,n8231);
and (n8184,n8185,n8188);
xor (n8185,n8186,n8187);
wire s0n8186,s1n8186,notn8186;
or (n8186,s0n8186,s1n8186);
not(notn8186,n7737);
and (s0n8186,notn8186,1'b0);
and (s1n8186,n7737,n8102);
wire s0n8187,s1n8187,notn8187;
or (n8187,s0n8187,s1n8187);
not(notn8187,n7883);
and (s0n8187,notn8187,1'b0);
and (s1n8187,n7883,n8087);
xor (n8188,n8189,n8084);
xor (n8189,n8081,n8082);
and (n8190,n8188,n8191);
or (n8191,n8192,n8198,n8230);
and (n8192,n8193,n8196);
xor (n8193,n8194,n8195);
wire s0n8194,s1n8194,notn8194;
or (n8194,s0n8194,s1n8194);
not(notn8194,n7737);
and (s0n8194,notn8194,1'b0);
and (s1n8194,n7737,n8117);
wire s0n8195,s1n8195,notn8195;
or (n8195,s0n8195,s1n8195);
not(notn8195,n7883);
and (s0n8195,notn8195,1'b0);
and (s1n8195,n7883,n8102);
xor (n8196,n8197,n8099);
xor (n8197,n8086,n8097);
and (n8198,n8196,n8199);
or (n8199,n8200,n8206,n8229);
and (n8200,n8201,n8204);
xor (n8201,n8202,n8203);
wire s0n8202,s1n8202,notn8202;
or (n8202,s0n8202,s1n8202);
not(notn8202,n7737);
and (s0n8202,notn8202,1'b0);
and (s1n8202,n7737,n8132);
wire s0n8203,s1n8203,notn8203;
or (n8203,s0n8203,s1n8203);
not(notn8203,n7883);
and (s0n8203,notn8203,1'b0);
and (s1n8203,n7883,n8117);
xor (n8204,n8205,n8114);
xor (n8205,n8101,n8112);
and (n8206,n8204,n8207);
or (n8207,n8208,n8214,n8228);
and (n8208,n8209,n8212);
xor (n8209,n8210,n8211);
wire s0n8210,s1n8210,notn8210;
or (n8210,s0n8210,s1n8210);
not(notn8210,n7737);
and (s0n8210,notn8210,1'b0);
and (s1n8210,n7737,n8147);
wire s0n8211,s1n8211,notn8211;
or (n8211,s0n8211,s1n8211);
not(notn8211,n7883);
and (s0n8211,notn8211,1'b0);
and (s1n8211,n7883,n8132);
xor (n8212,n8213,n8129);
xor (n8213,n8116,n8127);
and (n8214,n8212,n8215);
or (n8215,n8216,n8222,n8227);
and (n8216,n8217,n8220);
xor (n8217,n8218,n8219);
wire s0n8218,s1n8218,notn8218;
or (n8218,s0n8218,s1n8218);
not(notn8218,n7737);
and (s0n8218,notn8218,1'b0);
and (s1n8218,n7737,n8161);
wire s0n8219,s1n8219,notn8219;
or (n8219,s0n8219,s1n8219);
not(notn8219,n7883);
and (s0n8219,notn8219,1'b0);
and (s1n8219,n7883,n8147);
xor (n8220,n8221,n8144);
xor (n8221,n8131,n8142);
and (n8222,n8220,n8223);
and (n8223,n8224,n8225);
wire s0n8224,s1n8224,notn8224;
or (n8224,s0n8224,s1n8224);
not(notn8224,n7883);
and (s0n8224,notn8224,1'b0);
and (s1n8224,n7883,n8161);
xor (n8225,n8226,n8159);
xor (n8226,n8146,n8157);
and (n8227,n8217,n8223);
and (n8228,n8209,n8215);
and (n8229,n8201,n8207);
and (n8230,n8193,n8199);
and (n8231,n8185,n8191);
and (n8232,n8178,n8183);
wire s0n8233,s1n8233,notn8233;
or (n8233,s0n8233,s1n8233);
not(notn8233,n8236);
and (s0n8233,notn8233,1'b0);
and (s1n8233,n8236,n8234);
xor (n8234,n8235,n7990);
xor (n8235,n7870,n7888);
xor (n8236,n8237,n8238);
not (n8237,n7786);
and (n8238,n8049,n8050);
xor (n8239,n8240,n8635);
xor (n8240,n8241,n8619);
or (n8241,n8242,n8618);
and (n8242,n8243,n8486);
xor (n8243,n8244,n8474);
and (n8244,n8245,n8458);
xor (n8245,n8246,n8378);
wire s0n8246,s1n8246,notn8246;
or (n8246,s0n8246,s1n8246);
not(notn8246,n7785);
and (s0n8246,notn8246,1'b0);
and (s1n8246,n7785,n8247);
xor (n8247,n8248,n8350);
xor (n8248,n8249,n8261);
not (n8249,n8250);
nand (n8250,n7738,n8251);
nand (n8251,n8252,n8260);
or (n8252,n8253,n7982);
not (n8253,n8254);
or (n8254,1'b0,n8255,n8256,n8257,n8258);
and (n8255,n2397,n910);
and (n8256,n5709,n909);
and (n8257,n1429,n906);
and (n8258,n8259,n900);
nand (n8260,n7863,n8259);
xor (n8261,n8262,n8285);
xor (n8262,n8263,n8274);
wire s0n8263,s1n8263,notn8263;
or (n8263,s0n8263,s1n8263);
not(notn8263,n826);
and (s0n8263,notn8263,1'b0);
and (s1n8263,n826,n8264);
nand (n8264,n8265,n8273);
or (n8265,n8266,n7982);
not (n8266,n8267);
or (n8267,1'b0,n8268,n8269,n8270,n8271);
and (n8268,n2278,n910);
and (n8269,n5619,n909);
and (n8270,n1309,n906);
and (n8271,n8272,n900);
nand (n8273,n7863,n8272);
wire s0n8274,s1n8274,notn8274;
or (n8274,s0n8274,s1n8274);
not(notn8274,n753);
and (s0n8274,notn8274,1'b0);
and (s1n8274,n753,n8275);
nand (n8275,n8276,n8279);
or (n8276,n8277,n7862);
not (n8277,n8278);
nand (n8279,n7867,n8280);
or (n8280,1'b0,n8281,n8282,n8283,n8284);
and (n8281,n2157,n910);
and (n8282,n5553,n909);
and (n8283,n1181,n906);
and (n8284,n8278,n900);
or (n8285,n8286,n8289,n8349);
and (n8286,n8287,n8288);
wire s0n8287,s1n8287,notn8287;
or (n8287,s0n8287,s1n8287);
not(notn8287,n826);
and (s0n8287,notn8287,1'b0);
and (s1n8287,n826,n8251);
wire s0n8288,s1n8288,notn8288;
or (n8288,s0n8288,s1n8288);
not(notn8288,n753);
and (s0n8288,notn8288,1'b0);
and (s1n8288,n753,n8264);
and (n8289,n8288,n8290);
or (n8290,n8291,n8304,n8348);
and (n8291,n8292,n8303);
wire s0n8292,s1n8292,notn8292;
or (n8292,s0n8292,s1n8292);
not(notn8292,n826);
and (s0n8292,notn8292,1'b0);
and (s1n8292,n826,n8293);
nand (n8293,n8294,n8297);
or (n8294,n8295,n7862);
not (n8295,n8296);
nand (n8297,n7867,n8298);
or (n8298,1'b0,n8299,n8300,n8301,n8302);
and (n8299,n2525,n910);
and (n8300,n5788,n909);
and (n8301,n1548,n906);
and (n8302,n8296,n900);
wire s0n8303,s1n8303,notn8303;
or (n8303,s0n8303,s1n8303);
not(notn8303,n753);
and (s0n8303,notn8303,1'b0);
and (s1n8303,n753,n8251);
and (n8304,n8303,n8305);
or (n8305,n8306,n8319,n8321);
and (n8306,n8307,n8318);
wire s0n8307,s1n8307,notn8307;
or (n8307,s0n8307,s1n8307);
not(notn8307,n826);
and (s0n8307,notn8307,1'b0);
and (s1n8307,n826,n8308);
nand (n8308,n8309,n8317);
or (n8309,n8310,n7982);
not (n8310,n8311);
or (n8311,1'b0,n8312,n8313,n8314,n8315);
and (n8312,n2642,n910);
and (n8313,n5828,n909);
and (n8314,n1672,n906);
and (n8315,n8316,n900);
nand (n8317,n7863,n8316);
wire s0n8318,s1n8318,notn8318;
or (n8318,s0n8318,s1n8318);
not(notn8318,n753);
and (s0n8318,notn8318,1'b0);
and (s1n8318,n753,n8293);
and (n8319,n8318,n8320);
or (n8320,n8321,n8334,n8335);
and (n8321,n8322,n8333);
wire s0n8322,s1n8322,notn8322;
or (n8322,s0n8322,s1n8322);
not(notn8322,n826);
and (s0n8322,notn8322,1'b0);
and (s1n8322,n826,n8323);
nand (n8323,n8324,n8327);
or (n8324,n8325,n7862);
not (n8325,n8326);
nand (n8327,n7867,n8328);
or (n8328,1'b0,n8329,n8330,n8331,n8332);
and (n8329,n2762,n910);
and (n8330,n5927,n909);
and (n8331,n1795,n906);
and (n8332,n8326,n900);
wire s0n8333,s1n8333,notn8333;
or (n8333,s0n8333,s1n8333);
not(notn8333,n753);
and (s0n8333,notn8333,1'b0);
and (s1n8333,n753,n8308);
and (n8334,n8333,n8335);
and (n8335,n8336,n8347);
wire s0n8336,s1n8336,notn8336;
or (n8336,s0n8336,s1n8336);
not(notn8336,n826);
and (s0n8336,notn8336,1'b0);
and (s1n8336,n826,n8337);
nand (n8337,n8338,n8341);
or (n8338,n8339,n7862);
not (n8339,n8340);
nand (n8341,n7867,n8342);
or (n8342,1'b0,n8343,n8344,n8345,n8346);
and (n8343,n2885,n910);
and (n8344,n5999,n909);
and (n8345,n1915,n906);
and (n8346,n8340,n900);
wire s0n8347,s1n8347,notn8347;
or (n8347,s0n8347,s1n8347);
not(notn8347,n753);
and (s0n8347,notn8347,1'b0);
and (s1n8347,n753,n8323);
and (n8348,n8292,n8305);
and (n8349,n8287,n8290);
or (n8350,n8351,n8356,n8377);
and (n8351,n8352,n8354);
not (n8352,n8353);
nand (n8353,n7738,n8293);
xor (n8354,n8355,n8290);
xor (n8355,n8287,n8288);
and (n8356,n8354,n8357);
or (n8357,n8358,n8363,n8376);
and (n8358,n8359,n8361);
not (n8359,n8360);
nand (n8360,n7738,n8308);
xor (n8361,n8362,n8305);
xor (n8362,n8292,n8303);
and (n8363,n8361,n8364);
or (n8364,n8365,n8370,n8375);
and (n8365,n8366,n8368);
not (n8366,n8367);
nand (n8367,n7738,n8323);
xor (n8368,n8369,n8320);
xor (n8369,n8307,n8318);
and (n8370,n8368,n8371);
and (n8371,n8372,n8373);
and (n8372,n7738,n8337);
xor (n8373,n8374,n8335);
xor (n8374,n8322,n8333);
and (n8375,n8366,n8371);
and (n8376,n8359,n8364);
and (n8377,n8352,n8357);
xor (n8378,n8379,n8420);
xor (n8379,n8380,n8408);
xor (n8380,n8381,n8406);
xor (n8381,n8382,n8394);
nor (n8382,n8383,n8050);
nand (n8383,n7738,n8384);
nand (n8384,n8385,n8393);
or (n8385,n8386,n7982);
not (n8386,n8387);
or (n8387,1'b0,n8388,n8389,n8390,n8391);
and (n8388,n2102,n910);
and (n8389,n5459,n909);
and (n8390,n3077,n906);
and (n8391,n8392,n900);
nand (n8393,n7863,n8392);
and (n8394,n8395,n35);
and (n8395,n7738,n8396);
nand (n8396,n8397,n8400);
or (n8397,n8398,n7862);
not (n8398,n8399);
nand (n8400,n7867,n8401);
or (n8401,1'b0,n8402,n8403,n8404,n8405);
and (n8402,n2052,n910);
and (n8403,n5458,n909);
and (n8404,n1026,n906);
and (n8405,n8399,n900);
and (n8406,n8394,n8407);
wire s0n8407,s1n8407,notn8407;
or (n8407,s0n8407,s1n8407);
not(notn8407,n826);
and (s0n8407,notn8407,1'b0);
and (s1n8407,n826,n8275);
and (n8408,n8382,n8409);
wire s0n8409,s1n8409,notn8409;
or (n8409,s0n8409,s1n8409);
not(notn8409,n826);
and (s0n8409,notn8409,1'b0);
and (s1n8409,n826,n8410);
nand (n8410,n8411,n8419);
or (n8411,n8412,n7982);
not (n8412,n8413);
or (n8413,1'b0,n8414,n8415,n8416,n8417);
and (n8414,n2221,n910);
and (n8415,n5554,n909);
and (n8416,n3009,n906);
and (n8417,n8418,n900);
nand (n8419,n7863,n8418);
or (n8420,n8421,n8457);
and (n8421,n8422,n8436);
xor (n8422,n8423,n8428);
nor (n8423,n8424,n8050);
xnor (n8424,n8425,n8426);
nand (n8425,n7738,n8410);
not (n8426,n8427);
wire s0n8427,s1n8427,notn8427;
or (n8427,s0n8427,s1n8427);
not(notn8427,n826);
and (s0n8427,notn8427,1'b0);
and (s1n8427,n826,n8384);
and (n8428,n8429,n35);
nand (n8429,n8430,n8435);
or (n8430,n8431,n8433);
not (n8431,n8432);
wire s0n8432,s1n8432,notn8432;
or (n8432,s0n8432,s1n8432);
not(notn8432,n826);
and (s0n8432,notn8432,1'b0);
and (s1n8432,n826,n8396);
not (n8433,n8434);
nand (n8434,n7738,n8275);
or (n8435,n8434,n8432);
and (n8436,n8437,n35);
or (n8437,n8438,n8454);
nor (n8438,n8439,n8453);
and (n8439,n8440,n8451);
nand (n8440,n7738,n8441);
nand (n8441,n8442,n8450);
or (n8442,n8443,n7982);
not (n8443,n8444);
or (n8444,1'b0,n8445,n8446,n8447,n8448);
and (n8445,n2332,n910);
and (n8446,n5620,n909);
and (n8447,n3449,n906);
and (n8448,n8449,n900);
nand (n8450,n7863,n8449);
not (n8451,n8452);
wire s0n8452,s1n8452,notn8452;
or (n8452,s0n8452,s1n8452);
not(notn8452,n753);
and (s0n8452,notn8452,1'b0);
and (s1n8452,n753,n8384);
not (n8453,n8409);
nor (n8454,n8455,n8383);
not (n8455,n8456);
wire s0n8456,s1n8456,notn8456;
or (n8456,s0n8456,s1n8456);
not(notn8456,n753);
and (s0n8456,notn8456,1'b0);
and (s1n8456,n753,n8441);
and (n8457,n8423,n8428);
wire s0n8458,s1n8458,notn8458;
or (n8458,s0n8458,s1n8458);
not(notn8458,n8236);
and (s0n8458,notn8458,1'b0);
and (s1n8458,n8236,n8459);
xor (n8459,n8460,n8470);
xor (n8460,n8461,n8463);
not (n8461,n8462);
nand (n8462,n7738,n8264);
xor (n8463,n8464,n8466);
xor (n8464,n8407,n8465);
wire s0n8465,s1n8465,notn8465;
or (n8465,s0n8465,s1n8465);
not(notn8465,n753);
and (s0n8465,notn8465,1'b0);
and (s1n8465,n753,n8396);
or (n8466,n8467,n8468,n8469);
and (n8467,n8263,n8274);
and (n8468,n8274,n8285);
and (n8469,n8263,n8285);
or (n8470,n8471,n8472,n8473);
and (n8471,n8249,n8261);
and (n8472,n8261,n8350);
and (n8473,n8249,n8350);
wire s0n8474,s1n8474,notn8474;
or (n8474,s0n8474,s1n8474);
not(notn8474,n8236);
and (s0n8474,notn8474,1'b0);
and (s1n8474,n8236,n8475);
xor (n8475,n8476,n8482);
xor (n8476,n8433,n8477);
xor (n8477,n8432,n8478);
or (n8478,n8479,n8480,n8481);
and (n8479,n8407,n8465);
and (n8480,n8465,n8466);
and (n8481,n8407,n8466);
or (n8482,n8483,n8484,n8485);
and (n8483,n8461,n8463);
and (n8484,n8463,n8470);
and (n8485,n8461,n8470);
wire s0n8486,s1n8486,notn8486;
or (n8486,s0n8486,s1n8486);
not(notn8486,n7786);
and (s0n8486,notn8486,1'b0);
and (s1n8486,n7786,n8487);
xor (n8487,n8488,n8575);
xor (n8488,n8489,n8490);
not (n8489,n8425);
xor (n8490,n8427,n8491);
or (n8491,n8492,n8493,n8574);
and (n8492,n8409,n8452);
and (n8493,n8452,n8494);
or (n8494,n8495,n8498,n8573);
and (n8495,n8496,n8497);
wire s0n8496,s1n8496,notn8496;
or (n8496,s0n8496,s1n8496);
not(notn8496,n826);
and (s0n8496,notn8496,1'b0);
and (s1n8496,n826,n8441);
wire s0n8497,s1n8497,notn8497;
or (n8497,s0n8497,s1n8497);
not(notn8497,n753);
and (s0n8497,notn8497,1'b0);
and (s1n8497,n753,n8410);
and (n8498,n8497,n8499);
or (n8499,n8500,n8512,n8572);
and (n8500,n8501,n8456);
wire s0n8501,s1n8501,notn8501;
or (n8501,s0n8501,s1n8501);
not(notn8501,n826);
and (s0n8501,notn8501,1'b0);
and (s1n8501,n826,n8502);
nand (n8502,n8503,n8511);
or (n8503,n8504,n7982);
not (n8504,n8505);
or (n8505,1'b0,n8506,n8507,n8508,n8509);
and (n8506,n2457,n910);
and (n8507,n5710,n909);
and (n8508,n3516,n906);
and (n8509,n8510,n900);
nand (n8511,n7863,n8510);
and (n8512,n8456,n8513);
or (n8513,n8514,n8527,n8571);
and (n8514,n8515,n8526);
wire s0n8515,s1n8515,notn8515;
or (n8515,s0n8515,s1n8515);
not(notn8515,n826);
and (s0n8515,notn8515,1'b0);
and (s1n8515,n826,n8516);
nand (n8516,n8517,n8525);
or (n8517,n8518,n7982);
not (n8518,n8519);
or (n8519,1'b0,n8520,n8521,n8522,n8523);
and (n8520,n2582,n910);
and (n8521,n5789,n909);
and (n8522,n3376,n906);
and (n8523,n8524,n900);
nand (n8525,n7863,n8524);
wire s0n8526,s1n8526,notn8526;
or (n8526,s0n8526,s1n8526);
not(notn8526,n753);
and (s0n8526,notn8526,1'b0);
and (s1n8526,n753,n8502);
and (n8527,n8526,n8528);
or (n8528,n8529,n8542,n8544);
and (n8529,n8530,n8541);
wire s0n8530,s1n8530,notn8530;
or (n8530,s0n8530,s1n8530);
not(notn8530,n826);
and (s0n8530,notn8530,1'b0);
and (s1n8530,n826,n8531);
nand (n8531,n8532,n8535);
or (n8532,n8533,n7862);
not (n8533,n8534);
nand (n8535,n7867,n8536);
or (n8536,1'b0,n8537,n8538,n8539,n8540);
and (n8537,n2699,n910);
and (n8538,n5829,n909);
and (n8539,n3167,n906);
and (n8540,n8534,n900);
wire s0n8541,s1n8541,notn8541;
or (n8541,s0n8541,s1n8541);
not(notn8541,n753);
and (s0n8541,notn8541,1'b0);
and (s1n8541,n753,n8516);
and (n8542,n8541,n8543);
or (n8543,n8544,n8557,n8558);
and (n8544,n8545,n8556);
wire s0n8545,s1n8545,notn8545;
or (n8545,s0n8545,s1n8545);
not(notn8545,n826);
and (s0n8545,notn8545,1'b0);
and (s1n8545,n826,n8546);
nand (n8546,n8547,n8555);
or (n8547,n8548,n7982);
not (n8548,n8549);
or (n8549,1'b0,n8550,n8551,n8552,n8553);
and (n8550,n2823,n910);
and (n8551,n5928,n909);
and (n8552,n3234,n906);
and (n8553,n8554,n900);
nand (n8555,n7863,n8554);
wire s0n8556,s1n8556,notn8556;
or (n8556,s0n8556,s1n8556);
not(notn8556,n753);
and (s0n8556,notn8556,1'b0);
and (s1n8556,n753,n8531);
and (n8557,n8556,n8558);
and (n8558,n8559,n8570);
wire s0n8559,s1n8559,notn8559;
or (n8559,s0n8559,s1n8559);
not(notn8559,n826);
and (s0n8559,notn8559,1'b0);
and (s1n8559,n826,n8560);
nand (n8560,n8561,n8569);
or (n8561,n8562,n7982);
not (n8562,n8563);
or (n8563,1'b0,n8564,n8565,n8566,n8567);
and (n8564,n2948,n910);
and (n8565,n6000,n909);
and (n8566,n3303,n906);
and (n8567,n8568,n900);
nand (n8569,n7863,n8568);
wire s0n8570,s1n8570,notn8570;
or (n8570,s0n8570,s1n8570);
not(notn8570,n753);
and (s0n8570,notn8570,1'b0);
and (s1n8570,n753,n8546);
and (n8571,n8515,n8528);
and (n8572,n8501,n8513);
and (n8573,n8496,n8499);
and (n8574,n8409,n8494);
or (n8575,n8576,n8580,n8617);
and (n8576,n8577,n8578);
not (n8577,n8440);
xor (n8578,n8579,n8494);
xor (n8579,n8409,n8452);
and (n8580,n8578,n8581);
or (n8581,n8582,n8587,n8616);
and (n8582,n8583,n8585);
not (n8583,n8584);
nand (n8584,n7738,n8502);
xor (n8585,n8586,n8499);
xor (n8586,n8496,n8497);
and (n8587,n8585,n8588);
or (n8588,n8589,n8593,n8615);
and (n8589,n8590,n8591);
and (n8590,n7738,n8516);
xor (n8591,n8592,n8513);
xor (n8592,n8501,n8456);
and (n8593,n8591,n8594);
or (n8594,n8595,n8600,n8614);
and (n8595,n8596,n8598);
not (n8596,n8597);
nand (n8597,n7738,n8531);
xor (n8598,n8599,n8528);
xor (n8599,n8515,n8526);
and (n8600,n8598,n8601);
or (n8601,n8602,n8607,n8613);
and (n8602,n8603,n8605);
not (n8603,n8604);
nand (n8604,n7738,n8546);
xor (n8605,n8606,n8543);
xor (n8606,n8530,n8541);
and (n8607,n8605,n8608);
and (n8608,n8609,n8611);
not (n8609,n8610);
nand (n8610,n7738,n8560);
xor (n8611,n8612,n8558);
xor (n8612,n8545,n8556);
and (n8613,n8603,n8608);
and (n8614,n8596,n8601);
and (n8615,n8590,n8594);
and (n8616,n8583,n8588);
and (n8617,n8577,n8581);
and (n8618,n8244,n8474);
xor (n8619,n8620,n8632);
xor (n8620,n8621,n8631);
wire s0n8621,s1n8621,notn8621;
or (n8621,s0n8621,s1n8621);
not(notn8621,n8048);
and (s0n8621,notn8621,1'b0);
and (s1n8621,n8048,n8622);
or (n8622,n8623,n8625,n8630);
and (n8623,n8395,n8624);
and (n8624,n8432,n8478);
and (n8625,n8624,n8626);
or (n8626,n8627,n8628,n8629);
and (n8627,n8433,n8477);
and (n8628,n8477,n8482);
and (n8629,n8433,n8482);
and (n8630,n8395,n8626);
wire s0n8631,s1n8631,notn8631;
or (n8631,s0n8631,s1n8631);
not(notn8631,n7785);
and (s0n8631,notn8631,1'b0);
and (s1n8631,n7785,n8475);
wire s0n8632,s1n8632,notn8632;
or (n8632,s0n8632,s1n8632);
not(notn8632,n8236);
and (s0n8632,notn8632,1'b0);
and (s1n8632,n8236,n8633);
xor (n8633,n8634,n8626);
xor (n8634,n8395,n8624);
wire s0n8635,s1n8635,notn8635;
or (n8635,s0n8635,s1n8635);
not(notn8635,n679);
and (s0n8635,notn8635,1'b0);
and (s1n8635,n679,n8636);
or (n8636,n8637,n8640,n8645);
and (n8637,n8638,n8639);
not (n8638,n8383);
and (n8639,n8427,n8491);
and (n8640,n8639,n8641);
or (n8641,n8642,n8643,n8644);
and (n8642,n8489,n8490);
and (n8643,n8490,n8575);
and (n8644,n8489,n8575);
and (n8645,n8638,n8641);
or (n8646,n8647,n8791);
and (n8647,n8648,n8712);
xor (n8648,n8649,n8711);
or (n8649,n8650,n8710);
and (n8650,n8651,n8658);
xor (n8651,n8652,n8655);
wire s0n8652,s1n8652,notn8652;
or (n8652,s0n8652,s1n8652);
not(notn8652,n679);
and (s0n8652,notn8652,1'b0);
and (s1n8652,n679,n8653);
xor (n8653,n8654,n8183);
xor (n8654,n8178,n8181);
wire s0n8655,s1n8655,notn8655;
or (n8655,s0n8655,s1n8655);
not(notn8655,n7786);
and (s0n8655,notn8655,1'b0);
and (s1n8655,n7786,n8656);
xor (n8656,n8657,n8191);
xor (n8657,n8185,n8188);
and (n8658,n8659,n8236);
xor (n8659,n8660,n8672);
nor (n8660,n8661,n8671);
not (n8661,n8662);
or (n8662,n8663,n8666);
xor (n8663,n8664,n7897);
xor (n8664,n8001,n8665);
xor (n8665,n8003,n8000);
or (n8666,n8667,n8670);
and (n8667,n8668,n7912);
xor (n8668,n8009,n8669);
xor (n8669,n8011,n8008);
and (n8670,n8009,n8669);
and (n8671,n8663,n8666);
nand (n8672,n8673,n8709);
or (n8673,n8674,n8682);
not (n8674,n8675);
or (n8675,n8676,n8677);
xor (n8676,n8668,n7912);
or (n8677,n8678,n8681);
and (n8678,n8679,n7927);
xor (n8679,n8017,n8680);
xor (n8680,n8019,n8016);
and (n8681,n8017,n8680);
not (n8682,n8683);
nand (n8683,n8684,n8705,n8708);
nand (n8684,n8685,n8692,n8702);
or (n8685,n8686,n8687);
xor (n8686,n8679,n7927);
or (n8687,n8688,n8691);
and (n8688,n8689,n8690);
xor (n8689,n8025,n7942);
xor (n8690,n8027,n8024);
and (n8691,n8025,n7942);
or (n8692,n8693,n8701);
and (n8693,n8694,n8699);
xor (n8694,n7957,n8695);
or (n8695,n8696,n8698);
and (n8696,n8697,n8040);
xor (n8697,n7971,n8038);
and (n8698,n7971,n8038);
xor (n8699,n8700,n8033);
xor (n8700,n8032,n8035);
and (n8701,n7957,n8695);
or (n8702,n8703,n8704);
xor (n8703,n8689,n8690);
and (n8704,n8700,n8033);
nand (n8705,n8706,n8685);
not (n8706,n8707);
nand (n8707,n8703,n8704);
nand (n8708,n8686,n8687);
nand (n8709,n8676,n8677);
and (n8710,n8652,n8655);
xor (n8711,n8243,n8486);
and (n8712,n8713,n8788);
xor (n8713,n8714,n8717);
and (n8714,n8715,n7785);
xnor (n8715,n8683,n8716);
nand (n8716,n8675,n8709);
or (n8717,n8718,n8787);
and (n8718,n8719,n8755);
xor (n8719,n8720,n8723);
wire s0n8720,s1n8720,notn8720;
or (n8720,s0n8720,s1n8720);
not(notn8720,n7786);
and (s0n8720,notn8720,1'b0);
and (s1n8720,n7786,n8721);
xor (n8721,n8722,n8588);
xor (n8722,n8583,n8585);
and (n8723,n8724,n8749);
or (n8724,n8725,n8748);
and (n8725,n8726,n8740);
xor (n8726,n8727,n8734);
and (n8727,n8728,n35);
nand (n8728,n8729,n8731,n8733);
or (n8729,n8730,n8440);
not (n8730,n8541);
or (n8731,n8584,n8732);
not (n8732,n8515);
not (n8733,n8500);
nor (n8734,n8050,n8735);
nor (n8735,n8286,n8736);
nor (n8736,n8737,n8353);
and (n8737,n8738,n8739);
not (n8738,n8288);
not (n8739,n8287);
nor (n8740,n8741,n8050);
nor (n8741,n8742,n8746);
and (n8742,n8743,n8263);
not (n8743,n8744);
xor (n8744,n8250,n8745);
not (n8745,n8274);
and (n8746,n8744,n8747);
not (n8747,n8263);
and (n8748,n8727,n8734);
and (n8749,n8750,n35);
nor (n8750,n8751,n8753);
and (n8751,n8752,n8409);
xor (n8752,n8440,n8451);
and (n8753,n8754,n8453);
not (n8754,n8752);
or (n8755,n8756,n8786);
and (n8756,n8757,n8783);
xor (n8757,n8758,n8761);
wire s0n8758,s1n8758,notn8758;
or (n8758,s0n8758,s1n8758);
not(notn8758,n8236);
and (s0n8758,notn8758,1'b0);
and (s1n8758,n8236,n8759);
xor (n8759,n8760,n8357);
xor (n8760,n8352,n8354);
xor (n8761,n8762,n8775);
xor (n8762,n8763,n8768);
and (n8763,n8764,n35);
nand (n8764,n8765,n8766,n8767);
or (n8765,n8462,n8739);
not (n8766,n8467);
or (n8767,n8250,n8745);
and (n8768,n8769,n35);
nand (n8769,n8770,n8774);
or (n8770,n8771,n8584);
and (n8771,n8772,n8773);
not (n8772,n8496);
not (n8773,n8497);
not (n8774,n8495);
and (n8775,n8776,n35);
nor (n8776,n8777,n8780);
and (n8777,n8778,n8407);
xor (n8778,n8779,n8462);
not (n8779,n8465);
and (n8780,n8781,n8782);
not (n8781,n8778);
not (n8782,n8407);
wire s0n8783,s1n8783,notn8783;
or (n8783,s0n8783,s1n8783);
not(notn8783,n7786);
and (s0n8783,notn8783,1'b0);
and (s1n8783,n7786,n8784);
xor (n8784,n8785,n8594);
xor (n8785,n8590,n8591);
and (n8786,n8758,n8761);
and (n8787,n8720,n8723);
wire s0n8788,s1n8788,notn8788;
or (n8788,s0n8788,s1n8788);
not(notn8788,n8048);
and (s0n8788,notn8788,1'b0);
and (s1n8788,n8048,n8789);
xor (n8789,n8790,n7997);
xor (n8790,n7992,n7995);
and (n8791,n8649,n8711);
xor (n8792,n8793,n8824);
xor (n8793,n8794,n8807);
xor (n8794,n8795,n8804);
xor (n8795,n8796,n8797);
wire s0n8796,s1n8796,notn8796;
or (n8796,s0n8796,s1n8796);
not(notn8796,n7785);
and (s0n8796,notn8796,1'b0);
and (s1n8796,n7785,n8789);
and (n8797,n8798,n8801);
or (n8798,n8799,n8800);
and (n8799,n8379,n8420);
and (n8800,n8380,n8408);
or (n8801,n8802,n8803);
and (n8802,n8381,n8406);
and (n8803,n8382,n8394);
wire s0n8804,s1n8804,notn8804;
or (n8804,s0n8804,s1n8804);
not(notn8804,n7786);
and (s0n8804,notn8804,1'b0);
and (s1n8804,n7786,n8805);
xor (n8805,n8806,n8641);
xor (n8806,n8638,n8639);
or (n8807,n8808,n8823);
and (n8808,n8809,n8822);
xor (n8809,n8810,n8821);
or (n8810,n8811,n8820);
and (n8811,n8812,n8819);
xor (n8812,n8813,n8814);
xor (n8813,n8245,n8458);
and (n8814,n8815,n8818);
xor (n8815,n8816,n8817);
wire s0n8816,s1n8816,notn8816;
or (n8816,s0n8816,s1n8816);
not(notn8816,n7785);
and (s0n8816,notn8816,1'b0);
and (s1n8816,n7785,n8759);
wire s0n8817,s1n8817,notn8817;
or (n8817,s0n8817,s1n8817);
not(notn8817,n8236);
and (s0n8817,notn8817,1'b0);
and (s1n8817,n8236,n8247);
wire s0n8818,s1n8818,notn8818;
or (n8818,s0n8818,s1n8818);
not(notn8818,n8048);
and (s0n8818,notn8818,1'b0);
and (s1n8818,n8048,n8459);
wire s0n8819,s1n8819,notn8819;
or (n8819,s0n8819,s1n8819);
not(notn8819,n679);
and (s0n8819,notn8819,1'b0);
and (s1n8819,n679,n8487);
and (n8820,n8813,n8814);
wire s0n8821,s1n8821,notn8821;
or (n8821,s0n8821,s1n8821);
not(notn8821,n7786);
and (s0n8821,notn8821,1'b0);
and (s1n8821,n7786,n8653);
wire s0n8822,s1n8822,notn8822;
or (n8822,s0n8822,s1n8822);
not(notn8822,n8236);
and (s0n8822,notn8822,1'b0);
and (s1n8822,n8236,n8789);
and (n8823,n8810,n8821);
or (n8824,n8825,n8836);
and (n8825,n8826,n8835);
xor (n8826,n8827,n8828);
wire s0n8827,s1n8827,notn8827;
or (n8827,s0n8827,s1n8827);
not(notn8827,n35);
and (s0n8827,notn8827,1'b0);
and (s1n8827,n35,n7857);
wire s0n8828,s1n8828,notn8828;
or (n8828,s0n8828,s1n8828);
not(notn8828,n35);
and (s0n8828,notn8828,1'b0);
and (s1n8828,n35,n8829);
xor (n8829,n8830,n8831);
wire s0n8830,s1n8830,notn8830;
or (n8830,s0n8830,s1n8830);
not(notn8830,n7737);
and (s0n8830,notn8830,1'b0);
and (s1n8830,n7737,n8067);
or (n8831,n8832,n8833,n8834);
and (n8832,n8054,n8077);
and (n8833,n8077,n8176);
and (n8834,n8054,n8176);
wire s0n8835,s1n8835,notn8835;
or (n8835,s0n8835,s1n8835);
not(notn8835,n8048);
and (s0n8835,notn8835,1'b0);
and (s1n8835,n8048,n8234);
and (n8836,n8827,n8828);
or (n8837,n8838,n9030);
and (n8838,n8839,n8880);
xor (n8839,n8840,n8841);
xor (n8840,n8648,n8712);
or (n8841,n8842,n8879);
and (n8842,n8843,n8852);
xor (n8843,n8844,n8845);
xor (n8844,n8713,n8788);
or (n8845,n8846,n8851);
and (n8846,n8847,n8850);
xor (n8847,n8848,n8849);
and (n8848,n8715,n8236);
xor (n8849,n8719,n8755);
wire s0n8850,s1n8850,notn8850;
or (n8850,s0n8850,s1n8850);
not(notn8850,n35);
and (s0n8850,notn8850,1'b0);
and (s1n8850,n35,n8653);
and (n8851,n8848,n8849);
or (n8852,n8853,n8878);
and (n8853,n8854,n8877);
xor (n8854,n8855,n8856);
wire s0n8855,s1n8855,notn8855;
or (n8855,s0n8855,s1n8855);
not(notn8855,n679);
and (s0n8855,notn8855,1'b0);
and (s1n8855,n679,n8656);
or (n8856,n8857,n8876);
and (n8857,n8858,n8873);
xor (n8858,n8859,n8864);
xor (n8859,n8860,n8861);
xor (n8860,n8724,n8749);
wire s0n8861,s1n8861,notn8861;
or (n8861,s0n8861,s1n8861);
not(notn8861,n7785);
and (s0n8861,notn8861,1'b0);
and (s1n8861,n7785,n8862);
xor (n8862,n8863,n8364);
xor (n8863,n8359,n8361);
and (n8864,n8865,n8870);
xor (n8865,n8866,n8867);
xor (n8866,n8726,n8740);
wire s0n8867,s1n8867,notn8867;
or (n8867,s0n8867,s1n8867);
not(notn8867,n7785);
and (s0n8867,notn8867,1'b0);
and (s1n8867,n7785,n8868);
xor (n8868,n8869,n8371);
xor (n8869,n8366,n8368);
wire s0n8870,s1n8870,notn8870;
or (n8870,s0n8870,s1n8870);
not(notn8870,n7786);
and (s0n8870,notn8870,1'b0);
and (s1n8870,n7786,n8871);
xor (n8871,n8872,n8601);
xor (n8872,n8596,n8598);
wire s0n8873,s1n8873,notn8873;
or (n8873,s0n8873,s1n8873);
not(notn8873,n7785);
and (s0n8873,notn8873,1'b0);
and (s1n8873,n7785,n8874);
xor (n8874,n8875,n8029);
xor (n8875,n8023,n8026);
and (n8876,n8859,n8864);
and (n8877,n8659,n8048);
and (n8878,n8855,n8856);
and (n8879,n8844,n8845);
or (n8880,n8881,n9029);
and (n8881,n8882,n9005);
xor (n8882,n8883,n9004);
or (n8883,n8884,n9003);
and (n8884,n8885,n9002);
xor (n8885,n8886,n8919);
or (n8886,n8887,n8918);
and (n8887,n8888,n8915);
xor (n8888,n8889,n8890);
xor (n8889,n8757,n8783);
or (n8890,n8891,n8914);
and (n8891,n8892,n8913);
xor (n8892,n8893,n8894);
wire s0n8893,s1n8893,notn8893;
or (n8893,s0n8893,s1n8893);
not(notn8893,n8048);
and (s0n8893,notn8893,1'b0);
and (s1n8893,n8048,n8759);
or (n8894,n8895,n8912);
and (n8895,n8896,n8911);
xor (n8896,n8897,n8907);
and (n8897,n8898,n35);
nand (n8898,n8899,n8905);
or (n8899,n8501,n8900);
not (n8900,n8901);
nand (n8901,n8902,n8904);
or (n8902,n8456,n8903);
not (n8903,n8590);
or (n8904,n8590,n8455);
or (n8905,n8901,n8906);
not (n8906,n8501);
and (n8907,n8908,n35);
nand (n8908,n8909,n8910);
or (n8909,n8353,n8355);
nand (n8910,n8355,n8353);
wire s0n8911,s1n8911,notn8911;
or (n8911,s0n8911,s1n8911);
not(notn8911,n8236);
and (s0n8911,notn8911,1'b0);
and (s1n8911,n8236,n8868);
and (n8912,n8897,n8907);
wire s0n8913,s1n8913,notn8913;
or (n8913,s0n8913,s1n8913);
not(notn8913,n679);
and (s0n8913,notn8913,1'b0);
and (s1n8913,n679,n8784);
and (n8914,n8893,n8894);
wire s0n8915,s1n8915,notn8915;
or (n8915,s0n8915,s1n8915);
not(notn8915,n7786);
and (s0n8915,notn8915,1'b0);
and (s1n8915,n7786,n8916);
xor (n8916,n8917,n8207);
xor (n8917,n8201,n8204);
and (n8918,n8889,n8890);
or (n8919,n8920,n9001);
and (n8920,n8921,n8998);
xor (n8921,n8922,n8946);
xor (n8922,n8923,n8945);
xor (n8923,n8924,n8925);
wire s0n8924,s1n8924,notn8924;
or (n8924,s0n8924,s1n8924);
not(notn8924,n8048);
and (s0n8924,notn8924,1'b0);
and (s1n8924,n8048,n8247);
or (n8925,n8926,n8944);
and (n8926,n8927,n8943);
xor (n8927,n8928,n8941);
or (n8928,n8929,n8936);
and (n8929,n8930,n35);
nand (n8930,n8931,n8933,n8935);
or (n8931,n8250,n8932);
not (n8932,n8333);
or (n8933,n8353,n8934);
not (n8934,n8307);
not (n8935,n8291);
and (n8936,n8937,n35);
or (n8937,n8938,n8514);
nor (n8938,n8939,n8597);
and (n8939,n8940,n8732);
not (n8940,n8526);
nor (n8941,n8942,n8050);
xor (n8942,n8586,n8584);
wire s0n8943,s1n8943,notn8943;
or (n8943,s0n8943,s1n8943);
not(notn8943,n8236);
and (s0n8943,notn8943,1'b0);
and (s1n8943,n8236,n8862);
and (n8944,n8928,n8941);
wire s0n8945,s1n8945,notn8945;
or (n8945,s0n8945,s1n8945);
not(notn8945,n679);
and (s0n8945,notn8945,1'b0);
and (s1n8945,n679,n8721);
and (n8946,n8947,n8997);
xor (n8947,n8948,n8991);
or (n8948,n8949,n8990);
and (n8949,n8950,n8987);
xor (n8950,n8951,n8965);
and (n8951,n8952,n8963);
xor (n8952,n8953,n8961);
and (n8953,n8954,n8958);
nor (n8954,n8955,n8597);
not (n8955,n8956);
wire s0n8956,s1n8956,notn8956;
or (n8956,s0n8956,s1n8956);
not(notn8956,n35);
and (s0n8956,notn8956,1'b0);
and (s1n8956,n35,n8957);
wire s0n8957,s1n8957,notn8957;
or (n8957,s0n8957,s1n8957);
not(notn8957,n753);
and (s0n8957,notn8957,1'b0);
and (s1n8957,n753,n8560);
and (n8958,n8959,n35);
nor (n8959,n8960,n8932);
not (n8960,n8372);
wire s0n8961,s1n8961,notn8961;
or (n8961,s0n8961,s1n8961);
not(notn8961,n7785);
and (s0n8961,notn8961,1'b0);
and (s1n8961,n7785,n8962);
xor (n8962,n8336,n8347);
and (n8963,n8964,n35);
xnor (n8964,n8597,n8599);
or (n8965,n8966,n8986);
and (n8966,n8967,n8981);
xor (n8967,n8968,n8974);
and (n8968,n8969,n35);
nand (n8969,n8970,n8971,n8973);
or (n8970,n8367,n8934);
or (n8971,n8353,n8972);
not (n8972,n8347);
not (n8973,n8306);
and (n8974,n8975,n35);
not (n8975,n8976);
nor (n8976,n8977,n8978);
and (n8977,n8596,n8545);
nor (n8978,n8979,n8730);
and (n8979,n8604,n8980);
not (n8980,n8530);
and (n8981,n8982,n35);
xor (n8982,n8983,n8984);
not (n8983,n8292);
xnor (n8984,n8360,n8985);
not (n8985,n8303);
and (n8986,n8968,n8974);
wire s0n8987,s1n8987,notn8987;
or (n8987,s0n8987,s1n8987);
not(notn8987,n7786);
and (s0n8987,notn8987,1'b0);
and (s1n8987,n7786,n8988);
xor (n8988,n8989,n8608);
xor (n8989,n8603,n8605);
and (n8990,n8951,n8965);
and (n8991,n8992,n8996);
xor (n8992,n8993,n8994);
wire s0n8993,s1n8993,notn8993;
or (n8993,s0n8993,s1n8993);
not(notn8993,n679);
and (s0n8993,notn8993,1'b0);
and (s1n8993,n679,n8871);
wire s0n8994,s1n8994,notn8994;
or (n8994,s0n8994,s1n8994);
not(notn8994,n7785);
and (s0n8994,notn8994,1'b0);
and (s1n8994,n7785,n8995);
xor (n8995,n8372,n8373);
wire s0n8996,s1n8996,notn8996;
or (n8996,s0n8996,s1n8996);
not(notn8996,n8048);
and (s0n8996,notn8996,1'b0);
and (s1n8996,n8048,n8862);
xor (n8997,n8865,n8870);
wire s0n8998,s1n8998,notn8998;
or (n8998,s0n8998,s1n8998);
not(notn8998,n8236);
and (s0n8998,notn8998,1'b0);
and (s1n8998,n8236,n8999);
xor (n8999,n9000,n8021);
xor (n9000,n8015,n8018);
and (n9001,n8922,n8946);
wire s0n9002,s1n9002,notn9002;
or (n9002,s0n9002,s1n9002);
not(notn9002,n35);
and (s0n9002,notn9002,1'b0);
and (s1n9002,n35,n8789);
and (n9003,n8886,n8919);
xor (n9004,n8651,n8658);
xor (n9005,n9006,n9028);
xor (n9006,n9007,n9008);
wire s0n9007,s1n9007,notn9007;
or (n9007,s0n9007,s1n9007);
not(notn9007,n35);
and (s0n9007,notn9007,1'b0);
and (s1n9007,n35,n8052);
xor (n9008,n9009,n9025);
xor (n9009,n9010,n9011);
wire s0n9010,s1n9010,notn9010;
or (n9010,s0n9010,s1n9010);
not(notn9010,n8048);
and (s0n9010,notn9010,1'b0);
and (s1n9010,n8048,n8475);
or (n9011,n9012,n9024);
and (n9012,n9013,n9021);
xor (n9013,n9014,n9015);
xor (n9014,n8422,n8436);
and (n9015,n9016,n35);
nand (n9016,n9017,n9019);
or (n9017,n9018,n8782);
and (n9018,n8779,n8462);
or (n9019,n8738,n9020);
not (n9020,n8395);
or (n9021,n9022,n9023);
and (n9022,n8762,n8775);
and (n9023,n8763,n8768);
and (n9024,n9014,n9015);
wire s0n9025,s1n9025,notn9025;
or (n9025,s0n9025,s1n9025);
not(notn9025,n7786);
and (s0n9025,notn9025,1'b0);
and (s1n9025,n7786,n9026);
xor (n9026,n9027,n8581);
xor (n9027,n8577,n8578);
wire s0n9028,s1n9028,notn9028;
or (n9028,s0n9028,s1n9028);
not(notn9028,n35);
and (s0n9028,notn9028,1'b0);
and (s1n9028,n35,n8234);
and (n9029,n8883,n9004);
and (n9030,n8840,n8841);
and (n9031,n7852,n8792);
xor (n9032,n9033,n9056);
xor (n9033,n9034,n9037);
or (n9034,n9035,n9036);
and (n9035,n8793,n8824);
and (n9036,n8794,n8807);
and (n9037,n9038,n9049);
xor (n9038,n9039,n9048);
or (n9039,n9040,n9047);
and (n9040,n9041,n9046);
xor (n9041,n9042,n9043);
wire s0n9042,s1n9042,notn9042;
or (n9042,s0n9042,s1n9042);
not(notn9042,n8048);
and (s0n9042,notn9042,1'b0);
and (s1n9042,n8048,n8633);
xor (n9043,n9044,n9045);
xor (n9044,n8798,n8801);
wire s0n9045,s1n9045,notn9045;
or (n9045,s0n9045,s1n9045);
not(notn9045,n7785);
and (s0n9045,notn9045,1'b0);
and (s1n9045,n7785,n8459);
wire s0n9046,s1n9046,notn9046;
or (n9046,s0n9046,s1n9046);
not(notn9046,n679);
and (s0n9046,notn9046,1'b0);
and (s1n9046,n679,n8052);
and (n9047,n9042,n9043);
wire s0n9048,s1n9048,notn9048;
or (n9048,s0n9048,s1n9048);
not(notn9048,n679);
and (s0n9048,notn9048,1'b0);
and (s1n9048,n679,n8829);
and (n9049,n9050,n9055);
xor (n9050,n9051,n9052);
and (n9051,n8659,n7785);
or (n9052,n9053,n9054);
and (n9053,n9009,n9025);
and (n9054,n9010,n9011);
wire s0n9055,s1n9055,notn9055;
or (n9055,s0n9055,s1n9055);
not(notn9055,n679);
and (s0n9055,notn9055,1'b0);
and (s1n9055,n679,n8805);
xor (n9056,n9057,n9060);
xor (n9057,n9058,n9059);
and (n9058,n8795,n8804);
and (n9059,n8620,n8632);
or (n9060,n9061,n9062);
and (n9061,n7855,n8233);
and (n9062,n7856,n8051);
xor (n9063,n9064,n9083);
xor (n9064,n9065,n9068);
or (n9065,n9066,n9067);
and (n9066,n7853,n8646);
and (n9067,n7854,n8239);
xor (n9068,n9069,n9078);
xor (n9069,n9070,n9073);
or (n9070,n9071,n9072);
and (n9071,n8240,n8635);
and (n9072,n8241,n8619);
xor (n9073,n9074,n9077);
xor (n9074,n9075,n9076);
wire s0n9075,s1n9075,notn9075;
or (n9075,s0n9075,s1n9075);
not(notn9075,n7785);
and (s0n9075,notn9075,1'b0);
and (s1n9075,n7785,n8633);
wire s0n9076,s1n9076,notn9076;
or (n9076,s0n9076,s1n9076);
not(notn9076,n8236);
and (s0n9076,notn9076,1'b0);
and (s1n9076,n8236,n8622);
wire s0n9077,s1n9077,notn9077;
or (n9077,s0n9077,s1n9077);
not(notn9077,n7785);
and (s0n9077,notn9077,1'b0);
and (s1n9077,n7785,n8234);
xor (n9078,n9079,n9082);
xor (n9079,n9080,n9081);
wire s0n9080,s1n9080,notn9080;
or (n9080,s0n9080,s1n9080);
not(notn9080,n7786);
and (s0n9080,notn9080,1'b0);
and (s1n9080,n7786,n8829);
wire s0n9081,s1n9081,notn9081;
or (n9081,s0n9081,s1n9081);
not(notn9081,n7786);
and (s0n9081,notn9081,1'b0);
and (s1n9081,n7786,n8636);
wire s0n9082,s1n9082,notn9082;
or (n9082,s0n9082,s1n9082);
not(notn9082,n8236);
and (s0n9082,notn9082,1'b0);
and (s1n9082,n8236,n7857);
or (n9083,n9084,n9125);
and (n9084,n9085,n9096);
xor (n9085,n9086,n9095);
or (n9086,n9087,n9094);
and (n9087,n9088,n9091);
xor (n9088,n9089,n9090);
xor (n9089,n8809,n8822);
xor (n9090,n9041,n9046);
or (n9091,n9092,n9093);
and (n9092,n9006,n9028);
and (n9093,n9007,n9008);
and (n9094,n9089,n9090);
xor (n9095,n9038,n9049);
or (n9096,n9097,n9124);
and (n9097,n9098,n9123);
xor (n9098,n9099,n9100);
xor (n9099,n9050,n9055);
or (n9100,n9101,n9122);
and (n9101,n9102,n9113);
xor (n9102,n9103,n9104);
xor (n9103,n8812,n8819);
or (n9104,n9105,n9112);
and (n9105,n9106,n9111);
xor (n9106,n9107,n9110);
or (n9107,n9108,n9109);
and (n9108,n8923,n8945);
and (n9109,n8924,n8925);
xor (n9110,n9013,n9021);
wire s0n9111,s1n9111,notn9111;
or (n9111,s0n9111,s1n9111);
not(notn9111,n679);
and (s0n9111,notn9111,1'b0);
and (s1n9111,n679,n9026);
and (n9112,n9107,n9110);
or (n9113,n9114,n9121);
and (n9114,n9115,n9118);
xor (n9115,n9116,n9117);
wire s0n9116,s1n9116,notn9116;
or (n9116,s0n9116,s1n9116);
not(notn9116,n7785);
and (s0n9116,notn9116,1'b0);
and (s1n9116,n7785,n8999);
xor (n9117,n8815,n8818);
wire s0n9118,s1n9118,notn9118;
or (n9118,s0n9118,s1n9118);
not(notn9118,n7786);
and (s0n9118,notn9118,1'b0);
and (s1n9118,n7786,n9119);
xor (n9119,n9120,n8199);
xor (n9120,n8193,n8196);
and (n9121,n9116,n9117);
and (n9122,n9103,n9104);
xor (n9123,n8826,n8835);
and (n9124,n9099,n9100);
and (n9125,n9086,n9095);
or (n9126,n9127,n9198);
and (n9127,n9128,n9197);
xor (n9128,n9129,n9130);
xor (n9129,n9085,n9096);
or (n9130,n9131,n9196);
and (n9131,n9132,n9135);
xor (n9132,n9133,n9134);
xor (n9133,n9098,n9123);
xor (n9134,n9088,n9091);
or (n9135,n9136,n9195);
and (n9136,n9137,n9182);
xor (n9137,n9138,n9181);
or (n9138,n9139,n9180);
and (n9139,n9140,n9143);
xor (n9140,n9141,n9142);
xor (n9141,n9115,n9118);
xor (n9142,n9106,n9111);
or (n9143,n9144,n9179);
and (n9144,n9145,n9178);
xor (n9145,n9146,n9169);
or (n9146,n9147,n9168);
and (n9147,n9148,n9167);
xor (n9148,n9149,n9150);
xor (n9149,n8892,n8913);
or (n9150,n9151,n9166);
and (n9151,n9152,n9158);
xor (n9152,n9153,n9154);
xor (n9153,n8896,n8911);
nand (n9154,n9155,n8928);
or (n9155,n9156,n9157);
not (n9156,n8936);
not (n9157,n8929);
or (n9158,n9159,n9165);
and (n9159,n9160,n9164);
xor (n9160,n9161,n9162);
wire s0n9161,s1n9161,notn9161;
or (n9161,s0n9161,s1n9161);
not(notn9161,n8236);
and (s0n9161,notn9161,1'b0);
and (s1n9161,n8236,n8995);
wire s0n9162,s1n9162,notn9162;
or (n9162,s0n9162,s1n9162);
not(notn9162,n7786);
and (s0n9162,notn9162,1'b0);
and (s1n9162,n7786,n9163);
xor (n9163,n8609,n8611);
wire s0n9164,s1n9164,notn9164;
or (n9164,s0n9164,s1n9164);
not(notn9164,n8048);
and (s0n9164,notn9164,1'b0);
and (s1n9164,n8048,n8868);
and (n9165,n9161,n9162);
and (n9166,n9153,n9154);
wire s0n9167,s1n9167,notn9167;
or (n9167,s0n9167,s1n9167);
not(notn9167,n8236);
and (s0n9167,notn9167,1'b0);
and (s1n9167,n8236,n8874);
and (n9168,n9149,n9150);
and (n9169,n9170,n9175);
xor (n9170,n9171,n9174);
wire s0n9171,s1n9171,notn9171;
or (n9171,s0n9171,s1n9171);
not(notn9171,n7785);
and (s0n9171,notn9171,1'b0);
and (s1n9171,n7785,n9172);
xor (n9172,n9173,n8037);
xor (n9173,n8031,n8034);
xor (n9174,n8927,n8943);
wire s0n9175,s1n9175,notn9175;
or (n9175,s0n9175,s1n9175);
not(notn9175,n7786);
and (s0n9175,notn9175,1'b0);
and (s1n9175,n7786,n9176);
xor (n9176,n9177,n8215);
xor (n9177,n8209,n8212);
wire s0n9178,s1n9178,notn9178;
or (n9178,s0n9178,s1n9178);
not(notn9178,n35);
and (s0n9178,notn9178,1'b0);
and (s1n9178,n35,n8656);
and (n9179,n9146,n9169);
and (n9180,n9141,n9142);
xor (n9181,n9102,n9113);
or (n9182,n9183,n9194);
and (n9183,n9184,n9193);
xor (n9184,n9185,n9186);
xor (n9185,n8847,n8850);
or (n9186,n9187,n9192);
and (n9187,n9188,n9191);
xor (n9188,n9189,n9190);
and (n9189,n8715,n8048);
wire s0n9190,s1n9190,notn9190;
or (n9190,s0n9190,s1n9190);
not(notn9190,n679);
and (s0n9190,notn9190,1'b0);
and (s1n9190,n679,n9119);
and (n9191,n8659,n35);
and (n9192,n9189,n9190);
xor (n9193,n8854,n8877);
and (n9194,n9185,n9186);
and (n9195,n9138,n9181);
and (n9196,n9133,n9134);
xor (n9197,n7851,n8837);
and (n9198,n9129,n9130);
or (n9199,n9200,n9673);
and (n9200,n9201,n9278);
xor (n9201,n9202,n9203);
xor (n9202,n9128,n9197);
or (n9203,n9204,n9277);
and (n9204,n9205,n9276);
xor (n9205,n9206,n9207);
xor (n9206,n8839,n8880);
or (n9207,n9208,n9275);
and (n9208,n9209,n9212);
xor (n9209,n9210,n9211);
xor (n9210,n8843,n8852);
xor (n9211,n8882,n9005);
or (n9212,n9213,n9274);
and (n9213,n9214,n9253);
xor (n9214,n9215,n9216);
xor (n9215,n8885,n9002);
or (n9216,n9217,n9252);
and (n9217,n9218,n9221);
xor (n9218,n9219,n9220);
xor (n9219,n8888,n8915);
xor (n9220,n8858,n8873);
or (n9221,n9222,n9251);
and (n9222,n9223,n9250);
xor (n9223,n9224,n9249);
and (n9224,n9225,n9226);
xor (n9225,n8950,n8987);
or (n9226,n9227,n9248);
and (n9227,n9228,n9247);
xor (n9228,n9229,n9246);
or (n9229,n9230,n9245);
and (n9230,n9231,n9238);
xor (n9231,n9232,n9234);
wire s0n9232,s1n9232,notn9232;
or (n9232,s0n9232,s1n9232);
not(notn9232,n7786);
and (s0n9232,notn9232,1'b0);
and (s1n9232,n7786,n9233);
xor (n9233,n8559,n8570);
and (n9234,n9235,n9236);
wire s0n9235,s1n9235,notn9235;
or (n9235,s0n9235,s1n9235);
not(notn9235,n7786);
and (s0n9235,notn9235,1'b0);
and (s1n9235,n7786,n8957);
wire s0n9236,s1n9236,notn9236;
or (n9236,s0n9236,s1n9236);
not(notn9236,n7786);
and (s0n9236,notn9236,1'b0);
and (s1n9236,n7786,n9237);
wire s0n9237,s1n9237,notn9237;
or (n9237,s0n9237,s1n9237);
not(notn9237,n753);
and (s0n9237,notn9237,1'b0);
and (s1n9237,n753,n8161);
and (n9238,n9239,n35);
nand (n9239,n9240,n9244);
or (n9240,n8980,n9241);
nand (n9241,n9242,n9243);
or (n9242,n8541,n8604);
nand (n9243,n8541,n8604);
nand (n9244,n9241,n8980);
and (n9245,n9232,n9234);
xor (n9246,n8967,n8981);
wire s0n9247,s1n9247,notn9247;
or (n9247,s0n9247,s1n9247);
not(notn9247,n679);
and (s0n9247,notn9247,1'b0);
and (s1n9247,n679,n8988);
and (n9248,n9229,n9246);
wire s0n9249,s1n9249,notn9249;
or (n9249,s0n9249,s1n9249);
not(notn9249,n8048);
and (s0n9249,notn9249,1'b0);
and (s1n9249,n8048,n8999);
wire s0n9250,s1n9250,notn9250;
or (n9250,s0n9250,s1n9250);
not(notn9250,n679);
and (s0n9250,notn9250,1'b0);
and (s1n9250,n679,n8916);
and (n9251,n9224,n9249);
and (n9252,n9219,n9220);
or (n9253,n9254,n9273);
and (n9254,n9255,n9272);
xor (n9255,n9256,n9257);
xor (n9256,n8921,n8998);
or (n9257,n9258,n9271);
and (n9258,n9259,n9270);
xor (n9259,n9260,n9269);
or (n9260,n9261,n9268);
and (n9261,n9262,n9267);
xor (n9262,n9263,n9264);
xor (n9263,n8992,n8996);
wire s0n9264,s1n9264,notn9264;
or (n9264,s0n9264,s1n9264);
not(notn9264,n7786);
and (s0n9264,notn9264,1'b0);
and (s1n9264,n7786,n9265);
xor (n9265,n9266,n8223);
xor (n9266,n8217,n8220);
wire s0n9267,s1n9267,notn9267;
or (n9267,s0n9267,s1n9267);
not(notn9267,n8236);
and (s0n9267,notn9267,1'b0);
and (s1n9267,n8236,n9172);
and (n9268,n9263,n9264);
xor (n9269,n8947,n8997);
and (n9270,n8715,n35);
and (n9271,n9260,n9269);
xor (n9272,n9188,n9191);
and (n9273,n9256,n9257);
and (n9274,n9215,n9216);
and (n9275,n9210,n9211);
xor (n9276,n9132,n9135);
and (n9277,n9206,n9207);
or (n9278,n9279,n9672);
and (n9279,n9280,n9410);
xor (n9280,n9281,n9282);
xor (n9281,n9205,n9276);
or (n9282,n9283,n9409);
and (n9283,n9284,n9408);
xor (n9284,n9285,n9286);
xor (n9285,n9137,n9182);
or (n9286,n9287,n9407);
and (n9287,n9288,n9406);
xor (n9288,n9289,n9290);
xor (n9289,n9140,n9143);
or (n9290,n9291,n9405);
and (n9291,n9292,n9337);
xor (n9292,n9293,n9336);
or (n9293,n9294,n9335);
and (n9294,n9295,n9298);
xor (n9295,n9296,n9297);
xor (n9296,n9170,n9175);
wire s0n9297,s1n9297,notn9297;
or (n9297,s0n9297,s1n9297);
not(notn9297,n35);
and (s0n9297,notn9297,1'b0);
and (s1n9297,n35,n9119);
or (n9298,n9299,n9334);
and (n9299,n9300,n9333);
xor (n9300,n9301,n9315);
or (n9301,n9302,n9314);
and (n9302,n9303,n9312);
xor (n9303,n9304,n9306);
wire s0n9304,s1n9304,notn9304;
or (n9304,s0n9304,s1n9304);
not(notn9304,n7786);
and (s0n9304,notn9304,1'b0);
and (s1n9304,n7786,n9305);
xor (n9305,n8224,n8225);
and (n9306,n9307,n9311);
xor (n9307,n9308,n9309);
xor (n9308,n8954,n8958);
wire s0n9309,s1n9309,notn9309;
or (n9309,s0n9309,s1n9309);
not(notn9309,n7785);
and (s0n9309,notn9309,1'b0);
and (s1n9309,n7785,n9310);
wire s0n9310,s1n9310,notn9310;
or (n9310,s0n9310,s1n9310);
not(notn9310,n753);
and (s0n9310,notn9310,1'b0);
and (s1n9310,n753,n8337);
wire s0n9311,s1n9311,notn9311;
or (n9311,s0n9311,s1n9311);
not(notn9311,n679);
and (s0n9311,notn9311,1'b0);
and (s1n9311,n679,n9163);
wire s0n9312,s1n9312,notn9312;
or (n9312,s0n9312,s1n9312);
not(notn9312,n8236);
and (s0n9312,notn9312,1'b0);
and (s1n9312,n8236,n9313);
xor (n9313,n8038,n8039);
and (n9314,n9304,n9306);
or (n9315,n9316,n9332);
and (n9316,n9317,n9330);
xor (n9317,n9318,n9319);
xor (n9318,n8952,n8963);
and (n9319,n9320,n9329);
xor (n9320,n9321,n9327);
and (n9321,n9322,n35);
xnor (n9322,n9323,n8934);
nand (n9323,n9324,n9326);
or (n9324,n8366,n9325);
not (n9325,n8318);
nand (n9326,n8366,n9325);
wire s0n9327,s1n9327,notn9327;
or (n9327,s0n9327,s1n9327);
not(notn9327,n7785);
and (s0n9327,notn9327,1'b0);
and (s1n9327,n7785,n9328);
wire s0n9328,s1n9328,notn9328;
or (n9328,s0n9328,s1n9328);
not(notn9328,n753);
and (s0n9328,notn9328,1'b0);
and (s1n9328,n753,n7973);
wire s0n9329,s1n9329,notn9329;
or (n9329,s0n9329,s1n9329);
not(notn9329,n8236);
and (s0n9329,notn9329,1'b0);
and (s1n9329,n8236,n8962);
wire s0n9330,s1n9330,notn9330;
or (n9330,s0n9330,s1n9330);
not(notn9330,n7785);
and (s0n9330,notn9330,1'b0);
and (s1n9330,n7785,n9331);
xor (n9331,n7972,n7984);
and (n9332,n9318,n9319);
wire s0n9333,s1n9333,notn9333;
or (n9333,s0n9333,s1n9333);
not(notn9333,n8048);
and (s0n9333,notn9333,1'b0);
and (s1n9333,n8048,n8874);
and (n9334,n9301,n9315);
and (n9335,n9296,n9297);
xor (n9336,n9145,n9178);
or (n9337,n9338,n9404);
and (n9338,n9339,n9403);
xor (n9339,n9340,n9402);
or (n9340,n9341,n9401);
and (n9341,n9342,n9400);
xor (n9342,n9343,n9344);
xor (n9343,n9152,n9158);
or (n9344,n9345,n9399);
and (n9345,n9346,n9374);
xor (n9346,n9347,n9348);
xor (n9347,n9160,n9164);
or (n9348,n9349,n9373);
and (n9349,n9350,n9372);
xor (n9350,n9351,n9361);
or (n9351,n9352,n9360);
and (n9352,n9353,n9356);
xor (n9353,n9354,n9355);
wire s0n9354,s1n9354,notn9354;
or (n9354,s0n9354,s1n9354);
not(notn9354,n679);
and (s0n9354,notn9354,1'b0);
and (s1n9354,n679,n9233);
xor (n9355,n9235,n9236);
and (n9356,n9357,n35);
nand (n9357,n9358,n9359);
or (n9358,n8333,n8960);
or (n9359,n8372,n8932);
and (n9360,n9354,n9355);
or (n9361,n9362,n9371);
and (n9362,n9363,n9366);
xor (n9363,n9364,n9365);
and (n9364,n8322,n35);
and (n9365,n8545,n35);
and (n9366,n9367,n35);
nand (n9367,n9368,n9370);
or (n9368,n8609,n9369);
not (n9369,n8556);
nand (n9370,n8609,n9369);
and (n9371,n9364,n9365);
wire s0n9372,s1n9372,notn9372;
or (n9372,s0n9372,s1n9372);
not(notn9372,n8048);
and (s0n9372,notn9372,1'b0);
and (s1n9372,n8048,n8995);
and (n9373,n9351,n9361);
or (n9374,n9375,n9398);
and (n9375,n9376,n9396);
xor (n9376,n9377,n9378);
xor (n9377,n9231,n9238);
or (n9378,n9379,n9395);
and (n9379,n9380,n9394);
xor (n9380,n9381,n9389);
or (n9381,n9382,n9388);
and (n9382,n9383,n9386);
xor (n9383,n9384,n9385);
nor (n9384,n8972,n8050);
wire s0n9385,s1n9385,notn9385;
or (n9385,s0n9385,s1n9385);
not(notn9385,n679);
and (s0n9385,notn9385,1'b0);
and (s1n9385,n679,n8957);
nor (n9386,n9387,n8050);
not (n9387,n8570);
and (n9388,n9384,n9385);
and (n9389,n9390,n9392);
nor (n9390,n9391,n8050);
not (n9391,n8336);
nor (n9392,n9393,n8050);
not (n9393,n8559);
wire s0n9394,s1n9394,notn9394;
or (n9394,s0n9394,s1n9394);
not(notn9394,n8236);
and (s0n9394,notn9394,1'b0);
and (s1n9394,n8236,n9328);
and (n9395,n9381,n9389);
wire s0n9396,s1n9396,notn9396;
or (n9396,s0n9396,s1n9396);
not(notn9396,n7786);
and (s0n9396,notn9396,1'b0);
and (s1n9396,n7786,n9397);
xor (n9397,n8160,n8171);
and (n9398,n9377,n9378);
and (n9399,n9347,n9348);
wire s0n9400,s1n9400,notn9400;
or (n9400,s0n9400,s1n9400);
not(notn9400,n679);
and (s0n9400,notn9400,1'b0);
and (s1n9400,n679,n9176);
and (n9401,n9343,n9344);
xor (n9402,n9148,n9167);
xor (n9403,n9223,n9250);
and (n9404,n9340,n9402);
and (n9405,n9293,n9336);
xor (n9406,n9184,n9193);
and (n9407,n9289,n9290);
xor (n9408,n9209,n9212);
and (n9409,n9285,n9286);
or (n9410,n9411,n9671);
and (n9411,n9412,n9471);
xor (n9412,n9413,n9414);
xor (n9413,n9284,n9408);
or (n9414,n9415,n9470);
and (n9415,n9416,n9469);
xor (n9416,n9417,n9418);
xor (n9417,n9214,n9253);
or (n9418,n9419,n9468);
and (n9419,n9420,n9467);
xor (n9420,n9421,n9422);
xor (n9421,n9218,n9221);
or (n9422,n9423,n9466);
and (n9423,n9424,n9465);
xor (n9424,n9425,n9434);
or (n9425,n9426,n9433);
and (n9426,n9427,n9432);
xor (n9427,n9428,n9431);
xor (n9428,n9429,n9430);
xor (n9429,n9225,n9226);
wire s0n9430,s1n9430,notn9430;
or (n9430,s0n9430,s1n9430);
not(notn9430,n7785);
and (s0n9430,notn9430,1'b0);
and (s1n9430,n7785,n9313);
wire s0n9431,s1n9431,notn9431;
or (n9431,s0n9431,s1n9431);
not(notn9431,n35);
and (s0n9431,notn9431,1'b0);
and (s1n9431,n35,n8999);
wire s0n9432,s1n9432,notn9432;
or (n9432,s0n9432,s1n9432);
not(notn9432,n35);
and (s0n9432,notn9432,1'b0);
and (s1n9432,n35,n8916);
and (n9433,n9428,n9431);
or (n9434,n9435,n9464);
and (n9435,n9436,n9457);
xor (n9436,n9437,n9456);
or (n9437,n9438,n9455);
and (n9438,n9439,n9454);
xor (n9439,n9440,n9441);
xor (n9440,n9317,n9330);
or (n9441,n9442,n9453);
and (n9442,n9443,n9452);
xor (n9443,n9444,n9445);
wire s0n9444,s1n9444,notn9444;
or (n9444,s0n9444,s1n9444);
not(notn9444,n8236);
and (s0n9444,notn9444,1'b0);
and (s1n9444,n8236,n9331);
or (n9445,n9446,n9451);
and (n9446,n9447,n9450);
xor (n9447,n9448,n9449);
xor (n9448,n9363,n9366);
wire s0n9449,s1n9449,notn9449;
or (n9449,s0n9449,s1n9449);
not(notn9449,n8048);
and (s0n9449,notn9449,1'b0);
and (s1n9449,n8048,n8962);
wire s0n9450,s1n9450,notn9450;
or (n9450,s0n9450,s1n9450);
not(notn9450,n8236);
and (s0n9450,notn9450,1'b0);
and (s1n9450,n8236,n9310);
and (n9451,n9448,n9449);
xor (n9452,n9307,n9311);
and (n9453,n9444,n9445);
wire s0n9454,s1n9454,notn9454;
or (n9454,s0n9454,s1n9454);
not(notn9454,n8048);
and (s0n9454,notn9454,1'b0);
and (s1n9454,n8048,n9172);
and (n9455,n9440,n9441);
xor (n9456,n9262,n9267);
or (n9457,n9458,n9463);
and (n9458,n9459,n9462);
xor (n9459,n9460,n9461);
wire s0n9460,s1n9460,notn9460;
or (n9460,s0n9460,s1n9460);
not(notn9460,n679);
and (s0n9460,notn9460,1'b0);
and (s1n9460,n679,n9265);
xor (n9461,n9228,n9247);
wire s0n9462,s1n9462,notn9462;
or (n9462,s0n9462,s1n9462);
not(notn9462,n35);
and (s0n9462,notn9462,1'b0);
and (s1n9462,n35,n8874);
and (n9463,n9460,n9461);
and (n9464,n9437,n9456);
xor (n9465,n9259,n9270);
and (n9466,n9425,n9434);
xor (n9467,n9255,n9272);
and (n9468,n9421,n9422);
xor (n9469,n9288,n9406);
and (n9470,n9417,n9418);
or (n9471,n9472,n9670);
and (n9472,n9473,n9506);
xor (n9473,n9474,n9505);
or (n9474,n9475,n9504);
and (n9475,n9476,n9503);
xor (n9476,n9477,n9502);
or (n9477,n9478,n9501);
and (n9478,n9479,n9500);
xor (n9479,n9480,n9499);
or (n9480,n9481,n9498);
and (n9481,n9482,n9485);
xor (n9482,n9483,n9484);
xor (n9483,n9300,n9333);
xor (n9484,n9342,n9400);
or (n9485,n9486,n9497);
and (n9486,n9487,n9496);
xor (n9487,n9488,n9489);
xor (n9488,n9303,n9312);
or (n9489,n9490,n9495);
and (n9490,n9491,n9494);
xor (n9491,n9492,n9493);
xor (n9492,n9320,n9329);
wire s0n9493,s1n9493,notn9493;
or (n9493,s0n9493,s1n9493);
not(notn9493,n679);
and (s0n9493,notn9493,1'b0);
and (s1n9493,n679,n9305);
wire s0n9494,s1n9494,notn9494;
or (n9494,s0n9494,s1n9494);
not(notn9494,n8048);
and (s0n9494,notn9494,1'b0);
and (s1n9494,n8048,n9313);
and (n9495,n9492,n9493);
wire s0n9496,s1n9496,notn9496;
or (n9496,s0n9496,s1n9496);
not(notn9496,n35);
and (s0n9496,notn9496,1'b0);
and (s1n9496,n35,n9176);
and (n9497,n9488,n9489);
and (n9498,n9483,n9484);
xor (n9499,n9295,n9298);
xor (n9500,n9339,n9403);
and (n9501,n9480,n9499);
xor (n9502,n9292,n9337);
xor (n9503,n9420,n9467);
and (n9504,n9477,n9502);
xor (n9505,n9416,n9469);
or (n9506,n9507,n9669);
and (n9507,n9508,n9573);
xor (n9508,n9509,n9572);
or (n9509,n9510,n9571);
and (n9510,n9511,n9570);
xor (n9511,n9512,n9569);
or (n9512,n9513,n9568);
and (n9513,n9514,n9561);
xor (n9514,n9515,n9560);
or (n9515,n9516,n9559);
and (n9516,n9517,n9540);
xor (n9517,n9518,n9539);
or (n9518,n9519,n9538);
and (n9519,n9520,n9537);
xor (n9520,n9521,n9536);
or (n9521,n9522,n9535);
and (n9522,n9523,n9534);
xor (n9523,n9524,n9525);
xor (n9524,n9353,n9356);
or (n9525,n9526,n9533);
and (n9526,n9527,n9532);
xor (n9527,n9528,n9531);
and (n9528,n9529,n9530);
wire s0n9529,s1n9529,notn9529;
or (n9529,s0n9529,s1n9529);
not(notn9529,n35);
and (s0n9529,notn9529,1'b0);
and (s1n9529,n35,n9310);
wire s0n9530,s1n9530,notn9530;
or (n9530,s0n9530,s1n9530);
not(notn9530,n35);
and (s0n9530,notn9530,1'b0);
and (s1n9530,n35,n9237);
wire s0n9531,s1n9531,notn9531;
or (n9531,s0n9531,s1n9531);
not(notn9531,n679);
and (s0n9531,notn9531,1'b0);
and (s1n9531,n679,n9237);
xor (n9532,n9390,n9392);
and (n9533,n9528,n9531);
wire s0n9534,s1n9534,notn9534;
or (n9534,s0n9534,s1n9534);
not(notn9534,n8048);
and (s0n9534,notn9534,1'b0);
and (s1n9534,n8048,n9331);
and (n9535,n9524,n9525);
xor (n9536,n9350,n9372);
xor (n9537,n9376,n9396);
and (n9538,n9521,n9536);
xor (n9539,n9346,n9374);
or (n9540,n9541,n9558);
and (n9541,n9542,n9557);
xor (n9542,n9543,n9556);
or (n9543,n9544,n9555);
and (n9544,n9545,n9554);
xor (n9545,n9546,n9547);
wire s0n9546,s1n9546,notn9546;
or (n9546,s0n9546,s1n9546);
not(notn9546,n679);
and (s0n9546,notn9546,1'b0);
and (s1n9546,n679,n9397);
or (n9547,n9548,n9553);
and (n9548,n9549,n9552);
xor (n9549,n9550,n9551);
wire s0n9550,s1n9550,notn9550;
or (n9550,s0n9550,s1n9550);
not(notn9550,n8048);
and (s0n9550,notn9550,1'b0);
and (s1n9550,n8048,n9328);
xor (n9551,n9383,n9386);
wire s0n9552,s1n9552,notn9552;
or (n9552,s0n9552,s1n9552);
not(notn9552,n8048);
and (s0n9552,notn9552,1'b0);
and (s1n9552,n8048,n9310);
and (n9553,n9550,n9551);
xor (n9554,n9447,n9450);
and (n9555,n9546,n9547);
wire s0n9556,s1n9556,notn9556;
or (n9556,s0n9556,s1n9556);
not(notn9556,n35);
and (s0n9556,notn9556,1'b0);
and (s1n9556,n35,n9265);
wire s0n9557,s1n9557,notn9557;
or (n9557,s0n9557,s1n9557);
not(notn9557,n35);
and (s0n9557,notn9557,1'b0);
and (s1n9557,n35,n9172);
and (n9558,n9543,n9556);
and (n9559,n9518,n9539);
xor (n9560,n9427,n9432);
or (n9561,n9562,n9567);
and (n9562,n9563,n9566);
xor (n9563,n9564,n9565);
xor (n9564,n9439,n9454);
xor (n9565,n9459,n9462);
xor (n9566,n9487,n9496);
and (n9567,n9564,n9565);
and (n9568,n9515,n9560);
xor (n9569,n9424,n9465);
xor (n9570,n9479,n9500);
and (n9571,n9512,n9569);
xor (n9572,n9476,n9503);
or (n9573,n9574,n9668);
and (n9574,n9575,n9667);
xor (n9575,n9576,n9619);
or (n9576,n9577,n9618);
and (n9577,n9578,n9617);
xor (n9578,n9579,n9616);
or (n9579,n9580,n9615);
and (n9580,n9581,n9596);
xor (n9581,n9582,n9595);
or (n9582,n9583,n9594);
and (n9583,n9584,n9593);
xor (n9584,n9585,n9592);
or (n9585,n9586,n9591);
and (n9586,n9587,n9590);
xor (n9587,n9588,n9589);
wire s0n9588,s1n9588,notn9588;
or (n9588,s0n9588,s1n9588);
not(notn9588,n35);
and (s0n9588,notn9588,1'b0);
and (s1n9588,n35,n9305);
xor (n9589,n9380,n9394);
wire s0n9590,s1n9590,notn9590;
or (n9590,s0n9590,s1n9590);
not(notn9590,n35);
and (s0n9590,notn9590,1'b0);
and (s1n9590,n35,n9313);
and (n9591,n9588,n9589);
xor (n9592,n9443,n9452);
xor (n9593,n9491,n9494);
and (n9594,n9585,n9592);
xor (n9595,n9517,n9540);
or (n9596,n9597,n9614);
and (n9597,n9598,n9613);
xor (n9598,n9599,n9600);
xor (n9599,n9520,n9537);
or (n9600,n9601,n9612);
and (n9601,n9602,n9611);
xor (n9602,n9603,n9610);
or (n9603,n9604,n9609);
and (n9604,n9605,n9608);
xor (n9605,n9606,n9607);
wire s0n9606,s1n9606,notn9606;
or (n9606,s0n9606,s1n9606);
not(notn9606,n35);
and (s0n9606,notn9606,1'b0);
and (s1n9606,n35,n9331);
xor (n9607,n9527,n9532);
wire s0n9608,s1n9608,notn9608;
or (n9608,s0n9608,s1n9608);
not(notn9608,n35);
and (s0n9608,notn9608,1'b0);
and (s1n9608,n35,n9397);
and (n9609,n9606,n9607);
xor (n9610,n9523,n9534);
xor (n9611,n9545,n9554);
and (n9612,n9603,n9610);
xor (n9613,n9542,n9557);
and (n9614,n9599,n9600);
and (n9615,n9582,n9595);
xor (n9616,n9436,n9457);
xor (n9617,n9482,n9485);
and (n9618,n9579,n9616);
nand (n9619,n9620,n9663);
or (n9620,n9621,n9661);
not (n9621,n9622);
nand (n9622,n9623,n9625,n9660);
not (n9623,n9624);
xor (n9624,n9514,n9561);
nand (n9625,n9626,n9659);
or (n9626,n9627,n9628);
xor (n9627,n9581,n9596);
nand (n9628,n9629,n9656);
or (n9629,n9630,n9654);
not (n9630,n9631);
nand (n9631,n9632,n9651);
or (n9632,n9633,n9649);
not (n9633,n9634);
nand (n9634,n9635,n9646);
or (n9635,n9636,n9644);
not (n9636,n9637);
nand (n9637,n9638,n9641);
or (n9638,n8955,n9639);
not (n9639,n9640);
wire s0n9640,s1n9640,notn9640;
or (n9640,s0n9640,s1n9640);
not(notn9640,n35);
and (s0n9640,notn9640,1'b0);
and (s1n9640,n35,n9328);
nand (n9641,n9642,n9643);
or (n9642,n9640,n8956);
xor (n9643,n9529,n9530);
not (n9644,n9645);
xor (n9645,n9549,n9552);
nand (n9646,n9647,n9648);
or (n9647,n9645,n9637);
xor (n9648,n9605,n9608);
not (n9649,n9650);
xor (n9650,n9587,n9590);
nand (n9651,n9652,n9653);
or (n9652,n9650,n9634);
xor (n9653,n9602,n9611);
not (n9654,n9655);
xor (n9655,n9584,n9593);
nand (n9656,n9657,n9658);
or (n9657,n9655,n9631);
xor (n9658,n9598,n9613);
xor (n9659,n9563,n9566);
nand (n9660,n9627,n9628);
not (n9661,n9662);
xor (n9662,n9578,n9617);
nand (n9663,n9664,n9624);
or (n9664,n9665,n9666);
not (n9665,n9660);
not (n9666,n9625);
xor (n9667,n9511,n9570);
and (n9668,n9576,n9619);
and (n9669,n9509,n9572);
and (n9670,n9474,n9505);
and (n9671,n9413,n9414);
and (n9672,n9281,n9282);
and (n9673,n9202,n9203);
and (n9674,n7847,n9126);
nor (n9675,n9676,n9701);
not (n9676,n9677);
nor (n9677,n9678,n9698);
not (n9678,n9679);
nor (n9679,n9680,n9695);
not (n9680,n9681);
nor (n9681,n9682,n9692);
not (n9682,n9683);
nor (n9683,n9684,n9685);
and (n9684,n9079,n9082);
not (n9685,n9686);
nor (n9686,n9687,n9688);
and (n9687,n9074,n9077);
not (n9688,n9689);
xnor (n9689,n9690,n9691);
wire s0n9690,s1n9690,notn9690;
or (n9690,s0n9690,s1n9690);
not(notn9690,n7785);
and (s0n9690,notn9690,1'b0);
and (s1n9690,n7785,n7857);
wire s0n9691,s1n9691,notn9691;
or (n9691,s0n9691,s1n9691);
not(notn9691,n7785);
and (s0n9691,notn9691,1'b0);
and (s1n9691,n7785,n8622);
or (n9692,n9693,n9694);
and (n9693,n9069,n9078);
and (n9694,n9070,n9073);
or (n9695,n9696,n9697);
and (n9696,n9033,n9056);
and (n9697,n9034,n9037);
or (n9698,n9699,n9700);
and (n9699,n9064,n9083);
and (n9700,n9065,n9068);
or (n9701,n9702,n9703);
and (n9702,n7848,n9063);
and (n9703,n7849,n9032);
nor (n9704,n9705,n7735);
not (n9705,n9706);
and (n9706,n626,n4651);
wire s0n9707,s1n9707,notn9707;
or (n9707,s0n9707,s1n9707);
not(notn9707,n7196);
and (s0n9707,notn9707,n9708);
and (s1n9707,n7196,n10448);
wire s0n9708,s1n9708,notn9708;
or (n9708,s0n9708,s1n9708);
not(notn9708,n7735);
and (s0n9708,notn9708,n9709);
and (s1n9708,n7735,n7725);
xor (n9709,n9710,n10425);
xor (n9710,n9711,n10326);
xor (n9711,n9712,n10029);
xor (n9712,n9713,n9936);
xor (n9713,n9714,n9821);
xor (n9714,n9690,n9715);
or (n9715,n9716,n9754,n9820);
and (n9716,n9717,n9718);
xor (n9717,n9077,n9082);
and (n9718,n7856,n9719);
or (n9719,n9720,n9721,n9753);
and (n9720,n8835,n8827);
and (n9721,n8827,n9722);
or (n9722,n9723,n9724,n9752);
and (n9723,n8788,n9028);
and (n9724,n9028,n9725);
or (n9725,n9726,n9727,n9751);
and (n9726,n8877,n9002);
and (n9727,n9002,n9728);
or (n9728,n9729,n9730,n9750);
and (n9729,n9189,n9191);
and (n9730,n9191,n9731);
or (n9731,n9732,n9733,n9749);
and (n9732,n9249,n9270);
and (n9733,n9270,n9734);
or (n9734,n9735,n9736,n9748);
and (n9735,n9333,n9431);
and (n9736,n9431,n9737);
or (n9737,n9738,n9739,n9747);
and (n9738,n9454,n9462);
and (n9739,n9462,n9740);
or (n9740,n9741,n9742,n9744);
and (n9741,n9494,n9557);
and (n9742,n9557,n9743);
or (n9743,n9744,n9745,n9746);
and (n9744,n9534,n9590);
and (n9745,n9590,n9746);
and (n9746,n9550,n9606);
and (n9747,n9454,n9740);
and (n9748,n9333,n9737);
and (n9749,n9249,n9734);
and (n9750,n9189,n9731);
and (n9751,n8877,n9728);
and (n9752,n8788,n9725);
and (n9753,n8835,n9722);
and (n9754,n9718,n9755);
or (n9755,n9756,n9759,n9819);
and (n9756,n9757,n9758);
xor (n9757,n8796,n8233);
xor (n9758,n7856,n9719);
and (n9759,n9758,n9760);
or (n9760,n9761,n9765,n9818);
and (n9761,n9762,n9763);
xor (n9762,n9051,n8822);
xor (n9763,n9764,n9722);
xor (n9764,n8835,n8827);
and (n9765,n9763,n9766);
or (n9766,n9767,n9771,n9817);
and (n9767,n9768,n9769);
xor (n9768,n8714,n8658);
xor (n9769,n9770,n9725);
xor (n9770,n8788,n9028);
and (n9771,n9769,n9772);
or (n9772,n9773,n9777,n9816);
and (n9773,n9774,n9775);
xor (n9774,n9116,n8848);
xor (n9775,n9776,n9728);
xor (n9776,n8877,n9002);
and (n9777,n9775,n9778);
or (n9778,n9779,n9783,n9815);
and (n9779,n9780,n9781);
xor (n9780,n8873,n8998);
xor (n9781,n9782,n9731);
xor (n9782,n9189,n9191);
and (n9783,n9781,n9784);
or (n9784,n9785,n9789,n9814);
and (n9785,n9786,n9787);
xor (n9786,n9171,n9167);
xor (n9787,n9788,n9734);
xor (n9788,n9249,n9270);
and (n9789,n9787,n9790);
or (n9790,n9791,n9795,n9813);
and (n9791,n9792,n9793);
xor (n9792,n9430,n9267);
xor (n9793,n9794,n9737);
xor (n9794,n9333,n9431);
and (n9795,n9793,n9796);
or (n9796,n9797,n9801,n9812);
and (n9797,n9798,n9799);
xor (n9798,n9330,n9312);
xor (n9799,n9800,n9740);
xor (n9800,n9454,n9462);
and (n9801,n9799,n9802);
or (n9802,n9803,n9807,n9811);
and (n9803,n9804,n9805);
xor (n9804,n9327,n9444);
xor (n9805,n9806,n9743);
xor (n9806,n9494,n9557);
and (n9807,n9805,n9808);
and (n9808,n9394,n9809);
xor (n9809,n9810,n9746);
xor (n9810,n9534,n9590);
and (n9811,n9804,n9808);
and (n9812,n9798,n9802);
and (n9813,n9792,n9796);
and (n9814,n9786,n9790);
and (n9815,n9780,n9784);
and (n9816,n9774,n9778);
and (n9817,n9768,n9772);
and (n9818,n9762,n9766);
and (n9819,n9757,n9760);
and (n9820,n9717,n9755);
xor (n9821,n9691,n9822);
or (n9822,n9823,n9870,n9935);
and (n9823,n9074,n9824);
and (n9824,n8621,n9825);
or (n9825,n9826,n9828,n9869);
and (n9826,n9042,n9827);
wire s0n9827,s1n9827,notn9827;
or (n9827,s0n9827,s1n9827);
not(notn9827,n35);
and (s0n9827,notn9827,1'b0);
and (s1n9827,n35,n8622);
and (n9828,n9827,n9829);
or (n9829,n9830,n9832,n9868);
and (n9830,n9010,n9831);
wire s0n9831,s1n9831,notn9831;
or (n9831,s0n9831,s1n9831);
not(notn9831,n35);
and (s0n9831,notn9831,1'b0);
and (s1n9831,n35,n8633);
and (n9832,n9831,n9833);
or (n9833,n9834,n9836,n9867);
and (n9834,n8818,n9835);
wire s0n9835,s1n9835,notn9835;
or (n9835,s0n9835,s1n9835);
not(notn9835,n35);
and (s0n9835,notn9835,1'b0);
and (s1n9835,n35,n8475);
and (n9836,n9835,n9837);
or (n9837,n9838,n9840,n9866);
and (n9838,n8924,n9839);
wire s0n9839,s1n9839,notn9839;
or (n9839,s0n9839,s1n9839);
not(notn9839,n35);
and (s0n9839,notn9839,1'b0);
and (s1n9839,n35,n8459);
and (n9840,n9839,n9841);
or (n9841,n9842,n9844,n9865);
and (n9842,n8893,n9843);
wire s0n9843,s1n9843,notn9843;
or (n9843,s0n9843,s1n9843);
not(notn9843,n35);
and (s0n9843,notn9843,1'b0);
and (s1n9843,n35,n8247);
and (n9844,n9843,n9845);
or (n9845,n9846,n9848,n9864);
and (n9846,n8996,n9847);
wire s0n9847,s1n9847,notn9847;
or (n9847,s0n9847,s1n9847);
not(notn9847,n35);
and (s0n9847,notn9847,1'b0);
and (s1n9847,n35,n8759);
and (n9848,n9847,n9849);
or (n9849,n9850,n9852,n9863);
and (n9850,n9164,n9851);
wire s0n9851,s1n9851,notn9851;
or (n9851,s0n9851,s1n9851);
not(notn9851,n35);
and (s0n9851,notn9851,1'b0);
and (s1n9851,n35,n8862);
and (n9852,n9851,n9853);
or (n9853,n9854,n9856,n9858);
and (n9854,n9372,n9855);
wire s0n9855,s1n9855,notn9855;
or (n9855,s0n9855,s1n9855);
not(notn9855,n35);
and (s0n9855,notn9855,1'b0);
and (s1n9855,n35,n8868);
and (n9856,n9855,n9857);
or (n9857,n9858,n9860,n9861);
and (n9858,n9449,n9859);
wire s0n9859,s1n9859,notn9859;
or (n9859,s0n9859,s1n9859);
not(notn9859,n35);
and (s0n9859,notn9859,1'b0);
and (s1n9859,n35,n8995);
and (n9860,n9859,n9861);
and (n9861,n9552,n9862);
wire s0n9862,s1n9862,notn9862;
or (n9862,s0n9862,s1n9862);
not(notn9862,n35);
and (s0n9862,notn9862,1'b0);
and (s1n9862,n35,n8962);
and (n9863,n9164,n9853);
and (n9864,n8996,n9849);
and (n9865,n8893,n9845);
and (n9866,n8924,n9841);
and (n9867,n8818,n9837);
and (n9868,n9010,n9833);
and (n9869,n9042,n9829);
and (n9870,n9824,n9871);
or (n9871,n9872,n9875,n9934);
and (n9872,n9873,n9874);
xor (n9873,n8631,n8632);
xor (n9874,n8621,n9825);
and (n9875,n9874,n9876);
or (n9876,n9877,n9881,n9933);
and (n9877,n9878,n9879);
xor (n9878,n9045,n8474);
xor (n9879,n9880,n9829);
xor (n9880,n9042,n9827);
and (n9881,n9879,n9882);
or (n9882,n9883,n9887,n9932);
and (n9883,n9884,n9885);
xor (n9884,n8246,n8458);
xor (n9885,n9886,n9833);
xor (n9886,n9010,n9831);
and (n9887,n9885,n9888);
or (n9888,n9889,n9892,n9931);
and (n9889,n8815,n9890);
xor (n9890,n9891,n9837);
xor (n9891,n8818,n9835);
and (n9892,n9890,n9893);
or (n9893,n9894,n9898,n9930);
and (n9894,n9895,n9896);
xor (n9895,n8861,n8758);
xor (n9896,n9897,n9841);
xor (n9897,n8924,n9839);
and (n9898,n9896,n9899);
or (n9899,n9900,n9904,n9929);
and (n9900,n9901,n9902);
xor (n9901,n8867,n8943);
xor (n9902,n9903,n9845);
xor (n9903,n8893,n9843);
and (n9904,n9902,n9905);
or (n9905,n9906,n9910,n9928);
and (n9906,n9907,n9908);
xor (n9907,n8994,n8911);
xor (n9908,n9909,n9849);
xor (n9909,n8996,n9847);
and (n9910,n9908,n9911);
or (n9911,n9912,n9916,n9927);
and (n9912,n9913,n9914);
xor (n9913,n8961,n9161);
xor (n9914,n9915,n9853);
xor (n9915,n9164,n9851);
and (n9916,n9914,n9917);
or (n9917,n9918,n9922,n9926);
and (n9918,n9919,n9920);
xor (n9919,n9309,n9329);
xor (n9920,n9921,n9857);
xor (n9921,n9372,n9855);
and (n9922,n9920,n9923);
and (n9923,n9450,n9924);
xor (n9924,n9925,n9861);
xor (n9925,n9449,n9859);
and (n9926,n9919,n9923);
and (n9927,n9913,n9917);
and (n9928,n9907,n9911);
and (n9929,n9901,n9905);
and (n9930,n9895,n9899);
and (n9931,n8815,n9893);
and (n9932,n9884,n9888);
and (n9933,n9878,n9882);
and (n9934,n9873,n9876);
and (n9935,n9074,n9871);
or (n9936,n9937,n9942,n10028);
and (n9937,n9938,n9940);
xor (n9938,n9939,n9755);
xor (n9939,n9717,n9718);
xor (n9940,n9941,n9871);
xor (n9941,n9074,n9824);
and (n9942,n9940,n9943);
or (n9943,n9944,n9949,n10027);
and (n9944,n9945,n9947);
xor (n9945,n9946,n9760);
xor (n9946,n9757,n9758);
xor (n9947,n9948,n9876);
xor (n9948,n9873,n9874);
and (n9949,n9947,n9950);
or (n9950,n9951,n9956,n10026);
and (n9951,n9952,n9954);
xor (n9952,n9953,n9766);
xor (n9953,n9762,n9763);
xor (n9954,n9955,n9882);
xor (n9955,n9878,n9879);
and (n9956,n9954,n9957);
or (n9957,n9958,n9963,n10025);
and (n9958,n9959,n9961);
xor (n9959,n9960,n9772);
xor (n9960,n9768,n9769);
xor (n9961,n9962,n9888);
xor (n9962,n9884,n9885);
and (n9963,n9961,n9964);
or (n9964,n9965,n9970,n10024);
and (n9965,n9966,n9968);
xor (n9966,n9967,n9778);
xor (n9967,n9774,n9775);
xor (n9968,n9969,n9893);
xor (n9969,n8815,n9890);
and (n9970,n9968,n9971);
or (n9971,n9972,n9977,n10023);
and (n9972,n9973,n9975);
xor (n9973,n9974,n9784);
xor (n9974,n9780,n9781);
xor (n9975,n9976,n9899);
xor (n9976,n9895,n9896);
and (n9977,n9975,n9978);
or (n9978,n9979,n9984,n10022);
and (n9979,n9980,n9982);
xor (n9980,n9981,n9790);
xor (n9981,n9786,n9787);
xor (n9982,n9983,n9905);
xor (n9983,n9901,n9902);
and (n9984,n9982,n9985);
or (n9985,n9986,n9991,n10021);
and (n9986,n9987,n9989);
xor (n9987,n9988,n9796);
xor (n9988,n9792,n9793);
xor (n9989,n9990,n9911);
xor (n9990,n9907,n9908);
and (n9991,n9989,n9992);
or (n9992,n9993,n9998,n10020);
and (n9993,n9994,n9996);
xor (n9994,n9995,n9802);
xor (n9995,n9798,n9799);
xor (n9996,n9997,n9917);
xor (n9997,n9913,n9914);
and (n9998,n9996,n9999);
or (n9999,n10000,n10005,n10019);
and (n10000,n10001,n10003);
xor (n10001,n10002,n9808);
xor (n10002,n9804,n9805);
xor (n10003,n10004,n9923);
xor (n10004,n9919,n9920);
and (n10005,n10003,n10006);
or (n10006,n10007,n10010,n10018);
and (n10007,n10008,n10009);
xor (n10008,n9394,n9809);
xor (n10009,n9450,n9924);
and (n10010,n10009,n10011);
or (n10011,n10012,n10015,n10017);
and (n10012,n10013,n10014);
xor (n10013,n9550,n9606);
xor (n10014,n9552,n9862);
and (n10015,n10014,n10016);
and (n10016,n9640,n9529);
and (n10017,n10013,n10016);
and (n10018,n10008,n10011);
and (n10019,n10001,n10006);
and (n10020,n9994,n9999);
and (n10021,n9987,n9992);
and (n10022,n9980,n9985);
and (n10023,n9973,n9978);
and (n10024,n9966,n9971);
and (n10025,n9959,n9964);
and (n10026,n9952,n9957);
and (n10027,n9945,n9950);
and (n10028,n9938,n9943);
xor (n10029,n10030,n10233);
xor (n10030,n10031,n10127);
or (n10031,n10032,n10069,n10126);
and (n10032,n9080,n10033);
and (n10033,n9048,n10034);
or (n10034,n10035,n10036,n10068);
and (n10035,n9046,n8828);
and (n10036,n8828,n10037);
or (n10037,n10038,n10039,n10067);
and (n10038,n8652,n9007);
and (n10039,n9007,n10040);
or (n10040,n10041,n10042,n10066);
and (n10041,n8855,n8850);
and (n10042,n8850,n10043);
or (n10043,n10044,n10045,n10065);
and (n10044,n9190,n9178);
and (n10045,n9178,n10046);
or (n10046,n10047,n10048,n10064);
and (n10047,n9250,n9297);
and (n10048,n9297,n10049);
or (n10049,n10050,n10051,n10063);
and (n10050,n9400,n9432);
and (n10051,n9432,n10052);
or (n10052,n10053,n10054,n10062);
and (n10053,n9460,n9496);
and (n10054,n9496,n10055);
or (n10055,n10056,n10057,n10059);
and (n10056,n9493,n9556);
and (n10057,n9556,n10058);
or (n10058,n10059,n10060,n10061);
and (n10059,n9546,n9588);
and (n10060,n9588,n10061);
and (n10061,n9531,n9608);
and (n10062,n9460,n10055);
and (n10063,n9400,n10052);
and (n10064,n9250,n10049);
and (n10065,n9190,n10046);
and (n10066,n8855,n10043);
and (n10067,n8652,n10040);
and (n10068,n9046,n10037);
and (n10069,n10033,n10070);
or (n10070,n10071,n10073,n10125);
and (n10071,n8051,n10072);
xor (n10072,n9048,n10034);
and (n10073,n10072,n10074);
or (n10074,n10075,n10078,n10124);
and (n10075,n8821,n10076);
xor (n10076,n10077,n10037);
xor (n10077,n9046,n8828);
and (n10078,n10076,n10079);
or (n10079,n10080,n10083,n10123);
and (n10080,n8655,n10081);
xor (n10081,n10082,n10040);
xor (n10082,n8652,n9007);
and (n10083,n10081,n10084);
or (n10084,n10085,n10088,n10122);
and (n10085,n9118,n10086);
xor (n10086,n10087,n10043);
xor (n10087,n8855,n8850);
and (n10088,n10086,n10089);
or (n10089,n10090,n10093,n10121);
and (n10090,n8915,n10091);
xor (n10091,n10092,n10046);
xor (n10092,n9190,n9178);
and (n10093,n10091,n10094);
or (n10094,n10095,n10098,n10120);
and (n10095,n9175,n10096);
xor (n10096,n10097,n10049);
xor (n10097,n9250,n9297);
and (n10098,n10096,n10099);
or (n10099,n10100,n10103,n10119);
and (n10100,n9264,n10101);
xor (n10101,n10102,n10052);
xor (n10102,n9400,n9432);
and (n10103,n10101,n10104);
or (n10104,n10105,n10108,n10118);
and (n10105,n9304,n10106);
xor (n10106,n10107,n10055);
xor (n10107,n9460,n9496);
and (n10108,n10106,n10109);
or (n10109,n10110,n10113,n10117);
and (n10110,n9396,n10111);
xor (n10111,n10112,n10058);
xor (n10112,n9493,n9556);
and (n10113,n10111,n10114);
and (n10114,n9236,n10115);
xor (n10115,n10116,n10061);
xor (n10116,n9546,n9588);
and (n10117,n9396,n10114);
and (n10118,n9304,n10109);
and (n10119,n9264,n10104);
and (n10120,n9175,n10099);
and (n10121,n8915,n10094);
and (n10122,n9118,n10089);
and (n10123,n8655,n10084);
and (n10124,n8821,n10079);
and (n10125,n8051,n10074);
and (n10126,n9080,n10070);
or (n10127,n10128,n10175,n10232);
and (n10128,n9081,n10129);
and (n10129,n8635,n10130);
or (n10130,n10131,n10133,n10174);
and (n10131,n9055,n10132);
wire s0n10132,s1n10132,notn10132;
or (n10132,s0n10132,s1n10132);
not(notn10132,n35);
and (s0n10132,notn10132,1'b0);
and (s1n10132,n35,n8636);
and (n10133,n10132,n10134);
or (n10134,n10135,n10137,n10173);
and (n10135,n8819,n10136);
wire s0n10136,s1n10136,notn10136;
or (n10136,s0n10136,s1n10136);
not(notn10136,n35);
and (s0n10136,notn10136,1'b0);
and (s1n10136,n35,n8805);
and (n10137,n10136,n10138);
or (n10138,n10139,n10141,n10172);
and (n10139,n9111,n10140);
wire s0n10140,s1n10140,notn10140;
or (n10140,s0n10140,s1n10140);
not(notn10140,n35);
and (s0n10140,notn10140,1'b0);
and (s1n10140,n35,n8487);
and (n10141,n10140,n10142);
or (n10142,n10143,n10145,n10171);
and (n10143,n8945,n10144);
wire s0n10144,s1n10144,notn10144;
or (n10144,s0n10144,s1n10144);
not(notn10144,n35);
and (s0n10144,notn10144,1'b0);
and (s1n10144,n35,n9026);
and (n10145,n10144,n10146);
or (n10146,n10147,n10149,n10170);
and (n10147,n8913,n10148);
wire s0n10148,s1n10148,notn10148;
or (n10148,s0n10148,s1n10148);
not(notn10148,n35);
and (s0n10148,notn10148,1'b0);
and (s1n10148,n35,n8721);
and (n10149,n10148,n10150);
or (n10150,n10151,n10153,n10169);
and (n10151,n8993,n10152);
wire s0n10152,s1n10152,notn10152;
or (n10152,s0n10152,s1n10152);
not(notn10152,n35);
and (s0n10152,notn10152,1'b0);
and (s1n10152,n35,n8784);
and (n10153,n10152,n10154);
or (n10154,n10155,n10157,n10168);
and (n10155,n9247,n10156);
wire s0n10156,s1n10156,notn10156;
or (n10156,s0n10156,s1n10156);
not(notn10156,n35);
and (s0n10156,notn10156,1'b0);
and (s1n10156,n35,n8871);
and (n10157,n10156,n10158);
or (n10158,n10159,n10161,n10163);
and (n10159,n9311,n10160);
wire s0n10160,s1n10160,notn10160;
or (n10160,s0n10160,s1n10160);
not(notn10160,n35);
and (s0n10160,notn10160,1'b0);
and (s1n10160,n35,n8988);
and (n10161,n10160,n10162);
or (n10162,n10163,n10165,n10166);
and (n10163,n9354,n10164);
wire s0n10164,s1n10164,notn10164;
or (n10164,s0n10164,s1n10164);
not(notn10164,n35);
and (s0n10164,notn10164,1'b0);
and (s1n10164,n35,n9163);
and (n10165,n10164,n10166);
and (n10166,n9385,n10167);
wire s0n10167,s1n10167,notn10167;
or (n10167,s0n10167,s1n10167);
not(notn10167,n35);
and (s0n10167,notn10167,1'b0);
and (s1n10167,n35,n9233);
and (n10168,n9247,n10158);
and (n10169,n8993,n10154);
and (n10170,n8913,n10150);
and (n10171,n8945,n10146);
and (n10172,n9111,n10142);
and (n10173,n8819,n10138);
and (n10174,n9055,n10134);
and (n10175,n10129,n10176);
or (n10176,n10177,n10179,n10231);
and (n10177,n8804,n10178);
xor (n10178,n8635,n10130);
and (n10179,n10178,n10180);
or (n10180,n10181,n10184,n10230);
and (n10181,n8486,n10182);
xor (n10182,n10183,n10134);
xor (n10183,n9055,n10132);
and (n10184,n10182,n10185);
or (n10185,n10186,n10189,n10229);
and (n10186,n9025,n10187);
xor (n10187,n10188,n10138);
xor (n10188,n8819,n10136);
and (n10189,n10187,n10190);
or (n10190,n10191,n10194,n10228);
and (n10191,n8720,n10192);
xor (n10192,n10193,n10142);
xor (n10193,n9111,n10140);
and (n10194,n10192,n10195);
or (n10195,n10196,n10199,n10227);
and (n10196,n8783,n10197);
xor (n10197,n10198,n10146);
xor (n10198,n8945,n10144);
and (n10199,n10197,n10200);
or (n10200,n10201,n10204,n10226);
and (n10201,n8870,n10202);
xor (n10202,n10203,n10150);
xor (n10203,n8913,n10148);
and (n10204,n10202,n10205);
or (n10205,n10206,n10209,n10225);
and (n10206,n8987,n10207);
xor (n10207,n10208,n10154);
xor (n10208,n8993,n10152);
and (n10209,n10207,n10210);
or (n10210,n10211,n10214,n10224);
and (n10211,n9162,n10212);
xor (n10212,n10213,n10158);
xor (n10213,n9247,n10156);
and (n10214,n10212,n10215);
or (n10215,n10216,n10219,n10223);
and (n10216,n9232,n10217);
xor (n10217,n10218,n10162);
xor (n10218,n9311,n10160);
and (n10219,n10217,n10220);
and (n10220,n9235,n10221);
xor (n10221,n10222,n10166);
xor (n10222,n9354,n10164);
and (n10223,n9232,n10220);
and (n10224,n9162,n10215);
and (n10225,n8987,n10210);
and (n10226,n8870,n10205);
and (n10227,n8783,n10200);
and (n10228,n8720,n10195);
and (n10229,n9025,n10190);
and (n10230,n8486,n10185);
and (n10231,n8804,n10180);
and (n10232,n9081,n10176);
or (n10233,n10234,n10239,n10325);
and (n10234,n10235,n10237);
xor (n10235,n10236,n10070);
xor (n10236,n9080,n10033);
xor (n10237,n10238,n10176);
xor (n10238,n9081,n10129);
and (n10239,n10237,n10240);
or (n10240,n10241,n10246,n10324);
and (n10241,n10242,n10244);
xor (n10242,n10243,n10074);
xor (n10243,n8051,n10072);
xor (n10244,n10245,n10180);
xor (n10245,n8804,n10178);
and (n10246,n10244,n10247);
or (n10247,n10248,n10253,n10323);
and (n10248,n10249,n10251);
xor (n10249,n10250,n10079);
xor (n10250,n8821,n10076);
xor (n10251,n10252,n10185);
xor (n10252,n8486,n10182);
and (n10253,n10251,n10254);
or (n10254,n10255,n10260,n10322);
and (n10255,n10256,n10258);
xor (n10256,n10257,n10084);
xor (n10257,n8655,n10081);
xor (n10258,n10259,n10190);
xor (n10259,n9025,n10187);
and (n10260,n10258,n10261);
or (n10261,n10262,n10267,n10321);
and (n10262,n10263,n10265);
xor (n10263,n10264,n10089);
xor (n10264,n9118,n10086);
xor (n10265,n10266,n10195);
xor (n10266,n8720,n10192);
and (n10267,n10265,n10268);
or (n10268,n10269,n10274,n10320);
and (n10269,n10270,n10272);
xor (n10270,n10271,n10094);
xor (n10271,n8915,n10091);
xor (n10272,n10273,n10200);
xor (n10273,n8783,n10197);
and (n10274,n10272,n10275);
or (n10275,n10276,n10281,n10319);
and (n10276,n10277,n10279);
xor (n10277,n10278,n10099);
xor (n10278,n9175,n10096);
xor (n10279,n10280,n10205);
xor (n10280,n8870,n10202);
and (n10281,n10279,n10282);
or (n10282,n10283,n10288,n10318);
and (n10283,n10284,n10286);
xor (n10284,n10285,n10104);
xor (n10285,n9264,n10101);
xor (n10286,n10287,n10210);
xor (n10287,n8987,n10207);
and (n10288,n10286,n10289);
or (n10289,n10290,n10295,n10317);
and (n10290,n10291,n10293);
xor (n10291,n10292,n10109);
xor (n10292,n9304,n10106);
xor (n10293,n10294,n10215);
xor (n10294,n9162,n10212);
and (n10295,n10293,n10296);
or (n10296,n10297,n10302,n10316);
and (n10297,n10298,n10300);
xor (n10298,n10299,n10114);
xor (n10299,n9396,n10111);
xor (n10300,n10301,n10220);
xor (n10301,n9232,n10217);
and (n10302,n10300,n10303);
or (n10303,n10304,n10307,n10315);
and (n10304,n10305,n10306);
xor (n10305,n9236,n10115);
xor (n10306,n9235,n10221);
and (n10307,n10306,n10308);
or (n10308,n10309,n10312,n10314);
and (n10309,n10310,n10311);
xor (n10310,n9531,n9608);
xor (n10311,n9385,n10167);
and (n10312,n10311,n10313);
and (n10313,n9530,n8956);
and (n10314,n10310,n10313);
and (n10315,n10305,n10308);
and (n10316,n10298,n10303);
and (n10317,n10291,n10296);
and (n10318,n10284,n10289);
and (n10319,n10277,n10282);
and (n10320,n10270,n10275);
and (n10321,n10263,n10268);
and (n10322,n10256,n10261);
and (n10323,n10249,n10254);
and (n10324,n10242,n10247);
and (n10325,n10235,n10240);
or (n10326,n10327,n10332,n10424);
and (n10327,n10328,n10330);
xor (n10328,n10329,n9943);
xor (n10329,n9938,n9940);
xor (n10330,n10331,n10240);
xor (n10331,n10235,n10237);
and (n10332,n10330,n10333);
or (n10333,n10334,n10339,n10423);
and (n10334,n10335,n10337);
xor (n10335,n10336,n9950);
xor (n10336,n9945,n9947);
xor (n10337,n10338,n10247);
xor (n10338,n10242,n10244);
and (n10339,n10337,n10340);
or (n10340,n10341,n10346,n10422);
and (n10341,n10342,n10344);
xor (n10342,n10343,n9957);
xor (n10343,n9952,n9954);
xor (n10344,n10345,n10254);
xor (n10345,n10249,n10251);
and (n10346,n10344,n10347);
or (n10347,n10348,n10353,n10421);
and (n10348,n10349,n10351);
xor (n10349,n10350,n9964);
xor (n10350,n9959,n9961);
xor (n10351,n10352,n10261);
xor (n10352,n10256,n10258);
and (n10353,n10351,n10354);
or (n10354,n10355,n10360,n10420);
and (n10355,n10356,n10358);
xor (n10356,n10357,n9971);
xor (n10357,n9966,n9968);
xor (n10358,n10359,n10268);
xor (n10359,n10263,n10265);
and (n10360,n10358,n10361);
or (n10361,n10362,n10367,n10419);
and (n10362,n10363,n10365);
xor (n10363,n10364,n9978);
xor (n10364,n9973,n9975);
xor (n10365,n10366,n10275);
xor (n10366,n10270,n10272);
and (n10367,n10365,n10368);
or (n10368,n10369,n10374,n10418);
and (n10369,n10370,n10372);
xor (n10370,n10371,n9985);
xor (n10371,n9980,n9982);
xor (n10372,n10373,n10282);
xor (n10373,n10277,n10279);
and (n10374,n10372,n10375);
or (n10375,n10376,n10381,n10417);
and (n10376,n10377,n10379);
xor (n10377,n10378,n9992);
xor (n10378,n9987,n9989);
xor (n10379,n10380,n10289);
xor (n10380,n10284,n10286);
and (n10381,n10379,n10382);
or (n10382,n10383,n10388,n10416);
and (n10383,n10384,n10386);
xor (n10384,n10385,n9999);
xor (n10385,n9994,n9996);
xor (n10386,n10387,n10296);
xor (n10387,n10291,n10293);
and (n10388,n10386,n10389);
or (n10389,n10390,n10395,n10415);
and (n10390,n10391,n10393);
xor (n10391,n10392,n10006);
xor (n10392,n10001,n10003);
xor (n10393,n10394,n10303);
xor (n10394,n10298,n10300);
and (n10395,n10393,n10396);
or (n10396,n10397,n10402,n10414);
and (n10397,n10398,n10400);
xor (n10398,n10399,n10011);
xor (n10399,n10008,n10009);
xor (n10400,n10401,n10308);
xor (n10401,n10305,n10306);
and (n10402,n10400,n10403);
or (n10403,n10404,n10409,n10413);
and (n10404,n10405,n10407);
xor (n10405,n10406,n10016);
xor (n10406,n10013,n10014);
xor (n10407,n10408,n10313);
xor (n10408,n10310,n10311);
and (n10409,n10407,n10410);
and (n10410,n10411,n10412);
xor (n10411,n9640,n9529);
xor (n10412,n9530,n8956);
and (n10413,n10405,n10410);
and (n10414,n10398,n10403);
and (n10415,n10391,n10396);
and (n10416,n10384,n10389);
and (n10417,n10377,n10382);
and (n10418,n10370,n10375);
and (n10419,n10363,n10368);
and (n10420,n10356,n10361);
and (n10421,n10349,n10354);
and (n10422,n10342,n10347);
and (n10423,n10335,n10340);
and (n10424,n10328,n10333);
and (n10425,n10426,n10428);
xor (n10426,n10427,n10333);
xor (n10427,n10328,n10330);
and (n10428,n10429,n10431);
xor (n10429,n10430,n10340);
xor (n10430,n10335,n10337);
and (n10431,n10432,n10434);
xor (n10432,n10433,n10347);
xor (n10433,n10342,n10344);
and (n10434,n10435,n10437);
xor (n10435,n10436,n10354);
xor (n10436,n10349,n10351);
and (n10437,n10438,n10440);
xor (n10438,n10439,n10361);
xor (n10439,n10356,n10358);
and (n10440,n10441,n10443);
xor (n10441,n10442,n10368);
xor (n10442,n10363,n10365);
and (n10443,n10444,n10446);
xor (n10444,n10445,n10375);
xor (n10445,n10370,n10372);
xor (n10446,n10447,n10382);
xor (n10447,n10377,n10379);
or (n10448,n10449,n10454,n7725);
and (n10449,n10450,n10451);
wire s0n10450,s1n10450,notn10450;
or (n10450,s0n10450,s1n10450);
not(notn10450,n897);
and (s0n10450,notn10450,1'b0);
and (s1n10450,n897,n2);
nor (n10451,n7839,n10452,n1071);
not (n10452,n10453);
nand (n10453,n32,n677,n751,n914);
and (n10454,n10455,n917);
wire s0n10455,s1n10455,notn10455;
or (n10455,s0n10455,s1n10455);
not(notn10455,n918);
and (s0n10455,notn10455,1'b0);
and (s1n10455,n918,n2);
endmodule
