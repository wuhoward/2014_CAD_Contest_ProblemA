module top (out,n19,n20,n24,n26,n28,n29,n30,n33,n34
        ,n35,n39,n40,n44,n46,n48,n49,n52,n54,n56
        ,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67
        ,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77
        ,n78,n79,n80,n81,n82,n83,n84,n85,n86,n94
        ,n95,n96,n100,n101,n102,n110,n111,n112,n116,n117
        ,n118,n129,n130,n131,n141,n142,n143,n146,n147,n148
        ,n154,n155,n156,n163,n164,n165,n179,n180,n181,n190
        ,n191,n192,n195,n196,n197,n206,n207,n208,n222,n223
        ,n224,n235,n236,n237,n243,n244,n245,n251,n252,n253
        ,n260,n261,n262,n275,n276,n277,n286,n287,n288,n291
        ,n292,n293,n305,n306,n307,n318,n319,n320,n331,n332
        ,n333,n347,n348,n349,n358,n359,n360,n386,n387,n388
        ,n414,n415,n416,n522,n523,n524,n1144,n1145,n1149,n1151
        ,n1153,n1156,n1157,n1161,n1163,n1165,n1166,n1169,n1171,n1173
        ,n1175,n1176,n1177,n1178,n1179,n1180,n1181,n1182,n1183,n1184
        ,n1185,n1186,n1187,n1188,n1189,n1190,n1191,n1192,n1193,n1194
        ,n1195,n1196,n1197,n1198,n1199,n1200,n1201,n1202,n1203,n1206
        ,n1207,n1210,n1211,n1212);
output out;
input n19;
input n20;
input n24;
input n26;
input n28;
input n29;
input n30;
input n33;
input n34;
input n35;
input n39;
input n40;
input n44;
input n46;
input n48;
input n49;
input n52;
input n54;
input n56;
input n58;
input n59;
input n60;
input n61;
input n62;
input n63;
input n64;
input n65;
input n66;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n81;
input n82;
input n83;
input n84;
input n85;
input n86;
input n94;
input n95;
input n96;
input n100;
input n101;
input n102;
input n110;
input n111;
input n112;
input n116;
input n117;
input n118;
input n129;
input n130;
input n131;
input n141;
input n142;
input n143;
input n146;
input n147;
input n148;
input n154;
input n155;
input n156;
input n163;
input n164;
input n165;
input n179;
input n180;
input n181;
input n190;
input n191;
input n192;
input n195;
input n196;
input n197;
input n206;
input n207;
input n208;
input n222;
input n223;
input n224;
input n235;
input n236;
input n237;
input n243;
input n244;
input n245;
input n251;
input n252;
input n253;
input n260;
input n261;
input n262;
input n275;
input n276;
input n277;
input n286;
input n287;
input n288;
input n291;
input n292;
input n293;
input n305;
input n306;
input n307;
input n318;
input n319;
input n320;
input n331;
input n332;
input n333;
input n347;
input n348;
input n349;
input n358;
input n359;
input n360;
input n386;
input n387;
input n388;
input n414;
input n415;
input n416;
input n522;
input n523;
input n524;
input n1144;
input n1145;
input n1149;
input n1151;
input n1153;
input n1156;
input n1157;
input n1161;
input n1163;
input n1165;
input n1166;
input n1169;
input n1171;
input n1173;
input n1175;
input n1176;
input n1177;
input n1178;
input n1179;
input n1180;
input n1181;
input n1182;
input n1183;
input n1184;
input n1185;
input n1186;
input n1187;
input n1188;
input n1189;
input n1190;
input n1191;
input n1192;
input n1193;
input n1194;
input n1195;
input n1196;
input n1197;
input n1198;
input n1199;
input n1200;
input n1201;
input n1202;
input n1203;
input n1206;
input n1207;
input n1210;
input n1211;
input n1212;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n31;
wire n32;
wire n36;
wire n37;
wire n38;
wire n41;
wire n42;
wire n43;
wire n45;
wire n47;
wire n50;
wire n51;
wire n53;
wire n55;
wire n57;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n97;
wire n98;
wire n99;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n113;
wire n114;
wire n115;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n144;
wire n145;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n193;
wire n194;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n289;
wire n290;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1146;
wire n1147;
wire n1148;
wire n1150;
wire n1152;
wire n1154;
wire n1155;
wire n1158;
wire n1159;
wire n1160;
wire n1162;
wire n1164;
wire n1167;
wire n1168;
wire n1170;
wire n1172;
wire n1174;
wire n1204;
wire n1205;
wire n1208;
wire n1209;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
xor (out,n0,n1221);
and (n0,n1,n1139);
nand (n1,n2,n1138);
or (n2,n3,n662);
nand (n3,n4,n661);
nand (n4,n5,n594);
not (n5,n6);
xor (n6,n7,n507);
xor (n7,n8,n373);
xor (n8,n9,n265);
xor (n9,n10,n168);
or (n10,n11,n167);
and (n11,n12,n133);
xor (n12,n13,n87);
and (n13,n14,n37);
nand (n14,n15,n36);
or (n15,n16,n31);
not (n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n30);
and (s0n17,notn17,n18);
and (s1n17,n30,n29);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,n19);
and (s1n18,n21,n20);
and (n21,n22,n27);
and (n22,n23,n25);
not (n23,n24);
not (n25,n26);
not (n27,n28);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n30);
and (s0n31,notn31,n32);
and (s1n31,n30,n35);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n21);
and (s0n32,notn32,n33);
and (s1n32,n21,n34);
nand (n36,n31,n16);
wire s0n37,s1n37,notn37;
or (n37,s0n37,s1n37);
not(notn37,n50);
and (s0n37,notn37,n38);
and (s1n37,n50,n49);
wire s0n38,s1n38,notn38;
or (n38,s0n38,s1n38);
not(notn38,n41);
and (s0n38,notn38,n39);
and (s1n38,n41,n40);
and (n41,n42,n47);
and (n42,n43,n45);
not (n43,n44);
not (n45,n46);
not (n47,n48);
and (n50,n51,n53);
not (n51,n52);
or (n53,n54,n55);
and (n55,n56,n57);
or (n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86);
nand (n87,n88,n123);
or (n88,n89,n104);
not (n89,n90);
nand (n90,n91,n103);
or (n91,n92,n97);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n30);
and (s0n92,notn92,n93);
and (s1n92,n30,n96);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n21);
and (s0n93,notn93,n94);
and (s1n93,n21,n95);
not (n97,n98);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n50);
and (s0n98,notn98,n99);
and (s1n98,n50,n102);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n41);
and (s0n99,notn99,n100);
and (s1n99,n41,n101);
nand (n103,n97,n92);
nand (n104,n105,n120);
not (n105,n106);
nand (n106,n107,n119);
or (n107,n108,n113);
wire s0n108,s1n108,notn108;
or (n108,s0n108,s1n108);
not(notn108,n30);
and (s0n108,notn108,n109);
and (s1n108,n30,n112);
wire s0n109,s1n109,notn109;
or (n109,s0n109,s1n109);
not(notn109,n21);
and (s0n109,notn109,n110);
and (s1n109,n21,n111);
not (n113,n114);
wire s0n114,s1n114,notn114;
or (n114,s0n114,s1n114);
not(notn114,n30);
and (s0n114,notn114,n115);
and (s1n114,n30,n118);
wire s0n115,s1n115,notn115;
or (n115,s0n115,s1n115);
not(notn115,n21);
and (s0n115,notn115,n116);
and (s1n115,n21,n117);
nand (n119,n113,n108);
nand (n120,n121,n122);
or (n121,n113,n92);
nand (n122,n92,n113);
nand (n123,n124,n106);
nand (n124,n125,n132);
or (n125,n126,n127);
not (n126,n92);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n50);
and (s0n127,notn127,n128);
and (s1n127,n50,n131);
wire s0n128,s1n128,notn128;
or (n128,s0n128,s1n128);
not(notn128,n41);
and (s0n128,notn128,n129);
and (s1n128,n41,n130);
nand (n132,n127,n126);
nand (n133,n134,n157);
or (n134,n135,n150);
not (n135,n136);
nand (n136,n137,n149);
or (n137,n138,n144);
not (n138,n139);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n30);
and (s0n139,notn139,n140);
and (s1n139,n30,n143);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n21);
and (s0n140,notn140,n141);
and (s1n140,n21,n142);
wire s0n144,s1n144,notn144;
or (n144,s0n144,s1n144);
not(notn144,n50);
and (s0n144,notn144,n145);
and (s1n144,n50,n148);
wire s0n145,s1n145,notn145;
or (n145,s0n145,s1n145);
not(notn145,n41);
and (s0n145,notn145,n146);
and (s1n145,n41,n147);
nand (n149,n144,n138);
not (n150,n151);
nor (n151,n138,n152);
wire s0n152,s1n152,notn152;
or (n152,s0n152,s1n152);
not(notn152,n30);
and (s0n152,notn152,n153);
and (s1n152,n30,n156);
wire s0n153,s1n153,notn153;
or (n153,s0n153,s1n153);
not(notn153,n21);
and (s0n153,notn153,n154);
and (s1n153,n21,n155);
nand (n157,n158,n152);
nor (n158,n159,n166);
and (n159,n138,n160);
not (n160,n161);
wire s0n161,s1n161,notn161;
or (n161,s0n161,s1n161);
not(notn161,n50);
and (s0n161,notn161,n162);
and (s1n161,n50,n165);
wire s0n162,s1n162,notn162;
or (n162,s0n162,s1n162);
not(notn162,n41);
and (s0n162,notn162,n163);
and (s1n162,n41,n164);
and (n166,n161,n139);
and (n167,n13,n87);
xor (n168,n169,n226);
xor (n169,n170,n183);
nand (n170,n171,n173);
or (n171,n172,n150);
not (n172,n158);
nand (n173,n174,n152);
nand (n174,n175,n182);
or (n175,n139,n176);
not (n176,n177);
wire s0n177,s1n177,notn177;
or (n177,s0n177,s1n177);
not(notn177,n50);
and (s0n177,notn177,n178);
and (s1n177,n50,n181);
wire s0n178,s1n178,notn178;
or (n178,s0n178,s1n178);
not(notn178,n41);
and (s0n178,notn178,n179);
and (s1n178,n41,n180);
nand (n182,n176,n139);
nand (n183,n184,n210);
or (n184,n185,n200);
nor (n185,n186,n198);
and (n186,n187,n193);
not (n187,n188);
wire s0n188,s1n188,notn188;
or (n188,s0n188,s1n188);
not(notn188,n30);
and (s0n188,notn188,n189);
and (s1n188,n30,n192);
wire s0n189,s1n189,notn189;
or (n189,s0n189,s1n189);
not(notn189,n21);
and (s0n189,notn189,n190);
and (s1n189,n21,n191);
wire s0n193,s1n193,notn193;
or (n193,s0n193,s1n193);
not(notn193,n30);
and (s0n193,notn193,n194);
and (s1n193,n30,n197);
wire s0n194,s1n194,notn194;
or (n194,s0n194,s1n194);
not(notn194,n21);
and (s0n194,notn194,n195);
and (s1n194,n21,n196);
and (n198,n188,n199);
not (n199,n193);
not (n200,n201);
nand (n201,n202,n209);
or (n202,n203,n204);
not (n203,n31);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n50);
and (s0n204,notn204,n205);
and (s1n204,n50,n208);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n41);
and (s0n205,notn205,n206);
and (s1n205,n41,n207);
nand (n209,n204,n203);
nand (n210,n211,n218);
not (n211,n212);
nand (n212,n213,n185);
or (n213,n214,n216);
not (n214,n215);
nand (n215,n31,n199);
not (n216,n217);
nand (n217,n203,n193);
nand (n218,n219,n225);
or (n219,n203,n220);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n50);
and (s0n220,notn220,n221);
and (s1n220,n50,n224);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n41);
and (s0n221,notn221,n222);
and (s1n221,n41,n223);
nand (n225,n220,n203);
nand (n226,n227,n255);
or (n227,n228,n246);
nand (n228,n229,n240);
or (n229,n230,n238);
not (n230,n231);
nand (n231,n188,n232);
not (n232,n233);
wire s0n233,s1n233,notn233;
or (n233,s0n233,s1n233);
not(notn233,n30);
and (s0n233,notn233,n234);
and (s1n233,n30,n237);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n21);
and (s0n234,notn234,n235);
and (s1n234,n21,n236);
not (n238,n239);
nand (n239,n187,n233);
xnor (n240,n241,n233);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n30);
and (s0n241,notn241,n242);
and (s1n241,n30,n245);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n21);
and (s0n242,notn242,n243);
and (s1n242,n21,n244);
not (n246,n247);
nand (n247,n248,n254);
or (n248,n187,n249);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n50);
and (s0n249,notn249,n250);
and (s1n249,n50,n253);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n41);
and (s0n250,notn250,n251);
and (s1n250,n41,n252);
nand (n254,n249,n187);
nand (n255,n256,n264);
nand (n256,n257,n263);
or (n257,n187,n258);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n50);
and (s0n258,notn258,n259);
and (s1n258,n50,n262);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n41);
and (s0n259,notn259,n260);
and (s1n259,n41,n261);
nand (n263,n258,n187);
not (n264,n240);
xor (n265,n266,n339);
xor (n266,n267,n309);
nand (n267,n268,n299);
or (n268,n269,n279);
not (n269,n270);
nand (n270,n271,n278);
or (n271,n108,n272);
not (n272,n273);
wire s0n273,s1n273,notn273;
or (n273,s0n273,s1n273);
not(notn273,n50);
and (s0n273,notn273,n274);
and (s1n273,n50,n277);
wire s0n274,s1n274,notn274;
or (n274,s0n274,s1n274);
not(notn274,n41);
and (s0n274,notn274,n275);
and (s1n274,n41,n276);
nand (n278,n272,n108);
nand (n279,n280,n295);
not (n280,n281);
nand (n281,n282,n294);
or (n282,n283,n289);
not (n283,n284);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n30);
and (s0n284,notn284,n285);
and (s1n284,n30,n288);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n21);
and (s0n285,notn285,n286);
and (s1n285,n21,n287);
wire s0n289,s1n289,notn289;
or (n289,s0n289,s1n289);
not(notn289,n30);
and (s0n289,notn289,n290);
and (s1n289,n30,n293);
wire s0n290,s1n290,notn290;
or (n290,s0n290,s1n290);
not(notn290,n21);
and (s0n290,notn290,n291);
and (s1n290,n21,n292);
nand (n294,n289,n283);
nand (n295,n296,n298);
or (n296,n297,n284);
not (n297,n108);
nand (n298,n297,n284);
nand (n299,n300,n281);
nor (n300,n301,n308);
and (n301,n297,n302);
not (n302,n303);
wire s0n303,s1n303,notn303;
or (n303,s0n303,s1n303);
not(notn303,n50);
and (s0n303,notn303,n304);
and (s1n303,n50,n307);
wire s0n304,s1n304,notn304;
or (n304,s0n304,s1n304);
not(notn304,n41);
and (s0n304,notn304,n305);
and (s1n304,n41,n306);
and (n308,n303,n108);
nand (n309,n310,n335);
or (n310,n311,n326);
not (n311,n312);
nor (n312,n313,n323);
nor (n313,n314,n321);
and (n314,n315,n316);
not (n315,n241);
wire s0n316,s1n316,notn316;
or (n316,s0n316,s1n316);
not(notn316,n30);
and (s0n316,notn316,n317);
and (s1n316,n30,n320);
wire s0n317,s1n317,notn317;
or (n317,s0n317,s1n317);
not(notn317,n21);
and (s0n317,notn317,n318);
and (s1n317,n21,n319);
and (n321,n241,n322);
not (n322,n316);
nand (n323,n324,n325);
or (n324,n322,n92);
nand (n325,n92,n322);
not (n326,n327);
nand (n327,n328,n334);
or (n328,n315,n329);
wire s0n329,s1n329,notn329;
or (n329,s0n329,s1n329);
not(notn329,n50);
and (s0n329,notn329,n330);
and (s1n329,n50,n333);
wire s0n330,s1n330,notn330;
or (n330,s0n330,s1n330);
not(notn330,n41);
and (s0n330,notn330,n331);
and (s1n330,n41,n332);
nand (n334,n329,n315);
nand (n335,n336,n323);
nand (n336,n337,n338);
or (n337,n315,n98);
nand (n338,n98,n315);
nand (n339,n340,n368);
or (n340,n341,n351);
not (n341,n342);
nand (n342,n343,n350);
or (n343,n289,n344);
not (n344,n345);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n50);
and (s0n345,notn345,n346);
and (s1n345,n50,n349);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n41);
and (s0n346,notn346,n347);
and (s1n346,n41,n348);
nand (n350,n344,n289);
nand (n351,n352,n364);
or (n352,n353,n361);
not (n353,n354);
nand (n354,n289,n355);
not (n355,n356);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n30);
and (s0n356,notn356,n357);
and (s1n356,n30,n360);
wire s0n357,s1n357,notn357;
or (n357,s0n357,s1n357);
not(notn357,n21);
and (s0n357,notn357,n358);
and (s1n357,n21,n359);
not (n361,n362);
nand (n362,n363,n356);
not (n363,n289);
not (n364,n365);
nand (n365,n366,n367);
or (n366,n139,n355);
nand (n367,n355,n139);
nand (n368,n365,n369);
nor (n369,n370,n371);
and (n370,n144,n289);
and (n371,n363,n372);
not (n372,n144);
or (n373,n374,n506);
and (n374,n375,n442);
xor (n375,n376,n405);
xor (n376,n377,n398);
xor (n377,n378,n391);
nand (n378,n379,n390);
or (n379,n380,n279);
not (n380,n381);
nand (n381,n382,n389);
or (n382,n108,n383);
not (n383,n384);
wire s0n384,s1n384,notn384;
or (n384,s0n384,s1n384);
not(notn384,n50);
and (s0n384,notn384,n385);
and (s1n384,n50,n388);
wire s0n385,s1n385,notn385;
or (n385,s0n385,s1n385);
not(notn385,n41);
and (s0n385,notn385,n386);
and (s1n385,n41,n387);
nand (n389,n383,n108);
nand (n390,n270,n281);
nand (n391,n392,n397);
or (n392,n311,n393);
not (n393,n394);
nand (n394,n395,n396);
or (n395,n315,n258);
nand (n396,n258,n315);
nand (n397,n327,n323);
nand (n398,n399,n404);
or (n399,n228,n400);
not (n400,n401);
nand (n401,n402,n403);
or (n402,n187,n204);
nand (n403,n204,n187);
nand (n404,n247,n264);
xor (n405,n406,n427);
xor (n406,n407,n420);
nand (n407,n408,n418);
or (n408,n409,n212);
not (n409,n410);
nand (n410,n411,n417);
or (n411,n203,n412);
wire s0n412,s1n412,notn412;
or (n412,s0n412,s1n412);
not(notn412,n50);
and (s0n412,notn412,n413);
and (s1n412,n50,n416);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n41);
and (s0n413,notn413,n414);
and (s1n413,n41,n415);
nand (n417,n412,n203);
nand (n418,n218,n419);
not (n419,n185);
nand (n420,n421,n426);
or (n421,n422,n351);
not (n422,n423);
nand (n423,n424,n425);
or (n424,n363,n303);
nand (n425,n303,n363);
nand (n426,n342,n365);
and (n427,n428,n435);
nor (n428,n429,n203);
and (n429,n430,n433);
nand (n430,n431,n187);
not (n431,n432);
and (n432,n37,n193);
nand (n433,n434,n199);
not (n434,n37);
nand (n435,n436,n441);
or (n436,n104,n437);
not (n437,n438);
nand (n438,n439,n440);
or (n439,n126,n329);
nand (n440,n329,n126);
nand (n441,n90,n106);
or (n442,n443,n505);
and (n443,n444,n470);
xor (n444,n445,n446);
xor (n445,n428,n435);
or (n446,n447,n469);
and (n447,n448,n461);
xor (n448,n449,n450);
nor (n449,n434,n185);
nand (n450,n451,n456);
or (n451,n452,n279);
not (n452,n453);
nand (n453,n454,n455);
or (n454,n297,n98);
nand (n455,n98,n297);
nand (n456,n457,n281);
nand (n457,n458,n460);
or (n458,n108,n459);
not (n459,n127);
nand (n460,n459,n108);
nand (n461,n462,n468);
or (n462,n463,n104);
not (n463,n464);
nand (n464,n465,n467);
or (n465,n92,n466);
not (n466,n258);
nand (n467,n466,n92);
nand (n468,n438,n106);
and (n469,n449,n450);
or (n470,n471,n504);
and (n471,n472,n494);
xor (n472,n473,n483);
nand (n473,n474,n479);
or (n474,n475,n228);
not (n475,n476);
nand (n476,n477,n478);
or (n477,n187,n412);
nand (n478,n187,n412);
nand (n479,n480,n264);
nand (n480,n481,n482);
or (n481,n187,n220);
nand (n482,n220,n187);
nand (n483,n484,n490);
or (n484,n485,n486);
not (n485,n323);
not (n486,n487);
nand (n487,n488,n489);
or (n488,n315,n249);
nand (n489,n249,n315);
nand (n490,n491,n312);
nand (n491,n492,n493);
or (n492,n315,n204);
nand (n493,n204,n315);
nand (n494,n495,n500);
or (n495,n150,n496);
not (n496,n497);
nand (n497,n498,n499);
or (n498,n139,n302);
nand (n499,n302,n139);
nand (n500,n501,n152);
nand (n501,n502,n503);
or (n502,n138,n345);
nand (n503,n345,n138);
and (n504,n473,n483);
and (n505,n445,n446);
and (n506,n376,n405);
xor (n507,n508,n553);
xor (n508,n509,n512);
or (n509,n510,n511);
and (n510,n406,n427);
and (n511,n407,n420);
xor (n512,n513,n550);
xor (n513,n514,n536);
nand (n514,n515,n528);
or (n515,n516,n517);
not (n516,n14);
not (n517,n518);
nor (n518,n519,n525);
and (n519,n412,n520);
wire s0n520,s1n520,notn520;
or (n520,s0n520,s1n520);
not(notn520,n30);
and (s0n520,notn520,n521);
and (s1n520,n30,n524);
wire s0n521,s1n521,notn521;
or (n521,s0n521,s1n521);
not(notn521,n21);
and (s0n521,notn521,n522);
and (s1n521,n21,n523);
and (n525,n526,n527);
not (n526,n520);
not (n527,n412);
nand (n528,n529,n532);
nor (n529,n530,n531);
and (n530,n37,n520);
and (n531,n526,n434);
nor (n532,n14,n533);
nor (n533,n534,n535);
and (n534,n17,n526);
and (n535,n16,n520);
xor (n536,n537,n543);
nor (n537,n538,n526);
and (n538,n539,n542);
nand (n539,n540,n203);
not (n540,n541);
and (n541,n37,n17);
nand (n542,n434,n16);
nand (n543,n544,n546);
or (n544,n545,n104);
not (n545,n124);
nand (n546,n547,n106);
nand (n547,n548,n549);
or (n548,n92,n383);
nand (n549,n383,n92);
or (n550,n551,n552);
and (n551,n377,n398);
and (n552,n378,n391);
or (n553,n554,n593);
and (n554,n555,n592);
xor (n555,n556,n577);
or (n556,n557,n576);
and (n557,n558,n569);
xor (n558,n559,n563);
nand (n559,n560,n562);
or (n560,n561,n228);
not (n561,n480);
nand (n562,n264,n401);
nand (n563,n564,n568);
or (n564,n565,n212);
nor (n565,n566,n567);
and (n566,n31,n434);
and (n567,n203,n37);
nand (n568,n410,n419);
nand (n569,n570,n575);
or (n570,n571,n351);
not (n571,n572);
nand (n572,n573,n574);
or (n573,n363,n273);
nand (n574,n273,n363);
nand (n575,n423,n365);
and (n576,n559,n563);
or (n577,n578,n591);
and (n578,n579,n588);
xor (n579,n580,n584);
nand (n580,n581,n583);
or (n581,n582,n150);
not (n582,n501);
nand (n583,n136,n152);
nand (n584,n585,n587);
nand (n585,n586,n457);
not (n586,n279);
nand (n587,n281,n381);
nand (n588,n589,n590);
or (n589,n311,n486);
nand (n590,n394,n323);
and (n591,n580,n584);
xor (n592,n12,n133);
and (n593,n556,n577);
not (n594,n595);
or (n595,n596,n660);
and (n596,n597,n600);
xor (n597,n598,n599);
xor (n598,n555,n592);
xor (n599,n375,n442);
or (n600,n601,n659);
and (n601,n602,n605);
xor (n602,n603,n604);
xor (n603,n558,n569);
xor (n604,n579,n588);
or (n605,n606,n658);
and (n606,n607,n633);
xor (n607,n608,n615);
nand (n608,n609,n614);
or (n609,n610,n351);
not (n610,n611);
nand (n611,n612,n613);
or (n612,n363,n384);
nand (n613,n384,n363);
nand (n614,n572,n365);
nor (n615,n616,n625);
not (n616,n617);
nand (n617,n618,n624);
or (n618,n619,n279);
not (n619,n620);
nand (n620,n621,n623);
or (n621,n108,n622);
not (n622,n329);
nand (n623,n622,n108);
nand (n624,n453,n281);
nand (n625,n626,n188);
or (n626,n627,n629);
not (n627,n628);
nand (n628,n434,n232);
not (n629,n630);
nand (n630,n631,n315);
not (n631,n632);
and (n632,n37,n233);
or (n633,n634,n657);
and (n634,n635,n650);
xor (n635,n636,n643);
nand (n636,n637,n638);
or (n637,n105,n463);
nand (n638,n639,n642);
nand (n639,n640,n641);
or (n640,n126,n249);
nand (n641,n249,n126);
not (n642,n104);
nand (n643,n644,n649);
or (n644,n645,n228);
not (n645,n646);
nor (n646,n647,n648);
and (n647,n187,n434);
and (n648,n37,n188);
nand (n649,n476,n264);
nand (n650,n651,n653);
or (n651,n485,n652);
not (n652,n491);
nand (n653,n654,n312);
nand (n654,n655,n656);
or (n655,n315,n220);
nand (n656,n220,n315);
and (n657,n636,n643);
and (n658,n608,n615);
and (n659,n603,n604);
and (n660,n598,n599);
nand (n661,n6,n595);
nand (n662,n663,n1128);
or (n663,n664,n814);
not (n664,n665);
nor (n665,n666,n809);
nand (n666,n667,n757);
not (n667,n668);
nor (n668,n669,n701);
xor (n669,n670,n700);
xor (n670,n671,n672);
xor (n671,n444,n470);
or (n672,n673,n699);
and (n673,n674,n677);
xor (n674,n675,n676);
xor (n675,n472,n494);
xor (n676,n448,n461);
or (n677,n678,n698);
and (n678,n679,n694);
xor (n679,n680,n687);
nand (n680,n681,n686);
or (n681,n682,n351);
not (n682,n683);
nand (n683,n684,n685);
or (n684,n363,n127);
nand (n685,n127,n363);
nand (n686,n365,n611);
nand (n687,n688,n693);
or (n688,n689,n150);
not (n689,n690);
nand (n690,n691,n692);
or (n691,n139,n272);
nand (n692,n272,n139);
nand (n693,n497,n152);
nand (n694,n695,n697);
or (n695,n696,n616);
not (n696,n625);
or (n697,n625,n617);
and (n698,n680,n687);
and (n699,n675,n676);
xor (n700,n602,n605);
or (n701,n702,n756);
and (n702,n703,n755);
xor (n703,n704,n705);
xor (n704,n607,n633);
or (n705,n706,n754);
and (n706,n707,n753);
xor (n707,n708,n734);
or (n708,n709,n733);
and (n709,n710,n726);
xor (n710,n711,n718);
nand (n711,n712,n717);
or (n712,n713,n311);
not (n713,n714);
nand (n714,n715,n716);
or (n715,n241,n527);
nand (n716,n527,n241);
nand (n717,n654,n323);
nand (n718,n719,n721);
or (n719,n105,n720);
not (n720,n639);
nand (n721,n642,n722);
nand (n722,n723,n725);
or (n723,n92,n724);
not (n724,n204);
nand (n725,n724,n92);
nand (n726,n727,n732);
or (n727,n728,n351);
not (n728,n729);
nor (n729,n730,n731);
and (n730,n98,n289);
and (n731,n363,n97);
nand (n732,n683,n365);
and (n733,n711,n718);
or (n734,n735,n752);
and (n735,n736,n745);
xor (n736,n737,n738);
nor (n737,n434,n240);
nand (n738,n739,n744);
or (n739,n279,n740);
not (n740,n741);
nand (n741,n742,n743);
or (n742,n108,n466);
nand (n743,n466,n108);
nand (n744,n620,n281);
nand (n745,n746,n751);
or (n746,n747,n150);
not (n747,n748);
nand (n748,n749,n750);
or (n749,n139,n383);
nand (n750,n383,n139);
nand (n751,n690,n152);
and (n752,n737,n738);
xor (n753,n635,n650);
and (n754,n708,n734);
xor (n755,n674,n677);
and (n756,n704,n705);
or (n757,n758,n759);
xor (n758,n703,n755);
or (n759,n760,n808);
and (n760,n761,n764);
xor (n761,n762,n763);
xor (n762,n679,n694);
xor (n763,n707,n753);
or (n764,n765,n807);
and (n765,n766,n806);
xor (n766,n767,n781);
and (n767,n768,n774);
nor (n768,n769,n315);
and (n769,n770,n773);
nand (n770,n771,n126);
not (n771,n772);
and (n772,n37,n316);
nand (n773,n434,n322);
nand (n774,n775,n780);
or (n775,n279,n776);
not (n776,n777);
nand (n777,n778,n779);
or (n778,n297,n249);
nand (n779,n249,n297);
nand (n780,n741,n281);
or (n781,n782,n805);
and (n782,n783,n798);
xor (n783,n784,n791);
nand (n784,n785,n790);
or (n785,n150,n786);
not (n786,n787);
nand (n787,n788,n789);
or (n788,n139,n459);
nand (n789,n459,n139);
nand (n790,n748,n152);
nand (n791,n792,n797);
or (n792,n793,n351);
not (n793,n794);
nand (n794,n795,n796);
or (n795,n363,n329);
nand (n796,n329,n363);
nand (n797,n729,n365);
nand (n798,n799,n804);
or (n799,n800,n104);
not (n800,n801);
nand (n801,n802,n803);
or (n802,n126,n220);
nand (n803,n220,n126);
nand (n804,n722,n106);
and (n805,n784,n791);
xor (n806,n736,n745);
and (n807,n767,n781);
and (n808,n762,n763);
nor (n809,n810,n811);
xor (n810,n597,n600);
or (n811,n812,n813);
and (n812,n670,n700);
and (n813,n671,n672);
not (n814,n815);
nand (n815,n816,n1112,n1118);
nand (n816,n817,n858,n965);
nand (n817,n818,n820);
not (n818,n819);
xor (n819,n761,n764);
not (n820,n821);
or (n821,n822,n857);
and (n822,n823,n856);
xor (n823,n824,n825);
xor (n824,n710,n726);
or (n825,n826,n855);
and (n826,n827,n836);
xor (n827,n828,n835);
nand (n828,n829,n834);
or (n829,n311,n830);
not (n830,n831);
nor (n831,n832,n833);
and (n832,n37,n241);
and (n833,n315,n434);
nand (n834,n323,n714);
xor (n835,n768,n774);
or (n836,n837,n854);
and (n837,n838,n847);
xor (n838,n839,n840);
and (n839,n323,n37);
nand (n840,n841,n846);
or (n841,n351,n842);
not (n842,n843);
nand (n843,n844,n845);
or (n844,n289,n466);
nand (n845,n466,n289);
nand (n846,n794,n365);
nand (n847,n848,n853);
or (n848,n150,n849);
not (n849,n850);
nor (n850,n851,n852);
and (n851,n98,n139);
and (n852,n138,n97);
nand (n853,n787,n152);
and (n854,n839,n840);
and (n855,n828,n835);
xor (n856,n766,n806);
and (n857,n824,n825);
not (n858,n859);
nand (n859,n860,n958);
nor (n860,n861,n928);
nor (n861,n862,n898);
xor (n862,n863,n897);
xor (n863,n864,n865);
xor (n864,n783,n798);
or (n865,n866,n896);
and (n866,n867,n882);
xor (n867,n868,n875);
nand (n868,n869,n874);
or (n869,n870,n104);
not (n870,n871);
nand (n871,n872,n873);
or (n872,n126,n412);
nand (n873,n412,n126);
nand (n874,n801,n106);
nand (n875,n876,n881);
or (n876,n877,n279);
not (n877,n878);
nand (n878,n879,n880);
or (n879,n297,n204);
nand (n880,n204,n297);
nand (n881,n777,n281);
and (n882,n883,n890);
nand (n883,n884,n889);
or (n884,n885,n351);
not (n885,n886);
nand (n886,n887,n888);
or (n887,n363,n249);
nand (n888,n249,n363);
nand (n889,n843,n365);
nor (n890,n891,n126);
and (n891,n892,n895);
nand (n892,n893,n297);
not (n893,n894);
and (n894,n37,n114);
nand (n895,n434,n113);
and (n896,n868,n875);
xor (n897,n827,n836);
or (n898,n899,n927);
and (n899,n900,n926);
xor (n900,n901,n925);
or (n901,n902,n924);
and (n902,n903,n917);
xor (n903,n904,n910);
nand (n904,n905,n909);
nand (n905,n906,n151);
nand (n906,n907,n908);
or (n907,n138,n329);
nand (n908,n329,n138);
nand (n909,n850,n152);
nand (n910,n911,n916);
or (n911,n912,n104);
not (n912,n913);
nand (n913,n914,n915);
or (n914,n92,n434);
or (n915,n37,n126);
nand (n916,n871,n106);
nand (n917,n918,n923);
or (n918,n919,n279);
not (n919,n920);
nand (n920,n921,n922);
or (n921,n297,n220);
nand (n922,n220,n297);
nand (n923,n878,n281);
and (n924,n904,n910);
xor (n925,n838,n847);
xor (n926,n867,n882);
and (n927,n901,n925);
nor (n928,n929,n930);
xor (n929,n900,n926);
or (n930,n931,n957);
and (n931,n932,n956);
xor (n932,n933,n937);
nand (n933,n934,n936);
or (n934,n890,n935);
not (n935,n883);
nand (n936,n935,n890);
or (n937,n938,n955);
and (n938,n939,n948);
xor (n939,n940,n941);
nor (n940,n434,n105);
nand (n941,n942,n947);
or (n942,n943,n351);
not (n943,n944);
nand (n944,n945,n946);
or (n945,n289,n724);
nand (n946,n724,n289);
nand (n947,n886,n365);
nand (n948,n949,n954);
or (n949,n950,n279);
not (n950,n951);
nand (n951,n952,n953);
or (n952,n297,n412);
nand (n953,n412,n297);
nand (n954,n920,n281);
and (n955,n940,n941);
xor (n956,n903,n917);
and (n957,n933,n937);
nand (n958,n959,n961);
not (n959,n960);
xor (n960,n823,n856);
not (n961,n962);
or (n962,n963,n964);
and (n963,n863,n897);
and (n964,n864,n865);
nand (n965,n966,n1111);
or (n966,n967,n998);
not (n967,n968);
nand (n968,n969,n971);
not (n969,n970);
xor (n970,n932,n956);
not (n971,n972);
or (n972,n973,n997);
and (n973,n974,n996);
xor (n974,n975,n982);
nand (n975,n976,n981);
or (n976,n150,n977);
not (n977,n978);
nand (n978,n979,n980);
or (n979,n139,n466);
nand (n980,n139,n466);
nand (n981,n906,n152);
and (n982,n983,n990);
nand (n983,n984,n985);
or (n984,n364,n943);
nand (n985,n986,n987);
not (n986,n351);
nand (n987,n988,n989);
or (n988,n363,n220);
nand (n989,n220,n363);
nor (n990,n991,n297);
and (n991,n992,n995);
nand (n992,n993,n363);
not (n993,n994);
and (n994,n37,n284);
nand (n995,n434,n283);
xor (n996,n939,n948);
and (n997,n975,n982);
not (n998,n999);
nand (n999,n1000,n1110);
or (n1000,n1001,n1029);
not (n1001,n1002);
nand (n1002,n1003,n1005);
not (n1003,n1004);
xor (n1004,n974,n996);
not (n1005,n1006);
or (n1006,n1007,n1028);
and (n1007,n1008,n1024);
xor (n1008,n1009,n1016);
nand (n1009,n1010,n1015);
or (n1010,n1011,n279);
not (n1011,n1012);
nor (n1012,n1013,n1014);
and (n1013,n297,n434);
and (n1014,n37,n108);
nand (n1015,n281,n951);
nand (n1016,n1017,n1019);
or (n1017,n1018,n977);
not (n1018,n152);
nand (n1019,n1020,n151);
nand (n1020,n1021,n1023);
or (n1021,n139,n1022);
not (n1022,n249);
nand (n1023,n139,n1022);
nand (n1024,n1025,n1027);
or (n1025,n990,n1026);
not (n1026,n983);
nand (n1027,n1026,n990);
and (n1028,n1009,n1016);
not (n1029,n1030);
nand (n1030,n1031,n1109);
or (n1031,n1032,n1104);
nor (n1032,n1033,n1103);
and (n1033,n1034,n1070);
nand (n1034,n1035,n1053);
not (n1035,n1036);
xor (n1036,n1037,n1046);
xor (n1037,n1038,n1039);
and (n1038,n281,n37);
nand (n1039,n1040,n1042);
or (n1040,n1018,n1041);
not (n1041,n1020);
nand (n1042,n1043,n151);
nand (n1043,n1044,n1045);
or (n1044,n139,n724);
nand (n1045,n724,n139);
nand (n1046,n1047,n1052);
or (n1047,n1048,n351);
not (n1048,n1049);
nand (n1049,n1050,n1051);
or (n1050,n363,n412);
nand (n1051,n412,n363);
nand (n1052,n987,n365);
nand (n1053,n1054,n1063);
not (n1054,n1055);
nand (n1055,n1056,n289);
or (n1056,n1057,n1059);
not (n1057,n1058);
nand (n1058,n355,n434);
not (n1059,n1060);
nand (n1060,n1061,n138);
not (n1061,n1062);
and (n1062,n37,n356);
nand (n1063,n1064,n1066);
or (n1064,n1018,n1065);
not (n1065,n1043);
nand (n1066,n1067,n151);
nand (n1067,n1068,n1069);
or (n1068,n138,n220);
nand (n1069,n220,n138);
nand (n1070,n1071,n1102);
nand (n1071,n1072,n1083);
or (n1072,n1073,n1076);
nand (n1073,n1074,n1075);
or (n1074,n1055,n1063);
nand (n1075,n1063,n1055);
nand (n1076,n1077,n1082);
or (n1077,n1078,n351);
not (n1078,n1079);
nor (n1079,n1080,n1081);
and (n1080,n363,n434);
and (n1081,n37,n289);
nand (n1082,n365,n1049);
or (n1083,n1084,n1101);
and (n1084,n1085,n1094);
xor (n1085,n1086,n1087);
and (n1086,n37,n365);
nand (n1087,n1088,n1090);
or (n1088,n1018,n1089);
not (n1089,n1067);
nand (n1090,n1091,n151);
nand (n1091,n1092,n1093);
or (n1092,n138,n412);
nand (n1093,n412,n138);
nor (n1094,n1095,n1098);
nor (n1095,n1096,n1097);
and (n1096,n151,n434);
and (n1097,n1091,n152);
nand (n1098,n1099,n139);
not (n1099,n1100);
and (n1100,n37,n152);
and (n1101,n1086,n1087);
nand (n1102,n1073,n1076);
nor (n1103,n1035,n1053);
nor (n1104,n1105,n1106);
xor (n1105,n1008,n1024);
or (n1106,n1107,n1108);
and (n1107,n1037,n1046);
and (n1108,n1038,n1039);
nand (n1109,n1105,n1106);
nand (n1110,n1004,n1006);
nand (n1111,n970,n972);
nand (n1112,n1113,n817);
or (n1113,n1114,n1116);
not (n1114,n1115);
nand (n1115,n960,n962);
not (n1116,n1117);
nand (n1117,n819,n821);
nand (n1118,n817,n1119);
nor (n1119,n1120,n1127);
nand (n1120,n1121,n1126);
or (n1121,n1122,n1124);
not (n1122,n1123);
nand (n1123,n929,n930);
not (n1124,n1125);
nand (n1125,n862,n898);
not (n1126,n861);
not (n1127,n958);
nor (n1128,n1129,n1135);
and (n1129,n1130,n1134);
nand (n1130,n1131,n1133);
or (n1131,n668,n1132);
nand (n1132,n758,n759);
nand (n1133,n669,n701);
not (n1134,n809);
nor (n1135,n1136,n1137);
not (n1136,n810);
not (n1137,n811);
nand (n1138,n662,n3);
xor (n1139,n1140,n1217);
xor (n1140,n1141,n1213);
xor (n1141,n1142,n1204);
and (n1142,n1143,n1154);
wire s0n1143,s1n1143,notn1143;
or (n1143,s0n1143,s1n1143);
not(notn1143,n1146);
and (s0n1143,notn1143,n1144);
and (s1n1143,n1146,n1145);
and (n1146,n1147,n1152);
and (n1147,n1148,n1150);
not (n1148,n1149);
not (n1150,n1151);
not (n1152,n1153);
wire s0n1154,s1n1154,notn1154;
or (n1154,s0n1154,s1n1154);
not(notn1154,n1167);
and (s0n1154,notn1154,n1155);
and (s1n1154,n1167,n1166);
wire s0n1155,s1n1155,notn1155;
or (n1155,s0n1155,s1n1155);
not(notn1155,n1158);
and (s0n1155,notn1155,n1156);
and (s1n1155,n1158,n1157);
and (n1158,n1159,n1164);
and (n1159,n1160,n1162);
not (n1160,n1161);
not (n1162,n1163);
not (n1164,n1165);
and (n1167,n1168,n1170);
not (n1168,n1169);
or (n1170,n1171,n1172);
and (n1172,n1173,n1174);
or (n1174,n1175,n1176,n1177,n1178,n1179,n1180,n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,n1190,n1191,n1192,n1193,n1194,n1195,n1196,n1197,n1198,n1199,n1200,n1201,n1202,n1203);
and (n1204,n1205,n1208);
wire s0n1205,s1n1205,notn1205;
or (n1205,s0n1205,s1n1205);
not(notn1205,n1146);
and (s0n1205,notn1205,n1206);
and (s1n1205,n1146,n1207);
wire s0n1208,s1n1208,notn1208;
or (n1208,s0n1208,s1n1208);
not(notn1208,n1167);
and (s0n1208,notn1208,n1209);
and (s1n1208,n1167,n1212);
wire s0n1209,s1n1209,notn1209;
or (n1209,s0n1209,s1n1209);
not(notn1209,n1158);
and (s0n1209,notn1209,n1210);
and (s1n1209,n1158,n1211);
not (n1213,n1214);
xor (n1214,n1215,n1216);
and (n1215,n140,n37);
and (n1216,n153,n412);
or (n1217,n1218,n1219);
and (n1218,n1205,n1154);
not (n1219,n1220);
and (n1220,n153,n37);
and (n1221,n1139,n1222);
xor (n1222,n1223,n530);
xor (n1223,n1224,n1838);
xor (n1224,n1225,n1837);
xor (n1225,n1226,n1828);
xor (n1226,n1227,n1827);
xor (n1227,n1228,n1813);
xor (n1228,n1229,n1812);
xor (n1229,n1230,n1792);
xor (n1230,n1231,n1791);
xor (n1231,n1232,n1765);
xor (n1232,n1233,n1764);
xor (n1233,n1234,n1732);
xor (n1234,n1235,n1731);
xor (n1235,n1236,n1693);
xor (n1236,n1237,n1692);
xor (n1237,n1238,n1647);
xor (n1238,n1239,n1646);
xor (n1239,n1240,n1596);
xor (n1240,n1241,n1595);
xor (n1241,n1242,n1539);
xor (n1242,n1243,n1538);
xor (n1243,n1244,n1476);
xor (n1244,n1245,n1475);
xor (n1245,n1246,n1408);
xor (n1246,n1247,n1407);
xor (n1247,n1248,n1333);
xor (n1248,n1249,n1332);
xor (n1249,n1250,n1252);
xor (n1250,n1251,n166);
and (n1251,n177,n152);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
and (n1254,n161,n152);
and (n1255,n144,n139);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
and (n1260,n144,n152);
and (n1261,n345,n139);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
and (n1266,n345,n152);
and (n1267,n303,n139);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
and (n1272,n303,n152);
and (n1273,n273,n139);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
and (n1278,n273,n152);
and (n1279,n384,n139);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
and (n1284,n384,n152);
and (n1285,n127,n139);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1291);
and (n1289,n1290,n851);
and (n1290,n127,n152);
and (n1291,n1292,n1293);
xor (n1292,n1290,n851);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
and (n1295,n98,n152);
and (n1296,n329,n139);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
and (n1301,n329,n152);
and (n1302,n258,n139);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
and (n1307,n258,n152);
and (n1308,n249,n139);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
and (n1313,n249,n152);
and (n1314,n204,n139);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
and (n1319,n204,n152);
and (n1320,n220,n139);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
and (n1325,n220,n152);
and (n1326,n412,n139);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
and (n1329,n1330,n1331);
and (n1330,n412,n152);
and (n1331,n37,n139);
and (n1332,n144,n356);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
xor (n1335,n1257,n1258);
and (n1336,n345,n356);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1263,n1264);
and (n1342,n303,n356);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
xor (n1347,n1269,n1270);
and (n1348,n273,n356);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
xor (n1353,n1275,n1276);
and (n1354,n384,n356);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1281,n1282);
and (n1360,n127,n356);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1287,n1288);
and (n1366,n98,n356);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1292,n1293);
and (n1372,n329,n356);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1298,n1299);
and (n1378,n258,n356);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1304,n1305);
and (n1384,n249,n356);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1310,n1311);
and (n1390,n204,n356);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1316,n1317);
and (n1396,n220,n356);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1322,n1323);
and (n1402,n412,n356);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
and (n1405,n1406,n1062);
xor (n1406,n1328,n1329);
and (n1407,n345,n289);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1338,n1339);
and (n1411,n303,n289);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1344,n1345);
and (n1417,n273,n289);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1350,n1351);
and (n1423,n384,n289);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1356,n1357);
and (n1429,n127,n289);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
or (n1432,n1433,n1435);
and (n1433,n1434,n730);
xor (n1434,n1362,n1363);
and (n1435,n1436,n1437);
xor (n1436,n1434,n730);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1368,n1369);
and (n1440,n329,n289);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
or (n1443,n1444,n1447);
and (n1444,n1445,n1446);
xor (n1445,n1374,n1375);
and (n1446,n258,n289);
and (n1447,n1448,n1449);
xor (n1448,n1445,n1446);
or (n1449,n1450,n1453);
and (n1450,n1451,n1452);
xor (n1451,n1380,n1381);
and (n1452,n249,n289);
and (n1453,n1454,n1455);
xor (n1454,n1451,n1452);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1386,n1387);
and (n1458,n204,n289);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1392,n1393);
and (n1464,n220,n289);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1398,n1399);
and (n1470,n412,n289);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
and (n1473,n1474,n1081);
xor (n1474,n1404,n1405);
and (n1475,n303,n284);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1413,n1414);
and (n1479,n273,n284);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1419,n1420);
and (n1485,n384,n284);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1425,n1426);
and (n1491,n127,n284);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1431,n1432);
and (n1497,n98,n284);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1436,n1437);
and (n1503,n329,n284);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1442,n1443);
and (n1509,n258,n284);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1448,n1449);
and (n1515,n249,n284);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1454,n1455);
and (n1521,n204,n284);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1460,n1461);
and (n1527,n220,n284);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1466,n1467);
and (n1533,n412,n284);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
and (n1536,n1537,n994);
xor (n1537,n1472,n1473);
and (n1538,n273,n108);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1481,n1482);
and (n1542,n384,n108);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1487,n1488);
and (n1548,n127,n108);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1493,n1494);
and (n1554,n98,n108);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1499,n1500);
and (n1560,n329,n108);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1505,n1506);
and (n1566,n258,n108);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
or (n1569,n1570,n1573);
and (n1570,n1571,n1572);
xor (n1571,n1511,n1512);
and (n1572,n249,n108);
and (n1573,n1574,n1575);
xor (n1574,n1571,n1572);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1517,n1518);
and (n1578,n204,n108);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1523,n1524);
and (n1584,n220,n108);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1591);
and (n1588,n1589,n1590);
xor (n1589,n1529,n1530);
and (n1590,n412,n108);
and (n1591,n1592,n1593);
xor (n1592,n1589,n1590);
and (n1593,n1594,n1014);
xor (n1594,n1535,n1536);
and (n1595,n384,n114);
or (n1596,n1597,n1600);
and (n1597,n1598,n1599);
xor (n1598,n1544,n1545);
and (n1599,n127,n114);
and (n1600,n1601,n1602);
xor (n1601,n1598,n1599);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1550,n1551);
and (n1605,n98,n114);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1556,n1557);
and (n1611,n329,n114);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1562,n1563);
and (n1617,n258,n114);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
or (n1620,n1621,n1624);
and (n1621,n1622,n1623);
xor (n1622,n1568,n1569);
and (n1623,n249,n114);
and (n1624,n1625,n1626);
xor (n1625,n1622,n1623);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1574,n1575);
and (n1629,n204,n114);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1580,n1581);
and (n1635,n220,n114);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1586,n1587);
and (n1641,n412,n114);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
and (n1644,n1645,n894);
xor (n1645,n1592,n1593);
and (n1646,n127,n92);
or (n1647,n1648,n1651);
and (n1648,n1649,n1650);
xor (n1649,n1601,n1602);
and (n1650,n98,n92);
and (n1651,n1652,n1653);
xor (n1652,n1649,n1650);
or (n1653,n1654,n1657);
and (n1654,n1655,n1656);
xor (n1655,n1607,n1608);
and (n1656,n329,n92);
and (n1657,n1658,n1659);
xor (n1658,n1655,n1656);
or (n1659,n1660,n1663);
and (n1660,n1661,n1662);
xor (n1661,n1613,n1614);
and (n1662,n258,n92);
and (n1663,n1664,n1665);
xor (n1664,n1661,n1662);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n1619,n1620);
and (n1668,n249,n92);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1625,n1626);
and (n1674,n204,n92);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1631,n1632);
and (n1680,n220,n92);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1637,n1638);
and (n1686,n412,n92);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
and (n1689,n1690,n1691);
xor (n1690,n1643,n1644);
and (n1691,n37,n92);
and (n1692,n98,n316);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1652,n1653);
and (n1696,n329,n316);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1658,n1659);
and (n1702,n258,n316);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
or (n1705,n1706,n1709);
and (n1706,n1707,n1708);
xor (n1707,n1664,n1665);
and (n1708,n249,n316);
and (n1709,n1710,n1711);
xor (n1710,n1707,n1708);
or (n1711,n1712,n1715);
and (n1712,n1713,n1714);
xor (n1713,n1670,n1671);
and (n1714,n204,n316);
and (n1715,n1716,n1717);
xor (n1716,n1713,n1714);
or (n1717,n1718,n1721);
and (n1718,n1719,n1720);
xor (n1719,n1676,n1677);
and (n1720,n220,n316);
and (n1721,n1722,n1723);
xor (n1722,n1719,n1720);
or (n1723,n1724,n1727);
and (n1724,n1725,n1726);
xor (n1725,n1682,n1683);
and (n1726,n412,n316);
and (n1727,n1728,n1729);
xor (n1728,n1725,n1726);
and (n1729,n1730,n772);
xor (n1730,n1688,n1689);
and (n1731,n329,n241);
or (n1732,n1733,n1736);
and (n1733,n1734,n1735);
xor (n1734,n1698,n1699);
and (n1735,n258,n241);
and (n1736,n1737,n1738);
xor (n1737,n1734,n1735);
or (n1738,n1739,n1742);
and (n1739,n1740,n1741);
xor (n1740,n1704,n1705);
and (n1741,n249,n241);
and (n1742,n1743,n1744);
xor (n1743,n1740,n1741);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1710,n1711);
and (n1747,n204,n241);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
or (n1750,n1751,n1754);
and (n1751,n1752,n1753);
xor (n1752,n1716,n1717);
and (n1753,n220,n241);
and (n1754,n1755,n1756);
xor (n1755,n1752,n1753);
or (n1756,n1757,n1760);
and (n1757,n1758,n1759);
xor (n1758,n1722,n1723);
and (n1759,n412,n241);
and (n1760,n1761,n1762);
xor (n1761,n1758,n1759);
and (n1762,n1763,n832);
xor (n1763,n1728,n1729);
and (n1764,n258,n233);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1737,n1738);
and (n1768,n249,n233);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1743,n1744);
and (n1774,n204,n233);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1749,n1750);
and (n1780,n220,n233);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1755,n1756);
and (n1786,n412,n233);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
and (n1789,n1790,n632);
xor (n1790,n1761,n1762);
and (n1791,n249,n188);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1770,n1771);
and (n1795,n204,n188);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1776,n1777);
and (n1801,n220,n188);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1782,n1783);
and (n1807,n412,n188);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
and (n1810,n1811,n648);
xor (n1811,n1788,n1789);
and (n1812,n204,n193);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1797,n1798);
and (n1816,n220,n193);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1803,n1804);
and (n1822,n412,n193);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
and (n1825,n1826,n432);
xor (n1826,n1809,n1810);
and (n1827,n220,n31);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1818,n1819);
and (n1831,n412,n31);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
and (n1834,n1835,n1836);
xor (n1835,n1824,n1825);
and (n1836,n37,n31);
and (n1837,n412,n17);
and (n1838,n1839,n541);
xor (n1839,n1833,n1834);
endmodule
