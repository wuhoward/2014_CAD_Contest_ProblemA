module top (out,n6,n25,n28,n29,n37,n38,n44,n45,n50
        ,n58,n60,n61,n70,n71,n81,n96,n97,n100,n106
        ,n128,n129,n136,n244,n245,n253,n310,n316,n365,n376
        ,n382,n392,n398,n405,n410,n774);
output out;
input n6;
input n25;
input n28;
input n29;
input n37;
input n38;
input n44;
input n45;
input n50;
input n58;
input n60;
input n61;
input n70;
input n71;
input n81;
input n96;
input n97;
input n100;
input n106;
input n128;
input n129;
input n136;
input n244;
input n245;
input n253;
input n310;
input n316;
input n365;
input n376;
input n382;
input n392;
input n398;
input n405;
input n410;
input n774;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n406;
wire n407;
wire n408;
wire n409;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
xor (out,n0,n776);
nor (n0,n1,n775);
not (n1,n2);
nand (n2,n3,n774);
nand (n3,n4,n346);
or (n4,n5,n7);
not (n5,n6);
not (n7,n8);
nand (n8,n9,n345);
or (n9,n10,n292);
not (n10,n11);
nor (n11,n12,n290);
and (n12,n13,n233);
or (n13,n14,n232);
and (n14,n15,n148);
xor (n15,n16,n111);
or (n16,n17,n110);
and (n17,n18,n84);
xor (n18,n19,n53);
nand (n19,n20,n47);
or (n20,n21,n31);
not (n21,n22);
nor (n22,n23,n30);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
wire s0n27,s1n27,notn27;
or (n27,s0n27,s1n27);
not(notn27,n6);
and (s0n27,notn27,n28);
and (s1n27,n6,n29);
and (n30,n25,n27);
not (n31,n32);
and (n32,n33,n40);
nand (n33,n34,n39);
or (n34,n35,n27);
not (n35,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n6);
and (s0n36,notn36,n37);
and (s1n36,n6,n38);
nand (n39,n27,n35);
not (n40,n41);
nand (n41,n42,n46);
or (n42,n35,n43);
wire s0n43,s1n43,notn43;
or (n43,s0n43,s1n43);
not(notn43,n6);
and (s0n43,notn43,n44);
and (s1n43,n6,n45);
nand (n46,n43,n35);
nand (n47,n41,n48);
nor (n48,n49,n51);
and (n49,n50,n27);
and (n51,n26,n52);
not (n52,n50);
nand (n53,n54,n73);
or (n54,n55,n65);
not (n55,n56);
nor (n56,n57,n62);
and (n57,n58,n59);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n6);
and (s0n59,notn59,n60);
and (s1n59,n6,n61);
and (n62,n63,n64);
not (n63,n58);
not (n64,n59);
not (n65,n66);
nand (n66,n67,n72);
or (n67,n68,n27);
not (n68,n69);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n6);
and (s0n69,notn69,n70);
and (s1n69,n6,n71);
nand (n72,n27,n68);
nand (n73,n74,n79);
not (n74,n75);
nand (n75,n65,n76);
nand (n76,n77,n78);
or (n77,n68,n59);
nand (n78,n59,n68);
nand (n79,n80,n82);
or (n80,n64,n81);
or (n82,n59,n83);
not (n83,n81);
xor (n84,n85,n90);
and (n85,n86,n59);
nand (n86,n87,n89);
or (n87,n27,n88);
and (n88,n81,n69);
or (n89,n69,n81);
nand (n90,n91,n103);
or (n91,n92,n98);
not (n92,n93);
nor (n93,n94,n95);
not (n94,n43);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n6);
and (s0n95,notn95,n96);
and (s1n95,n6,n97);
nor (n98,n99,n101);
and (n99,n94,n100);
and (n101,n43,n102);
not (n102,n100);
or (n103,n104,n109);
nor (n104,n105,n107);
and (n105,n106,n94);
and (n107,n108,n43);
not (n108,n106);
not (n109,n95);
and (n110,n19,n53);
xor (n111,n112,n120);
xor (n112,n113,n119);
nand (n113,n114,n115);
or (n114,n55,n75);
or (n115,n65,n116);
nor (n116,n117,n118);
and (n117,n64,n25);
and (n118,n59,n24);
and (n119,n85,n90);
xor (n120,n121,n141);
xor (n121,n122,n131);
and (n122,n123,n81);
not (n123,n124);
nor (n124,n125,n130);
and (n125,n126,n59);
not (n126,n127);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n6);
and (s0n127,notn127,n128);
and (s1n127,n6,n129);
and (n130,n127,n64);
nand (n131,n132,n139);
or (n132,n109,n133);
not (n133,n134);
nor (n134,n135,n137);
and (n135,n136,n43);
and (n137,n138,n94);
not (n138,n136);
nand (n139,n140,n93);
not (n140,n104);
nand (n141,n142,n144);
or (n142,n143,n31);
not (n143,n48);
nand (n144,n41,n145);
nand (n145,n146,n147);
or (n146,n27,n102);
or (n147,n26,n100);
or (n148,n149,n231);
and (n149,n150,n171);
xor (n150,n151,n170);
or (n151,n152,n169);
and (n152,n153,n162);
xor (n153,n154,n155);
and (n154,n66,n81);
nand (n155,n156,n161);
or (n156,n157,n31);
not (n157,n158);
nor (n158,n159,n160);
and (n159,n58,n27);
and (n160,n63,n26);
nand (n161,n22,n41);
nand (n162,n163,n168);
or (n163,n92,n164);
not (n164,n165);
nor (n165,n166,n167);
and (n166,n52,n94);
and (n167,n50,n43);
or (n168,n98,n109);
and (n169,n154,n155);
xor (n170,n18,n84);
or (n171,n172,n230);
and (n172,n173,n229);
xor (n173,n174,n188);
nor (n174,n175,n183);
not (n175,n176);
nand (n176,n177,n182);
or (n177,n178,n92);
not (n178,n179);
nand (n179,n180,n181);
or (n180,n24,n43);
nand (n181,n43,n24);
nand (n182,n165,n95);
nand (n183,n184,n27);
nand (n184,n185,n187);
or (n185,n43,n186);
and (n186,n81,n36);
or (n187,n36,n81);
nand (n188,n189,n227);
or (n189,n190,n213);
not (n190,n191);
nand (n191,n192,n212);
or (n192,n193,n202);
nor (n193,n194,n201);
nand (n194,n195,n200);
or (n195,n196,n92);
not (n196,n197);
nand (n197,n198,n199);
or (n198,n63,n43);
nand (n199,n43,n63);
nand (n200,n179,n95);
nor (n201,n40,n83);
nand (n202,n203,n210);
nand (n203,n204,n209);
or (n204,n205,n92);
not (n205,n206);
nand (n206,n207,n208);
or (n207,n94,n81);
or (n208,n43,n83);
nand (n209,n197,n95);
nor (n210,n211,n94);
and (n211,n81,n95);
nand (n212,n194,n201);
not (n213,n214);
nand (n214,n215,n223);
not (n215,n216);
nand (n216,n217,n222);
or (n217,n218,n31);
not (n218,n219);
nand (n219,n220,n221);
or (n220,n26,n81);
or (n221,n27,n83);
nand (n222,n41,n158);
nor (n223,n224,n226);
and (n224,n175,n225);
not (n225,n183);
and (n226,n176,n183);
nand (n227,n228,n216);
not (n228,n223);
xor (n229,n153,n162);
and (n230,n174,n188);
and (n231,n151,n170);
and (n232,n16,n111);
or (n233,n234,n287);
xor (n234,n235,n258);
xor (n235,n236,n255);
xor (n236,n237,n246);
nor (n237,n238,n242);
nor (n238,n239,n241);
and (n239,n64,n240);
nand (n240,n127,n81);
and (n241,n126,n83);
not (n242,n243);
wire s0n243,s1n243,notn243;
or (n243,s0n243,s1n243);
not(notn243,n6);
and (s0n243,notn243,n244);
and (s1n243,n6,n245);
nand (n246,n247,n248);
or (n247,n133,n92);
nand (n248,n249,n95);
not (n249,n250);
nor (n250,n251,n254);
and (n251,n252,n43);
not (n252,n253);
and (n254,n253,n94);
or (n255,n256,n257);
and (n256,n121,n141);
and (n257,n122,n131);
xor (n258,n259,n281);
xor (n259,n260,n274);
nand (n260,n261,n270);
or (n261,n262,n266);
not (n262,n263);
nand (n263,n264,n265);
or (n264,n242,n81);
or (n265,n243,n83);
nand (n266,n124,n267);
nand (n267,n268,n269);
or (n268,n126,n243);
nand (n269,n243,n126);
or (n270,n124,n271);
nor (n271,n272,n273);
and (n272,n58,n242);
and (n273,n63,n243);
nand (n274,n275,n277);
or (n275,n276,n31);
not (n276,n145);
nand (n277,n41,n278);
nor (n278,n279,n280);
and (n279,n106,n27);
and (n280,n108,n26);
nand (n281,n282,n283);
or (n282,n75,n116);
or (n283,n65,n284);
nor (n284,n285,n286);
and (n285,n64,n50);
and (n286,n59,n52);
or (n287,n288,n289);
and (n288,n112,n120);
and (n289,n113,n119);
not (n290,n291);
nand (n291,n234,n287);
not (n292,n293);
nor (n293,n294,n344);
not (n294,n295);
nand (n295,n296,n341);
xor (n296,n297,n325);
xor (n297,n298,n301);
or (n298,n299,n300);
and (n299,n259,n281);
and (n300,n260,n274);
xor (n301,n302,n319);
xor (n302,n303,n311);
and (n303,n304,n81);
not (n304,n305);
nand (n305,n243,n306);
not (n306,n307);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n6);
and (s0n307,notn307,1'b0);
and (s1n307,n6,n309);
and (n309,n310,n245);
nand (n311,n312,n313);
or (n312,n92,n250);
or (n313,n314,n109);
nor (n314,n315,n317);
and (n315,n94,n316);
and (n317,n43,n318);
not (n318,n316);
nand (n319,n320,n321);
or (n320,n266,n271);
or (n321,n124,n322);
nor (n322,n323,n324);
and (n323,n25,n242);
and (n324,n24,n243);
xor (n325,n326,n340);
xor (n326,n327,n334);
nand (n327,n328,n330);
or (n328,n31,n329);
not (n329,n278);
or (n330,n40,n331);
nor (n331,n332,n333);
and (n332,n26,n136);
and (n333,n27,n138);
nand (n334,n335,n336);
or (n335,n75,n284);
or (n336,n65,n337);
nor (n337,n338,n339);
and (n338,n64,n100);
and (n339,n59,n102);
and (n340,n237,n246);
or (n341,n342,n343);
and (n342,n235,n258);
and (n343,n236,n255);
nor (n344,n296,n341);
or (n345,n293,n11);
nand (n346,n347,n5);
xor (n347,n348,n531);
and (n348,n349,n529);
not (n349,n350);
nor (n350,n351,n484);
or (n351,n352,n483);
and (n352,n353,n445);
xor (n353,n354,n385);
xor (n354,n355,n372);
xor (n355,n356,n368);
nand (n356,n357,n362);
or (n357,n358,n266);
not (n358,n359);
nor (n359,n360,n361);
and (n360,n316,n243);
and (n361,n318,n242);
nand (n362,n123,n363);
nor (n363,n364,n366);
and (n364,n365,n243);
and (n366,n367,n242);
not (n367,n365);
nor (n368,n305,n369);
nor (n369,n370,n371);
and (n370,n307,n252);
and (n371,n306,n253);
nand (n372,n373,n379);
or (n373,n75,n374);
nor (n374,n375,n377);
and (n375,n64,n376);
and (n377,n59,n378);
not (n378,n376);
or (n379,n65,n380);
nor (n380,n381,n383);
and (n381,n64,n382);
and (n383,n59,n384);
not (n384,n382);
xor (n385,n386,n425);
xor (n386,n387,n411);
xor (n387,n388,n401);
nand (n388,n389,n395);
or (n389,n92,n390);
nor (n390,n391,n393);
and (n391,n94,n392);
and (n393,n43,n394);
not (n394,n392);
or (n395,n396,n109);
nor (n396,n397,n399);
and (n397,n94,n398);
and (n399,n43,n400);
not (n400,n398);
nand (n401,n402,n408);
or (n402,n31,n403);
nor (n403,n404,n406);
and (n404,n26,n405);
and (n406,n27,n407);
not (n407,n405);
or (n408,n409,n40);
xor (n409,n410,n26);
and (n411,n412,n419);
nand (n412,n413,n418);
or (n413,n92,n414);
nor (n414,n415,n416);
and (n415,n94,n410);
and (n416,n43,n417);
not (n417,n410);
or (n418,n390,n109);
nand (n419,n420,n424);
or (n420,n31,n421);
nor (n421,n422,n423);
and (n422,n26,n382);
and (n423,n27,n384);
or (n424,n40,n403);
or (n425,n426,n444);
and (n426,n427,n438);
xor (n427,n428,n434);
nand (n428,n429,n433);
or (n429,n430,n266);
nor (n430,n431,n432);
and (n431,n253,n242);
and (n432,n252,n243);
nand (n433,n123,n359);
nor (n434,n305,n435);
nor (n435,n436,n437);
and (n436,n307,n138);
and (n437,n306,n136);
nand (n438,n439,n443);
or (n439,n75,n440);
nor (n440,n441,n442);
and (n441,n64,n365);
and (n442,n59,n367);
or (n443,n65,n374);
and (n444,n428,n434);
or (n445,n446,n482);
and (n446,n447,n462);
xor (n447,n448,n449);
xor (n448,n412,n419);
and (n449,n450,n456);
nand (n450,n451,n455);
or (n451,n92,n452);
nor (n452,n453,n454);
and (n453,n94,n405);
and (n454,n43,n407);
or (n455,n414,n109);
nand (n456,n457,n461);
or (n457,n31,n458);
nor (n458,n459,n460);
and (n459,n26,n376);
and (n460,n27,n378);
or (n461,n421,n40);
or (n462,n463,n481);
and (n463,n464,n475);
xor (n464,n465,n471);
nand (n465,n466,n470);
or (n466,n266,n467);
nor (n467,n468,n469);
and (n468,n242,n136);
and (n469,n243,n138);
or (n470,n124,n430);
nor (n471,n305,n472);
nor (n472,n473,n474);
and (n473,n307,n108);
and (n474,n306,n106);
nand (n475,n476,n477);
or (n476,n440,n65);
or (n477,n75,n478);
nor (n478,n479,n480);
and (n479,n64,n316);
and (n480,n59,n318);
and (n481,n465,n471);
and (n482,n448,n449);
and (n483,n354,n385);
xor (n484,n485,n526);
xor (n485,n486,n505);
xor (n486,n487,n499);
xor (n487,n488,n495);
nand (n488,n489,n491);
or (n489,n490,n266);
not (n490,n363);
or (n491,n124,n492);
nor (n492,n493,n494);
and (n493,n242,n376);
and (n494,n243,n378);
nor (n495,n305,n496);
nor (n496,n497,n498);
and (n497,n307,n318);
and (n498,n306,n316);
nand (n499,n500,n501);
or (n500,n75,n380);
or (n501,n65,n502);
nor (n502,n503,n504);
and (n503,n64,n405);
and (n504,n59,n407);
xor (n505,n506,n523);
xor (n506,n507,n522);
xor (n507,n508,n516);
nand (n508,n509,n510);
or (n509,n92,n396);
or (n510,n511,n109);
nor (n511,n512,n514);
and (n512,n94,n513);
and (n513,n310,n398);
and (n514,n43,n515);
not (n515,n513);
nand (n516,n517,n518);
or (n517,n409,n31);
nand (n518,n41,n519);
nand (n519,n520,n521);
or (n520,n27,n394);
or (n521,n26,n392);
and (n522,n388,n401);
or (n523,n524,n525);
and (n524,n355,n372);
and (n525,n356,n368);
or (n526,n527,n528);
and (n527,n386,n425);
and (n528,n387,n411);
not (n529,n530);
and (n530,n351,n484);
nand (n531,n532,n763,n773);
nand (n532,n533,n684);
nand (n533,n534,n678,n683);
nand (n534,n535,n631);
nand (n535,n536,n630);
or (n536,n537,n585);
nor (n537,n538,n584);
and (n538,n539,n294);
not (n539,n540);
nor (n540,n541,n544);
or (n541,n542,n543);
and (n542,n297,n325);
and (n543,n298,n301);
xor (n544,n545,n567);
xor (n545,n546,n564);
xor (n546,n547,n558);
xor (n547,n548,n554);
nand (n548,n549,n550);
or (n549,n322,n266);
nand (n550,n551,n123);
nor (n551,n552,n553);
and (n552,n50,n243);
and (n553,n52,n242);
nor (n554,n305,n555);
nor (n555,n556,n557);
and (n556,n307,n63);
and (n557,n306,n58);
nand (n558,n559,n560);
or (n559,n92,n314);
or (n560,n561,n109);
nor (n561,n562,n563);
and (n562,n94,n365);
and (n563,n43,n367);
or (n564,n565,n566);
and (n565,n326,n340);
and (n566,n327,n334);
xor (n567,n568,n581);
xor (n568,n569,n575);
nand (n569,n570,n571);
or (n570,n75,n337);
or (n571,n65,n572);
nor (n572,n573,n574);
and (n573,n64,n106);
and (n574,n59,n108);
nand (n575,n576,n577);
or (n576,n31,n331);
or (n577,n578,n40);
nor (n578,n579,n580);
and (n579,n26,n253);
and (n580,n27,n252);
or (n581,n582,n583);
and (n582,n302,n319);
and (n583,n303,n311);
and (n584,n541,n544);
nor (n585,n586,n627);
xor (n586,n587,n624);
xor (n587,n588,n607);
xor (n588,n589,n601);
xor (n589,n590,n597);
nand (n590,n591,n593);
or (n591,n592,n266);
not (n592,n551);
nand (n593,n123,n594);
nor (n594,n595,n596);
and (n595,n100,n243);
and (n596,n102,n242);
nor (n597,n305,n598);
nor (n598,n599,n600);
and (n599,n307,n24);
and (n600,n306,n25);
nand (n601,n602,n603);
or (n602,n75,n572);
or (n603,n65,n604);
nor (n604,n605,n606);
and (n605,n64,n136);
and (n606,n59,n138);
xor (n607,n608,n621);
xor (n608,n609,n615);
nand (n609,n610,n611);
or (n610,n92,n561);
or (n611,n612,n109);
nor (n612,n613,n614);
and (n613,n94,n376);
and (n614,n43,n378);
nand (n615,n616,n617);
or (n616,n31,n578);
or (n617,n618,n40);
nor (n618,n619,n620);
and (n619,n26,n316);
and (n620,n27,n318);
or (n621,n622,n623);
and (n622,n547,n558);
and (n623,n548,n554);
or (n624,n625,n626);
and (n625,n568,n581);
and (n626,n569,n575);
or (n627,n628,n629);
and (n628,n545,n567);
and (n629,n546,n564);
nand (n630,n586,n627);
nand (n631,n632,n674);
not (n632,n633);
xor (n633,n634,n673);
xor (n634,n635,n654);
xor (n635,n636,n648);
xor (n636,n637,n644);
nand (n637,n638,n640);
or (n638,n639,n266);
not (n639,n594);
nand (n640,n123,n641);
nor (n641,n642,n643);
and (n642,n106,n243);
and (n643,n108,n242);
nor (n644,n305,n645);
nor (n645,n646,n647);
and (n646,n307,n52);
and (n647,n306,n50);
nand (n648,n649,n650);
or (n649,n75,n604);
or (n650,n65,n651);
nor (n651,n652,n653);
and (n652,n64,n253);
and (n653,n59,n252);
xor (n654,n655,n670);
xor (n655,n656,n669);
xor (n656,n657,n663);
nand (n657,n658,n659);
or (n658,n92,n612);
or (n659,n660,n109);
nor (n660,n661,n662);
and (n661,n94,n382);
and (n662,n43,n384);
nand (n663,n664,n665);
or (n664,n31,n618);
or (n665,n40,n666);
nor (n666,n667,n668);
and (n667,n26,n365);
and (n668,n27,n367);
and (n669,n609,n615);
or (n670,n671,n672);
and (n671,n589,n601);
and (n672,n590,n597);
and (n673,n608,n621);
not (n674,n675);
or (n675,n676,n677);
and (n676,n587,n624);
and (n677,n588,n607);
nand (n678,n631,n679,n682);
nor (n679,n11,n680);
nand (n680,n681,n539);
not (n681,n344);
not (n682,n585);
nand (n683,n633,n675);
nor (n684,n685,n742);
nand (n685,n686,n735);
not (n686,n687);
nor (n687,n688,n726);
xor (n688,n689,n717);
xor (n689,n690,n691);
xor (n690,n464,n475);
xor (n691,n692,n701);
xor (n692,n693,n694);
xor (n693,n450,n456);
and (n694,n695,n698);
nand (n695,n696,n697);
or (n696,n92,n660);
or (n697,n452,n109);
nand (n698,n699,n700);
or (n699,n31,n666);
or (n700,n458,n40);
or (n701,n702,n716);
and (n702,n703,n713);
xor (n703,n704,n709);
nand (n704,n705,n707);
or (n705,n706,n266);
not (n706,n641);
nand (n707,n708,n123);
not (n708,n467);
nor (n709,n305,n710);
nor (n710,n711,n712);
and (n711,n307,n102);
and (n712,n306,n100);
nand (n713,n714,n715);
or (n714,n75,n651);
or (n715,n65,n478);
and (n716,n704,n709);
or (n717,n718,n725);
and (n718,n719,n722);
xor (n719,n720,n721);
xor (n720,n695,n698);
and (n721,n657,n663);
or (n722,n723,n724);
and (n723,n636,n648);
and (n724,n637,n644);
and (n725,n720,n721);
or (n726,n727,n734);
and (n727,n728,n731);
xor (n728,n729,n730);
xor (n729,n703,n713);
xor (n730,n719,n722);
or (n731,n732,n733);
and (n732,n655,n670);
and (n733,n656,n669);
and (n734,n729,n730);
nand (n735,n736,n738);
not (n736,n737);
xor (n737,n728,n731);
not (n738,n739);
or (n739,n740,n741);
and (n740,n634,n673);
and (n741,n635,n654);
nand (n742,n743,n756);
nand (n743,n744,n752);
not (n744,n745);
xor (n745,n746,n749);
xor (n746,n747,n748);
xor (n747,n427,n438);
xor (n748,n447,n462);
or (n749,n750,n751);
and (n750,n692,n701);
and (n751,n693,n694);
not (n752,n753);
or (n753,n754,n755);
and (n754,n689,n717);
and (n755,n690,n691);
nand (n756,n757,n759);
not (n757,n758);
xor (n758,n353,n445);
not (n759,n760);
or (n760,n761,n762);
and (n761,n746,n749);
and (n762,n747,n748);
nand (n763,n764,n756);
nand (n764,n765,n772);
or (n765,n766,n767);
not (n766,n743);
not (n767,n768);
nand (n768,n769,n771);
or (n769,n687,n770);
nand (n770,n737,n739);
nand (n771,n688,n726);
nand (n772,n745,n753);
nand (n773,n760,n758);
nor (n775,n3,n774);
xor (n776,n774,n777);
wire s0n777,s1n777,notn777;
or (n777,s0n777,s1n777);
not(notn777,n6);
and (s0n777,notn777,n778);
and (s1n777,n6,n1451);
xor (n778,n779,n1331);
xor (n779,n780,n1449);
xor (n780,n781,n1326);
xor (n781,n782,n1442);
xor (n782,n783,n1320);
xor (n783,n784,n1430);
xor (n784,n785,n1314);
xor (n785,n786,n1413);
xor (n786,n787,n1308);
xor (n787,n788,n1391);
xor (n788,n789,n1302);
xor (n789,n790,n1364);
xor (n790,n791,n1296);
xor (n791,n792,n1332);
xor (n792,n793,n1290);
xor (n793,n794,n1287);
xor (n794,n795,n1286);
xor (n795,n796,n1239);
xor (n796,n797,n364);
xor (n797,n798,n1182);
xor (n798,n799,n1181);
xor (n799,n800,n1119);
xor (n800,n801,n1118);
xor (n801,n802,n1050);
xor (n802,n803,n1049);
xor (n803,n804,n978);
xor (n804,n805,n977);
xor (n805,n806,n897);
xor (n806,n807,n896);
xor (n807,n808,n811);
xor (n808,n809,n810);
and (n809,n513,n95);
and (n810,n398,n43);
or (n811,n812,n815);
and (n812,n813,n814);
and (n813,n398,n95);
and (n814,n392,n43);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n821);
and (n818,n819,n820);
and (n819,n392,n95);
and (n820,n410,n43);
and (n821,n822,n823);
xor (n822,n819,n820);
or (n823,n824,n827);
and (n824,n825,n826);
and (n825,n410,n95);
and (n826,n405,n43);
and (n827,n828,n829);
xor (n828,n825,n826);
or (n829,n830,n833);
and (n830,n831,n832);
and (n831,n405,n95);
and (n832,n382,n43);
and (n833,n834,n835);
xor (n834,n831,n832);
or (n835,n836,n839);
and (n836,n837,n838);
and (n837,n382,n95);
and (n838,n376,n43);
and (n839,n840,n841);
xor (n840,n837,n838);
or (n841,n842,n845);
and (n842,n843,n844);
and (n843,n376,n95);
and (n844,n365,n43);
and (n845,n846,n847);
xor (n846,n843,n844);
or (n847,n848,n851);
and (n848,n849,n850);
and (n849,n365,n95);
and (n850,n316,n43);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n857);
and (n854,n855,n856);
and (n855,n316,n95);
and (n856,n253,n43);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n862);
and (n860,n861,n135);
and (n861,n253,n95);
and (n862,n863,n864);
xor (n863,n861,n135);
or (n864,n865,n868);
and (n865,n866,n867);
and (n866,n136,n95);
and (n867,n106,n43);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n874);
and (n871,n872,n873);
and (n872,n106,n95);
and (n873,n100,n43);
and (n874,n875,n876);
xor (n875,n872,n873);
or (n876,n877,n879);
and (n877,n878,n167);
and (n878,n100,n95);
and (n879,n880,n881);
xor (n880,n878,n167);
or (n881,n882,n885);
and (n882,n883,n884);
and (n883,n50,n95);
and (n884,n25,n43);
and (n885,n886,n887);
xor (n886,n883,n884);
or (n887,n888,n891);
and (n888,n889,n890);
and (n889,n25,n95);
and (n890,n58,n43);
and (n891,n892,n893);
xor (n892,n889,n890);
and (n893,n894,n895);
and (n894,n58,n95);
and (n895,n81,n43);
and (n896,n392,n36);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n816,n817);
and (n900,n410,n36);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n822,n823);
and (n906,n405,n36);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n828,n829);
and (n912,n382,n36);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
xor (n917,n834,n835);
and (n918,n376,n36);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n925);
and (n922,n923,n924);
xor (n923,n840,n841);
and (n924,n365,n36);
and (n925,n926,n927);
xor (n926,n923,n924);
or (n927,n928,n931);
and (n928,n929,n930);
xor (n929,n846,n847);
and (n930,n316,n36);
and (n931,n932,n933);
xor (n932,n929,n930);
or (n933,n934,n937);
and (n934,n935,n936);
xor (n935,n852,n853);
and (n936,n253,n36);
and (n937,n938,n939);
xor (n938,n935,n936);
or (n939,n940,n943);
and (n940,n941,n942);
xor (n941,n858,n859);
and (n942,n136,n36);
and (n943,n944,n945);
xor (n944,n941,n942);
or (n945,n946,n949);
and (n946,n947,n948);
xor (n947,n863,n864);
and (n948,n106,n36);
and (n949,n950,n951);
xor (n950,n947,n948);
or (n951,n952,n955);
and (n952,n953,n954);
xor (n953,n869,n870);
and (n954,n100,n36);
and (n955,n956,n957);
xor (n956,n953,n954);
or (n957,n958,n961);
and (n958,n959,n960);
xor (n959,n875,n876);
and (n960,n50,n36);
and (n961,n962,n963);
xor (n962,n959,n960);
or (n963,n964,n967);
and (n964,n965,n966);
xor (n965,n880,n881);
and (n966,n25,n36);
and (n967,n968,n969);
xor (n968,n965,n966);
or (n969,n970,n973);
and (n970,n971,n972);
xor (n971,n886,n887);
and (n972,n58,n36);
and (n973,n974,n975);
xor (n974,n971,n972);
and (n975,n976,n186);
xor (n976,n892,n893);
and (n977,n410,n27);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n902,n903);
and (n981,n405,n27);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n908,n909);
and (n987,n382,n27);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n914,n915);
and (n993,n376,n27);
and (n994,n995,n996);
xor (n995,n992,n993);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n920,n921);
and (n999,n365,n27);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n926,n927);
and (n1005,n316,n27);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n932,n933);
and (n1011,n253,n27);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
xor (n1016,n938,n939);
and (n1017,n136,n27);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1023);
and (n1021,n1022,n279);
xor (n1022,n944,n945);
and (n1023,n1024,n1025);
xor (n1024,n1022,n279);
or (n1025,n1026,n1029);
and (n1026,n1027,n1028);
xor (n1027,n950,n951);
and (n1028,n100,n27);
and (n1029,n1030,n1031);
xor (n1030,n1027,n1028);
or (n1031,n1032,n1034);
and (n1032,n1033,n49);
xor (n1033,n956,n957);
and (n1034,n1035,n1036);
xor (n1035,n1033,n49);
or (n1036,n1037,n1039);
and (n1037,n1038,n30);
xor (n1038,n962,n963);
and (n1039,n1040,n1041);
xor (n1040,n1038,n30);
or (n1041,n1042,n1044);
and (n1042,n1043,n159);
xor (n1043,n968,n969);
and (n1044,n1045,n1046);
xor (n1045,n1043,n159);
and (n1046,n1047,n1048);
xor (n1047,n974,n975);
and (n1048,n81,n27);
and (n1049,n405,n69);
or (n1050,n1051,n1054);
and (n1051,n1052,n1053);
xor (n1052,n983,n984);
and (n1053,n382,n69);
and (n1054,n1055,n1056);
xor (n1055,n1052,n1053);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n989,n990);
and (n1059,n376,n69);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
xor (n1064,n995,n996);
and (n1065,n365,n69);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
or (n1068,n1069,n1072);
and (n1069,n1070,n1071);
xor (n1070,n1001,n1002);
and (n1071,n316,n69);
and (n1072,n1073,n1074);
xor (n1073,n1070,n1071);
or (n1074,n1075,n1078);
and (n1075,n1076,n1077);
xor (n1076,n1007,n1008);
and (n1077,n253,n69);
and (n1078,n1079,n1080);
xor (n1079,n1076,n1077);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
xor (n1082,n1013,n1014);
and (n1083,n136,n69);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
xor (n1088,n1019,n1020);
and (n1089,n106,n69);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
xor (n1094,n1024,n1025);
and (n1095,n100,n69);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
xor (n1100,n1030,n1031);
and (n1101,n50,n69);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
xor (n1106,n1035,n1036);
and (n1107,n25,n69);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1114);
and (n1111,n1112,n1113);
xor (n1112,n1040,n1041);
and (n1113,n58,n69);
and (n1114,n1115,n1116);
xor (n1115,n1112,n1113);
and (n1116,n1117,n88);
xor (n1117,n1045,n1046);
and (n1118,n382,n59);
or (n1119,n1120,n1123);
and (n1120,n1121,n1122);
xor (n1121,n1055,n1056);
and (n1122,n376,n59);
and (n1123,n1124,n1125);
xor (n1124,n1121,n1122);
or (n1125,n1126,n1129);
and (n1126,n1127,n1128);
xor (n1127,n1061,n1062);
and (n1128,n365,n59);
and (n1129,n1130,n1131);
xor (n1130,n1127,n1128);
or (n1131,n1132,n1135);
and (n1132,n1133,n1134);
xor (n1133,n1067,n1068);
and (n1134,n316,n59);
and (n1135,n1136,n1137);
xor (n1136,n1133,n1134);
or (n1137,n1138,n1141);
and (n1138,n1139,n1140);
xor (n1139,n1073,n1074);
and (n1140,n253,n59);
and (n1141,n1142,n1143);
xor (n1142,n1139,n1140);
or (n1143,n1144,n1147);
and (n1144,n1145,n1146);
xor (n1145,n1079,n1080);
and (n1146,n136,n59);
and (n1147,n1148,n1149);
xor (n1148,n1145,n1146);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
xor (n1151,n1085,n1086);
and (n1152,n106,n59);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
xor (n1157,n1091,n1092);
and (n1158,n100,n59);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n1097,n1098);
and (n1164,n50,n59);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1103,n1104);
and (n1170,n25,n59);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1176);
and (n1174,n1175,n57);
xor (n1175,n1109,n1110);
and (n1176,n1177,n1178);
xor (n1177,n1175,n57);
and (n1178,n1179,n1180);
xor (n1179,n1115,n1116);
and (n1180,n81,n59);
and (n1181,n376,n127);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1124,n1125);
and (n1185,n365,n127);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1130,n1131);
and (n1191,n316,n127);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1136,n1137);
and (n1197,n253,n127);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1142,n1143);
and (n1203,n136,n127);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1148,n1149);
and (n1209,n106,n127);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1154,n1155);
and (n1215,n100,n127);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1160,n1161);
and (n1221,n50,n127);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1166,n1167);
and (n1227,n25,n127);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1172,n1173);
and (n1233,n58,n127);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
and (n1236,n1237,n1238);
xor (n1237,n1177,n1178);
not (n1238,n240);
or (n1239,n1240,n1242);
and (n1240,n1241,n360);
xor (n1241,n1187,n1188);
and (n1242,n1243,n1244);
xor (n1243,n1241,n360);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1193,n1194);
and (n1247,n253,n243);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1254);
and (n1251,n1252,n1253);
xor (n1252,n1199,n1200);
and (n1253,n136,n243);
and (n1254,n1255,n1256);
xor (n1255,n1252,n1253);
or (n1256,n1257,n1259);
and (n1257,n1258,n642);
xor (n1258,n1205,n1206);
and (n1259,n1260,n1261);
xor (n1260,n1258,n642);
or (n1261,n1262,n1264);
and (n1262,n1263,n595);
xor (n1263,n1211,n1212);
and (n1264,n1265,n1266);
xor (n1265,n1263,n595);
or (n1266,n1267,n1269);
and (n1267,n1268,n552);
xor (n1268,n1217,n1218);
and (n1269,n1270,n1271);
xor (n1270,n1268,n552);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1223,n1224);
and (n1274,n25,n243);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1229,n1230);
and (n1280,n58,n243);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
and (n1283,n1284,n1285);
xor (n1284,n1235,n1236);
and (n1285,n81,n243);
and (n1286,n316,n307);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1243,n1244);
and (n1290,n253,n307);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1249,n1250);
and (n1296,n136,n307);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1255,n1256);
and (n1302,n106,n307);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1260,n1261);
and (n1308,n100,n307);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1265,n1266);
and (n1314,n50,n307);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1270,n1271);
and (n1320,n25,n307);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1276,n1277);
and (n1326,n58,n307);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
and (n1329,n1330,n1331);
xor (n1330,n1282,n1283);
and (n1331,n81,n307);
or (n1332,n1333,n1335);
and (n1333,n1334,n1296);
xor (n1334,n1292,n1293);
and (n1335,n1336,n1337);
xor (n1336,n1334,n1296);
or (n1337,n1338,n1340);
and (n1338,n1339,n1302);
xor (n1339,n1298,n1299);
and (n1340,n1341,n1342);
xor (n1341,n1339,n1302);
or (n1342,n1343,n1345);
and (n1343,n1344,n1308);
xor (n1344,n1304,n1305);
and (n1345,n1346,n1347);
xor (n1346,n1344,n1308);
or (n1347,n1348,n1350);
and (n1348,n1349,n1314);
xor (n1349,n1310,n1311);
and (n1350,n1351,n1352);
xor (n1351,n1349,n1314);
or (n1352,n1353,n1355);
and (n1353,n1354,n1320);
xor (n1354,n1316,n1317);
and (n1355,n1356,n1357);
xor (n1356,n1354,n1320);
or (n1357,n1358,n1360);
and (n1358,n1359,n1326);
xor (n1359,n1322,n1323);
and (n1360,n1361,n1362);
xor (n1361,n1359,n1326);
and (n1362,n1363,n1331);
xor (n1363,n1328,n1329);
or (n1364,n1365,n1367);
and (n1365,n1366,n1302);
xor (n1366,n1336,n1337);
and (n1367,n1368,n1369);
xor (n1368,n1366,n1302);
or (n1369,n1370,n1372);
and (n1370,n1371,n1308);
xor (n1371,n1341,n1342);
and (n1372,n1373,n1374);
xor (n1373,n1371,n1308);
or (n1374,n1375,n1377);
and (n1375,n1376,n1314);
xor (n1376,n1346,n1347);
and (n1377,n1378,n1379);
xor (n1378,n1376,n1314);
or (n1379,n1380,n1382);
and (n1380,n1381,n1320);
xor (n1381,n1351,n1352);
and (n1382,n1383,n1384);
xor (n1383,n1381,n1320);
or (n1384,n1385,n1387);
and (n1385,n1386,n1326);
xor (n1386,n1356,n1357);
and (n1387,n1388,n1389);
xor (n1388,n1386,n1326);
and (n1389,n1390,n1331);
xor (n1390,n1361,n1362);
or (n1391,n1392,n1394);
and (n1392,n1393,n1308);
xor (n1393,n1368,n1369);
and (n1394,n1395,n1396);
xor (n1395,n1393,n1308);
or (n1396,n1397,n1399);
and (n1397,n1398,n1314);
xor (n1398,n1373,n1374);
and (n1399,n1400,n1401);
xor (n1400,n1398,n1314);
or (n1401,n1402,n1404);
and (n1402,n1403,n1320);
xor (n1403,n1378,n1379);
and (n1404,n1405,n1406);
xor (n1405,n1403,n1320);
or (n1406,n1407,n1409);
and (n1407,n1408,n1326);
xor (n1408,n1383,n1384);
and (n1409,n1410,n1411);
xor (n1410,n1408,n1326);
and (n1411,n1412,n1331);
xor (n1412,n1388,n1389);
or (n1413,n1414,n1416);
and (n1414,n1415,n1314);
xor (n1415,n1395,n1396);
and (n1416,n1417,n1418);
xor (n1417,n1415,n1314);
or (n1418,n1419,n1421);
and (n1419,n1420,n1320);
xor (n1420,n1400,n1401);
and (n1421,n1422,n1423);
xor (n1422,n1420,n1320);
or (n1423,n1424,n1426);
and (n1424,n1425,n1326);
xor (n1425,n1405,n1406);
and (n1426,n1427,n1428);
xor (n1427,n1425,n1326);
and (n1428,n1429,n1331);
xor (n1429,n1410,n1411);
or (n1430,n1431,n1433);
and (n1431,n1432,n1320);
xor (n1432,n1417,n1418);
and (n1433,n1434,n1435);
xor (n1434,n1432,n1320);
or (n1435,n1436,n1438);
and (n1436,n1437,n1326);
xor (n1437,n1422,n1423);
and (n1438,n1439,n1440);
xor (n1439,n1437,n1326);
and (n1440,n1441,n1331);
xor (n1441,n1427,n1428);
or (n1442,n1443,n1445);
and (n1443,n1444,n1326);
xor (n1444,n1434,n1435);
and (n1445,n1446,n1447);
xor (n1446,n1444,n1326);
and (n1447,n1448,n1331);
xor (n1448,n1439,n1440);
and (n1449,n1450,n1331);
xor (n1450,n1446,n1447);
xor (n1451,n1330,n1331);
endmodule
