module top (out,n18,n20,n27,n28,n37,n45,n47,n54,n55
        ,n64,n69,n74,n78,n88,n94,n95,n106,n115,n124
        ,n132,n134,n140,n149,n154,n164,n175,n184,n242,n243
        ,n273,n367,n430,n490,n575);
output out;
input n18;
input n20;
input n27;
input n28;
input n37;
input n45;
input n47;
input n54;
input n55;
input n64;
input n69;
input n74;
input n78;
input n88;
input n94;
input n95;
input n106;
input n115;
input n124;
input n132;
input n134;
input n140;
input n149;
input n154;
input n164;
input n175;
input n184;
input n242;
input n243;
input n273;
input n367;
input n430;
input n490;
input n575;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
xor (out,n0,n1542);
nand (n0,n1,n1541);
or (n1,n2,n503);
nand (n2,n3,n502);
not (n3,n4);
nor (n4,n5,n381);
xor (n5,n6,n323);
xor (n6,n7,n190);
xor (n7,n8,n126);
xor (n8,n9,n80);
or (n9,n10,n79);
and (n10,n11,n66);
xor (n11,n12,n39);
nand (n12,n13,n34);
or (n13,n14,n22);
not (n14,n15);
nor (n15,n16,n21);
and (n16,n17,n19);
not (n17,n18);
not (n19,n20);
and (n21,n18,n20);
not (n22,n23);
nor (n23,n24,n30);
nand (n24,n25,n29);
or (n25,n26,n28);
not (n26,n27);
nand (n29,n26,n28);
nor (n30,n31,n32);
and (n31,n19,n28);
and (n32,n20,n33);
not (n33,n28);
nand (n34,n24,n35);
nand (n35,n36,n38);
or (n36,n37,n19);
nand (n38,n19,n37);
nand (n39,n40,n60);
or (n40,n41,n49);
not (n41,n42);
nor (n42,n43,n48);
and (n43,n44,n46);
not (n44,n45);
not (n46,n47);
and (n48,n45,n47);
nand (n49,n50,n57);
not (n50,n51);
nand (n51,n52,n56);
or (n52,n53,n55);
not (n53,n54);
nand (n56,n55,n53);
nand (n57,n58,n59);
or (n58,n55,n46);
nand (n59,n46,n55);
nand (n60,n51,n61);
nor (n61,n62,n65);
and (n62,n63,n46);
not (n63,n64);
and (n65,n64,n47);
nand (n66,n67,n77);
or (n67,n68,n70);
not (n68,n69);
not (n70,n71);
nor (n71,n72,n76);
nand (n72,n73,n75);
or (n73,n46,n74);
nand (n75,n74,n46);
not (n76,n74);
nand (n77,n72,n78);
and (n79,n12,n39);
xor (n80,n81,n117);
xor (n81,n82,n108);
nand (n82,n83,n101);
or (n83,n84,n90);
not (n84,n85);
nand (n85,n86,n89);
or (n86,n87,n54);
not (n87,n88);
or (n89,n88,n53);
nand (n90,n91,n98);
nor (n91,n92,n96);
and (n92,n93,n95);
not (n93,n94);
and (n96,n94,n97);
not (n97,n95);
nor (n98,n99,n100);
and (n99,n93,n53);
and (n100,n94,n54);
nand (n101,n102,n103);
not (n102,n91);
nor (n103,n104,n107);
and (n104,n53,n105);
not (n105,n106);
and (n107,n106,n54);
nand (n108,n109,n111);
or (n109,n110,n22);
not (n110,n35);
nand (n111,n24,n112);
nor (n112,n113,n116);
and (n113,n114,n19);
not (n114,n115);
and (n116,n115,n20);
nand (n117,n118,n120);
or (n118,n49,n119);
not (n119,n61);
or (n120,n50,n121);
nor (n121,n122,n125);
and (n122,n123,n47);
not (n123,n124);
and (n125,n124,n46);
xor (n126,n127,n167);
xor (n127,n128,n143);
nand (n128,n129,n140);
or (n129,n130,n136);
nand (n130,n131,n135);
or (n131,n132,n133);
not (n133,n134);
nand (n135,n132,n133);
nor (n136,n130,n137);
nor (n137,n138,n141);
and (n138,n139,n140);
not (n139,n132);
and (n141,n132,n142);
not (n142,n140);
nand (n143,n144,n160);
or (n144,n145,n151);
not (n145,n146);
nor (n146,n147,n150);
and (n147,n148,n26);
not (n148,n149);
and (n150,n149,n27);
nand (n151,n152,n156);
nand (n152,n153,n155);
or (n153,n154,n26);
nand (n155,n26,n154);
not (n156,n157);
nand (n157,n158,n159);
or (n158,n142,n154);
nand (n159,n154,n142);
nand (n160,n161,n157);
not (n161,n162);
nor (n162,n163,n165);
and (n163,n26,n164);
and (n165,n27,n166);
not (n166,n164);
nand (n167,n168,n186);
or (n168,n169,n180);
not (n169,n170);
and (n170,n171,n177);
not (n171,n172);
nand (n172,n173,n176);
or (n173,n174,n20);
not (n174,n175);
nand (n176,n20,n174);
nand (n177,n178,n179);
nand (n178,n95,n174);
nand (n179,n175,n97);
not (n180,n181);
nor (n181,n182,n185);
and (n182,n183,n97);
not (n183,n184);
and (n185,n184,n95);
or (n186,n171,n187);
nor (n187,n188,n189);
and (n188,n97,n18);
and (n189,n95,n17);
xor (n190,n191,n292);
xor (n191,n192,n231);
xor (n192,n193,n206);
xor (n193,n194,n199);
nand (n194,n195,n197);
or (n195,n196,n70);
not (n196,n78);
or (n197,n198,n44);
not (n198,n72);
not (n199,n200);
nor (n200,n201,n205);
and (n201,n136,n202);
nor (n202,n203,n204);
and (n203,n166,n142);
and (n204,n164,n140);
and (n205,n130,n140);
or (n206,n207,n230);
and (n207,n208,n223);
xor (n208,n209,n216);
nand (n209,n210,n215);
or (n210,n211,n151);
not (n211,n212);
nor (n212,n213,n214);
and (n213,n114,n26);
and (n214,n115,n27);
nand (n215,n157,n146);
nand (n216,n217,n222);
or (n217,n218,n169);
not (n218,n219);
nor (n219,n220,n221);
and (n220,n105,n97);
and (n221,n106,n95);
nand (n222,n172,n181);
nand (n223,n224,n225);
or (n224,n84,n91);
nand (n225,n226,n227);
not (n226,n90);
nor (n227,n228,n229);
and (n228,n123,n53);
and (n229,n124,n54);
and (n230,n209,n216);
or (n231,n232,n291);
and (n232,n233,n267);
xor (n233,n200,n234);
or (n234,n235,n266);
and (n235,n236,n259);
xor (n236,n237,n251);
nand (n237,n238,n134);
or (n238,n239,n245);
nand (n239,n240,n244);
or (n240,n241,n243);
not (n241,n242);
nand (n244,n243,n241);
not (n245,n246);
nand (n246,n247,n248);
not (n247,n239);
nand (n248,n249,n250);
or (n249,n241,n134);
nand (n250,n241,n134);
nand (n251,n252,n258);
or (n252,n253,n257);
not (n253,n254);
nand (n254,n255,n256);
or (n255,n149,n142);
nand (n256,n142,n149);
not (n257,n136);
nand (n258,n202,n130);
nand (n259,n260,n265);
or (n260,n261,n22);
not (n261,n262);
nor (n262,n263,n264);
and (n263,n183,n19);
and (n264,n184,n20);
nand (n265,n24,n15);
and (n266,n237,n251);
or (n267,n268,n290);
and (n268,n269,n282);
xor (n269,n270,n275);
nand (n270,n271,n274);
or (n271,n272,n70);
not (n272,n273);
nand (n274,n72,n69);
nand (n275,n276,n281);
or (n276,n277,n169);
not (n277,n278);
nor (n278,n279,n280);
and (n279,n87,n97);
and (n280,n88,n95);
nand (n281,n172,n219);
nand (n282,n283,n284);
or (n283,n211,n156);
or (n284,n151,n285);
not (n285,n286);
nor (n286,n287,n289);
and (n287,n288,n26);
not (n288,n37);
and (n289,n37,n27);
and (n290,n270,n275);
and (n291,n200,n234);
or (n292,n293,n322);
and (n293,n294,n297);
xor (n294,n295,n296);
xor (n295,n11,n66);
xor (n296,n208,n223);
or (n297,n298,n321);
and (n298,n299,n314);
xor (n299,n300,n307);
nand (n300,n301,n306);
or (n301,n302,n90);
not (n302,n303);
nor (n303,n304,n305);
and (n304,n53,n63);
and (n305,n64,n54);
nand (n306,n102,n227);
nand (n307,n308,n313);
or (n308,n309,n49);
not (n309,n310);
nor (n310,n311,n312);
and (n311,n196,n46);
and (n312,n78,n47);
nand (n313,n51,n42);
not (n314,n315);
nor (n315,n316,n320);
and (n316,n245,n317);
nor (n317,n318,n319);
and (n318,n166,n133);
and (n319,n164,n134);
nor (n320,n247,n133);
and (n321,n300,n307);
and (n322,n295,n296);
or (n323,n324,n380);
and (n324,n325,n379);
xor (n325,n326,n327);
xor (n326,n233,n267);
or (n327,n328,n378);
and (n328,n329,n377);
xor (n329,n330,n354);
or (n330,n331,n353);
and (n331,n332,n347);
xor (n332,n333,n340);
nand (n333,n334,n339);
or (n334,n335,n169);
not (n335,n336);
nand (n336,n337,n338);
or (n337,n124,n97);
nand (n338,n97,n124);
nand (n339,n278,n172);
nand (n340,n341,n346);
or (n341,n342,n151);
not (n342,n343);
nor (n343,n344,n345);
and (n344,n17,n26);
and (n345,n18,n27);
nand (n346,n157,n286);
nand (n347,n348,n349);
or (n348,n91,n302);
or (n349,n90,n350);
nor (n350,n351,n352);
and (n351,n45,n53);
and (n352,n54,n44);
and (n353,n333,n340);
or (n354,n355,n376);
and (n355,n356,n369);
xor (n356,n357,n364);
nand (n357,n358,n363);
or (n358,n359,n257);
not (n359,n360);
nor (n360,n361,n362);
and (n361,n114,n142);
and (n362,n115,n140);
nand (n363,n130,n254);
nand (n364,n365,n368);
or (n365,n366,n70);
not (n366,n367);
nand (n368,n72,n273);
nand (n369,n370,n375);
or (n370,n371,n22);
not (n371,n372);
nor (n372,n373,n374);
and (n373,n105,n19);
and (n374,n106,n20);
nand (n375,n24,n262);
and (n376,n357,n364);
xor (n377,n236,n259);
and (n378,n330,n354);
xor (n379,n294,n297);
and (n380,n326,n327);
or (n381,n382,n501);
and (n382,n383,n410);
xor (n383,n384,n409);
or (n384,n385,n408);
and (n385,n386,n389);
xor (n386,n387,n388);
xor (n387,n269,n282);
xor (n388,n299,n314);
or (n389,n390,n407);
and (n390,n391,n399);
xor (n391,n392,n315);
nand (n392,n393,n398);
or (n393,n394,n49);
not (n394,n395);
nor (n395,n396,n397);
and (n396,n68,n46);
and (n397,n69,n47);
nand (n398,n51,n310);
nand (n399,n400,n243);
nor (n400,n401,n406);
and (n401,n402,n403);
not (n402,n151);
nand (n403,n404,n405);
or (n404,n184,n26);
nand (n405,n26,n184);
and (n406,n157,n343);
and (n407,n392,n315);
and (n408,n387,n388);
xor (n409,n325,n379);
or (n410,n411,n500);
and (n411,n412,n464);
xor (n412,n413,n414);
xor (n413,n329,n377);
or (n414,n415,n463);
and (n415,n416,n462);
xor (n416,n417,n439);
or (n417,n418,n438);
and (n418,n419,n432);
xor (n419,n420,n427);
nand (n420,n421,n426);
or (n421,n422,n49);
not (n422,n423);
nand (n423,n424,n425);
or (n424,n272,n47);
nand (n425,n47,n272);
nand (n426,n395,n51);
nand (n427,n428,n431);
or (n428,n429,n70);
not (n429,n430);
nand (n431,n72,n367);
nand (n432,n433,n435);
or (n433,n434,n247);
not (n434,n317);
or (n435,n246,n436);
not (n436,n437);
xor (n437,n148,n133);
and (n438,n420,n427);
or (n439,n440,n461);
and (n440,n441,n455);
xor (n441,n442,n449);
nand (n442,n443,n448);
or (n443,n444,n22);
not (n444,n445);
nor (n445,n446,n447);
and (n446,n87,n19);
and (n447,n88,n20);
nand (n448,n24,n372);
nand (n449,n450,n454);
or (n450,n451,n257);
nor (n451,n452,n453);
and (n452,n288,n140);
and (n453,n37,n142);
nand (n454,n360,n130);
nand (n455,n456,n460);
or (n456,n169,n457);
nor (n457,n458,n459);
and (n458,n63,n95);
and (n459,n64,n97);
or (n460,n171,n335);
and (n461,n442,n449);
xor (n462,n332,n347);
and (n463,n417,n439);
or (n464,n465,n499);
and (n465,n466,n469);
xor (n466,n467,n468);
xor (n467,n356,n369);
xor (n468,n391,n399);
and (n469,n470,n493);
or (n470,n471,n492);
and (n471,n472,n487);
xor (n472,n473,n480);
nand (n473,n474,n479);
or (n474,n475,n151);
not (n475,n476);
nor (n476,n477,n478);
and (n477,n105,n26);
and (n478,n106,n27);
nand (n479,n403,n157);
nand (n480,n481,n486);
or (n481,n482,n49);
not (n482,n483);
nand (n483,n484,n485);
or (n484,n367,n46);
nand (n485,n367,n46);
nand (n486,n51,n423);
nand (n487,n488,n491);
or (n488,n489,n70);
not (n489,n490);
nand (n491,n72,n430);
and (n492,n473,n480);
nand (n493,n494,n498);
or (n494,n90,n495);
nor (n495,n496,n497);
and (n496,n53,n78);
and (n497,n54,n196);
or (n498,n91,n350);
and (n499,n467,n468);
and (n500,n413,n414);
and (n501,n384,n409);
nand (n502,n5,n381);
nand (n503,n504,n1536);
or (n504,n505,n680);
not (n505,n506);
nor (n506,n507,n587);
nor (n507,n508,n509);
xor (n508,n383,n410);
or (n509,n510,n586);
and (n510,n511,n514);
xor (n511,n512,n513);
xor (n512,n386,n389);
xor (n513,n412,n464);
or (n514,n515,n585);
and (n515,n516,n549);
xor (n516,n517,n518);
xor (n517,n416,n462);
or (n518,n519,n548);
and (n519,n520,n546);
xor (n520,n521,n545);
or (n521,n522,n544);
and (n522,n523,n538);
xor (n523,n524,n531);
nand (n524,n525,n530);
or (n525,n526,n246);
not (n526,n527);
nor (n527,n528,n529);
and (n528,n114,n133);
and (n529,n115,n134);
nand (n530,n239,n437);
nand (n531,n532,n537);
or (n532,n533,n22);
not (n533,n534);
nor (n534,n535,n536);
and (n535,n123,n19);
and (n536,n124,n20);
nand (n537,n24,n445);
nand (n538,n539,n542);
or (n539,n257,n540);
not (n540,n541);
xor (n541,n17,n142);
or (n542,n451,n543);
not (n543,n130);
and (n544,n524,n531);
xor (n545,n441,n455);
nand (n546,n547,n399);
or (n547,n243,n400);
and (n548,n521,n545);
or (n549,n550,n584);
and (n550,n551,n583);
xor (n551,n552,n553);
xor (n552,n419,n432);
or (n553,n554,n582);
and (n554,n555,n571);
xor (n555,n556,n564);
nand (n556,n557,n562);
or (n557,n558,n169);
not (n558,n559);
nand (n559,n560,n561);
or (n560,n95,n44);
or (n561,n97,n45);
nand (n562,n563,n172);
not (n563,n457);
nand (n564,n565,n570);
or (n565,n566,n90);
not (n566,n567);
nand (n567,n568,n569);
or (n568,n54,n68);
or (n569,n53,n69);
or (n570,n91,n495);
nand (n571,n572,n581);
or (n572,n573,n576);
nand (n573,n574,n243);
not (n574,n575);
not (n576,n577);
nor (n577,n578,n580);
and (n578,n166,n579);
not (n579,n243);
and (n580,n164,n243);
or (n581,n579,n574);
and (n582,n556,n564);
xor (n583,n493,n470);
and (n584,n552,n553);
and (n585,n517,n518);
and (n586,n512,n513);
nor (n587,n588,n589);
xor (n588,n511,n514);
or (n589,n590,n679);
and (n590,n591,n678);
xor (n591,n592,n593);
xor (n592,n466,n469);
or (n593,n594,n677);
and (n594,n595,n676);
xor (n595,n596,n669);
or (n596,n597,n668);
and (n597,n598,n642);
xor (n598,n599,n617);
or (n599,n600,n616);
and (n600,n601,n609);
xor (n601,n602,n603);
and (n602,n72,n490);
nand (n603,n604,n608);
or (n604,n573,n605);
nor (n605,n606,n607);
and (n606,n148,n243);
and (n607,n149,n579);
nand (n608,n577,n575);
nand (n609,n610,n615);
or (n610,n611,n246);
not (n611,n612);
nor (n612,n613,n614);
and (n613,n288,n133);
and (n614,n37,n134);
nand (n615,n239,n527);
and (n616,n602,n603);
or (n617,n618,n641);
and (n618,n619,n634);
xor (n619,n620,n627);
nand (n620,n621,n626);
or (n621,n622,n257);
not (n622,n623);
nor (n623,n624,n625);
and (n624,n183,n142);
and (n625,n184,n140);
nand (n626,n541,n130);
nand (n627,n628,n629);
or (n628,n171,n558);
nand (n629,n630,n170);
not (n630,n631);
nor (n631,n632,n633);
and (n632,n78,n97);
and (n633,n196,n95);
nand (n634,n635,n636);
or (n635,n566,n91);
nand (n636,n637,n226);
not (n637,n638);
nor (n638,n639,n640);
and (n639,n273,n53);
and (n640,n54,n272);
and (n641,n620,n627);
or (n642,n643,n667);
and (n643,n644,n659);
xor (n644,n645,n652);
nand (n645,n646,n651);
or (n646,n647,n49);
not (n647,n648);
nor (n648,n649,n650);
and (n649,n429,n46);
and (n650,n430,n47);
nand (n651,n483,n51);
nand (n652,n653,n658);
or (n653,n654,n151);
not (n654,n655);
nand (n655,n656,n657);
or (n656,n27,n87);
or (n657,n26,n88);
nand (n658,n157,n476);
nand (n659,n660,n665);
or (n660,n22,n661);
not (n661,n662);
nor (n662,n663,n664);
and (n663,n63,n19);
and (n664,n64,n20);
or (n665,n666,n533);
not (n666,n24);
and (n667,n645,n652);
and (n668,n599,n617);
or (n669,n670,n675);
and (n670,n671,n674);
xor (n671,n672,n673);
xor (n672,n472,n487);
xor (n673,n523,n538);
xor (n674,n555,n571);
and (n675,n672,n673);
xor (n676,n520,n546);
and (n677,n596,n669);
xor (n678,n516,n549);
and (n679,n592,n593);
not (n680,n681);
nand (n681,n682,n1521);
or (n682,n683,n1451);
not (n683,n684);
nand (n684,n685,n1438);
or (n685,n686,n1139);
not (n686,n687);
nand (n687,n688,n1128,n1138);
nand (n688,n689,n916,n994);
nor (n689,n690,n854);
not (n690,n691);
or (n691,n692,n817);
xor (n692,n693,n777);
xor (n693,n694,n724);
xor (n694,n695,n715);
xor (n695,n696,n706);
nand (n696,n697,n702);
or (n697,n698,n22);
not (n698,n699);
nor (n699,n700,n701);
and (n700,n429,n19);
and (n701,n430,n20);
nand (n702,n24,n703);
nand (n703,n704,n705);
or (n704,n20,n366);
or (n705,n19,n367);
nand (n706,n707,n711);
or (n707,n708,n573);
nor (n708,n709,n710);
and (n709,n579,n88);
and (n710,n243,n87);
or (n711,n712,n574);
nor (n712,n713,n714);
and (n713,n579,n106);
and (n714,n243,n105);
nand (n715,n716,n720);
or (n716,n257,n717);
nor (n717,n718,n719);
and (n718,n142,n78);
and (n719,n140,n196);
or (n720,n721,n543);
nor (n721,n722,n723);
and (n722,n142,n45);
and (n723,n140,n44);
or (n724,n725,n776);
and (n725,n726,n751);
xor (n726,n727,n733);
nand (n727,n728,n732);
or (n728,n257,n729);
nor (n729,n730,n731);
and (n730,n142,n69);
and (n731,n140,n68);
or (n732,n543,n717);
xor (n733,n734,n740);
and (n734,n735,n20);
nand (n735,n736,n737);
or (n736,n490,n28);
nand (n737,n738,n26);
not (n738,n739);
and (n739,n490,n28);
nand (n740,n741,n746);
or (n741,n742,n247);
not (n742,n743);
nand (n743,n744,n745);
or (n744,n134,n63);
or (n745,n133,n64);
nand (n746,n747,n245);
not (n747,n748);
nor (n748,n749,n750);
and (n749,n133,n45);
and (n750,n134,n44);
or (n751,n752,n775);
and (n752,n753,n765);
xor (n753,n754,n755);
and (n754,n24,n490);
nand (n755,n756,n761);
or (n756,n574,n757);
not (n757,n758);
nor (n758,n759,n760);
and (n759,n123,n579);
and (n760,n124,n243);
or (n761,n762,n573);
nor (n762,n763,n764);
and (n763,n579,n64);
and (n764,n243,n63);
nand (n765,n766,n770);
or (n766,n151,n767);
nor (n767,n768,n769);
and (n768,n26,n430);
and (n769,n27,n429);
or (n770,n156,n771);
not (n771,n772);
nor (n772,n773,n774);
and (n773,n367,n27);
and (n774,n366,n26);
and (n775,n754,n755);
and (n776,n727,n733);
xor (n777,n778,n800);
xor (n778,n779,n780);
and (n779,n734,n740);
or (n780,n781,n799);
and (n781,n782,n796);
xor (n782,n783,n789);
nand (n783,n784,n785);
or (n784,n771,n151);
nand (n785,n157,n786);
nor (n786,n787,n788);
and (n787,n272,n26);
and (n788,n273,n27);
nand (n789,n790,n795);
or (n790,n791,n22);
not (n791,n792);
nand (n792,n793,n794);
or (n793,n19,n490);
or (n794,n489,n20);
nand (n795,n24,n699);
nand (n796,n797,n798);
or (n797,n573,n757);
or (n798,n708,n574);
and (n799,n783,n789);
xor (n800,n801,n809);
xor (n801,n802,n803);
and (n802,n172,n490);
nand (n803,n804,n805);
or (n804,n742,n246);
nand (n805,n239,n806);
nand (n806,n807,n808);
or (n807,n134,n123);
or (n808,n133,n124);
nand (n809,n810,n812);
or (n810,n811,n151);
not (n811,n786);
nand (n812,n813,n157);
not (n813,n814);
nor (n814,n815,n816);
and (n815,n26,n69);
and (n816,n27,n68);
or (n817,n818,n853);
and (n818,n819,n852);
xor (n819,n820,n821);
xor (n820,n782,n796);
or (n821,n822,n851);
and (n822,n823,n836);
xor (n823,n824,n830);
nand (n824,n825,n829);
or (n825,n246,n826);
nor (n826,n827,n828);
and (n827,n133,n78);
and (n828,n134,n196);
or (n829,n247,n748);
nand (n830,n831,n835);
or (n831,n257,n832);
nor (n832,n833,n834);
and (n833,n142,n273);
and (n834,n140,n272);
or (n835,n729,n543);
and (n836,n837,n844);
nor (n837,n838,n26);
nor (n838,n839,n842);
and (n839,n840,n142);
not (n840,n841);
and (n841,n490,n154);
and (n842,n489,n843);
not (n843,n154);
nand (n844,n845,n850);
or (n845,n846,n573);
not (n846,n847);
nor (n847,n848,n849);
and (n848,n44,n579);
and (n849,n45,n243);
or (n850,n762,n574);
and (n851,n824,n830);
xor (n852,n726,n751);
and (n853,n820,n821);
nand (n854,n855,n910);
not (n855,n856);
nor (n856,n857,n885);
xor (n857,n858,n884);
xor (n858,n859,n883);
or (n859,n860,n882);
and (n860,n861,n876);
xor (n861,n862,n870);
nand (n862,n863,n868);
or (n863,n864,n151);
not (n864,n865);
nand (n865,n866,n867);
or (n866,n26,n490);
or (n867,n27,n489);
nand (n868,n869,n157);
not (n869,n767);
nand (n870,n871,n875);
or (n871,n246,n872);
nor (n872,n873,n874);
and (n873,n133,n69);
and (n874,n134,n68);
or (n875,n826,n247);
nand (n876,n877,n881);
or (n877,n257,n878);
nor (n878,n879,n880);
and (n879,n142,n367);
and (n880,n140,n366);
or (n881,n832,n543);
and (n882,n862,n870);
xor (n883,n753,n765);
xor (n884,n823,n836);
or (n885,n886,n909);
and (n886,n887,n908);
xor (n887,n888,n889);
xor (n888,n837,n844);
or (n889,n890,n907);
and (n890,n891,n900);
xor (n891,n892,n893);
and (n892,n157,n490);
nand (n893,n894,n899);
or (n894,n573,n895);
not (n895,n896);
nor (n896,n897,n898);
and (n897,n78,n243);
and (n898,n196,n579);
nand (n899,n847,n575);
nand (n900,n901,n906);
or (n901,n246,n902);
not (n902,n903);
nor (n903,n904,n905);
and (n904,n272,n133);
and (n905,n273,n134);
or (n906,n247,n872);
and (n907,n892,n893);
xor (n908,n861,n876);
and (n909,n888,n889);
not (n910,n911);
nor (n911,n912,n913);
xor (n912,n819,n852);
or (n913,n914,n915);
and (n914,n858,n884);
and (n915,n859,n883);
nand (n916,n917,n990);
not (n917,n918);
xor (n918,n919,n987);
xor (n919,n920,n957);
xor (n920,n921,n939);
xor (n921,n922,n933);
nand (n922,n923,n928);
or (n923,n924,n171);
not (n924,n925);
nand (n925,n926,n927);
or (n926,n95,n429);
or (n927,n97,n430);
nand (n928,n929,n170);
not (n929,n930);
nor (n930,n931,n932);
and (n931,n489,n95);
and (n932,n97,n490);
nand (n933,n934,n935);
or (n934,n257,n721);
or (n935,n543,n936);
nor (n936,n937,n938);
and (n937,n142,n64);
and (n938,n140,n63);
nand (n939,n940,n956);
or (n940,n941,n948);
not (n941,n942);
nand (n942,n943,n95);
nand (n943,n944,n945);
or (n944,n490,n175);
nand (n945,n946,n19);
not (n946,n947);
and (n947,n490,n175);
not (n948,n949);
nand (n949,n950,n952);
or (n950,n951,n246);
not (n951,n806);
nand (n952,n239,n953);
nor (n953,n954,n955);
and (n954,n87,n133);
and (n955,n88,n134);
or (n956,n949,n942);
xor (n957,n958,n965);
xor (n958,n959,n962);
or (n959,n960,n961);
and (n960,n801,n809);
and (n961,n802,n803);
or (n962,n963,n964);
and (n963,n695,n715);
and (n964,n696,n706);
xor (n965,n966,n980);
xor (n966,n967,n973);
nand (n967,n968,n969);
or (n968,n151,n814);
or (n969,n970,n156);
nor (n970,n971,n972);
and (n971,n26,n78);
and (n972,n27,n196);
nand (n973,n974,n979);
or (n974,n975,n666);
not (n975,n976);
nand (n976,n977,n978);
or (n977,n272,n20);
or (n978,n19,n273);
nand (n979,n23,n703);
nand (n980,n981,n982);
or (n981,n712,n573);
or (n982,n983,n574);
not (n983,n984);
nor (n984,n985,n986);
and (n985,n183,n579);
and (n986,n184,n243);
or (n987,n988,n989);
and (n988,n778,n800);
and (n989,n779,n780);
not (n990,n991);
or (n991,n992,n993);
and (n992,n693,n777);
and (n993,n694,n724);
or (n994,n995,n1127);
and (n995,n996,n1024);
xor (n996,n997,n1023);
or (n997,n998,n1022);
and (n998,n999,n1021);
xor (n999,n1000,n1007);
nand (n1000,n1001,n1006);
or (n1001,n257,n1002);
not (n1002,n1003);
nor (n1003,n1004,n1005);
and (n1004,n430,n140);
and (n1005,n429,n142);
or (n1006,n878,n543);
and (n1007,n1008,n1014);
nor (n1008,n1009,n142);
nor (n1009,n1010,n1013);
and (n1010,n1011,n133);
not (n1011,n1012);
and (n1012,n490,n132);
and (n1013,n489,n139);
nand (n1014,n1015,n1016);
or (n1015,n574,n895);
nand (n1016,n1017,n1020);
nand (n1017,n1018,n1019);
or (n1018,n69,n579);
nand (n1019,n579,n69);
not (n1020,n573);
xor (n1021,n891,n900);
and (n1022,n1000,n1007);
xor (n1023,n887,n908);
or (n1024,n1025,n1126);
and (n1025,n1026,n1045);
xor (n1026,n1027,n1044);
or (n1027,n1028,n1043);
and (n1028,n1029,n1042);
xor (n1029,n1030,n1035);
nand (n1030,n1031,n1034);
or (n1031,n1032,n246);
not (n1032,n1033);
xor (n1033,n366,n133);
nand (n1034,n239,n903);
nand (n1035,n1036,n1041);
or (n1036,n1037,n257);
not (n1037,n1038);
nand (n1038,n1039,n1040);
or (n1039,n142,n490);
or (n1040,n489,n140);
nand (n1041,n1003,n130);
xor (n1042,n1008,n1014);
and (n1043,n1030,n1035);
xor (n1044,n999,n1021);
or (n1045,n1046,n1125);
and (n1046,n1047,n1069);
xor (n1047,n1048,n1068);
or (n1048,n1049,n1067);
and (n1049,n1050,n1059);
xor (n1050,n1051,n1052);
and (n1051,n130,n490);
nand (n1052,n1053,n1058);
or (n1053,n1054,n246);
not (n1054,n1055);
nor (n1055,n1056,n1057);
and (n1056,n429,n133);
and (n1057,n430,n134);
nand (n1058,n239,n1033);
nand (n1059,n1060,n1065);
or (n1060,n573,n1061);
not (n1061,n1062);
nand (n1062,n1063,n1064);
or (n1063,n273,n579);
nand (n1064,n579,n273);
or (n1065,n1066,n574);
not (n1066,n1017);
and (n1067,n1051,n1052);
xor (n1068,n1029,n1042);
nand (n1069,n1070,n1124);
or (n1070,n1071,n1086);
nor (n1071,n1072,n1073);
xor (n1072,n1050,n1059);
nor (n1073,n1074,n1081);
not (n1074,n1075);
nand (n1075,n1076,n1080);
or (n1076,n573,n1077);
nor (n1077,n1078,n1079);
and (n1078,n366,n243);
and (n1079,n367,n579);
nand (n1080,n1062,n575);
nand (n1081,n1082,n134);
nand (n1082,n1083,n1085);
or (n1083,n1084,n243);
and (n1084,n490,n242);
or (n1085,n490,n242);
nor (n1086,n1087,n1123);
and (n1087,n1088,n1099);
nand (n1088,n1089,n1093);
nor (n1089,n1090,n1091);
and (n1090,n1081,n1075);
and (n1091,n1092,n1074);
not (n1092,n1081);
nor (n1093,n1094,n1098);
and (n1094,n245,n1095);
nand (n1095,n1096,n1097);
or (n1096,n133,n490);
or (n1097,n489,n134);
and (n1098,n239,n1055);
nand (n1099,n1100,n1122);
or (n1100,n1101,n1116);
not (n1101,n1102);
nor (n1102,n1103,n1114);
not (n1103,n1104);
nand (n1104,n1105,n1110);
or (n1105,n574,n1106);
not (n1106,n1107);
nor (n1107,n1108,n1109);
and (n1108,n429,n579);
and (n1109,n430,n243);
nand (n1110,n1111,n1020);
nor (n1111,n1112,n1113);
and (n1112,n489,n579);
and (n1113,n490,n243);
nand (n1114,n1115,n243);
nand (n1115,n490,n575);
not (n1116,n1117);
nand (n1117,n1118,n1121);
nor (n1118,n1119,n1120);
nor (n1119,n1106,n573);
nor (n1120,n1077,n574);
nand (n1121,n490,n239);
or (n1122,n1118,n1121);
nor (n1123,n1093,n1089);
nand (n1124,n1072,n1073);
and (n1125,n1048,n1068);
and (n1126,n1027,n1044);
and (n1127,n997,n1023);
nand (n1128,n1129,n916);
or (n1129,n1130,n1132);
not (n1130,n1131);
nand (n1131,n692,n817);
not (n1132,n1133);
nand (n1133,n691,n1134);
nand (n1134,n1135,n1137);
or (n1135,n911,n1136);
nand (n1136,n857,n885);
nand (n1137,n912,n913);
nand (n1138,n918,n991);
not (n1139,n1140);
nor (n1140,n1141,n1401);
nor (n1141,n1142,n1378);
xor (n1142,n1143,n1298);
xor (n1143,n1144,n1215);
xor (n1144,n1145,n1195);
xor (n1145,n1146,n1180);
or (n1146,n1147,n1179);
and (n1147,n1148,n1168);
xor (n1148,n1149,n1159);
nand (n1149,n1150,n1155);
or (n1150,n1151,n151);
not (n1151,n1152);
nor (n1152,n1153,n1154);
and (n1153,n64,n27);
and (n1154,n63,n26);
nand (n1155,n157,n1156);
nor (n1156,n1157,n1158);
and (n1157,n123,n26);
and (n1158,n124,n27);
nand (n1159,n1160,n1164);
or (n1160,n22,n1161);
nor (n1161,n1162,n1163);
and (n1162,n196,n20);
and (n1163,n78,n19);
nand (n1164,n24,n1165);
nor (n1165,n1166,n1167);
and (n1166,n44,n19);
and (n1167,n45,n20);
nand (n1168,n1169,n1174);
or (n1169,n543,n1170);
not (n1170,n1171);
nand (n1171,n1172,n1173);
or (n1172,n140,n105);
or (n1173,n142,n106);
nand (n1174,n1175,n136);
not (n1175,n1176);
nor (n1176,n1177,n1178);
and (n1177,n142,n88);
and (n1178,n140,n87);
and (n1179,n1149,n1159);
xor (n1180,n1181,n1189);
xor (n1181,n1182,n1186);
nand (n1182,n1183,n1185);
or (n1183,n1184,n22);
not (n1184,n1165);
nand (n1185,n24,n662);
nand (n1186,n1187,n1188);
or (n1187,n1170,n257);
nand (n1188,n130,n623);
nand (n1189,n1190,n1194);
or (n1190,n169,n1191);
nor (n1191,n1192,n1193);
and (n1192,n97,n69);
and (n1193,n95,n68);
or (n1194,n171,n631);
xor (n1195,n1196,n1211);
xor (n1196,n1197,n1204);
nand (n1197,n1198,n1203);
or (n1198,n1199,n246);
not (n1199,n1200);
nor (n1200,n1201,n1202);
and (n1201,n17,n133);
and (n1202,n18,n134);
nand (n1203,n612,n239);
nand (n1204,n1205,n1210);
or (n1205,n1206,n49);
not (n1206,n1207);
nand (n1207,n1208,n1209);
or (n1208,n46,n490);
or (n1209,n47,n489);
nand (n1210,n648,n51);
nand (n1211,n1212,n1213);
or (n1212,n654,n156);
or (n1213,n151,n1214);
not (n1214,n1156);
or (n1215,n1216,n1297);
and (n1216,n1217,n1254);
xor (n1217,n1218,n1219);
xor (n1218,n1148,n1168);
xor (n1219,n1220,n1238);
xor (n1220,n1221,n1228);
nand (n1221,n1222,n1226);
or (n1222,n1223,n169);
nor (n1223,n1224,n1225);
and (n1224,n272,n95);
and (n1225,n273,n97);
nand (n1226,n1227,n172);
not (n1227,n1191);
nand (n1228,n1229,n1233);
or (n1229,n90,n1230);
nor (n1230,n1231,n1232);
and (n1231,n53,n430);
and (n1232,n54,n429);
nand (n1233,n1234,n102);
not (n1234,n1235);
nor (n1235,n1236,n1237);
and (n1236,n53,n367);
and (n1237,n54,n366);
and (n1238,n1239,n1244);
nor (n1239,n1240,n53);
nor (n1240,n1241,n1243);
and (n1241,n1242,n97);
nand (n1242,n490,n94);
and (n1243,n489,n93);
nand (n1244,n1245,n1250);
or (n1245,n573,n1246);
not (n1246,n1247);
nor (n1247,n1248,n1249);
and (n1248,n17,n579);
and (n1249,n18,n243);
nand (n1250,n1251,n575);
nor (n1251,n1252,n1253);
and (n1252,n288,n579);
and (n1253,n37,n243);
or (n1254,n1255,n1296);
and (n1255,n1256,n1277);
xor (n1256,n1257,n1258);
xor (n1257,n1239,n1244);
or (n1258,n1259,n1276);
and (n1259,n1260,n1269);
xor (n1260,n1261,n1262);
and (n1261,n102,n490);
nand (n1262,n1263,n1265);
or (n1263,n1264,n246);
not (n1264,n953);
nand (n1265,n239,n1266);
nor (n1266,n1267,n1268);
and (n1267,n105,n133);
and (n1268,n106,n134);
nand (n1269,n1270,n1275);
or (n1270,n1271,n156);
not (n1271,n1272);
nand (n1272,n1273,n1274);
or (n1273,n27,n44);
or (n1274,n26,n45);
or (n1275,n151,n970);
and (n1276,n1261,n1262);
or (n1277,n1278,n1295);
and (n1278,n1279,n1289);
xor (n1279,n1280,n1286);
nand (n1280,n1281,n1282);
or (n1281,n975,n22);
nand (n1282,n1283,n24);
nor (n1283,n1284,n1285);
and (n1284,n68,n19);
and (n1285,n69,n20);
nand (n1286,n1287,n1288);
or (n1287,n574,n1246);
nand (n1288,n984,n1020);
nand (n1289,n1290,n1291);
or (n1290,n924,n169);
nand (n1291,n1292,n172);
nor (n1292,n1293,n1294);
and (n1293,n366,n97);
and (n1294,n367,n95);
and (n1295,n1280,n1286);
and (n1296,n1257,n1258);
and (n1297,n1218,n1219);
xor (n1298,n1299,n1338);
xor (n1299,n1300,n1303);
or (n1300,n1301,n1302);
and (n1301,n1220,n1238);
and (n1302,n1221,n1228);
xor (n1303,n1304,n1322);
xor (n1304,n1305,n1308);
nand (n1305,n1306,n1307);
or (n1306,n90,n1235);
or (n1307,n91,n638);
xor (n1308,n1309,n1315);
nor (n1309,n1310,n46);
nor (n1310,n1311,n1313);
and (n1311,n1312,n53);
nand (n1312,n490,n55);
and (n1313,n489,n1314);
not (n1314,n55);
nand (n1315,n1316,n1321);
or (n1316,n1317,n573);
not (n1317,n1318);
nor (n1318,n1319,n1320);
and (n1319,n114,n579);
and (n1320,n115,n243);
or (n1321,n605,n574);
or (n1322,n1323,n1337);
and (n1323,n1324,n1330);
xor (n1324,n1325,n1326);
and (n1325,n51,n490);
nand (n1326,n1327,n1329);
or (n1327,n573,n1328);
not (n1328,n1251);
nand (n1329,n1318,n575);
nand (n1330,n1331,n1336);
or (n1331,n246,n1332);
not (n1332,n1333);
nor (n1333,n1334,n1335);
and (n1334,n133,n183);
and (n1335,n184,n134);
or (n1336,n247,n1199);
and (n1337,n1325,n1326);
or (n1338,n1339,n1377);
and (n1339,n1340,n1376);
xor (n1340,n1341,n1356);
or (n1341,n1342,n1355);
and (n1342,n1343,n1351);
xor (n1343,n1344,n1348);
nand (n1344,n1345,n1347);
or (n1345,n1346,n246);
not (n1346,n1266);
nand (n1347,n1333,n239);
nand (n1348,n1349,n1350);
or (n1349,n1271,n151);
nand (n1350,n157,n1152);
nand (n1351,n1352,n1354);
or (n1352,n22,n1353);
not (n1353,n1283);
or (n1354,n666,n1161);
and (n1355,n1344,n1348);
or (n1356,n1357,n1375);
and (n1357,n1358,n1369);
xor (n1358,n1359,n1365);
nand (n1359,n1360,n1364);
or (n1360,n257,n1361);
nor (n1361,n1362,n1363);
and (n1362,n124,n142);
and (n1363,n123,n140);
or (n1364,n1176,n543);
nand (n1365,n1366,n1368);
or (n1366,n169,n1367);
not (n1367,n1292);
or (n1368,n1223,n171);
nand (n1369,n1370,n1374);
or (n1370,n90,n1371);
nor (n1371,n1372,n1373);
and (n1372,n489,n54);
and (n1373,n490,n53);
or (n1374,n1230,n91);
and (n1375,n1359,n1365);
xor (n1376,n1324,n1330);
and (n1377,n1341,n1356);
or (n1378,n1379,n1400);
and (n1379,n1380,n1383);
xor (n1380,n1381,n1382);
xor (n1381,n1340,n1376);
xor (n1382,n1217,n1254);
or (n1383,n1384,n1399);
and (n1384,n1385,n1388);
xor (n1385,n1386,n1387);
xor (n1386,n1358,n1369);
xor (n1387,n1343,n1351);
or (n1388,n1389,n1398);
and (n1389,n1390,n1395);
xor (n1390,n1391,n1394);
nand (n1391,n1392,n1393);
or (n1392,n257,n936);
or (n1393,n1361,n543);
nor (n1394,n948,n942);
or (n1395,n1396,n1397);
and (n1396,n966,n980);
and (n1397,n967,n973);
and (n1398,n1391,n1394);
and (n1399,n1386,n1387);
and (n1400,n1381,n1382);
nand (n1401,n1402,n1431);
nor (n1402,n1403,n1426);
nor (n1403,n1404,n1417);
xor (n1404,n1405,n1416);
xor (n1405,n1406,n1407);
xor (n1406,n1256,n1277);
or (n1407,n1408,n1415);
and (n1408,n1409,n1412);
xor (n1409,n1410,n1411);
xor (n1410,n1279,n1289);
xor (n1411,n1260,n1269);
or (n1412,n1413,n1414);
and (n1413,n921,n939);
and (n1414,n922,n933);
and (n1415,n1410,n1411);
xor (n1416,n1385,n1388);
or (n1417,n1418,n1425);
and (n1418,n1419,n1424);
xor (n1419,n1420,n1421);
xor (n1420,n1390,n1395);
or (n1421,n1422,n1423);
and (n1422,n958,n965);
and (n1423,n959,n962);
xor (n1424,n1409,n1412);
and (n1425,n1420,n1421);
nor (n1426,n1427,n1430);
or (n1427,n1428,n1429);
and (n1428,n919,n987);
and (n1429,n920,n957);
xor (n1430,n1419,n1424);
nand (n1431,n1432,n1434);
not (n1432,n1433);
xor (n1433,n1380,n1383);
not (n1434,n1435);
or (n1435,n1436,n1437);
and (n1436,n1405,n1416);
and (n1437,n1406,n1407);
nor (n1438,n1439,n1450);
and (n1439,n1440,n1449);
nand (n1440,n1441,n1448);
or (n1441,n1442,n1443);
not (n1442,n1431);
not (n1443,n1444);
nand (n1444,n1445,n1447);
or (n1445,n1403,n1446);
nand (n1446,n1427,n1430);
nand (n1447,n1404,n1417);
nand (n1448,n1433,n1435);
not (n1449,n1141);
and (n1450,n1142,n1378);
not (n1451,n1452);
and (n1452,n1453,n1504);
nor (n1453,n1454,n1485);
nor (n1454,n1455,n1456);
xor (n1455,n591,n678);
or (n1456,n1457,n1484);
and (n1457,n1458,n1483);
xor (n1458,n1459,n1460);
xor (n1459,n551,n583);
or (n1460,n1461,n1482);
and (n1461,n1462,n1475);
xor (n1462,n1463,n1474);
or (n1463,n1464,n1473);
and (n1464,n1465,n1470);
xor (n1465,n1466,n1467);
and (n1466,n1309,n1315);
or (n1467,n1468,n1469);
and (n1468,n1196,n1211);
and (n1469,n1197,n1204);
or (n1470,n1471,n1472);
and (n1471,n1181,n1189);
and (n1472,n1182,n1186);
and (n1473,n1466,n1467);
xor (n1474,n598,n642);
or (n1475,n1476,n1481);
and (n1476,n1477,n1480);
xor (n1477,n1478,n1479);
xor (n1478,n619,n634);
xor (n1479,n601,n609);
xor (n1480,n644,n659);
and (n1481,n1478,n1479);
and (n1482,n1463,n1474);
xor (n1483,n595,n676);
and (n1484,n1459,n1460);
nor (n1485,n1486,n1487);
xor (n1486,n1458,n1483);
or (n1487,n1488,n1503);
and (n1488,n1489,n1502);
xor (n1489,n1490,n1491);
xor (n1490,n671,n674);
or (n1491,n1492,n1501);
and (n1492,n1493,n1498);
xor (n1493,n1494,n1497);
or (n1494,n1495,n1496);
and (n1495,n1304,n1322);
and (n1496,n1305,n1308);
xor (n1497,n1465,n1470);
or (n1498,n1499,n1500);
and (n1499,n1145,n1195);
and (n1500,n1146,n1180);
and (n1501,n1494,n1497);
xor (n1502,n1462,n1475);
and (n1503,n1490,n1491);
nor (n1504,n1505,n1516);
nor (n1505,n1506,n1507);
xor (n1506,n1489,n1502);
or (n1507,n1508,n1515);
and (n1508,n1509,n1514);
xor (n1509,n1510,n1511);
xor (n1510,n1477,n1480);
or (n1511,n1512,n1513);
and (n1512,n1299,n1338);
and (n1513,n1300,n1303);
xor (n1514,n1493,n1498);
and (n1515,n1510,n1511);
nor (n1516,n1517,n1518);
xor (n1517,n1509,n1514);
or (n1518,n1519,n1520);
and (n1519,n1143,n1298);
and (n1520,n1144,n1215);
not (n1521,n1522);
nand (n1522,n1523,n1530);
or (n1523,n1524,n1529);
not (n1524,n1525);
nor (n1525,n1526,n1505);
and (n1526,n1527,n1528);
nand (n1527,n1506,n1507);
nand (n1528,n1517,n1518);
not (n1529,n1453);
nor (n1530,n1531,n1535);
and (n1531,n1532,n1533);
not (n1532,n1454);
not (n1533,n1534);
nand (n1534,n1486,n1487);
and (n1535,n1455,n1456);
not (n1536,n1537);
nor (n1537,n1538,n507);
and (n1538,n1539,n1540);
nand (n1539,n509,n508);
nand (n1540,n588,n589);
nand (n1541,n503,n2);
xor (n1542,n1543,n2665);
xor (n1543,n1544,n2664);
xor (n1544,n1545,n2629);
xor (n1545,n1546,n65);
xor (n1546,n1547,n2584);
xor (n1547,n1548,n2583);
xor (n1548,n1549,n2534);
xor (n1549,n1550,n2533);
xor (n1550,n1551,n2476);
xor (n1551,n1552,n2475);
xor (n1552,n1553,n2415);
xor (n1553,n1554,n185);
xor (n1554,n1555,n2347);
xor (n1555,n1556,n2346);
xor (n1556,n1557,n2280);
xor (n1557,n1558,n2279);
xor (n1558,n1559,n2199);
xor (n1559,n1560,n2198);
xor (n1560,n1561,n2119);
xor (n1561,n1562,n150);
xor (n1562,n1563,n2027);
xor (n1563,n1564,n2026);
or (n1564,n1565,n1934);
and (n1565,n1566,n204);
or (n1566,n1567,n1840);
and (n1567,n1568,n1839);
or (n1568,n1569,n1752);
and (n1569,n1570,n319);
or (n1570,n1571,n1658);
and (n1571,n1572,n1657);
and (n1572,n580,n1573);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
and (n1575,n164,n575);
and (n1576,n149,n243);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1582);
and (n1580,n1581,n1320);
and (n1581,n149,n575);
and (n1582,n1583,n1584);
xor (n1583,n1581,n1320);
or (n1584,n1585,n1587);
and (n1585,n1586,n1253);
and (n1586,n115,n575);
and (n1587,n1588,n1589);
xor (n1588,n1586,n1253);
or (n1589,n1590,n1592);
and (n1590,n1591,n1249);
and (n1591,n37,n575);
and (n1592,n1593,n1594);
xor (n1593,n1591,n1249);
or (n1594,n1595,n1597);
and (n1595,n1596,n986);
and (n1596,n18,n575);
and (n1597,n1598,n1599);
xor (n1598,n1596,n986);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
and (n1601,n184,n575);
and (n1602,n106,n243);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
and (n1607,n106,n575);
and (n1608,n88,n243);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1614);
and (n1612,n1613,n760);
and (n1613,n88,n575);
and (n1614,n1615,n1616);
xor (n1615,n1613,n760);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
and (n1618,n124,n575);
and (n1619,n64,n243);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1625);
and (n1623,n1624,n849);
and (n1624,n64,n575);
and (n1625,n1626,n1627);
xor (n1626,n1624,n849);
or (n1627,n1628,n1630);
and (n1628,n1629,n897);
and (n1629,n45,n575);
and (n1630,n1631,n1632);
xor (n1631,n1629,n897);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
and (n1634,n78,n575);
and (n1635,n69,n243);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
and (n1640,n69,n575);
and (n1641,n273,n243);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
and (n1646,n273,n575);
and (n1647,n367,n243);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
or (n1650,n1651,n1653);
and (n1651,n1652,n1109);
and (n1652,n367,n575);
and (n1653,n1654,n1655);
xor (n1654,n1652,n1109);
and (n1655,n1656,n1113);
and (n1656,n430,n575);
and (n1657,n164,n242);
and (n1658,n1659,n1660);
xor (n1659,n1572,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n580,n1573);
and (n1663,n149,n242);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1578,n1579);
and (n1669,n115,n242);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1583,n1584);
and (n1675,n37,n242);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1588,n1589);
and (n1681,n18,n242);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1593,n1594);
and (n1687,n184,n242);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
or (n1690,n1691,n1694);
and (n1691,n1692,n1693);
xor (n1692,n1598,n1599);
and (n1693,n106,n242);
and (n1694,n1695,n1696);
xor (n1695,n1692,n1693);
or (n1696,n1697,n1700);
and (n1697,n1698,n1699);
xor (n1698,n1604,n1605);
and (n1699,n88,n242);
and (n1700,n1701,n1702);
xor (n1701,n1698,n1699);
or (n1702,n1703,n1706);
and (n1703,n1704,n1705);
xor (n1704,n1610,n1611);
and (n1705,n124,n242);
and (n1706,n1707,n1708);
xor (n1707,n1704,n1705);
or (n1708,n1709,n1712);
and (n1709,n1710,n1711);
xor (n1710,n1615,n1616);
and (n1711,n64,n242);
and (n1712,n1713,n1714);
xor (n1713,n1710,n1711);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
xor (n1716,n1621,n1622);
and (n1717,n45,n242);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
xor (n1722,n1626,n1627);
and (n1723,n78,n242);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
xor (n1728,n1631,n1632);
and (n1729,n69,n242);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1736);
and (n1733,n1734,n1735);
xor (n1734,n1637,n1638);
and (n1735,n273,n242);
and (n1736,n1737,n1738);
xor (n1737,n1734,n1735);
or (n1738,n1739,n1742);
and (n1739,n1740,n1741);
xor (n1740,n1643,n1644);
and (n1741,n367,n242);
and (n1742,n1743,n1744);
xor (n1743,n1740,n1741);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1649,n1650);
and (n1747,n430,n242);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
and (n1750,n1751,n1084);
xor (n1751,n1654,n1655);
and (n1752,n1753,n1754);
xor (n1753,n1570,n319);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1659,n1660);
and (n1757,n149,n134);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1763);
and (n1761,n1762,n529);
xor (n1762,n1665,n1666);
and (n1763,n1764,n1765);
xor (n1764,n1762,n529);
or (n1765,n1766,n1768);
and (n1766,n1767,n614);
xor (n1767,n1671,n1672);
and (n1768,n1769,n1770);
xor (n1769,n1767,n614);
or (n1770,n1771,n1773);
and (n1771,n1772,n1202);
xor (n1772,n1677,n1678);
and (n1773,n1774,n1775);
xor (n1774,n1772,n1202);
or (n1775,n1776,n1778);
and (n1776,n1777,n1335);
xor (n1777,n1683,n1684);
and (n1778,n1779,n1780);
xor (n1779,n1777,n1335);
or (n1780,n1781,n1783);
and (n1781,n1782,n1268);
xor (n1782,n1689,n1690);
and (n1783,n1784,n1785);
xor (n1784,n1782,n1268);
or (n1785,n1786,n1788);
and (n1786,n1787,n955);
xor (n1787,n1695,n1696);
and (n1788,n1789,n1790);
xor (n1789,n1787,n955);
or (n1790,n1791,n1794);
and (n1791,n1792,n1793);
xor (n1792,n1701,n1702);
and (n1793,n124,n134);
and (n1794,n1795,n1796);
xor (n1795,n1792,n1793);
or (n1796,n1797,n1800);
and (n1797,n1798,n1799);
xor (n1798,n1707,n1708);
and (n1799,n64,n134);
and (n1800,n1801,n1802);
xor (n1801,n1798,n1799);
or (n1802,n1803,n1806);
and (n1803,n1804,n1805);
xor (n1804,n1713,n1714);
and (n1805,n45,n134);
and (n1806,n1807,n1808);
xor (n1807,n1804,n1805);
or (n1808,n1809,n1812);
and (n1809,n1810,n1811);
xor (n1810,n1719,n1720);
and (n1811,n78,n134);
and (n1812,n1813,n1814);
xor (n1813,n1810,n1811);
or (n1814,n1815,n1818);
and (n1815,n1816,n1817);
xor (n1816,n1725,n1726);
and (n1817,n69,n134);
and (n1818,n1819,n1820);
xor (n1819,n1816,n1817);
or (n1820,n1821,n1823);
and (n1821,n1822,n905);
xor (n1822,n1731,n1732);
and (n1823,n1824,n1825);
xor (n1824,n1822,n905);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
xor (n1827,n1737,n1738);
and (n1828,n367,n134);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
or (n1831,n1832,n1834);
and (n1832,n1833,n1057);
xor (n1833,n1743,n1744);
and (n1834,n1835,n1836);
xor (n1835,n1833,n1057);
and (n1836,n1837,n1838);
xor (n1837,n1749,n1750);
and (n1838,n490,n134);
and (n1839,n164,n132);
and (n1840,n1841,n1842);
xor (n1841,n1568,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1753,n1754);
and (n1845,n149,n132);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1759,n1760);
and (n1851,n115,n132);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1764,n1765);
and (n1857,n37,n132);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1769,n1770);
and (n1863,n18,n132);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1774,n1775);
and (n1869,n184,n132);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1779,n1780);
and (n1875,n106,n132);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1784,n1785);
and (n1881,n88,n132);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1789,n1790);
and (n1887,n124,n132);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1795,n1796);
and (n1893,n64,n132);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1801,n1802);
and (n1899,n45,n132);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1807,n1808);
and (n1905,n78,n132);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
or (n1908,n1909,n1912);
and (n1909,n1910,n1911);
xor (n1910,n1813,n1814);
and (n1911,n69,n132);
and (n1912,n1913,n1914);
xor (n1913,n1910,n1911);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1819,n1820);
and (n1917,n273,n132);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
or (n1920,n1921,n1924);
and (n1921,n1922,n1923);
xor (n1922,n1824,n1825);
and (n1923,n367,n132);
and (n1924,n1925,n1926);
xor (n1925,n1922,n1923);
or (n1926,n1927,n1930);
and (n1927,n1928,n1929);
xor (n1928,n1830,n1831);
and (n1929,n430,n132);
and (n1930,n1931,n1932);
xor (n1931,n1928,n1929);
and (n1932,n1933,n1012);
xor (n1933,n1835,n1836);
and (n1934,n1935,n1936);
xor (n1935,n1566,n204);
or (n1936,n1937,n1940);
and (n1937,n1938,n1939);
xor (n1938,n1841,n1842);
and (n1939,n149,n140);
and (n1940,n1941,n1942);
xor (n1941,n1938,n1939);
or (n1942,n1943,n1945);
and (n1943,n1944,n362);
xor (n1944,n1847,n1848);
and (n1945,n1946,n1947);
xor (n1946,n1944,n362);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1853,n1854);
and (n1950,n37,n140);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1859,n1860);
and (n1956,n18,n140);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1962);
and (n1960,n1961,n625);
xor (n1961,n1865,n1866);
and (n1962,n1963,n1964);
xor (n1963,n1961,n625);
or (n1964,n1965,n1968);
and (n1965,n1966,n1967);
xor (n1966,n1871,n1872);
and (n1967,n106,n140);
and (n1968,n1969,n1970);
xor (n1969,n1966,n1967);
or (n1970,n1971,n1974);
and (n1971,n1972,n1973);
xor (n1972,n1877,n1878);
and (n1973,n88,n140);
and (n1974,n1975,n1976);
xor (n1975,n1972,n1973);
or (n1976,n1977,n1980);
and (n1977,n1978,n1979);
xor (n1978,n1883,n1884);
and (n1979,n124,n140);
and (n1980,n1981,n1982);
xor (n1981,n1978,n1979);
or (n1982,n1983,n1986);
and (n1983,n1984,n1985);
xor (n1984,n1889,n1890);
and (n1985,n64,n140);
and (n1986,n1987,n1988);
xor (n1987,n1984,n1985);
or (n1988,n1989,n1992);
and (n1989,n1990,n1991);
xor (n1990,n1895,n1896);
and (n1991,n45,n140);
and (n1992,n1993,n1994);
xor (n1993,n1990,n1991);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1901,n1902);
and (n1997,n78,n140);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
or (n2000,n2001,n2004);
and (n2001,n2002,n2003);
xor (n2002,n1907,n1908);
and (n2003,n69,n140);
and (n2004,n2005,n2006);
xor (n2005,n2002,n2003);
or (n2006,n2007,n2010);
and (n2007,n2008,n2009);
xor (n2008,n1913,n1914);
and (n2009,n273,n140);
and (n2010,n2011,n2012);
xor (n2011,n2008,n2009);
or (n2012,n2013,n2016);
and (n2013,n2014,n2015);
xor (n2014,n1919,n1920);
and (n2015,n367,n140);
and (n2016,n2017,n2018);
xor (n2017,n2014,n2015);
or (n2018,n2019,n2021);
and (n2019,n2020,n1004);
xor (n2020,n1925,n1926);
and (n2021,n2022,n2023);
xor (n2022,n2020,n1004);
and (n2023,n2024,n2025);
xor (n2024,n1931,n1932);
and (n2025,n490,n140);
and (n2026,n164,n154);
or (n2027,n2028,n2031);
and (n2028,n2029,n2030);
xor (n2029,n1935,n1936);
and (n2030,n149,n154);
and (n2031,n2032,n2033);
xor (n2032,n2029,n2030);
or (n2033,n2034,n2037);
and (n2034,n2035,n2036);
xor (n2035,n1941,n1942);
and (n2036,n115,n154);
and (n2037,n2038,n2039);
xor (n2038,n2035,n2036);
or (n2039,n2040,n2043);
and (n2040,n2041,n2042);
xor (n2041,n1946,n1947);
and (n2042,n37,n154);
and (n2043,n2044,n2045);
xor (n2044,n2041,n2042);
or (n2045,n2046,n2049);
and (n2046,n2047,n2048);
xor (n2047,n1952,n1953);
and (n2048,n18,n154);
and (n2049,n2050,n2051);
xor (n2050,n2047,n2048);
or (n2051,n2052,n2055);
and (n2052,n2053,n2054);
xor (n2053,n1958,n1959);
and (n2054,n184,n154);
and (n2055,n2056,n2057);
xor (n2056,n2053,n2054);
or (n2057,n2058,n2061);
and (n2058,n2059,n2060);
xor (n2059,n1963,n1964);
and (n2060,n106,n154);
and (n2061,n2062,n2063);
xor (n2062,n2059,n2060);
or (n2063,n2064,n2067);
and (n2064,n2065,n2066);
xor (n2065,n1969,n1970);
and (n2066,n88,n154);
and (n2067,n2068,n2069);
xor (n2068,n2065,n2066);
or (n2069,n2070,n2073);
and (n2070,n2071,n2072);
xor (n2071,n1975,n1976);
and (n2072,n124,n154);
and (n2073,n2074,n2075);
xor (n2074,n2071,n2072);
or (n2075,n2076,n2079);
and (n2076,n2077,n2078);
xor (n2077,n1981,n1982);
and (n2078,n64,n154);
and (n2079,n2080,n2081);
xor (n2080,n2077,n2078);
or (n2081,n2082,n2085);
and (n2082,n2083,n2084);
xor (n2083,n1987,n1988);
and (n2084,n45,n154);
and (n2085,n2086,n2087);
xor (n2086,n2083,n2084);
or (n2087,n2088,n2091);
and (n2088,n2089,n2090);
xor (n2089,n1993,n1994);
and (n2090,n78,n154);
and (n2091,n2092,n2093);
xor (n2092,n2089,n2090);
or (n2093,n2094,n2097);
and (n2094,n2095,n2096);
xor (n2095,n1999,n2000);
and (n2096,n69,n154);
and (n2097,n2098,n2099);
xor (n2098,n2095,n2096);
or (n2099,n2100,n2103);
and (n2100,n2101,n2102);
xor (n2101,n2005,n2006);
and (n2102,n273,n154);
and (n2103,n2104,n2105);
xor (n2104,n2101,n2102);
or (n2105,n2106,n2109);
and (n2106,n2107,n2108);
xor (n2107,n2011,n2012);
and (n2108,n367,n154);
and (n2109,n2110,n2111);
xor (n2110,n2107,n2108);
or (n2111,n2112,n2115);
and (n2112,n2113,n2114);
xor (n2113,n2017,n2018);
and (n2114,n430,n154);
and (n2115,n2116,n2117);
xor (n2116,n2113,n2114);
and (n2117,n2118,n841);
xor (n2118,n2022,n2023);
or (n2119,n2120,n2122);
and (n2120,n2121,n214);
xor (n2121,n2032,n2033);
and (n2122,n2123,n2124);
xor (n2123,n2121,n214);
or (n2124,n2125,n2127);
and (n2125,n2126,n289);
xor (n2126,n2038,n2039);
and (n2127,n2128,n2129);
xor (n2128,n2126,n289);
or (n2129,n2130,n2132);
and (n2130,n2131,n345);
xor (n2131,n2044,n2045);
and (n2132,n2133,n2134);
xor (n2133,n2131,n345);
or (n2134,n2135,n2138);
and (n2135,n2136,n2137);
xor (n2136,n2050,n2051);
and (n2137,n184,n27);
and (n2138,n2139,n2140);
xor (n2139,n2136,n2137);
or (n2140,n2141,n2143);
and (n2141,n2142,n478);
xor (n2142,n2056,n2057);
and (n2143,n2144,n2145);
xor (n2144,n2142,n478);
or (n2145,n2146,n2149);
and (n2146,n2147,n2148);
xor (n2147,n2062,n2063);
and (n2148,n88,n27);
and (n2149,n2150,n2151);
xor (n2150,n2147,n2148);
or (n2151,n2152,n2154);
and (n2152,n2153,n1158);
xor (n2153,n2068,n2069);
and (n2154,n2155,n2156);
xor (n2155,n2153,n1158);
or (n2156,n2157,n2159);
and (n2157,n2158,n1153);
xor (n2158,n2074,n2075);
and (n2159,n2160,n2161);
xor (n2160,n2158,n1153);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2080,n2081);
and (n2164,n45,n27);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
or (n2167,n2168,n2171);
and (n2168,n2169,n2170);
xor (n2169,n2086,n2087);
and (n2170,n78,n27);
and (n2171,n2172,n2173);
xor (n2172,n2169,n2170);
or (n2173,n2174,n2177);
and (n2174,n2175,n2176);
xor (n2175,n2092,n2093);
and (n2176,n69,n27);
and (n2177,n2178,n2179);
xor (n2178,n2175,n2176);
or (n2179,n2180,n2182);
and (n2180,n2181,n788);
xor (n2181,n2098,n2099);
and (n2182,n2183,n2184);
xor (n2183,n2181,n788);
or (n2184,n2185,n2187);
and (n2185,n2186,n773);
xor (n2186,n2104,n2105);
and (n2187,n2188,n2189);
xor (n2188,n2186,n773);
or (n2189,n2190,n2193);
and (n2190,n2191,n2192);
xor (n2191,n2110,n2111);
and (n2192,n430,n27);
and (n2193,n2194,n2195);
xor (n2194,n2191,n2192);
and (n2195,n2196,n2197);
xor (n2196,n2116,n2117);
and (n2197,n490,n27);
and (n2198,n115,n28);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2123,n2124);
and (n2202,n37,n28);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
xor (n2207,n2128,n2129);
and (n2208,n18,n28);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2215);
and (n2212,n2213,n2214);
xor (n2213,n2133,n2134);
and (n2214,n184,n28);
and (n2215,n2216,n2217);
xor (n2216,n2213,n2214);
or (n2217,n2218,n2221);
and (n2218,n2219,n2220);
xor (n2219,n2139,n2140);
and (n2220,n106,n28);
and (n2221,n2222,n2223);
xor (n2222,n2219,n2220);
or (n2223,n2224,n2227);
and (n2224,n2225,n2226);
xor (n2225,n2144,n2145);
and (n2226,n88,n28);
and (n2227,n2228,n2229);
xor (n2228,n2225,n2226);
or (n2229,n2230,n2233);
and (n2230,n2231,n2232);
xor (n2231,n2150,n2151);
and (n2232,n124,n28);
and (n2233,n2234,n2235);
xor (n2234,n2231,n2232);
or (n2235,n2236,n2239);
and (n2236,n2237,n2238);
xor (n2237,n2155,n2156);
and (n2238,n64,n28);
and (n2239,n2240,n2241);
xor (n2240,n2237,n2238);
or (n2241,n2242,n2245);
and (n2242,n2243,n2244);
xor (n2243,n2160,n2161);
and (n2244,n45,n28);
and (n2245,n2246,n2247);
xor (n2246,n2243,n2244);
or (n2247,n2248,n2251);
and (n2248,n2249,n2250);
xor (n2249,n2166,n2167);
and (n2250,n78,n28);
and (n2251,n2252,n2253);
xor (n2252,n2249,n2250);
or (n2253,n2254,n2257);
and (n2254,n2255,n2256);
xor (n2255,n2172,n2173);
and (n2256,n69,n28);
and (n2257,n2258,n2259);
xor (n2258,n2255,n2256);
or (n2259,n2260,n2263);
and (n2260,n2261,n2262);
xor (n2261,n2178,n2179);
and (n2262,n273,n28);
and (n2263,n2264,n2265);
xor (n2264,n2261,n2262);
or (n2265,n2266,n2269);
and (n2266,n2267,n2268);
xor (n2267,n2183,n2184);
and (n2268,n367,n28);
and (n2269,n2270,n2271);
xor (n2270,n2267,n2268);
or (n2271,n2272,n2275);
and (n2272,n2273,n2274);
xor (n2273,n2188,n2189);
and (n2274,n430,n28);
and (n2275,n2276,n2277);
xor (n2276,n2273,n2274);
and (n2277,n2278,n739);
xor (n2278,n2194,n2195);
and (n2279,n37,n20);
or (n2280,n2281,n2283);
and (n2281,n2282,n21);
xor (n2282,n2204,n2205);
and (n2283,n2284,n2285);
xor (n2284,n2282,n21);
or (n2285,n2286,n2288);
and (n2286,n2287,n264);
xor (n2287,n2210,n2211);
and (n2288,n2289,n2290);
xor (n2289,n2287,n264);
or (n2290,n2291,n2293);
and (n2291,n2292,n374);
xor (n2292,n2216,n2217);
and (n2293,n2294,n2295);
xor (n2294,n2292,n374);
or (n2295,n2296,n2298);
and (n2296,n2297,n447);
xor (n2297,n2222,n2223);
and (n2298,n2299,n2300);
xor (n2299,n2297,n447);
or (n2300,n2301,n2303);
and (n2301,n2302,n536);
xor (n2302,n2228,n2229);
and (n2303,n2304,n2305);
xor (n2304,n2302,n536);
or (n2305,n2306,n2308);
and (n2306,n2307,n664);
xor (n2307,n2234,n2235);
and (n2308,n2309,n2310);
xor (n2309,n2307,n664);
or (n2310,n2311,n2313);
and (n2311,n2312,n1167);
xor (n2312,n2240,n2241);
and (n2313,n2314,n2315);
xor (n2314,n2312,n1167);
or (n2315,n2316,n2319);
and (n2316,n2317,n2318);
xor (n2317,n2246,n2247);
and (n2318,n78,n20);
and (n2319,n2320,n2321);
xor (n2320,n2317,n2318);
or (n2321,n2322,n2324);
and (n2322,n2323,n1285);
xor (n2323,n2252,n2253);
and (n2324,n2325,n2326);
xor (n2325,n2323,n1285);
or (n2326,n2327,n2330);
and (n2327,n2328,n2329);
xor (n2328,n2258,n2259);
and (n2329,n273,n20);
and (n2330,n2331,n2332);
xor (n2331,n2328,n2329);
or (n2332,n2333,n2336);
and (n2333,n2334,n2335);
xor (n2334,n2264,n2265);
and (n2335,n367,n20);
and (n2336,n2337,n2338);
xor (n2337,n2334,n2335);
or (n2338,n2339,n2341);
and (n2339,n2340,n701);
xor (n2340,n2270,n2271);
and (n2341,n2342,n2343);
xor (n2342,n2340,n701);
and (n2343,n2344,n2345);
xor (n2344,n2276,n2277);
and (n2345,n490,n20);
and (n2346,n18,n175);
or (n2347,n2348,n2351);
and (n2348,n2349,n2350);
xor (n2349,n2284,n2285);
and (n2350,n184,n175);
and (n2351,n2352,n2353);
xor (n2352,n2349,n2350);
or (n2353,n2354,n2357);
and (n2354,n2355,n2356);
xor (n2355,n2289,n2290);
and (n2356,n106,n175);
and (n2357,n2358,n2359);
xor (n2358,n2355,n2356);
or (n2359,n2360,n2363);
and (n2360,n2361,n2362);
xor (n2361,n2294,n2295);
and (n2362,n88,n175);
and (n2363,n2364,n2365);
xor (n2364,n2361,n2362);
or (n2365,n2366,n2369);
and (n2366,n2367,n2368);
xor (n2367,n2299,n2300);
and (n2368,n124,n175);
and (n2369,n2370,n2371);
xor (n2370,n2367,n2368);
or (n2371,n2372,n2375);
and (n2372,n2373,n2374);
xor (n2373,n2304,n2305);
and (n2374,n64,n175);
and (n2375,n2376,n2377);
xor (n2376,n2373,n2374);
or (n2377,n2378,n2381);
and (n2378,n2379,n2380);
xor (n2379,n2309,n2310);
and (n2380,n45,n175);
and (n2381,n2382,n2383);
xor (n2382,n2379,n2380);
or (n2383,n2384,n2387);
and (n2384,n2385,n2386);
xor (n2385,n2314,n2315);
and (n2386,n78,n175);
and (n2387,n2388,n2389);
xor (n2388,n2385,n2386);
or (n2389,n2390,n2393);
and (n2390,n2391,n2392);
xor (n2391,n2320,n2321);
and (n2392,n69,n175);
and (n2393,n2394,n2395);
xor (n2394,n2391,n2392);
or (n2395,n2396,n2399);
and (n2396,n2397,n2398);
xor (n2397,n2325,n2326);
and (n2398,n273,n175);
and (n2399,n2400,n2401);
xor (n2400,n2397,n2398);
or (n2401,n2402,n2405);
and (n2402,n2403,n2404);
xor (n2403,n2331,n2332);
and (n2404,n367,n175);
and (n2405,n2406,n2407);
xor (n2406,n2403,n2404);
or (n2407,n2408,n2411);
and (n2408,n2409,n2410);
xor (n2409,n2337,n2338);
and (n2410,n430,n175);
and (n2411,n2412,n2413);
xor (n2412,n2409,n2410);
and (n2413,n2414,n947);
xor (n2414,n2342,n2343);
or (n2415,n2416,n2418);
and (n2416,n2417,n221);
xor (n2417,n2352,n2353);
and (n2418,n2419,n2420);
xor (n2419,n2417,n221);
or (n2420,n2421,n2423);
and (n2421,n2422,n280);
xor (n2422,n2358,n2359);
and (n2423,n2424,n2425);
xor (n2424,n2422,n280);
or (n2425,n2426,n2429);
and (n2426,n2427,n2428);
xor (n2427,n2364,n2365);
and (n2428,n124,n95);
and (n2429,n2430,n2431);
xor (n2430,n2427,n2428);
or (n2431,n2432,n2435);
and (n2432,n2433,n2434);
xor (n2433,n2370,n2371);
and (n2434,n64,n95);
and (n2435,n2436,n2437);
xor (n2436,n2433,n2434);
or (n2437,n2438,n2441);
and (n2438,n2439,n2440);
xor (n2439,n2376,n2377);
and (n2440,n45,n95);
and (n2441,n2442,n2443);
xor (n2442,n2439,n2440);
or (n2443,n2444,n2447);
and (n2444,n2445,n2446);
xor (n2445,n2382,n2383);
and (n2446,n78,n95);
and (n2447,n2448,n2449);
xor (n2448,n2445,n2446);
or (n2449,n2450,n2453);
and (n2450,n2451,n2452);
xor (n2451,n2388,n2389);
and (n2452,n69,n95);
and (n2453,n2454,n2455);
xor (n2454,n2451,n2452);
or (n2455,n2456,n2459);
and (n2456,n2457,n2458);
xor (n2457,n2394,n2395);
and (n2458,n273,n95);
and (n2459,n2460,n2461);
xor (n2460,n2457,n2458);
or (n2461,n2462,n2464);
and (n2462,n2463,n1294);
xor (n2463,n2400,n2401);
and (n2464,n2465,n2466);
xor (n2465,n2463,n1294);
or (n2466,n2467,n2470);
and (n2467,n2468,n2469);
xor (n2468,n2406,n2407);
and (n2469,n430,n95);
and (n2470,n2471,n2472);
xor (n2471,n2468,n2469);
and (n2472,n2473,n2474);
xor (n2473,n2412,n2413);
and (n2474,n490,n95);
and (n2475,n106,n94);
or (n2476,n2477,n2480);
and (n2477,n2478,n2479);
xor (n2478,n2419,n2420);
and (n2479,n88,n94);
and (n2480,n2481,n2482);
xor (n2481,n2478,n2479);
or (n2482,n2483,n2486);
and (n2483,n2484,n2485);
xor (n2484,n2424,n2425);
and (n2485,n124,n94);
and (n2486,n2487,n2488);
xor (n2487,n2484,n2485);
or (n2488,n2489,n2492);
and (n2489,n2490,n2491);
xor (n2490,n2430,n2431);
and (n2491,n64,n94);
and (n2492,n2493,n2494);
xor (n2493,n2490,n2491);
or (n2494,n2495,n2498);
and (n2495,n2496,n2497);
xor (n2496,n2436,n2437);
and (n2497,n45,n94);
and (n2498,n2499,n2500);
xor (n2499,n2496,n2497);
or (n2500,n2501,n2504);
and (n2501,n2502,n2503);
xor (n2502,n2442,n2443);
and (n2503,n78,n94);
and (n2504,n2505,n2506);
xor (n2505,n2502,n2503);
or (n2506,n2507,n2510);
and (n2507,n2508,n2509);
xor (n2508,n2448,n2449);
and (n2509,n69,n94);
and (n2510,n2511,n2512);
xor (n2511,n2508,n2509);
or (n2512,n2513,n2516);
and (n2513,n2514,n2515);
xor (n2514,n2454,n2455);
and (n2515,n273,n94);
and (n2516,n2517,n2518);
xor (n2517,n2514,n2515);
or (n2518,n2519,n2522);
and (n2519,n2520,n2521);
xor (n2520,n2460,n2461);
and (n2521,n367,n94);
and (n2522,n2523,n2524);
xor (n2523,n2520,n2521);
or (n2524,n2525,n2528);
and (n2525,n2526,n2527);
xor (n2526,n2465,n2466);
and (n2527,n430,n94);
and (n2528,n2529,n2530);
xor (n2529,n2526,n2527);
and (n2530,n2531,n2532);
xor (n2531,n2471,n2472);
not (n2532,n1242);
and (n2533,n88,n54);
or (n2534,n2535,n2537);
and (n2535,n2536,n229);
xor (n2536,n2481,n2482);
and (n2537,n2538,n2539);
xor (n2538,n2536,n229);
or (n2539,n2540,n2542);
and (n2540,n2541,n305);
xor (n2541,n2487,n2488);
and (n2542,n2543,n2544);
xor (n2543,n2541,n305);
or (n2544,n2545,n2548);
and (n2545,n2546,n2547);
xor (n2546,n2493,n2494);
and (n2547,n45,n54);
and (n2548,n2549,n2550);
xor (n2549,n2546,n2547);
or (n2550,n2551,n2554);
and (n2551,n2552,n2553);
xor (n2552,n2499,n2500);
and (n2553,n78,n54);
and (n2554,n2555,n2556);
xor (n2555,n2552,n2553);
or (n2556,n2557,n2560);
and (n2557,n2558,n2559);
xor (n2558,n2505,n2506);
and (n2559,n69,n54);
and (n2560,n2561,n2562);
xor (n2561,n2558,n2559);
or (n2562,n2563,n2566);
and (n2563,n2564,n2565);
xor (n2564,n2511,n2512);
and (n2565,n273,n54);
and (n2566,n2567,n2568);
xor (n2567,n2564,n2565);
or (n2568,n2569,n2572);
and (n2569,n2570,n2571);
xor (n2570,n2517,n2518);
and (n2571,n367,n54);
and (n2572,n2573,n2574);
xor (n2573,n2570,n2571);
or (n2574,n2575,n2578);
and (n2575,n2576,n2577);
xor (n2576,n2523,n2524);
and (n2577,n430,n54);
and (n2578,n2579,n2580);
xor (n2579,n2576,n2577);
and (n2580,n2581,n2582);
xor (n2581,n2529,n2530);
and (n2582,n490,n54);
and (n2583,n124,n55);
or (n2584,n2585,n2588);
and (n2585,n2586,n2587);
xor (n2586,n2538,n2539);
and (n2587,n64,n55);
and (n2588,n2589,n2590);
xor (n2589,n2586,n2587);
or (n2590,n2591,n2594);
and (n2591,n2592,n2593);
xor (n2592,n2543,n2544);
and (n2593,n45,n55);
and (n2594,n2595,n2596);
xor (n2595,n2592,n2593);
or (n2596,n2597,n2600);
and (n2597,n2598,n2599);
xor (n2598,n2549,n2550);
and (n2599,n78,n55);
and (n2600,n2601,n2602);
xor (n2601,n2598,n2599);
or (n2602,n2603,n2606);
and (n2603,n2604,n2605);
xor (n2604,n2555,n2556);
and (n2605,n69,n55);
and (n2606,n2607,n2608);
xor (n2607,n2604,n2605);
or (n2608,n2609,n2612);
and (n2609,n2610,n2611);
xor (n2610,n2561,n2562);
and (n2611,n273,n55);
and (n2612,n2613,n2614);
xor (n2613,n2610,n2611);
or (n2614,n2615,n2618);
and (n2615,n2616,n2617);
xor (n2616,n2567,n2568);
and (n2617,n367,n55);
and (n2618,n2619,n2620);
xor (n2619,n2616,n2617);
or (n2620,n2621,n2624);
and (n2621,n2622,n2623);
xor (n2622,n2573,n2574);
and (n2623,n430,n55);
and (n2624,n2625,n2626);
xor (n2625,n2622,n2623);
and (n2626,n2627,n2628);
xor (n2627,n2579,n2580);
not (n2628,n1312);
or (n2629,n2630,n2632);
and (n2630,n2631,n48);
xor (n2631,n2589,n2590);
and (n2632,n2633,n2634);
xor (n2633,n2631,n48);
or (n2634,n2635,n2637);
and (n2635,n2636,n312);
xor (n2636,n2595,n2596);
and (n2637,n2638,n2639);
xor (n2638,n2636,n312);
or (n2639,n2640,n2642);
and (n2640,n2641,n397);
xor (n2641,n2601,n2602);
and (n2642,n2643,n2644);
xor (n2643,n2641,n397);
or (n2644,n2645,n2648);
and (n2645,n2646,n2647);
xor (n2646,n2607,n2608);
and (n2647,n273,n47);
and (n2648,n2649,n2650);
xor (n2649,n2646,n2647);
or (n2650,n2651,n2654);
and (n2651,n2652,n2653);
xor (n2652,n2613,n2614);
and (n2653,n367,n47);
and (n2654,n2655,n2656);
xor (n2655,n2652,n2653);
or (n2656,n2657,n2659);
and (n2657,n2658,n650);
xor (n2658,n2619,n2620);
and (n2659,n2660,n2661);
xor (n2660,n2658,n650);
and (n2661,n2662,n2663);
xor (n2662,n2625,n2626);
and (n2663,n490,n47);
and (n2664,n45,n74);
or (n2665,n2666,n2669);
and (n2666,n2667,n2668);
xor (n2667,n2633,n2634);
and (n2668,n78,n74);
and (n2669,n2670,n2671);
xor (n2670,n2667,n2668);
or (n2671,n2672,n2675);
and (n2672,n2673,n2674);
xor (n2673,n2638,n2639);
and (n2674,n69,n74);
and (n2675,n2676,n2677);
xor (n2676,n2673,n2674);
or (n2677,n2678,n2681);
and (n2678,n2679,n2680);
xor (n2679,n2643,n2644);
and (n2680,n273,n74);
and (n2681,n2682,n2683);
xor (n2682,n2679,n2680);
or (n2683,n2684,n2687);
and (n2684,n2685,n2686);
xor (n2685,n2649,n2650);
and (n2686,n367,n74);
and (n2687,n2688,n2689);
xor (n2688,n2685,n2686);
or (n2689,n2690,n2693);
and (n2690,n2691,n2692);
xor (n2691,n2655,n2656);
and (n2692,n430,n74);
and (n2693,n2694,n2695);
xor (n2694,n2691,n2692);
and (n2695,n2696,n2697);
xor (n2696,n2660,n2661);
and (n2697,n490,n74);
endmodule
