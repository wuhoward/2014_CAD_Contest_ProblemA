module top (out,n12,n14,n15,n17,n20,n21,n27,n29,n30
        ,n32,n35,n39,n41,n42,n44,n47,n52,n54,n56
        ,n68,n77,n79,n81,n84,n96,n103,n105,n107,n110
        ,n118,n119,n131,n143,n181,n185,n187,n189,n217,n218
        ,n325,n342,n343,n495,n499,n501,n512,n524,n538);
output out;
input n12;
input n14;
input n15;
input n17;
input n20;
input n21;
input n27;
input n29;
input n30;
input n32;
input n35;
input n39;
input n41;
input n42;
input n44;
input n47;
input n52;
input n54;
input n56;
input n68;
input n77;
input n79;
input n81;
input n84;
input n96;
input n103;
input n105;
input n107;
input n110;
input n118;
input n119;
input n131;
input n143;
input n181;
input n185;
input n187;
input n189;
input n217;
input n218;
input n325;
input n342;
input n343;
input n495;
input n499;
input n501;
input n512;
input n524;
input n538;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n16;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n31;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n40;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n80;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n106;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n186;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n496;
wire n497;
wire n498;
wire n500;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
xor (out,n0,n2516);
xnor (n0,n1,n2436);
nand (n1,n2,n476);
nand (n2,n3,n396);
nand (n3,n4,n312,n395);
nand (n4,n5,n171);
xor (n5,n6,n135);
xor (n6,n7,n60);
xor (n7,n8,n22);
xor (n8,n9,n21);
xor (n9,n10,n20);
or (n10,n11,n16);
and (n11,n12,n13);
xor (n13,n14,n15);
and (n16,n17,n18);
nor (n18,n13,n19);
xnor (n19,n20,n14);
nand (n22,n23,n48,n59);
nand (n23,n24,n36);
xor (n24,n25,n35);
or (n25,n26,n31);
and (n26,n27,n28);
xor (n28,n29,n30);
and (n31,n32,n33);
nor (n33,n28,n34);
xnor (n34,n35,n29);
xor (n36,n37,n47);
or (n37,n38,n43);
and (n38,n39,n40);
xor (n40,n41,n42);
and (n43,n44,n45);
nor (n45,n40,n46);
xnor (n46,n47,n41);
nand (n48,n49,n36);
xor (n49,n50,n30);
or (n50,n51,n55);
and (n51,n52,n53);
xor (n53,n54,n47);
and (n55,n56,n57);
nor (n57,n53,n58);
xnor (n58,n30,n54);
nand (n59,n24,n49);
nand (n60,n61,n111,n134);
nand (n61,n62,n86);
nand (n62,n63,n73,n85);
nand (n63,n64,n69);
xor (n64,n65,n35);
or (n65,n66,n67);
and (n66,n32,n28);
and (n67,n68,n33);
xor (n69,n70,n47);
or (n70,n71,n72);
and (n71,n44,n40);
and (n72,n52,n45);
nand (n73,n74,n69);
xor (n74,n75,n84);
or (n75,n76,n80);
and (n76,n77,n78);
xor (n78,n79,n35);
and (n80,n81,n82);
nor (n82,n78,n83);
xnor (n83,n84,n79);
nand (n85,n64,n74);
xor (n86,n87,n100);
xor (n87,n88,n92);
xor (n88,n89,n84);
or (n89,n90,n91);
and (n90,n68,n78);
and (n91,n77,n82);
xor (n92,n93,n15);
or (n93,n94,n97);
and (n94,n81,n95);
xor (n95,n96,n84);
and (n97,n12,n98);
nor (n98,n95,n99);
xnor (n99,n15,n96);
xor (n100,n101,n110);
or (n101,n102,n106);
and (n102,n103,n104);
xor (n104,n105,n20);
and (n106,n107,n108);
nor (n108,n104,n109);
xnor (n109,n110,n105);
nand (n111,n112,n86);
nand (n112,n113,n127,n133);
nand (n113,n114,n123);
xor (n114,n115,n42);
or (n115,n116,n120);
and (n116,n39,n117);
xor (n117,n118,n119);
and (n120,n44,n121);
nor (n121,n117,n122);
xnor (n122,n42,n118);
xor (n123,n124,n15);
or (n124,n125,n126);
and (n125,n12,n95);
and (n126,n17,n98);
nand (n127,n128,n123);
xor (n128,n129,n20);
or (n129,n130,n132);
and (n130,n131,n13);
and (n132,n103,n18);
nand (n133,n114,n128);
nand (n134,n62,n112);
xor (n135,n136,n167);
xor (n136,n137,n153);
xor (n137,n138,n149);
xor (n138,n139,n145);
not (n139,n140);
xor (n140,n141,n42);
or (n141,n142,n144);
and (n142,n143,n117);
and (n144,n143,n121);
xor (n145,n146,n47);
or (n146,n147,n148);
and (n147,n143,n40);
and (n148,n39,n45);
xor (n149,n150,n35);
or (n150,n151,n152);
and (n151,n56,n28);
and (n152,n27,n33);
xor (n153,n154,n163);
xor (n154,n155,n159);
xor (n155,n156,n30);
or (n156,n157,n158);
and (n157,n44,n53);
and (n158,n52,n57);
xor (n159,n160,n84);
or (n160,n161,n162);
and (n161,n32,n78);
and (n162,n68,n82);
xor (n163,n164,n15);
or (n164,n165,n166);
and (n165,n77,n95);
and (n166,n81,n98);
nand (n167,n168,n169,n170);
nand (n168,n88,n92);
nand (n169,n100,n92);
nand (n170,n88,n100);
xor (n171,n172,n251);
xor (n172,n173,n231);
nand (n173,n174,n204,n230);
nand (n174,n175,n194);
nand (n175,n176,n192,n193);
nand (n176,n177,n182);
xor (n177,n178,n110);
or (n178,n179,n180);
and (n179,n107,n104);
and (n180,n181,n108);
xor (n182,n183,n21);
or (n183,n184,n188);
and (n184,n185,n186);
xor (n186,n187,n110);
and (n188,n189,n190);
nor (n190,n186,n191);
xnor (n191,n21,n187);
nand (n192,n21,n182);
nand (n193,n177,n21);
xor (n194,n195,n200);
xor (n195,n196,n139);
xor (n196,n197,n21);
or (n197,n198,n199);
and (n198,n181,n186);
and (n199,n185,n190);
xor (n200,n201,n20);
or (n201,n202,n203);
and (n202,n17,n13);
and (n203,n131,n18);
nand (n204,n205,n194);
xor (n205,n206,n228);
xor (n206,n21,n207);
nand (n207,n208,n222,n227);
nand (n208,n209,n212);
xor (n209,n210,n42);
or (n210,n142,n211);
and (n211,n39,n121);
not (n212,n213);
xor (n213,n214,n119);
or (n214,n215,n219);
and (n215,n143,n216);
xor (n216,n217,n218);
and (n219,n143,n220);
nor (n220,n216,n221);
xnor (n221,n119,n217);
nand (n222,n223,n212);
xor (n223,n224,n30);
or (n224,n225,n226);
and (n225,n56,n53);
and (n226,n27,n57);
nand (n227,n209,n223);
xor (n228,n229,n49);
xor (n229,n24,n36);
nand (n230,n175,n205);
xor (n231,n232,n247);
xor (n232,n233,n237);
nand (n233,n234,n235,n236);
nand (n234,n196,n139);
nand (n235,n200,n139);
nand (n236,n196,n200);
xor (n237,n238,n140);
xor (n238,n239,n243);
xor (n239,n240,n110);
or (n240,n241,n242);
and (n241,n131,n104);
and (n242,n103,n108);
xor (n243,n244,n21);
or (n244,n245,n246);
and (n245,n107,n186);
and (n246,n181,n190);
nand (n247,n248,n249,n250);
nand (n248,n21,n207);
nand (n249,n228,n207);
nand (n250,n21,n228);
nand (n251,n252,n308,n311);
nand (n252,n253,n273);
nand (n253,n254,n269,n272);
nand (n254,n255,n267);
nand (n255,n256,n261,n266);
nand (n256,n213,n257);
xor (n257,n258,n30);
or (n258,n259,n260);
and (n259,n27,n53);
and (n260,n32,n57);
nand (n261,n262,n257);
xor (n262,n263,n35);
or (n263,n264,n265);
and (n264,n68,n28);
and (n265,n77,n33);
nand (n266,n213,n262);
xor (n267,n268,n74);
xor (n268,n64,n69);
nand (n269,n270,n267);
xor (n270,n271,n223);
xor (n271,n209,n212);
nand (n272,n255,n270);
nand (n273,n274,n304,n307);
nand (n274,n275,n288);
nand (n275,n276,n282,n287);
nand (n276,n277,n281);
xor (n277,n278,n47);
or (n278,n279,n280);
and (n279,n52,n40);
and (n280,n56,n45);
not (n281,n114);
nand (n282,n283,n281);
xor (n283,n284,n84);
or (n284,n285,n286);
and (n285,n81,n78);
and (n286,n12,n82);
nand (n287,n277,n283);
nand (n288,n289,n298,n303);
nand (n289,n290,n294);
xor (n290,n291,n15);
or (n291,n292,n293);
and (n292,n17,n95);
and (n293,n131,n98);
xor (n294,n295,n20);
or (n295,n296,n297);
and (n296,n103,n13);
and (n297,n107,n18);
nand (n298,n299,n294);
xor (n299,n300,n110);
or (n300,n301,n302);
and (n301,n181,n104);
and (n302,n185,n108);
nand (n303,n290,n299);
nand (n304,n305,n288);
xor (n305,n306,n128);
xor (n306,n114,n123);
nand (n307,n275,n305);
nand (n308,n309,n273);
xor (n309,n310,n112);
xor (n310,n62,n86);
nand (n311,n253,n309);
nand (n312,n313,n171);
nand (n313,n314,n391,n394);
nand (n314,n315,n317);
xor (n315,n316,n205);
xor (n316,n175,n194);
nand (n317,n318,n351,n390);
nand (n318,n319,n349);
nand (n319,n320,n326,n348);
nand (n320,n321,n21);
xor (n321,n322,n21);
or (n322,n323,n324);
and (n323,n189,n186);
and (n324,n325,n190);
nand (n326,n327,n21);
nand (n327,n328,n336,n347);
nand (n328,n329,n332);
xor (n329,n330,n119);
or (n330,n215,n331);
and (n331,n39,n220);
xor (n332,n333,n42);
or (n333,n334,n335);
and (n334,n44,n117);
and (n335,n52,n121);
nand (n336,n337,n332);
not (n337,n338);
xor (n338,n339,n218);
or (n339,n340,n344);
and (n340,n143,n341);
xor (n341,n342,n343);
and (n344,n143,n345);
nor (n345,n341,n346);
xnor (n346,n218,n342);
nand (n347,n329,n337);
nand (n348,n321,n327);
xor (n349,n350,n21);
xor (n350,n177,n182);
nand (n351,n352,n349);
nand (n352,n353,n372,n389);
nand (n353,n354,n370);
nand (n354,n355,n364,n369);
nand (n355,n356,n360);
xor (n356,n357,n47);
or (n357,n358,n359);
and (n358,n56,n40);
and (n359,n27,n45);
xor (n360,n361,n30);
or (n361,n362,n363);
and (n362,n32,n53);
and (n363,n68,n57);
nand (n364,n365,n360);
xor (n365,n366,n35);
or (n366,n367,n368);
and (n367,n77,n28);
and (n368,n81,n33);
nand (n369,n356,n365);
xor (n370,n371,n262);
xor (n371,n213,n257);
nand (n372,n373,n370);
nand (n373,n374,n383,n388);
nand (n374,n375,n379);
xor (n375,n376,n15);
or (n376,n377,n378);
and (n377,n131,n95);
and (n378,n103,n98);
xor (n379,n380,n119);
or (n380,n381,n382);
and (n381,n39,n216);
and (n382,n44,n220);
nand (n383,n384,n379);
xor (n384,n385,n84);
or (n385,n386,n387);
and (n386,n12,n78);
and (n387,n17,n82);
nand (n388,n375,n384);
nand (n389,n354,n373);
nand (n390,n319,n352);
nand (n391,n392,n317);
xor (n392,n393,n309);
xor (n393,n253,n273);
nand (n394,n315,n392);
nand (n395,n5,n313);
xor (n396,n397,n472);
xor (n397,n398,n402);
nand (n398,n399,n400,n401);
nand (n399,n7,n60);
nand (n400,n135,n60);
nand (n401,n7,n135);
xor (n402,n403,n442);
xor (n403,n404,n408);
nand (n404,n405,n406,n407);
nand (n405,n233,n237);
nand (n406,n247,n237);
nand (n407,n233,n247);
xor (n408,n409,n428);
xor (n409,n410,n414);
nand (n410,n411,n412,n413);
nand (n411,n239,n243);
nand (n412,n140,n243);
nand (n413,n239,n140);
xor (n414,n415,n424);
xor (n415,n416,n420);
xor (n416,n417,n20);
or (n417,n418,n419);
and (n418,n81,n13);
and (n419,n12,n18);
xor (n420,n421,n110);
or (n421,n422,n423);
and (n422,n17,n104);
and (n423,n131,n108);
nand (n424,n425,n426,n427);
nand (n425,n139,n145);
nand (n426,n149,n145);
nand (n427,n139,n149);
xor (n428,n429,n438);
xor (n429,n430,n434);
xor (n430,n431,n15);
or (n431,n432,n433);
and (n432,n68,n95);
and (n433,n77,n98);
xor (n434,n435,n21);
or (n435,n436,n437);
and (n436,n103,n186);
and (n437,n107,n190);
not (n438,n439);
xor (n439,n440,n47);
or (n440,n147,n441);
and (n441,n143,n45);
xor (n442,n443,n468);
xor (n443,n444,n448);
nand (n444,n445,n446,n447);
nand (n445,n9,n21);
nand (n446,n22,n21);
nand (n447,n9,n22);
xor (n448,n449,n464);
xor (n449,n21,n450);
xor (n450,n451,n460);
xor (n451,n452,n456);
xor (n452,n453,n30);
or (n453,n454,n455);
and (n454,n39,n53);
and (n455,n44,n57);
xor (n456,n457,n35);
or (n457,n458,n459);
and (n458,n52,n28);
and (n459,n56,n33);
xor (n460,n461,n84);
or (n461,n462,n463);
and (n462,n27,n78);
and (n463,n32,n82);
nand (n464,n465,n466,n467);
nand (n465,n155,n159);
nand (n466,n163,n159);
nand (n467,n155,n163);
nand (n468,n469,n470,n471);
nand (n469,n137,n153);
nand (n470,n167,n153);
nand (n471,n137,n167);
nand (n472,n473,n474,n475);
nand (n473,n173,n231);
nand (n474,n251,n231);
nand (n475,n173,n251);
nand (n476,n477,n2434);
nand (n477,n478,n2008);
nor (n478,n479,n1976);
nor (n479,n480,n1449);
nor (n480,n481,n1434);
nor (n481,n482,n1155);
nand (n482,n483,n938);
nor (n483,n484,n837);
nor (n484,n485,n747);
nand (n485,n486,n662,n746);
nand (n486,n487,n564);
xor (n487,n488,n540);
xor (n488,n489,n514);
xor (n489,n490,n502);
xor (n490,n491,n496);
xor (n491,n492,n84);
or (n492,n493,n494);
and (n493,n325,n78);
and (n494,n495,n82);
xor (n496,n497,n15);
or (n497,n498,n500);
and (n498,n499,n95);
and (n500,n501,n98);
xor (n502,n503,n507);
xor (n503,n504,n218);
or (n504,n505,n506);
and (n505,n32,n341);
and (n506,n68,n345);
xnor (n507,n508,n343);
nor (n508,n509,n513);
and (n509,n27,n510);
and (n510,n511,n343);
not (n511,n512);
and (n513,n56,n512);
nand (n514,n515,n525,n539);
nand (n515,n516,n520);
xor (n516,n517,n84);
or (n517,n518,n519);
and (n518,n495,n78);
and (n519,n499,n82);
xor (n520,n521,n15);
or (n521,n522,n523);
and (n522,n501,n95);
and (n523,n524,n98);
nand (n525,n526,n520);
xor (n526,n527,n536);
xor (n527,n528,n532);
xor (n528,n529,n218);
or (n529,n530,n531);
and (n530,n68,n341);
and (n531,n77,n345);
xor (n532,n533,n42);
or (n533,n534,n535);
and (n534,n17,n117);
and (n535,n131,n121);
xnor (n536,n537,n20);
nand (n537,n538,n13);
nand (n539,n516,n526);
xor (n540,n541,n550);
xor (n541,n542,n546);
xor (n542,n543,n20);
or (n543,n544,n545);
and (n544,n524,n13);
and (n545,n538,n18);
nand (n546,n547,n548,n549);
nand (n547,n528,n532);
nand (n548,n536,n532);
nand (n549,n528,n536);
xor (n550,n551,n560);
xor (n551,n552,n556);
xor (n552,n553,n42);
or (n553,n554,n555);
and (n554,n12,n117);
and (n555,n17,n121);
xor (n556,n557,n119);
or (n557,n558,n559);
and (n558,n77,n216);
and (n559,n81,n220);
xor (n560,n561,n47);
or (n561,n562,n563);
and (n562,n131,n40);
and (n563,n103,n45);
nand (n564,n565,n619,n661);
nand (n565,n566,n568);
xor (n566,n567,n526);
xor (n567,n516,n520);
xor (n568,n569,n608);
xor (n569,n570,n586);
nand (n570,n571,n580,n585);
nand (n571,n572,n576);
xor (n572,n573,n42);
or (n573,n574,n575);
and (n574,n131,n117);
and (n575,n103,n121);
xor (n576,n577,n119);
or (n577,n578,n579);
and (n578,n12,n216);
and (n579,n17,n220);
nand (n580,n581,n576);
xor (n581,n582,n47);
or (n582,n583,n584);
and (n583,n107,n40);
and (n584,n181,n45);
nand (n585,n572,n581);
nand (n586,n587,n602,n607);
nand (n587,n588,n597);
xor (n588,n589,n593);
xnor (n589,n590,n343);
nor (n590,n591,n592);
and (n591,n68,n510);
and (n592,n32,n512);
xor (n593,n594,n218);
or (n594,n595,n596);
and (n595,n77,n341);
and (n596,n81,n345);
and (n597,n598,n15);
xnor (n598,n599,n343);
nor (n599,n600,n601);
and (n600,n77,n510);
and (n601,n68,n512);
nand (n602,n603,n597);
xor (n603,n604,n30);
or (n604,n605,n606);
and (n605,n185,n53);
and (n606,n189,n57);
nand (n607,n588,n603);
xor (n608,n609,n615);
xor (n609,n610,n614);
xor (n610,n611,n30);
or (n611,n612,n613);
and (n612,n181,n53);
and (n613,n185,n57);
and (n614,n589,n593);
xor (n615,n616,n35);
or (n616,n617,n618);
and (n617,n189,n28);
and (n618,n325,n33);
nand (n619,n620,n568);
nand (n620,n621,n645,n660);
nand (n621,n622,n643);
nand (n622,n623,n637,n642);
nand (n623,n624,n633);
and (n624,n625,n629);
xnor (n625,n626,n343);
nor (n626,n627,n628);
and (n627,n81,n510);
and (n628,n77,n512);
xor (n629,n630,n218);
or (n630,n631,n632);
and (n631,n12,n341);
and (n632,n17,n345);
xor (n633,n634,n30);
or (n634,n635,n636);
and (n635,n189,n53);
and (n636,n325,n57);
nand (n637,n638,n633);
xor (n638,n639,n35);
or (n639,n640,n641);
and (n640,n495,n28);
and (n641,n499,n33);
nand (n642,n624,n638);
xor (n643,n644,n603);
xor (n644,n588,n597);
nand (n645,n646,n643);
xor (n646,n647,n656);
xor (n647,n648,n652);
xor (n648,n649,n35);
or (n649,n650,n651);
and (n650,n325,n28);
and (n651,n495,n33);
xor (n652,n653,n84);
or (n653,n654,n655);
and (n654,n499,n78);
and (n655,n501,n82);
xor (n656,n657,n15);
or (n657,n658,n659);
and (n658,n524,n95);
and (n659,n538,n98);
nand (n660,n622,n646);
nand (n661,n566,n620);
nand (n662,n663,n564);
xor (n663,n664,n703);
xor (n664,n665,n669);
nand (n665,n666,n667,n668);
nand (n666,n570,n586);
nand (n667,n608,n586);
nand (n668,n570,n608);
xor (n669,n670,n692);
xor (n670,n671,n688);
nand (n671,n672,n682,n687);
nand (n672,n673,n677);
xor (n673,n674,n119);
or (n674,n675,n676);
and (n675,n81,n216);
and (n676,n12,n220);
xor (n677,n678,n20);
xnor (n678,n679,n343);
nor (n679,n680,n681);
and (n680,n32,n510);
and (n681,n27,n512);
nand (n682,n683,n677);
xor (n683,n684,n47);
or (n684,n685,n686);
and (n685,n103,n40);
and (n686,n107,n45);
nand (n687,n673,n683);
nand (n688,n689,n690,n691);
nand (n689,n610,n614);
nand (n690,n615,n614);
nand (n691,n610,n615);
xor (n692,n693,n699);
xor (n693,n694,n695);
and (n694,n678,n20);
xor (n695,n696,n30);
or (n696,n697,n698);
and (n697,n107,n53);
and (n698,n181,n57);
xor (n699,n700,n35);
or (n700,n701,n702);
and (n701,n185,n28);
and (n702,n189,n33);
nand (n703,n704,n711,n745);
nand (n704,n705,n709);
nand (n705,n706,n707,n708);
nand (n706,n648,n652);
nand (n707,n656,n652);
nand (n708,n648,n656);
xor (n709,n710,n683);
xor (n710,n673,n677);
nand (n711,n712,n709);
nand (n712,n713,n730,n744);
nand (n713,n714,n728);
nand (n714,n715,n724,n727);
nand (n715,n716,n720);
xor (n716,n717,n218);
or (n717,n718,n719);
and (n718,n81,n341);
and (n719,n12,n345);
xor (n720,n721,n42);
or (n721,n722,n723);
and (n722,n103,n117);
and (n723,n107,n121);
nand (n724,n725,n720);
xnor (n725,n726,n15);
nand (n726,n538,n95);
nand (n727,n716,n725);
xor (n728,n729,n581);
xor (n729,n572,n576);
nand (n730,n731,n728);
nand (n731,n732,n738,n743);
nand (n732,n733,n737);
xor (n733,n734,n119);
or (n734,n735,n736);
and (n735,n17,n216);
and (n736,n131,n220);
xor (n737,n598,n15);
nand (n738,n739,n737);
xor (n739,n740,n47);
or (n740,n741,n742);
and (n741,n181,n40);
and (n742,n185,n45);
nand (n743,n733,n739);
nand (n744,n714,n731);
nand (n745,n705,n712);
nand (n746,n487,n663);
xor (n747,n748,n833);
xor (n748,n749,n770);
xor (n749,n750,n766);
xor (n750,n751,n762);
xor (n751,n752,n758);
xor (n752,n753,n757);
xor (n753,n754,n15);
or (n754,n755,n756);
and (n755,n495,n95);
and (n756,n499,n98);
and (n757,n503,n507);
xor (n758,n759,n20);
or (n759,n760,n761);
and (n760,n501,n13);
and (n761,n524,n18);
nand (n762,n763,n764,n765);
nand (n763,n542,n546);
nand (n764,n550,n546);
nand (n765,n542,n550);
nand (n766,n767,n768,n769);
nand (n767,n671,n688);
nand (n768,n692,n688);
nand (n769,n671,n692);
xor (n770,n771,n829);
xor (n771,n772,n796);
xor (n772,n773,n792);
xor (n773,n774,n778);
nand (n774,n775,n776,n777);
nand (n775,n694,n695);
nand (n776,n699,n695);
nand (n777,n694,n699);
xor (n778,n779,n788);
xor (n779,n780,n784);
xnor (n780,n781,n343);
nor (n781,n782,n783);
and (n782,n56,n510);
and (n783,n52,n512);
xor (n784,n785,n42);
or (n785,n786,n787);
and (n786,n81,n117);
and (n787,n12,n121);
xor (n788,n789,n119);
or (n789,n790,n791);
and (n790,n68,n216);
and (n791,n77,n220);
nand (n792,n793,n794,n795);
nand (n793,n552,n556);
nand (n794,n560,n556);
nand (n795,n552,n560);
xor (n796,n797,n815);
xor (n797,n798,n802);
nand (n798,n799,n800,n801);
nand (n799,n491,n496);
nand (n800,n502,n496);
nand (n801,n491,n502);
xor (n802,n803,n813);
xor (n803,n804,n808);
xor (n804,n805,n47);
or (n805,n806,n807);
and (n806,n17,n40);
and (n807,n131,n45);
xor (n808,n110,n809);
xor (n809,n810,n218);
or (n810,n811,n812);
and (n811,n27,n341);
and (n812,n32,n345);
xnor (n813,n814,n110);
nand (n814,n538,n104);
xor (n815,n816,n825);
xor (n816,n817,n821);
xor (n817,n818,n30);
or (n818,n819,n820);
and (n819,n103,n53);
and (n820,n107,n57);
xor (n821,n822,n35);
or (n822,n823,n824);
and (n823,n181,n28);
and (n824,n185,n33);
xor (n825,n826,n84);
or (n826,n827,n828);
and (n827,n189,n78);
and (n828,n325,n82);
nand (n829,n830,n831,n832);
nand (n830,n489,n514);
nand (n831,n540,n514);
nand (n832,n489,n540);
nand (n833,n834,n835,n836);
nand (n834,n665,n669);
nand (n835,n703,n669);
nand (n836,n665,n703);
nor (n837,n838,n842);
nand (n838,n839,n840,n841);
nand (n839,n749,n770);
nand (n840,n833,n770);
nand (n841,n749,n833);
xor (n842,n843,n852);
xor (n843,n844,n848);
nand (n844,n845,n846,n847);
nand (n845,n751,n762);
nand (n846,n766,n762);
nand (n847,n751,n766);
nand (n848,n849,n850,n851);
nand (n849,n772,n796);
nand (n850,n829,n796);
nand (n851,n772,n829);
xor (n852,n853,n914);
xor (n853,n854,n885);
xor (n854,n855,n874);
xor (n855,n856,n870);
xor (n856,n857,n866);
xor (n857,n858,n862);
xor (n858,n859,n42);
or (n859,n860,n861);
and (n860,n77,n117);
and (n861,n81,n121);
xor (n862,n863,n119);
or (n863,n864,n865);
and (n864,n32,n216);
and (n865,n68,n220);
xor (n866,n867,n47);
or (n867,n868,n869);
and (n868,n12,n40);
and (n869,n17,n45);
nand (n870,n871,n872,n873);
nand (n871,n804,n808);
nand (n872,n813,n808);
nand (n873,n804,n813);
xor (n874,n875,n881);
xor (n875,n876,n880);
xor (n876,n877,n30);
or (n877,n878,n879);
and (n878,n131,n53);
and (n879,n103,n57);
and (n880,n110,n809);
xor (n881,n882,n35);
or (n882,n883,n884);
and (n883,n107,n28);
and (n884,n181,n33);
xor (n885,n886,n910);
xor (n886,n887,n891);
nand (n887,n888,n889,n890);
nand (n888,n817,n821);
nand (n889,n825,n821);
nand (n890,n817,n825);
xor (n891,n892,n901);
xor (n892,n893,n897);
xor (n893,n894,n84);
or (n894,n895,n896);
and (n895,n185,n78);
and (n896,n189,n82);
xor (n897,n898,n15);
or (n898,n899,n900);
and (n899,n325,n95);
and (n900,n495,n98);
xor (n901,n902,n906);
xnor (n902,n903,n343);
nor (n903,n904,n905);
and (n904,n52,n510);
and (n905,n44,n512);
xor (n906,n907,n218);
or (n907,n908,n909);
and (n908,n56,n341);
and (n909,n27,n345);
nand (n910,n911,n912,n913);
nand (n911,n753,n757);
nand (n912,n758,n757);
nand (n913,n753,n758);
xor (n914,n915,n934);
xor (n915,n916,n930);
xor (n916,n917,n926);
xor (n917,n918,n922);
xor (n918,n919,n20);
or (n919,n920,n921);
and (n920,n499,n13);
and (n921,n501,n18);
xor (n922,n923,n110);
or (n923,n924,n925);
and (n924,n524,n104);
and (n925,n538,n108);
nand (n926,n927,n928,n929);
nand (n927,n780,n784);
nand (n928,n788,n784);
nand (n929,n780,n788);
nand (n930,n931,n932,n933);
nand (n931,n774,n778);
nand (n932,n792,n778);
nand (n933,n774,n792);
nand (n934,n935,n936,n937);
nand (n935,n798,n802);
nand (n936,n815,n802);
nand (n937,n798,n815);
nor (n938,n939,n1044);
nor (n939,n940,n944);
nand (n940,n941,n942,n943);
nand (n941,n844,n848);
nand (n942,n852,n848);
nand (n943,n844,n852);
xor (n944,n945,n1040);
xor (n945,n946,n980);
xor (n946,n947,n976);
xor (n947,n948,n952);
nand (n948,n949,n950,n951);
nand (n949,n856,n870);
nand (n950,n874,n870);
nand (n951,n856,n874);
xor (n952,n953,n962);
xor (n953,n954,n958);
xor (n954,n955,n110);
or (n955,n956,n957);
and (n956,n501,n104);
and (n957,n524,n108);
nand (n958,n959,n960,n961);
nand (n959,n876,n880);
nand (n960,n881,n880);
nand (n961,n876,n881);
xor (n962,n963,n972);
xor (n963,n964,n968);
xor (n964,n965,n42);
or (n965,n966,n967);
and (n966,n68,n117);
and (n967,n77,n121);
xnor (n968,n969,n343);
nor (n969,n970,n971);
and (n970,n44,n510);
and (n971,n39,n512);
xor (n972,n973,n119);
or (n973,n974,n975);
and (n974,n27,n216);
and (n975,n32,n220);
nand (n976,n977,n978,n979);
nand (n977,n887,n891);
nand (n978,n910,n891);
nand (n979,n887,n910);
xor (n980,n981,n1036);
xor (n981,n982,n1004);
xor (n982,n983,n992);
xor (n983,n984,n988);
nand (n984,n985,n986,n987);
nand (n985,n858,n862);
nand (n986,n866,n862);
nand (n987,n858,n866);
nand (n988,n989,n990,n991);
nand (n989,n893,n897);
nand (n990,n901,n897);
nand (n991,n893,n901);
xor (n992,n993,n1000);
xor (n993,n994,n998);
xor (n994,n995,n47);
or (n995,n996,n997);
and (n996,n81,n40);
and (n997,n12,n45);
xnor (n998,n999,n21);
nand (n999,n538,n186);
xor (n1000,n1001,n30);
or (n1001,n1002,n1003);
and (n1002,n17,n53);
and (n1003,n131,n57);
xor (n1004,n1005,n1024);
xor (n1005,n1006,n1010);
nand (n1006,n1007,n1008,n1009);
nand (n1007,n918,n922);
nand (n1008,n926,n922);
nand (n1009,n918,n926);
xor (n1010,n1011,n1020);
xor (n1011,n1012,n1016);
xor (n1012,n1013,n35);
or (n1013,n1014,n1015);
and (n1014,n103,n28);
and (n1015,n107,n33);
xor (n1016,n1017,n84);
or (n1017,n1018,n1019);
and (n1018,n181,n78);
and (n1019,n185,n82);
xor (n1020,n1021,n15);
or (n1021,n1022,n1023);
and (n1022,n189,n95);
and (n1023,n325,n98);
xor (n1024,n1025,n1032);
xor (n1025,n1026,n1031);
xor (n1026,n21,n1027);
xor (n1027,n1028,n218);
or (n1028,n1029,n1030);
and (n1029,n52,n341);
and (n1030,n56,n345);
and (n1031,n902,n906);
xor (n1032,n1033,n20);
or (n1033,n1034,n1035);
and (n1034,n495,n13);
and (n1035,n499,n18);
nand (n1036,n1037,n1038,n1039);
nand (n1037,n916,n930);
nand (n1038,n934,n930);
nand (n1039,n916,n934);
nand (n1040,n1041,n1042,n1043);
nand (n1041,n854,n885);
nand (n1042,n914,n885);
nand (n1043,n854,n914);
nor (n1044,n1045,n1049);
nand (n1045,n1046,n1047,n1048);
nand (n1046,n946,n980);
nand (n1047,n1040,n980);
nand (n1048,n946,n1040);
xor (n1049,n1050,n1059);
xor (n1050,n1051,n1055);
nand (n1051,n1052,n1053,n1054);
nand (n1052,n948,n952);
nand (n1053,n976,n952);
nand (n1054,n948,n976);
nand (n1055,n1056,n1057,n1058);
nand (n1056,n982,n1004);
nand (n1057,n1036,n1004);
nand (n1058,n982,n1036);
xor (n1059,n1060,n1121);
xor (n1060,n1061,n1085);
xor (n1061,n1062,n1081);
xor (n1062,n1063,n1067);
nand (n1063,n1064,n1065,n1066);
nand (n1064,n1012,n1016);
nand (n1065,n1020,n1016);
nand (n1066,n1012,n1020);
xor (n1067,n1068,n1077);
xor (n1068,n1069,n1073);
xor (n1069,n1070,n30);
or (n1070,n1071,n1072);
and (n1071,n12,n53);
and (n1072,n17,n57);
xor (n1073,n1074,n35);
or (n1074,n1075,n1076);
and (n1075,n131,n28);
and (n1076,n103,n33);
xor (n1077,n1078,n84);
or (n1078,n1079,n1080);
and (n1079,n107,n78);
and (n1080,n181,n82);
nand (n1081,n1082,n1083,n1084);
nand (n1082,n1026,n1031);
nand (n1083,n1032,n1031);
nand (n1084,n1026,n1032);
xor (n1085,n1086,n1107);
xor (n1086,n1087,n1103);
xor (n1087,n1088,n1102);
xor (n1088,n1089,n1093);
xor (n1089,n1090,n15);
or (n1090,n1091,n1092);
and (n1091,n185,n95);
and (n1092,n189,n98);
xor (n1093,n1094,n1098);
xnor (n1094,n1095,n343);
nor (n1095,n1096,n1097);
and (n1096,n39,n510);
and (n1097,n143,n512);
xor (n1098,n1099,n218);
or (n1099,n1100,n1101);
and (n1100,n44,n341);
and (n1101,n52,n345);
and (n1102,n21,n1027);
nand (n1103,n1104,n1105,n1106);
nand (n1104,n954,n958);
nand (n1105,n962,n958);
nand (n1106,n954,n962);
xor (n1107,n1108,n1117);
xor (n1108,n1109,n1113);
xor (n1109,n1110,n20);
or (n1110,n1111,n1112);
and (n1111,n325,n13);
and (n1112,n495,n18);
xor (n1113,n1114,n21);
or (n1114,n1115,n1116);
and (n1115,n524,n186);
and (n1116,n538,n190);
xor (n1117,n1118,n110);
or (n1118,n1119,n1120);
and (n1119,n499,n104);
and (n1120,n501,n108);
xor (n1121,n1122,n1151);
xor (n1122,n1123,n1147);
xor (n1123,n1124,n1143);
xor (n1124,n1125,n1129);
nand (n1125,n1126,n1127,n1128);
nand (n1126,n964,n968);
nand (n1127,n972,n968);
nand (n1128,n964,n972);
xor (n1129,n1130,n1139);
xor (n1130,n1131,n1135);
xor (n1131,n1132,n42);
or (n1132,n1133,n1134);
and (n1133,n32,n117);
and (n1134,n68,n121);
xor (n1135,n1136,n119);
or (n1136,n1137,n1138);
and (n1137,n56,n216);
and (n1138,n27,n220);
xor (n1139,n1140,n47);
or (n1140,n1141,n1142);
and (n1141,n77,n40);
and (n1142,n81,n45);
nand (n1143,n1144,n1145,n1146);
nand (n1144,n994,n998);
nand (n1145,n1000,n998);
nand (n1146,n994,n1000);
nand (n1147,n1148,n1149,n1150);
nand (n1148,n984,n988);
nand (n1149,n992,n988);
nand (n1150,n984,n992);
nand (n1151,n1152,n1153,n1154);
nand (n1152,n1006,n1010);
nand (n1153,n1024,n1010);
nand (n1154,n1006,n1024);
nor (n1155,n1156,n1428);
nor (n1156,n1157,n1404);
nor (n1157,n1158,n1402);
nor (n1158,n1159,n1377);
nand (n1159,n1160,n1339);
nand (n1160,n1161,n1286,n1338);
nand (n1161,n1162,n1213);
xor (n1162,n1163,n1200);
xor (n1163,n1164,n1185);
nand (n1164,n1165,n1179,n1184);
nand (n1165,n1166,n1175);
and (n1166,n1167,n1171);
xnor (n1167,n1168,n343);
nor (n1168,n1169,n1170);
and (n1169,n17,n510);
and (n1170,n12,n512);
xor (n1171,n1172,n218);
or (n1172,n1173,n1174);
and (n1173,n131,n341);
and (n1174,n103,n345);
xor (n1175,n1176,n30);
or (n1176,n1177,n1178);
and (n1177,n495,n53);
and (n1178,n499,n57);
nand (n1179,n1180,n1175);
xor (n1180,n1181,n35);
or (n1181,n1182,n1183);
and (n1182,n501,n28);
and (n1183,n524,n33);
nand (n1184,n1166,n1180);
xor (n1185,n1186,n1195);
xor (n1186,n1187,n1191);
xor (n1187,n1188,n42);
or (n1188,n1189,n1190);
and (n1189,n107,n117);
and (n1190,n181,n121);
xor (n1191,n1192,n119);
or (n1192,n1193,n1194);
and (n1193,n131,n216);
and (n1194,n103,n220);
and (n1195,n1196,n84);
xnor (n1196,n1197,n343);
nor (n1197,n1198,n1199);
and (n1198,n12,n510);
and (n1199,n81,n512);
nand (n1200,n1201,n1207,n1212);
nand (n1201,n1202,n1206);
xor (n1202,n1203,n119);
or (n1203,n1204,n1205);
and (n1204,n103,n216);
and (n1205,n107,n220);
xor (n1206,n1196,n84);
nand (n1207,n1208,n1206);
xor (n1208,n1209,n47);
or (n1209,n1210,n1211);
and (n1210,n189,n40);
and (n1211,n325,n45);
nand (n1212,n1202,n1208);
xor (n1213,n1214,n1250);
xor (n1214,n1215,n1226);
xor (n1215,n1216,n1222);
xor (n1216,n1217,n1221);
xor (n1217,n1218,n47);
or (n1218,n1219,n1220);
and (n1219,n185,n40);
and (n1220,n189,n45);
xor (n1221,n625,n629);
xor (n1222,n1223,n30);
or (n1223,n1224,n1225);
and (n1224,n325,n53);
and (n1225,n495,n57);
xor (n1226,n1227,n1236);
xor (n1227,n1228,n1232);
xor (n1228,n1229,n35);
or (n1229,n1230,n1231);
and (n1230,n499,n28);
and (n1231,n501,n33);
xor (n1232,n1233,n84);
or (n1233,n1234,n1235);
and (n1234,n524,n78);
and (n1235,n538,n82);
nand (n1236,n1237,n1244,n1249);
nand (n1237,n1238,n1242);
xor (n1238,n1239,n218);
or (n1239,n1240,n1241);
and (n1240,n17,n341);
and (n1241,n131,n345);
xnor (n1242,n1243,n84);
nand (n1243,n538,n78);
nand (n1244,n1245,n1242);
xor (n1245,n1246,n42);
or (n1246,n1247,n1248);
and (n1247,n181,n117);
and (n1248,n185,n121);
nand (n1249,n1238,n1245);
nand (n1250,n1251,n1271,n1285);
nand (n1251,n1252,n1254);
xor (n1252,n1253,n1245);
xor (n1253,n1238,n1242);
nand (n1254,n1255,n1264,n1270);
nand (n1255,n1256,n1260);
xor (n1256,n1257,n42);
or (n1257,n1258,n1259);
and (n1258,n185,n117);
and (n1259,n189,n121);
xor (n1260,n1261,n119);
or (n1261,n1262,n1263);
and (n1262,n107,n216);
and (n1263,n181,n220);
nand (n1264,n1265,n1260);
and (n1265,n1266,n35);
xnor (n1266,n1267,n343);
nor (n1267,n1268,n1269);
and (n1268,n131,n510);
and (n1269,n17,n512);
nand (n1270,n1256,n1265);
nand (n1271,n1272,n1254);
nand (n1272,n1273,n1279,n1284);
nand (n1273,n1274,n1278);
xor (n1274,n1275,n47);
or (n1275,n1276,n1277);
and (n1276,n325,n40);
and (n1277,n495,n45);
xor (n1278,n1167,n1171);
nand (n1279,n1280,n1278);
xor (n1280,n1281,n30);
or (n1281,n1282,n1283);
and (n1282,n499,n53);
and (n1283,n501,n57);
nand (n1284,n1274,n1280);
nand (n1285,n1252,n1272);
nand (n1286,n1287,n1213);
nand (n1287,n1288,n1293,n1337);
nand (n1288,n1289,n1291);
xor (n1289,n1290,n1180);
xor (n1290,n1166,n1175);
xor (n1291,n1292,n1208);
xor (n1292,n1202,n1206);
nand (n1293,n1294,n1291);
nand (n1294,n1295,n1314,n1336);
nand (n1295,n1296,n1300);
xor (n1296,n1297,n35);
or (n1297,n1298,n1299);
and (n1298,n524,n28);
and (n1299,n538,n33);
nand (n1300,n1301,n1308,n1313);
nand (n1301,n1302,n1306);
xor (n1302,n1303,n218);
or (n1303,n1304,n1305);
and (n1304,n103,n341);
and (n1305,n107,n345);
xnor (n1306,n1307,n35);
nand (n1307,n538,n28);
nand (n1308,n1309,n1306);
xor (n1309,n1310,n42);
or (n1310,n1311,n1312);
and (n1311,n189,n117);
and (n1312,n325,n121);
nand (n1313,n1302,n1309);
nand (n1314,n1315,n1300);
nand (n1315,n1316,n1330,n1335);
nand (n1316,n1317,n1321);
xor (n1317,n1318,n119);
or (n1318,n1319,n1320);
and (n1319,n181,n216);
and (n1320,n185,n220);
and (n1321,n1322,n1326);
xnor (n1322,n1323,n343);
nor (n1323,n1324,n1325);
and (n1324,n103,n510);
and (n1325,n131,n512);
xor (n1326,n1327,n218);
or (n1327,n1328,n1329);
and (n1328,n107,n341);
and (n1329,n181,n345);
nand (n1330,n1331,n1321);
xor (n1331,n1332,n47);
or (n1332,n1333,n1334);
and (n1333,n495,n40);
and (n1334,n499,n45);
nand (n1335,n1317,n1331);
nand (n1336,n1296,n1315);
nand (n1337,n1289,n1294);
nand (n1338,n1162,n1287);
xor (n1339,n1340,n1355);
xor (n1340,n1341,n1351);
xor (n1341,n1342,n1349);
xor (n1342,n1343,n1347);
nand (n1343,n1344,n1345,n1346);
nand (n1344,n1187,n1191);
nand (n1345,n1195,n1191);
nand (n1346,n1187,n1195);
xor (n1347,n1348,n638);
xor (n1348,n624,n633);
xor (n1349,n1350,n739);
xor (n1350,n733,n737);
nand (n1351,n1352,n1353,n1354);
nand (n1352,n1215,n1226);
nand (n1353,n1250,n1226);
nand (n1354,n1215,n1250);
xor (n1355,n1356,n1365);
xor (n1356,n1357,n1361);
nand (n1357,n1358,n1359,n1360);
nand (n1358,n1228,n1232);
nand (n1359,n1236,n1232);
nand (n1360,n1228,n1236);
nand (n1361,n1362,n1363,n1364);
nand (n1362,n1164,n1185);
nand (n1363,n1200,n1185);
nand (n1364,n1164,n1200);
xor (n1365,n1366,n1375);
xor (n1366,n1367,n1371);
xor (n1367,n1368,n84);
or (n1368,n1369,n1370);
and (n1369,n501,n78);
and (n1370,n524,n82);
nand (n1371,n1372,n1373,n1374);
nand (n1372,n1217,n1221);
nand (n1373,n1222,n1221);
nand (n1374,n1217,n1222);
xor (n1375,n1376,n725);
xor (n1376,n716,n720);
nor (n1377,n1378,n1382);
nand (n1378,n1379,n1380,n1381);
nand (n1379,n1341,n1351);
nand (n1380,n1355,n1351);
nand (n1381,n1341,n1355);
xor (n1382,n1383,n1390);
xor (n1383,n1384,n1386);
xor (n1384,n1385,n646);
xor (n1385,n622,n643);
nand (n1386,n1387,n1388,n1389);
nand (n1387,n1357,n1361);
nand (n1388,n1365,n1361);
nand (n1389,n1357,n1365);
xor (n1390,n1391,n1400);
xor (n1391,n1392,n1396);
nand (n1392,n1393,n1394,n1395);
nand (n1393,n1367,n1371);
nand (n1394,n1375,n1371);
nand (n1395,n1367,n1375);
nand (n1396,n1397,n1398,n1399);
nand (n1397,n1343,n1347);
nand (n1398,n1349,n1347);
nand (n1399,n1343,n1349);
xor (n1400,n1401,n731);
xor (n1401,n714,n728);
not (n1402,n1403);
nand (n1403,n1378,n1382);
not (n1404,n1405);
nor (n1405,n1406,n1421);
nor (n1406,n1407,n1411);
nand (n1407,n1408,n1409,n1410);
nand (n1408,n1384,n1386);
nand (n1409,n1390,n1386);
nand (n1410,n1384,n1390);
xor (n1411,n1412,n1419);
xor (n1412,n1413,n1415);
xor (n1413,n1414,n712);
xor (n1414,n705,n709);
nand (n1415,n1416,n1417,n1418);
nand (n1416,n1392,n1396);
nand (n1417,n1400,n1396);
nand (n1418,n1392,n1400);
xor (n1419,n1420,n620);
xor (n1420,n566,n568);
nor (n1421,n1422,n1426);
nand (n1422,n1423,n1424,n1425);
nand (n1423,n1413,n1415);
nand (n1424,n1419,n1415);
nand (n1425,n1413,n1419);
xor (n1426,n1427,n663);
xor (n1427,n487,n564);
not (n1428,n1429);
nor (n1429,n1430,n1432);
nor (n1430,n1431,n1421);
nand (n1431,n1407,n1411);
not (n1432,n1433);
nand (n1433,n1422,n1426);
not (n1434,n1435);
nor (n1435,n1436,n1443);
nor (n1436,n1437,n1442);
nor (n1437,n1438,n1440);
nor (n1438,n1439,n837);
nand (n1439,n485,n747);
not (n1440,n1441);
nand (n1441,n838,n842);
not (n1442,n938);
not (n1443,n1444);
nor (n1444,n1445,n1447);
nor (n1445,n1446,n1044);
nand (n1446,n940,n944);
not (n1447,n1448);
nand (n1448,n1045,n1049);
not (n1449,n1450);
nor (n1450,n1451,n1866);
nand (n1451,n1452,n1679);
nor (n1452,n1453,n1565);
nor (n1453,n1454,n1458);
nand (n1454,n1455,n1456,n1457);
nand (n1455,n1051,n1055);
nand (n1456,n1059,n1055);
nand (n1457,n1051,n1059);
xor (n1458,n1459,n1561);
xor (n1459,n1460,n1493);
xor (n1460,n1461,n1489);
xor (n1461,n1462,n1485);
xor (n1462,n1463,n1481);
xor (n1463,n1464,n1477);
xor (n1464,n1465,n1474);
xor (n1465,n1466,n1470);
xor (n1466,n1467,n218);
or (n1467,n1468,n1469);
and (n1468,n39,n341);
and (n1469,n44,n345);
xor (n1470,n1471,n119);
or (n1471,n1472,n1473);
and (n1472,n52,n216);
and (n1473,n56,n220);
xnor (n1474,n1475,n343);
nor (n1475,n1476,n1097);
and (n1476,n143,n510);
nand (n1477,n1478,n1479,n1480);
nand (n1478,n1069,n1073);
nand (n1479,n1077,n1073);
nand (n1480,n1069,n1077);
nand (n1481,n1482,n1483,n1484);
nand (n1482,n1089,n1093);
nand (n1483,n1102,n1093);
nand (n1484,n1089,n1102);
nand (n1485,n1486,n1487,n1488);
nand (n1486,n1063,n1067);
nand (n1487,n1081,n1067);
nand (n1488,n1063,n1081);
nand (n1489,n1490,n1491,n1492);
nand (n1490,n1087,n1103);
nand (n1491,n1107,n1103);
nand (n1492,n1087,n1107);
xor (n1493,n1494,n1557);
xor (n1494,n1495,n1533);
xor (n1495,n1496,n1518);
xor (n1496,n1497,n1511);
xor (n1497,n1498,n1507);
xor (n1498,n1499,n1503);
xor (n1499,n1500,n47);
or (n1500,n1501,n1502);
and (n1501,n68,n40);
and (n1502,n77,n45);
xor (n1503,n1504,n30);
or (n1504,n1505,n1506);
and (n1505,n81,n53);
and (n1506,n12,n57);
xor (n1507,n1508,n35);
or (n1508,n1509,n1510);
and (n1509,n17,n28);
and (n1510,n131,n33);
xor (n1511,n1512,n1514);
xor (n1512,n21,n1513);
and (n1513,n1094,n1098);
xor (n1514,n1515,n20);
or (n1515,n1516,n1517);
and (n1516,n189,n13);
and (n1517,n325,n18);
xor (n1518,n1519,n1528);
xor (n1519,n1520,n1524);
xor (n1520,n1521,n84);
or (n1521,n1522,n1523);
and (n1522,n103,n78);
and (n1523,n107,n82);
xor (n1524,n1525,n15);
or (n1525,n1526,n1527);
and (n1526,n181,n95);
and (n1527,n185,n98);
xor (n1528,n21,n1529);
xor (n1529,n1530,n42);
or (n1530,n1531,n1532);
and (n1531,n27,n117);
and (n1532,n32,n121);
xor (n1533,n1534,n1543);
xor (n1534,n1535,n1539);
nand (n1535,n1536,n1537,n1538);
nand (n1536,n1109,n1113);
nand (n1537,n1117,n1113);
nand (n1538,n1109,n1117);
nand (n1539,n1540,n1541,n1542);
nand (n1540,n1125,n1129);
nand (n1541,n1143,n1129);
nand (n1542,n1125,n1143);
xor (n1543,n1544,n1553);
xor (n1544,n1545,n1549);
xor (n1545,n1546,n110);
or (n1546,n1547,n1548);
and (n1547,n495,n104);
and (n1548,n499,n108);
xor (n1549,n1550,n21);
or (n1550,n1551,n1552);
and (n1551,n501,n186);
and (n1552,n524,n190);
nand (n1553,n1554,n1555,n1556);
nand (n1554,n1131,n1135);
nand (n1555,n1139,n1135);
nand (n1556,n1131,n1139);
nand (n1557,n1558,n1559,n1560);
nand (n1558,n1123,n1147);
nand (n1559,n1151,n1147);
nand (n1560,n1123,n1151);
nand (n1561,n1562,n1563,n1564);
nand (n1562,n1061,n1085);
nand (n1563,n1121,n1085);
nand (n1564,n1061,n1121);
nor (n1565,n1566,n1570);
nand (n1566,n1567,n1568,n1569);
nand (n1567,n1460,n1493);
nand (n1568,n1561,n1493);
nand (n1569,n1460,n1561);
xor (n1570,n1571,n1580);
xor (n1571,n1572,n1576);
nand (n1572,n1573,n1574,n1575);
nand (n1573,n1462,n1485);
nand (n1574,n1489,n1485);
nand (n1575,n1462,n1489);
nand (n1576,n1577,n1578,n1579);
nand (n1577,n1495,n1533);
nand (n1578,n1557,n1533);
nand (n1579,n1495,n1557);
xor (n1580,n1581,n1638);
xor (n1581,n1582,n1613);
xor (n1582,n1583,n1599);
xor (n1583,n1584,n1588);
nand (n1584,n1585,n1586,n1587);
nand (n1585,n21,n1513);
nand (n1586,n1514,n1513);
nand (n1587,n21,n1514);
xor (n1588,n1589,n1595);
xor (n1589,n1590,n1594);
xor (n1590,n1591,n15);
or (n1591,n1592,n1593);
and (n1592,n107,n95);
and (n1593,n181,n98);
and (n1594,n21,n1529);
xor (n1595,n1596,n20);
or (n1596,n1597,n1598);
and (n1597,n185,n13);
and (n1598,n189,n18);
xor (n1599,n1600,n1609);
xor (n1600,n1601,n1605);
xor (n1601,n1602,n110);
or (n1602,n1603,n1604);
and (n1603,n325,n104);
and (n1604,n495,n108);
xor (n1605,n1606,n21);
or (n1606,n1607,n1608);
and (n1607,n499,n186);
and (n1608,n501,n190);
nand (n1609,n1610,n1611,n1612);
nand (n1610,n1466,n1470);
nand (n1611,n1474,n1470);
nand (n1612,n1466,n1474);
xor (n1613,n1614,n1623);
xor (n1614,n1615,n1619);
nand (n1615,n1616,n1617,n1618);
nand (n1616,n1545,n1549);
nand (n1617,n1553,n1549);
nand (n1618,n1545,n1553);
nand (n1619,n1620,n1621,n1622);
nand (n1620,n1464,n1477);
nand (n1621,n1481,n1477);
nand (n1622,n1464,n1481);
xor (n1623,n1624,n21);
xor (n1624,n1625,n1629);
nand (n1625,n1626,n1627,n1628);
nand (n1626,n1499,n1503);
nand (n1627,n1507,n1503);
nand (n1628,n1499,n1507);
xor (n1629,n1630,n1635);
not (n1630,n1631);
xor (n1631,n1632,n42);
or (n1632,n1633,n1634);
and (n1633,n56,n117);
and (n1634,n27,n121);
xor (n1635,n1636,n218);
or (n1636,n340,n1637);
and (n1637,n39,n345);
xor (n1638,n1639,n1675);
xor (n1639,n1640,n1644);
nand (n1640,n1641,n1642,n1643);
nand (n1641,n1497,n1511);
nand (n1642,n1518,n1511);
nand (n1643,n1497,n1518);
xor (n1644,n1645,n1664);
xor (n1645,n1646,n1650);
nand (n1646,n1647,n1648,n1649);
nand (n1647,n1520,n1524);
nand (n1648,n1528,n1524);
nand (n1649,n1520,n1528);
xor (n1650,n1651,n1660);
xor (n1651,n1652,n1656);
xor (n1652,n1653,n30);
or (n1653,n1654,n1655);
and (n1654,n77,n53);
and (n1655,n81,n57);
xor (n1656,n1657,n35);
or (n1657,n1658,n1659);
and (n1658,n12,n28);
and (n1659,n17,n33);
xor (n1660,n1661,n84);
or (n1661,n1662,n1663);
and (n1662,n131,n78);
and (n1663,n103,n82);
xor (n1664,n1665,n1671);
xor (n1665,n1666,n1670);
xor (n1666,n1667,n119);
or (n1667,n1668,n1669);
and (n1668,n44,n216);
and (n1669,n52,n220);
not (n1670,n1474);
xor (n1671,n1672,n47);
or (n1672,n1673,n1674);
and (n1673,n32,n40);
and (n1674,n68,n45);
nand (n1675,n1676,n1677,n1678);
nand (n1676,n1535,n1539);
nand (n1677,n1543,n1539);
nand (n1678,n1535,n1543);
nor (n1679,n1680,n1787);
nor (n1680,n1681,n1685);
nand (n1681,n1682,n1683,n1684);
nand (n1682,n1572,n1576);
nand (n1683,n1580,n1576);
nand (n1684,n1572,n1580);
xor (n1685,n1686,n1783);
xor (n1686,n1687,n1727);
xor (n1687,n1688,n1723);
xor (n1688,n1689,n1719);
xor (n1689,n1690,n1715);
xor (n1690,n1691,n1705);
xor (n1691,n1692,n1701);
xor (n1692,n1693,n1697);
xor (n1693,n1694,n30);
or (n1694,n1695,n1696);
and (n1695,n68,n53);
and (n1696,n77,n57);
xor (n1697,n1698,n35);
or (n1698,n1699,n1700);
and (n1699,n81,n28);
and (n1700,n12,n33);
xor (n1701,n1702,n15);
or (n1702,n1703,n1704);
and (n1703,n103,n95);
and (n1704,n107,n98);
xor (n1705,n1706,n1711);
xor (n1706,n1707,n338);
xor (n1707,n1708,n42);
or (n1708,n1709,n1710);
and (n1709,n52,n117);
and (n1710,n56,n121);
xor (n1711,n1712,n47);
or (n1712,n1713,n1714);
and (n1713,n27,n40);
and (n1714,n32,n45);
nand (n1715,n1716,n1717,n1718);
nand (n1716,n1590,n1594);
nand (n1717,n1595,n1594);
nand (n1718,n1590,n1595);
nand (n1719,n1720,n1721,n1722);
nand (n1720,n1584,n1588);
nand (n1721,n1599,n1588);
nand (n1722,n1584,n1599);
nand (n1723,n1724,n1725,n1726);
nand (n1724,n1615,n1619);
nand (n1725,n1623,n1619);
nand (n1726,n1615,n1623);
xor (n1727,n1728,n1779);
xor (n1728,n1729,n1750);
xor (n1729,n1730,n1746);
xor (n1730,n1731,n1742);
xor (n1731,n1732,n1738);
xor (n1732,n1733,n1734);
not (n1733,n379);
xor (n1734,n1735,n84);
or (n1735,n1736,n1737);
and (n1736,n17,n78);
and (n1737,n131,n82);
xor (n1738,n1739,n20);
or (n1739,n1740,n1741);
and (n1740,n181,n13);
and (n1741,n185,n18);
nand (n1742,n1743,n1744,n1745);
nand (n1743,n1601,n1605);
nand (n1744,n1609,n1605);
nand (n1745,n1601,n1609);
nand (n1746,n1747,n1748,n1749);
nand (n1747,n1625,n1629);
nand (n1748,n21,n1629);
nand (n1749,n1625,n21);
xor (n1750,n1751,n1775);
xor (n1751,n1752,n1765);
xor (n1752,n1753,n1762);
xor (n1753,n1754,n1758);
xor (n1754,n1755,n110);
or (n1755,n1756,n1757);
and (n1756,n189,n104);
and (n1757,n325,n108);
xor (n1758,n1759,n21);
or (n1759,n1760,n1761);
and (n1760,n495,n186);
and (n1761,n499,n190);
nand (n1762,n1630,n1763,n1764);
nand (n1763,n1635,n1631);
not (n1764,n1635);
xor (n1765,n1766,n1771);
xor (n1766,n21,n1767);
nand (n1767,n1768,n1769,n1770);
nand (n1768,n1666,n1670);
nand (n1769,n1671,n1670);
nand (n1770,n1666,n1671);
nand (n1771,n1772,n1773,n1774);
nand (n1772,n1652,n1656);
nand (n1773,n1660,n1656);
nand (n1774,n1652,n1660);
nand (n1775,n1776,n1777,n1778);
nand (n1776,n1646,n1650);
nand (n1777,n1664,n1650);
nand (n1778,n1646,n1664);
nand (n1779,n1780,n1781,n1782);
nand (n1780,n1640,n1644);
nand (n1781,n1675,n1644);
nand (n1782,n1640,n1675);
nand (n1783,n1784,n1785,n1786);
nand (n1784,n1582,n1613);
nand (n1785,n1638,n1613);
nand (n1786,n1582,n1638);
nor (n1787,n1788,n1792);
nand (n1788,n1789,n1790,n1791);
nand (n1789,n1687,n1727);
nand (n1790,n1783,n1727);
nand (n1791,n1687,n1783);
xor (n1792,n1793,n1802);
xor (n1793,n1794,n1798);
nand (n1794,n1795,n1796,n1797);
nand (n1795,n1689,n1719);
nand (n1796,n1723,n1719);
nand (n1797,n1689,n1723);
nand (n1798,n1799,n1800,n1801);
nand (n1799,n1729,n1750);
nand (n1800,n1779,n1750);
nand (n1801,n1729,n1779);
xor (n1802,n1803,n1834);
xor (n1803,n1804,n1808);
nand (n1804,n1805,n1806,n1807);
nand (n1805,n1752,n1765);
nand (n1806,n1775,n1765);
nand (n1807,n1752,n1775);
xor (n1808,n1809,n1822);
xor (n1809,n1810,n1814);
nand (n1810,n1811,n1812,n1813);
nand (n1811,n21,n1767);
nand (n1812,n1771,n1767);
nand (n1813,n21,n1771);
xor (n1814,n1815,n1818);
xor (n1815,n1816,n21);
xor (n1816,n1817,n337);
xor (n1817,n329,n332);
nand (n1818,n1819,n1820,n1821);
nand (n1819,n1707,n338);
nand (n1820,n1711,n338);
nand (n1821,n1707,n1711);
xor (n1822,n1823,n1830);
xor (n1823,n1824,n1826);
xor (n1824,n1825,n365);
xor (n1825,n356,n360);
nand (n1826,n1827,n1828,n1829);
nand (n1827,n1693,n1697);
nand (n1828,n1701,n1697);
nand (n1829,n1693,n1701);
nand (n1830,n1831,n1832,n1833);
nand (n1831,n1754,n1758);
nand (n1832,n1762,n1758);
nand (n1833,n1754,n1762);
xor (n1834,n1835,n1844);
xor (n1835,n1836,n1840);
nand (n1836,n1837,n1838,n1839);
nand (n1837,n1691,n1705);
nand (n1838,n1715,n1705);
nand (n1839,n1691,n1715);
nand (n1840,n1841,n1842,n1843);
nand (n1841,n1731,n1742);
nand (n1842,n1746,n1742);
nand (n1843,n1731,n1746);
xor (n1844,n1845,n1852);
xor (n1845,n1846,n1850);
nand (n1846,n1847,n1848,n1849);
nand (n1847,n1733,n1734);
nand (n1848,n1738,n1734);
nand (n1849,n1733,n1738);
xor (n1850,n1851,n384);
xor (n1851,n375,n379);
xor (n1852,n1853,n1862);
xor (n1853,n1854,n1858);
xor (n1854,n1855,n20);
or (n1855,n1856,n1857);
and (n1856,n107,n13);
and (n1857,n181,n18);
xor (n1858,n1859,n110);
or (n1859,n1860,n1861);
and (n1860,n185,n104);
and (n1861,n189,n108);
xor (n1862,n1863,n21);
or (n1863,n1864,n1865);
and (n1864,n325,n186);
and (n1865,n495,n190);
nand (n1866,n1867,n1951);
nor (n1867,n1868,n1918);
nor (n1868,n1869,n1873);
nand (n1869,n1870,n1871,n1872);
nand (n1870,n1794,n1798);
nand (n1871,n1802,n1798);
nand (n1872,n1794,n1802);
xor (n1873,n1874,n1914);
xor (n1874,n1875,n1895);
xor (n1875,n1876,n1883);
xor (n1876,n1877,n1879);
xor (n1877,n1878,n373);
xor (n1878,n354,n370);
nand (n1879,n1880,n1881,n1882);
nand (n1880,n1846,n1850);
nand (n1881,n1852,n1850);
nand (n1882,n1846,n1852);
xor (n1883,n1884,n1891);
xor (n1884,n1885,n1889);
nand (n1885,n1886,n1887,n1888);
nand (n1886,n1854,n1858);
nand (n1887,n1862,n1858);
nand (n1888,n1854,n1862);
xor (n1889,n1890,n283);
xor (n1890,n277,n281);
nand (n1891,n1892,n1893,n1894);
nand (n1892,n1816,n21);
nand (n1893,n1818,n21);
nand (n1894,n1816,n1818);
xor (n1895,n1896,n1910);
xor (n1896,n1897,n1901);
nand (n1897,n1898,n1899,n1900);
nand (n1898,n1810,n1814);
nand (n1899,n1822,n1814);
nand (n1900,n1810,n1822);
xor (n1901,n1902,n1906);
xor (n1902,n1903,n1905);
xor (n1903,n1904,n299);
xor (n1904,n290,n294);
xor (n1905,n322,n327);
nand (n1906,n1907,n1908,n1909);
nand (n1907,n1824,n1826);
nand (n1908,n1830,n1826);
nand (n1909,n1824,n1830);
nand (n1910,n1911,n1912,n1913);
nand (n1911,n1836,n1840);
nand (n1912,n1844,n1840);
nand (n1913,n1836,n1844);
nand (n1914,n1915,n1916,n1917);
nand (n1915,n1804,n1808);
nand (n1916,n1834,n1808);
nand (n1917,n1804,n1834);
nor (n1918,n1919,n1923);
nand (n1919,n1920,n1921,n1922);
nand (n1920,n1875,n1895);
nand (n1921,n1914,n1895);
nand (n1922,n1875,n1914);
xor (n1923,n1924,n1947);
xor (n1924,n1925,n1935);
xor (n1925,n1926,n1933);
xor (n1926,n1927,n1929);
xor (n1927,n1928,n270);
xor (n1928,n255,n267);
nand (n1929,n1930,n1931,n1932);
nand (n1930,n1885,n1889);
nand (n1931,n1891,n1889);
nand (n1932,n1885,n1891);
xor (n1933,n1934,n305);
xor (n1934,n275,n288);
xor (n1935,n1936,n1943);
xor (n1936,n1937,n1939);
xor (n1937,n1938,n352);
xor (n1938,n319,n349);
nand (n1939,n1940,n1941,n1942);
nand (n1940,n1903,n1905);
nand (n1941,n1906,n1905);
nand (n1942,n1903,n1906);
nand (n1943,n1944,n1945,n1946);
nand (n1944,n1877,n1879);
nand (n1945,n1883,n1879);
nand (n1946,n1877,n1883);
nand (n1947,n1948,n1949,n1950);
nand (n1948,n1897,n1901);
nand (n1949,n1910,n1901);
nand (n1950,n1897,n1910);
nor (n1951,n1952,n1969);
nor (n1952,n1953,n1957);
nand (n1953,n1954,n1955,n1956);
nand (n1954,n1925,n1935);
nand (n1955,n1947,n1935);
nand (n1956,n1925,n1947);
xor (n1957,n1958,n1965);
xor (n1958,n1959,n1963);
nand (n1959,n1960,n1961,n1962);
nand (n1960,n1927,n1929);
nand (n1961,n1933,n1929);
nand (n1962,n1927,n1933);
xor (n1963,n1964,n392);
xor (n1964,n315,n317);
nand (n1965,n1966,n1967,n1968);
nand (n1966,n1937,n1939);
nand (n1967,n1943,n1939);
nand (n1968,n1937,n1943);
nor (n1969,n1970,n1974);
nand (n1970,n1971,n1972,n1973);
nand (n1971,n1959,n1963);
nand (n1972,n1965,n1963);
nand (n1973,n1959,n1965);
xor (n1974,n1975,n313);
xor (n1975,n5,n171);
not (n1976,n1977);
nor (n1977,n1978,n1993);
nor (n1978,n1866,n1979);
nor (n1979,n1980,n1987);
nor (n1980,n1981,n1986);
nor (n1981,n1982,n1984);
nor (n1982,n1983,n1565);
nand (n1983,n1454,n1458);
not (n1984,n1985);
nand (n1985,n1566,n1570);
not (n1986,n1679);
not (n1987,n1988);
nor (n1988,n1989,n1991);
nor (n1989,n1990,n1787);
nand (n1990,n1681,n1685);
not (n1991,n1992);
nand (n1992,n1788,n1792);
not (n1993,n1994);
nor (n1994,n1995,n2002);
nor (n1995,n1996,n2001);
nor (n1996,n1997,n1999);
nor (n1997,n1998,n1918);
nand (n1998,n1869,n1873);
not (n1999,n2000);
nand (n2000,n1919,n1923);
not (n2001,n1951);
not (n2002,n2003);
nor (n2003,n2004,n2006);
nor (n2004,n2005,n1969);
nand (n2005,n1953,n1957);
not (n2006,n2007);
nand (n2007,n1970,n1974);
nand (n2008,n2009,n2428);
nand (n2009,n2010,n2321);
nor (n2010,n2011,n2306);
nor (n2011,n2012,n2177);
nand (n2012,n2013,n2154);
nor (n2013,n2014,n2131);
nor (n2014,n2015,n2104);
nand (n2015,n2016,n2061,n2103);
nand (n2016,n2017,n2029);
xor (n2017,n2018,n2024);
xor (n2018,n2019,n2020);
xor (n2019,n1322,n1326);
xor (n2020,n2021,n30);
or (n2021,n2022,n2023);
and (n2022,n524,n53);
and (n2023,n538,n57);
and (n2024,n30,n2025);
xor (n2025,n2026,n218);
or (n2026,n2027,n2028);
and (n2027,n181,n341);
and (n2028,n185,n345);
nand (n2029,n2030,n2047,n2060);
nand (n2030,n2031,n2032);
xor (n2031,n30,n2025);
nand (n2032,n2033,n2042,n2046);
nand (n2033,n2034,n2038);
xor (n2034,n2035,n42);
or (n2035,n2036,n2037);
and (n2036,n499,n117);
and (n2037,n501,n121);
xor (n2038,n2039,n119);
or (n2039,n2040,n2041);
and (n2040,n325,n216);
and (n2041,n495,n220);
nand (n2042,n2043,n2038);
and (n2043,n47,n2044);
xnor (n2044,n2045,n47);
nand (n2045,n538,n40);
nand (n2046,n2034,n2043);
nand (n2047,n2048,n2032);
xor (n2048,n2049,n2056);
xor (n2049,n2050,n2054);
xnor (n2050,n2051,n343);
nor (n2051,n2052,n2053);
and (n2052,n107,n510);
and (n2053,n103,n512);
xnor (n2054,n2055,n30);
nand (n2055,n538,n53);
xor (n2056,n2057,n42);
or (n2057,n2058,n2059);
and (n2058,n495,n117);
and (n2059,n499,n121);
nand (n2060,n2031,n2048);
nand (n2061,n2062,n2029);
xor (n2062,n2063,n2082);
xor (n2063,n2064,n2068);
nand (n2064,n2065,n2066,n2067);
nand (n2065,n2050,n2054);
nand (n2066,n2056,n2054);
nand (n2067,n2050,n2056);
xor (n2068,n2069,n2078);
xor (n2069,n2070,n2074);
xor (n2070,n2071,n42);
or (n2071,n2072,n2073);
and (n2072,n325,n117);
and (n2073,n495,n121);
xor (n2074,n2075,n119);
or (n2075,n2076,n2077);
and (n2076,n185,n216);
and (n2077,n189,n220);
xor (n2078,n2079,n47);
or (n2079,n2080,n2081);
and (n2080,n499,n40);
and (n2081,n501,n45);
nand (n2082,n2083,n2097,n2102);
nand (n2083,n2084,n2088);
xor (n2084,n2085,n119);
or (n2085,n2086,n2087);
and (n2086,n189,n216);
and (n2087,n325,n220);
and (n2088,n2089,n2093);
xnor (n2089,n2090,n343);
nor (n2090,n2091,n2092);
and (n2091,n181,n510);
and (n2092,n107,n512);
xor (n2093,n2094,n218);
or (n2094,n2095,n2096);
and (n2095,n185,n341);
and (n2096,n189,n345);
nand (n2097,n2098,n2088);
xor (n2098,n2099,n47);
or (n2099,n2100,n2101);
and (n2100,n501,n40);
and (n2101,n524,n45);
nand (n2102,n2084,n2098);
nand (n2103,n2017,n2062);
xor (n2104,n2105,n2119);
xor (n2105,n2106,n2115);
xor (n2106,n2107,n2113);
xor (n2107,n2108,n2112);
xor (n2108,n2109,n30);
or (n2109,n2110,n2111);
and (n2110,n501,n53);
and (n2111,n524,n57);
xor (n2112,n1266,n35);
xor (n2113,n2114,n1309);
xor (n2114,n1302,n1306);
nand (n2115,n2116,n2117,n2118);
nand (n2116,n2064,n2068);
nand (n2117,n2082,n2068);
nand (n2118,n2064,n2082);
xor (n2119,n2120,n2129);
xor (n2120,n2121,n2125);
nand (n2121,n2122,n2123,n2124);
nand (n2122,n2019,n2020);
nand (n2123,n2024,n2020);
nand (n2124,n2019,n2024);
nand (n2125,n2126,n2127,n2128);
nand (n2126,n2070,n2074);
nand (n2127,n2078,n2074);
nand (n2128,n2070,n2078);
xor (n2129,n2130,n1331);
xor (n2130,n1317,n1321);
nor (n2131,n2132,n2136);
nand (n2132,n2133,n2134,n2135);
nand (n2133,n2106,n2115);
nand (n2134,n2119,n2115);
nand (n2135,n2106,n2119);
xor (n2136,n2137,n2144);
xor (n2137,n2138,n2140);
xor (n2138,n2139,n1315);
xor (n2139,n1296,n1300);
nand (n2140,n2141,n2142,n2143);
nand (n2141,n2121,n2125);
nand (n2142,n2129,n2125);
nand (n2143,n2121,n2129);
xor (n2144,n2145,n2150);
xor (n2145,n2146,n2148);
xor (n2146,n2147,n1265);
xor (n2147,n1256,n1260);
xor (n2148,n2149,n1280);
xor (n2149,n1274,n1278);
nand (n2150,n2151,n2152,n2153);
nand (n2151,n2108,n2112);
nand (n2152,n2113,n2112);
nand (n2153,n2108,n2113);
nor (n2154,n2155,n2170);
nor (n2155,n2156,n2160);
nand (n2156,n2157,n2158,n2159);
nand (n2157,n2138,n2140);
nand (n2158,n2144,n2140);
nand (n2159,n2138,n2144);
xor (n2160,n2161,n2168);
xor (n2161,n2162,n2164);
xor (n2162,n2163,n1272);
xor (n2163,n1252,n1254);
nand (n2164,n2165,n2166,n2167);
nand (n2165,n2146,n2148);
nand (n2166,n2150,n2148);
nand (n2167,n2146,n2150);
xor (n2168,n2169,n1294);
xor (n2169,n1289,n1291);
nor (n2170,n2171,n2175);
nand (n2171,n2172,n2173,n2174);
nand (n2172,n2162,n2164);
nand (n2173,n2168,n2164);
nand (n2174,n2162,n2168);
xor (n2175,n2176,n1287);
xor (n2176,n1162,n1213);
nor (n2177,n2178,n2300);
nor (n2178,n2179,n2276);
nor (n2179,n2180,n2273);
nor (n2180,n2181,n2249);
nand (n2181,n2182,n2221);
or (n2182,n2183,n2207,n2220);
and (n2183,n2184,n2193);
xor (n2184,n2185,n2189);
xnor (n2185,n2186,n343);
nor (n2186,n2187,n2188);
and (n2187,n189,n510);
and (n2188,n185,n512);
xnor (n2189,n2190,n218);
nor (n2190,n2191,n2192);
and (n2191,n495,n345);
and (n2192,n325,n341);
or (n2193,n2194,n2201,n2206);
and (n2194,n2195,n2197);
not (n2195,n2196);
nand (n2196,n538,n117);
xnor (n2197,n2198,n343);
nor (n2198,n2199,n2200);
and (n2199,n325,n510);
and (n2200,n189,n512);
and (n2201,n2197,n2202);
xnor (n2202,n2203,n218);
nor (n2203,n2204,n2205);
and (n2204,n499,n345);
and (n2205,n495,n341);
and (n2206,n2195,n2202);
and (n2207,n2193,n2208);
xor (n2208,n2209,n2216);
xor (n2209,n2210,n2212);
and (n2210,n42,n2211);
xnor (n2211,n2196,n42);
xnor (n2212,n2213,n119);
nor (n2213,n2214,n2215);
and (n2214,n501,n220);
and (n2215,n499,n216);
xnor (n2216,n2217,n42);
nor (n2217,n2218,n2219);
and (n2218,n538,n121);
and (n2219,n524,n117);
and (n2220,n2184,n2208);
xor (n2221,n2222,n2238);
xor (n2222,n2223,n2227);
or (n2223,n2224,n2225,n2226);
and (n2224,n2210,n2212);
and (n2225,n2212,n2216);
and (n2226,n2210,n2216);
xor (n2227,n2228,n2234);
xor (n2228,n2229,n2230);
and (n2229,n2185,n2189);
xnor (n2230,n2231,n119);
nor (n2231,n2232,n2233);
and (n2232,n499,n220);
and (n2233,n495,n216);
xnor (n2234,n2235,n42);
nor (n2235,n2236,n2237);
and (n2236,n524,n121);
and (n2237,n501,n117);
xor (n2238,n2239,n2245);
xor (n2239,n2240,n2241);
not (n2240,n2045);
xnor (n2241,n2242,n343);
nor (n2242,n2243,n2244);
and (n2243,n185,n510);
and (n2244,n181,n512);
xnor (n2245,n2246,n218);
nor (n2246,n2247,n2248);
and (n2247,n325,n345);
and (n2248,n189,n341);
nor (n2249,n2250,n2254);
or (n2250,n2251,n2252,n2253);
and (n2251,n2223,n2227);
and (n2252,n2227,n2238);
and (n2253,n2223,n2238);
xor (n2254,n2255,n2262);
xor (n2255,n2256,n2260);
or (n2256,n2257,n2258,n2259);
and (n2257,n2229,n2230);
and (n2258,n2230,n2234);
and (n2259,n2229,n2234);
xor (n2260,n2261,n2043);
xor (n2261,n2034,n2038);
xor (n2262,n2263,n2269);
xor (n2263,n2264,n2268);
xor (n2264,n2265,n47);
or (n2265,n2266,n2267);
and (n2266,n524,n40);
and (n2267,n538,n45);
xor (n2268,n2089,n2093);
or (n2269,n2270,n2271,n2272);
and (n2270,n2240,n2241);
and (n2271,n2241,n2245);
and (n2272,n2240,n2245);
not (n2273,n2274);
not (n2274,n2275);
and (n2275,n2250,n2254);
not (n2276,n2277);
nor (n2277,n2278,n2293);
nor (n2278,n2279,n2283);
nand (n2279,n2280,n2281,n2282);
nand (n2280,n2256,n2260);
nand (n2281,n2262,n2260);
nand (n2282,n2256,n2262);
xor (n2283,n2284,n2291);
xor (n2284,n2285,n2287);
xor (n2285,n2286,n2098);
xor (n2286,n2084,n2088);
nand (n2287,n2288,n2289,n2290);
nand (n2288,n2264,n2268);
nand (n2289,n2269,n2268);
nand (n2290,n2264,n2269);
xor (n2291,n2292,n2048);
xor (n2292,n2031,n2032);
nor (n2293,n2294,n2298);
nand (n2294,n2295,n2296,n2297);
nand (n2295,n2285,n2287);
nand (n2296,n2291,n2287);
nand (n2297,n2285,n2291);
xor (n2298,n2299,n2062);
xor (n2299,n2017,n2029);
not (n2300,n2301);
nor (n2301,n2302,n2304);
nor (n2302,n2303,n2293);
nand (n2303,n2279,n2283);
not (n2304,n2305);
nand (n2305,n2294,n2298);
not (n2306,n2307);
nor (n2307,n2308,n2315);
nor (n2308,n2309,n2314);
nor (n2309,n2310,n2312);
nor (n2310,n2311,n2131);
nand (n2311,n2015,n2104);
not (n2312,n2313);
nand (n2313,n2132,n2136);
not (n2314,n2154);
not (n2315,n2316);
nor (n2316,n2317,n2319);
nor (n2317,n2318,n2170);
nand (n2318,n2156,n2160);
not (n2319,n2320);
nand (n2320,n2171,n2175);
nand (n2321,n2322,n2326);
nor (n2322,n2323,n2012);
nand (n2323,n2324,n2277);
nor (n2324,n2325,n2249);
nor (n2325,n2182,n2221);
or (n2326,n2327,n2349);
and (n2327,n2328,n2330);
xor (n2328,n2329,n2208);
xor (n2329,n2184,n2193);
or (n2330,n2331,n2345,n2348);
and (n2331,n2332,n2341);
and (n2332,n2333,n2337);
xnor (n2333,n2334,n343);
nor (n2334,n2335,n2336);
and (n2335,n495,n510);
and (n2336,n325,n512);
xnor (n2337,n2338,n218);
nor (n2338,n2339,n2340);
and (n2339,n501,n345);
and (n2340,n499,n341);
xnor (n2341,n2342,n119);
nor (n2342,n2343,n2344);
and (n2343,n524,n220);
and (n2344,n501,n216);
and (n2345,n2341,n2346);
xor (n2346,n2347,n2202);
xor (n2347,n2195,n2197);
and (n2348,n2332,n2346);
and (n2349,n2350,n2351);
xor (n2350,n2328,n2330);
or (n2351,n2352,n2367);
and (n2352,n2353,n2365);
or (n2353,n2354,n2359,n2364);
and (n2354,n2355,n2356);
xor (n2355,n2333,n2337);
and (n2356,n119,n2357);
xnor (n2357,n2358,n119);
nand (n2358,n538,n216);
and (n2359,n2356,n2360);
xnor (n2360,n2361,n119);
nor (n2361,n2362,n2363);
and (n2362,n538,n220);
and (n2363,n524,n216);
and (n2364,n2355,n2360);
xor (n2365,n2366,n2346);
xor (n2366,n2332,n2341);
and (n2367,n2368,n2369);
xor (n2368,n2353,n2365);
or (n2369,n2370,n2386);
and (n2370,n2371,n2373);
xor (n2371,n2372,n2360);
xor (n2372,n2355,n2356);
or (n2373,n2374,n2380,n2385);
and (n2374,n2375,n2376);
not (n2375,n2358);
xnor (n2376,n2377,n343);
nor (n2377,n2378,n2379);
and (n2378,n499,n510);
and (n2379,n495,n512);
and (n2380,n2376,n2381);
xnor (n2381,n2382,n218);
nor (n2382,n2383,n2384);
and (n2383,n524,n345);
and (n2384,n501,n341);
and (n2385,n2375,n2381);
and (n2386,n2387,n2388);
xor (n2387,n2371,n2373);
or (n2388,n2389,n2400);
and (n2389,n2390,n2392);
xor (n2390,n2391,n2381);
xor (n2391,n2375,n2376);
and (n2392,n2393,n2396);
and (n2393,n218,n2394);
xnor (n2394,n2395,n218);
nand (n2395,n538,n341);
xnor (n2396,n2397,n343);
nor (n2397,n2398,n2399);
and (n2398,n501,n510);
and (n2399,n499,n512);
and (n2400,n2401,n2402);
xor (n2401,n2390,n2392);
or (n2402,n2403,n2409);
and (n2403,n2404,n2408);
xnor (n2404,n2405,n218);
nor (n2405,n2406,n2407);
and (n2406,n538,n345);
and (n2407,n524,n341);
xor (n2408,n2393,n2396);
and (n2409,n2410,n2411);
xor (n2410,n2404,n2408);
or (n2411,n2412,n2418);
and (n2412,n2413,n2417);
xnor (n2413,n2414,n343);
nor (n2414,n2415,n2416);
and (n2415,n524,n510);
and (n2416,n501,n512);
not (n2417,n2395);
and (n2418,n2419,n2420);
xor (n2419,n2413,n2417);
and (n2420,n2421,n2425);
xnor (n2421,n2422,n343);
nor (n2422,n2423,n2424);
and (n2423,n538,n510);
and (n2424,n524,n512);
and (n2425,n2426,n343);
xnor (n2426,n2427,n343);
nand (n2427,n538,n512);
not (n2428,n2429);
nand (n2429,n2430,n1450);
nor (n2430,n2431,n482);
nand (n2431,n2432,n1405);
nor (n2432,n2433,n1377);
nor (n2433,n1160,n1339);
not (n2434,n2435);
nor (n2435,n3,n396);
nand (n2436,n2437,n2515);
not (n2437,n2438);
nor (n2438,n2439,n2443);
nand (n2439,n2440,n2441,n2442);
nand (n2440,n398,n402);
nand (n2441,n472,n402);
nand (n2442,n398,n472);
xor (n2443,n2444,n2511);
xor (n2444,n2445,n2471);
xor (n2445,n2446,n2455);
xor (n2446,n2447,n2451);
nand (n2447,n2448,n2449,n2450);
nand (n2448,n416,n420);
nand (n2449,n424,n420);
nand (n2450,n416,n424);
nand (n2451,n2452,n2453,n2454);
nand (n2452,n21,n450);
nand (n2453,n464,n450);
nand (n2454,n21,n464);
xor (n2455,n2456,n2467);
xor (n2456,n21,n2457);
xor (n2457,n2458,n2463);
xor (n2458,n438,n2459);
xor (n2459,n2460,n30);
or (n2460,n2461,n2462);
and (n2461,n143,n53);
and (n2462,n39,n57);
xor (n2463,n2464,n35);
or (n2464,n2465,n2466);
and (n2465,n44,n28);
and (n2466,n52,n33);
nand (n2467,n2468,n2469,n2470);
nand (n2468,n452,n456);
nand (n2469,n460,n456);
nand (n2470,n452,n460);
xor (n2471,n2472,n2507);
xor (n2472,n2473,n2503);
xor (n2473,n2474,n2493);
xor (n2474,n2475,n2479);
nand (n2475,n2476,n2477,n2478);
nand (n2476,n430,n434);
nand (n2477,n438,n434);
nand (n2478,n430,n438);
xor (n2479,n2480,n2489);
xor (n2480,n2481,n2485);
xor (n2481,n2482,n84);
or (n2482,n2483,n2484);
and (n2483,n56,n78);
and (n2484,n27,n82);
xor (n2485,n2486,n15);
or (n2486,n2487,n2488);
and (n2487,n32,n95);
and (n2488,n68,n98);
xor (n2489,n2490,n21);
or (n2490,n2491,n2492);
and (n2491,n131,n186);
and (n2492,n103,n190);
xor (n2493,n2494,n2499);
xor (n2494,n439,n2495);
xor (n2495,n2496,n20);
or (n2496,n2497,n2498);
and (n2497,n77,n13);
and (n2498,n81,n18);
xor (n2499,n2500,n110);
or (n2500,n2501,n2502);
and (n2501,n12,n104);
and (n2502,n17,n108);
nand (n2503,n2504,n2505,n2506);
nand (n2504,n410,n414);
nand (n2505,n428,n414);
nand (n2506,n410,n428);
nand (n2507,n2508,n2509,n2510);
nand (n2508,n444,n448);
nand (n2509,n468,n448);
nand (n2510,n444,n468);
nand (n2511,n2512,n2513,n2514);
nand (n2512,n404,n408);
nand (n2513,n442,n408);
nand (n2514,n404,n442);
nand (n2515,n2439,n2443);
xor (n2516,n2517,n2712);
xor (n2517,n2518,n2630);
xor (n2518,n2519,n2582);
xor (n2519,n2520,n2556);
or (n2520,n2521,n2537,n2555);
and (n2521,n2522,n2525);
xor (n2522,n2523,n424);
xor (n2523,n464,n2524);
not (n2524,n411);
or (n2525,n2526,n2533,n2536);
and (n2526,n137,n2527);
or (n2527,n2528,n2530,n2532);
and (n2528,n228,n2529);
not (n2529,n194);
and (n2530,n2529,n2531);
not (n2531,n176);
and (n2532,n228,n2531);
and (n2533,n2527,n2534);
xor (n2534,n2535,n238);
xor (n2535,n9,n153);
and (n2536,n137,n2534);
and (n2537,n2525,n2538);
xor (n2538,n2539,n2552);
xor (n2539,n2540,n2544);
or (n2540,n2541,n2542,n2543);
and (n2541,n9,n153);
and (n2542,n153,n238);
and (n2543,n9,n238);
or (n2544,n2545,n2546,n2551);
and (n2545,n22,n167);
and (n2546,n167,n2547);
or (n2547,n2548,n2549,n2550);
and (n2548,n140,n200);
not (n2549,n236);
and (n2550,n140,n196);
and (n2551,n22,n2547);
xor (n2552,n2553,n415);
xor (n2553,n450,n2554);
not (n2554,n428);
and (n2555,n2522,n2538);
xor (n2556,n2557,n2570);
xor (n2557,n2558,n2562);
or (n2558,n2559,n2560,n2561);
and (n2559,n2540,n2544);
and (n2560,n2544,n2552);
and (n2561,n2540,n2552);
xor (n2562,n2563,n2565);
xor (n2563,n2564,n2457);
not (n2564,n2448);
xor (n2565,n2566,n2479);
or (n2566,n2567,n2568,n2569);
and (n2567,n439,n430);
not (n2568,n2476);
and (n2569,n439,n434);
xor (n2570,n2571,n2580);
xor (n2571,n2572,n2576);
or (n2572,n2573,n2574,n2575);
and (n2573,n450,n2554);
and (n2574,n2554,n415);
and (n2575,n450,n415);
or (n2576,n2577,n2578,n2579);
and (n2577,n464,n2524);
and (n2578,n2524,n424);
and (n2579,n464,n424);
xor (n2580,n2581,n2467);
xor (n2581,n2495,n2499);
or (n2582,n2583,n2594,n2629);
and (n2583,n2584,n2592);
or (n2584,n2585,n2588,n2591);
and (n2585,n2586,n60);
xor (n2586,n2587,n2547);
xor (n2587,n22,n167);
and (n2588,n60,n2589);
xor (n2589,n2590,n2534);
xor (n2590,n137,n2527);
and (n2591,n2586,n2589);
xor (n2592,n2593,n2538);
xor (n2593,n2522,n2525);
and (n2594,n2592,n2595);
or (n2595,n2596,n2625,n2628);
and (n2596,n2597,n2610);
or (n2597,n2598,n2608,n2609);
and (n2598,n2599,n273);
or (n2599,n2600,n2605,n2607);
and (n2600,n2601,n267);
or (n2601,n2602,n2603,n2604);
and (n2602,n212,n257);
not (n2603,n261);
and (n2604,n212,n262);
and (n2605,n267,n2606);
not (n2606,n270);
and (n2607,n2601,n2606);
not (n2608,n308);
and (n2609,n2599,n309);
or (n2610,n2611,n2618,n2624);
and (n2611,n2612,n2616);
or (n2612,n2613,n2614,n2615);
and (n2613,n213,n209);
not (n2614,n227);
and (n2615,n213,n223);
xor (n2616,n2617,n2531);
xor (n2617,n228,n2529);
and (n2618,n2616,n2619);
or (n2619,n2620,n2621,n2623);
and (n2620,n212,n350);
and (n2621,n350,n2622);
not (n2622,n1930);
and (n2623,n212,n2622);
and (n2624,n2612,n2619);
and (n2625,n2610,n2626);
xor (n2626,n2627,n2589);
xor (n2627,n2586,n60);
and (n2628,n2597,n2626);
and (n2629,n2584,n2595);
or (n2630,n2631,n2633);
xor (n2631,n2632,n2595);
xor (n2632,n2584,n2592);
or (n2633,n2634,n2656,n2711);
and (n2634,n2635,n2654);
or (n2635,n2636,n2650,n2653);
and (n2636,n2637,n2639);
xor (n2637,n2638,n309);
xor (n2638,n2599,n273);
or (n2639,n2640,n2643,n2649);
and (n2640,n2641,n1933);
xor (n2641,n2642,n2606);
xor (n2642,n2601,n267);
and (n2643,n1933,n2644);
or (n2644,n2645,n2646,n2648);
not (n2645,n389);
and (n2646,n373,n2647);
not (n2647,n370);
and (n2648,n354,n2647);
and (n2649,n2641,n2644);
and (n2650,n2639,n2651);
xor (n2651,n2652,n2619);
xor (n2652,n2612,n2616);
and (n2653,n2637,n2651);
xor (n2654,n2655,n2626);
xor (n2655,n2597,n2610);
and (n2656,n2654,n2657);
or (n2657,n2658,n2673,n2710);
and (n2658,n2659,n2671);
or (n2659,n2660,n2667,n2670);
and (n2660,n2661,n2665);
or (n2661,n2662,n2663,n2664);
and (n2662,n321,n1903);
and (n2663,n1903,n1884);
and (n2664,n321,n1884);
xor (n2665,n2666,n2622);
xor (n2666,n212,n350);
and (n2667,n2665,n2668);
and (n2668,n1879,n2669);
not (n2669,n1877);
and (n2670,n2661,n2668);
xor (n2671,n2672,n2651);
xor (n2672,n2637,n2639);
and (n2673,n2671,n2674);
or (n2674,n2675,n2695,n2709);
and (n2675,n2676,n2693);
or (n2676,n2677,n2682,n2692);
and (n2677,n2678,n1906);
or (n2678,n2679,n2680,n2681);
and (n2679,n338,n329);
not (n2680,n328);
and (n2681,n338,n332);
and (n2682,n1906,n2683);
or (n2683,n2684,n2689,n2691);
and (n2684,n337,n2685);
or (n2685,n2686,n2687,n2688);
and (n2686,n337,n1707);
not (n2687,n1821);
and (n2688,n337,n1711);
and (n2689,n2685,n2690);
not (n2690,n1816);
and (n2691,n337,n2690);
and (n2692,n2678,n2683);
xor (n2693,n2694,n2644);
xor (n2694,n2641,n1933);
and (n2695,n2693,n2696);
or (n2696,n2697,n2701,n2708);
and (n2697,n2698,n2700);
xor (n2698,n2699,n1884);
xor (n2699,n321,n1903);
not (n2700,n1876);
and (n2701,n2700,n2702);
or (n2702,n2703,n2706,n2707);
and (n2703,n2704,n1822);
and (n2704,n1691,n2705);
not (n2705,n1705);
and (n2706,n1822,n1844);
and (n2707,n2704,n1844);
and (n2708,n2698,n2702);
and (n2709,n2676,n2696);
and (n2710,n2659,n2674);
and (n2711,n2635,n2657);
and (n2712,n2713,n2714);
xnor (n2713,n2631,n2633);
or (n2714,n2715,n2919);
and (n2715,n2716,n2718);
xor (n2716,n2717,n2657);
xor (n2717,n2635,n2654);
or (n2718,n2719,n2794,n2918);
and (n2719,n2720,n2792);
or (n2720,n2721,n2788,n2791);
and (n2721,n2722,n2724);
xor (n2722,n2723,n2668);
xor (n2723,n2661,n2665);
or (n2724,n2725,n2759,n2787);
and (n2725,n2726,n2757);
or (n2726,n2727,n2745,n2756);
and (n2727,n2728,n2737);
and (n2728,n2729,n1731);
or (n2729,n2730,n2735,n2736);
and (n2730,n2731,n1601);
or (n2731,n2732,n2733,n2734);
and (n2732,n1670,n1466);
not (n2733,n1610);
and (n2734,n1670,n1470);
not (n2735,n1743);
and (n2736,n2731,n1605);
or (n2737,n2738,n2743,n2744);
and (n2738,n1771,n2739);
or (n2739,n2740,n2741,n2742);
and (n2740,n1670,n1590);
not (n2741,n1718);
and (n2742,n1670,n1595);
and (n2743,n2739,n1752);
and (n2744,n1771,n1752);
and (n2745,n2737,n2746);
or (n2746,n2747,n2753,n2755);
and (n2747,n2748,n2749);
not (n2748,n1690);
or (n2749,n2750,n2751,n2752);
and (n2750,n1474,n1666);
not (n2751,n1770);
and (n2752,n1474,n1671);
and (n2753,n2749,n2754);
not (n2754,n1747);
and (n2755,n2748,n2754);
and (n2756,n2728,n2746);
xor (n2757,n2758,n2683);
xor (n2758,n2678,n1906);
and (n2759,n2757,n2760);
or (n2760,n2761,n2783,n2786);
and (n2761,n2762,n2764);
xor (n2762,n2763,n2690);
xor (n2763,n337,n2685);
or (n2764,n2765,n2774,n2782);
and (n2765,n2766,n2773);
or (n2766,n2767,n2769,n2772);
and (n2767,n1650,n2768);
not (n2768,n1647);
and (n2769,n2768,n2770);
xor (n2770,n2771,n1595);
xor (n2771,n1670,n1590);
and (n2772,n1650,n2770);
xor (n2773,n2729,n1731);
and (n2774,n2773,n2775);
or (n2775,n2776,n2780,n2781);
and (n2776,n2777,n2778);
not (n2777,n1664);
xor (n2778,n2779,n1605);
xor (n2779,n2731,n1601);
and (n2780,n2778,n1624);
and (n2781,n2777,n1624);
and (n2782,n2766,n2775);
and (n2783,n2764,n2784);
xor (n2784,n2785,n1844);
xor (n2785,n2704,n1822);
and (n2786,n2762,n2784);
and (n2787,n2726,n2760);
and (n2788,n2724,n2789);
xor (n2789,n2790,n2696);
xor (n2790,n2676,n2693);
and (n2791,n2722,n2789);
xor (n2792,n2793,n2674);
xor (n2793,n2659,n2671);
and (n2794,n2792,n2795);
or (n2795,n2796,n2829,n2917);
and (n2796,n2797,n2827);
or (n2797,n2798,n2823,n2826);
and (n2798,n2799,n2801);
xor (n2799,n2800,n2702);
xor (n2800,n2698,n2700);
or (n2801,n2802,n2819,n2822);
and (n2802,n2803,n2805);
xor (n2803,n2804,n2746);
xor (n2804,n2728,n2737);
or (n2805,n2806,n2811,n2818);
and (n2806,n2807,n2809);
xor (n2807,n2808,n1752);
xor (n2808,n1771,n2739);
xor (n2809,n2810,n2754);
xor (n2810,n2748,n2749);
and (n2811,n2809,n2812);
and (n2812,n1615,n2813);
or (n2813,n2814,n2815,n2817);
not (n2814,n1621);
and (n2815,n1481,n2816);
not (n2816,n1464);
and (n2817,n1477,n2816);
and (n2818,n2807,n2812);
and (n2819,n2805,n2820);
xor (n2820,n2821,n2784);
xor (n2821,n2762,n2764);
and (n2822,n2803,n2820);
and (n2823,n2801,n2824);
xor (n2824,n2825,n2760);
xor (n2825,n2726,n2757);
and (n2826,n2799,n2824);
xor (n2827,n2828,n2789);
xor (n2828,n2722,n2724);
and (n2829,n2827,n2830);
or (n2830,n2831,n2888,n2916);
and (n2831,n2832,n2834);
xor (n2832,n2833,n2824);
xor (n2833,n2799,n2801);
or (n2834,n2835,n2867,n2887);
and (n2835,n2836,n2865);
or (n2836,n2837,n2850,n2864);
and (n2837,n2838,n2848);
or (n2838,n2839,n2846,n2847);
and (n2839,n2840,n2844);
or (n2840,n2841,n2842,n2843);
and (n2841,n1529,n1514);
and (n2842,n1514,n1497);
and (n2843,n1529,n1497);
xor (n2844,n2845,n2770);
xor (n2845,n1650,n2768);
and (n2846,n2844,n1675);
and (n2847,n2840,n1675);
xor (n2848,n2849,n2775);
xor (n2849,n2766,n2773);
and (n2850,n2848,n2851);
or (n2851,n2852,n2861,n2863);
and (n2852,n2853,n2859);
or (n2853,n2854,n2855,n2858);
and (n2854,n1519,n1513);
and (n2855,n1513,n2856);
xor (n2856,n2857,n1497);
xor (n2857,n1529,n1514);
and (n2858,n1519,n2856);
xor (n2859,n2860,n1624);
xor (n2860,n2777,n2778);
and (n2861,n2859,n2862);
xor (n2862,n1615,n2813);
and (n2863,n2853,n2862);
and (n2864,n2838,n2851);
xor (n2865,n2866,n2820);
xor (n2866,n2803,n2805);
and (n2867,n2865,n2868);
or (n2868,n2869,n2883,n2886);
and (n2869,n2870,n2872);
xor (n2870,n2871,n2812);
xor (n2871,n2807,n2809);
or (n2872,n2873,n2881,n2882);
and (n2873,n2874,n2876);
xor (n2874,n2875,n1675);
xor (n2875,n2840,n2844);
or (n2876,n2877,n2878,n2880);
not (n2877,n1574);
and (n2878,n1489,n2879);
not (n2879,n1462);
and (n2880,n1485,n2879);
and (n2881,n2876,n1576);
and (n2882,n2874,n1576);
and (n2883,n2872,n2884);
xor (n2884,n2885,n2851);
xor (n2885,n2838,n2848);
and (n2886,n2870,n2884);
and (n2887,n2836,n2868);
and (n2888,n2834,n2889);
or (n2889,n2890,n2892);
xor (n2890,n2891,n2868);
xor (n2891,n2836,n2865);
or (n2892,n2893,n2909,n2915);
and (n2893,n2894,n2907);
or (n2894,n2895,n2903,n2906);
and (n2895,n2896,n2898);
xor (n2896,n2897,n2862);
xor (n2897,n2853,n2859);
or (n2898,n2899,n2901,n2902);
and (n2899,n2900,n1561);
not (n2900,n1460);
not (n2901,n1568);
and (n2902,n2900,n1493);
and (n2903,n2898,n2904);
xor (n2904,n2905,n1576);
xor (n2905,n2874,n2876);
and (n2906,n2896,n2904);
xor (n2907,n2908,n2884);
xor (n2908,n2870,n2872);
and (n2909,n2907,n2910);
or (n2910,n2911,n2913);
or (n2911,n1454,n2912);
not (n2912,n1458);
xor (n2913,n2914,n2904);
xor (n2914,n2896,n2898);
and (n2915,n2894,n2910);
and (n2916,n2832,n2889);
and (n2917,n2797,n2830);
and (n2918,n2720,n2795);
and (n2919,n2920,n2921);
xor (n2920,n2716,n2718);
and (n2921,n2922,n2924);
xor (n2922,n2923,n2795);
xor (n2923,n2720,n2792);
or (n2924,n2925,n2927);
xor (n2925,n2926,n2830);
xor (n2926,n2797,n2827);
and (n2927,n2928,n2929);
not (n2928,n2925);
and (n2929,n2930,n2932);
xor (n2930,n2931,n2889);
xor (n2931,n2832,n2834);
and (n2932,n2933,n2934);
xnor (n2933,n2890,n2892);
and (n2934,n2935,n2937);
xor (n2935,n2936,n2910);
xor (n2936,n2894,n2907);
and (n2937,n2938,n2939);
xnor (n2938,n2911,n2913);
and (n2939,n2940,n2943);
not (n2940,n2941);
nand (n2941,n2942,n1983);
not (n2942,n1453);
nand (n2943,n480,n2944);
nand (n2944,n2430,n2009);
endmodule
