module top (out,n3,n6,n7,n25,n27,n34,n35,n46,n57
        ,n58,n64,n70,n75,n83,n84,n91,n101,n108,n114
        ,n118,n137,n145,n157,n162,n187,n236,n287,n289,n325
        ,n384,n416,n417,n447,n575,n608,n668,n745);
output out;
input n3;
input n6;
input n7;
input n25;
input n27;
input n34;
input n35;
input n46;
input n57;
input n58;
input n64;
input n70;
input n75;
input n83;
input n84;
input n91;
input n101;
input n108;
input n114;
input n118;
input n137;
input n145;
input n157;
input n162;
input n187;
input n236;
input n287;
input n289;
input n325;
input n384;
input n416;
input n417;
input n447;
input n575;
input n608;
input n668;
input n745;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n288;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
xor (out,n0,n1736);
nand (n0,n1,n8);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nor (n5,n6,n7);
nand (n8,n9,n1733);
nand (n9,n10,n1732);
or (n10,n11,n393);
nand (n11,n12,n392);
not (n12,n13);
nor (n13,n14,n248);
xor (n14,n15,n226);
xor (n15,n16,n167);
or (n16,n17,n166);
and (n17,n18,n123);
xor (n18,n19,n48);
nand (n19,n20,n41);
or (n20,n21,n29);
not (n21,n22);
nor (n22,n23,n28);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
and (n28,n25,n27);
not (n29,n30);
nor (n30,n31,n37);
nand (n31,n32,n36);
or (n32,n33,n35);
not (n33,n34);
nand (n36,n33,n35);
nor (n37,n38,n39);
and (n38,n26,n35);
and (n39,n27,n40);
not (n40,n35);
nand (n41,n42,n31);
not (n42,n43);
nor (n43,n44,n47);
and (n44,n45,n27);
not (n45,n46);
and (n47,n46,n26);
or (n48,n49,n122);
and (n49,n50,n103);
xor (n50,n51,n78);
nand (n51,n52,n72);
or (n52,n53,n66);
nand (n53,n54,n61);
nor (n54,n55,n59);
and (n55,n56,n58);
not (n56,n57);
and (n59,n57,n60);
not (n60,n58);
nor (n61,n62,n65);
and (n62,n56,n63);
not (n63,n64);
and (n65,n57,n64);
not (n66,n67);
nor (n67,n68,n71);
and (n68,n63,n69);
not (n69,n70);
and (n71,n70,n64);
or (n72,n73,n54);
nor (n73,n74,n76);
and (n74,n75,n63);
and (n76,n64,n77);
not (n77,n75);
nand (n78,n79,n93);
or (n79,n80,n88);
not (n80,n81);
nor (n81,n82,n85);
and (n82,n83,n84);
and (n85,n86,n87);
not (n86,n83);
not (n87,n84);
not (n88,n89);
nand (n89,n90,n92);
or (n90,n63,n91);
nand (n92,n91,n63);
or (n93,n94,n98);
nand (n94,n88,n95);
nand (n95,n96,n97);
or (n96,n91,n87);
nand (n97,n87,n91);
nor (n98,n99,n102);
and (n99,n100,n84);
not (n100,n101);
and (n102,n101,n87);
nand (n103,n104,n121);
or (n104,n105,n116);
nand (n105,n106,n110);
nand (n106,n107,n109);
or (n107,n108,n33);
nand (n109,n33,n108);
not (n110,n111);
nand (n111,n112,n115);
or (n112,n113,n108);
not (n113,n114);
nand (n115,n108,n113);
nor (n116,n117,n119);
and (n117,n33,n118);
and (n119,n34,n120);
not (n120,n118);
or (n121,n110,n33);
and (n122,n51,n78);
xor (n123,n124,n154);
xor (n124,n125,n131);
nand (n125,n126,n127);
or (n126,n80,n94);
nand (n127,n89,n128);
nor (n128,n129,n130);
and (n129,n69,n87);
and (n130,n70,n84);
nand (n131,n132,n150);
or (n132,n133,n139);
not (n133,n134);
nor (n134,n135,n138);
and (n135,n136,n60);
not (n136,n137);
and (n138,n137,n58);
not (n139,n140);
and (n140,n141,n147);
not (n141,n142);
nand (n142,n143,n146);
or (n143,n144,n27);
not (n144,n145);
nand (n146,n27,n144);
nand (n147,n148,n149);
nand (n148,n58,n144);
nand (n149,n145,n60);
nand (n150,n142,n151);
nor (n151,n152,n153);
and (n152,n24,n60);
and (n153,n25,n58);
nand (n154,n155,n165);
or (n155,n156,n158);
not (n156,n157);
not (n158,n159);
nor (n159,n160,n164);
nand (n160,n161,n163);
or (n161,n87,n162);
nand (n163,n162,n87);
not (n164,n162);
nand (n165,n160,n101);
and (n166,n19,n48);
xor (n167,n168,n206);
xor (n168,n169,n191);
or (n169,n170,n190);
and (n170,n171,n182);
xor (n171,n172,n175);
nand (n172,n173,n34);
or (n173,n111,n174);
not (n174,n105);
nand (n175,n176,n177);
or (n176,n29,n43);
or (n177,n178,n179);
not (n178,n31);
nor (n179,n180,n181);
and (n180,n26,n118);
and (n181,n27,n120);
nand (n182,n183,n184);
or (n183,n53,n73);
or (n184,n54,n185);
nor (n185,n186,n188);
and (n186,n63,n187);
and (n188,n64,n189);
not (n189,n187);
and (n190,n172,n175);
xor (n191,n192,n203);
xor (n192,n193,n200);
nand (n193,n194,n196);
or (n194,n94,n195);
not (n195,n128);
or (n196,n88,n197);
nor (n197,n198,n199);
and (n198,n87,n75);
and (n199,n84,n77);
nand (n200,n201,n202);
or (n201,n100,n158);
nand (n202,n160,n83);
nand (n203,n204,n205);
or (n204,n29,n179);
or (n205,n178,n26);
xor (n206,n207,n223);
xor (n207,n208,n214);
nand (n208,n209,n210);
or (n209,n53,n185);
or (n210,n54,n211);
nor (n211,n212,n213);
and (n212,n63,n137);
and (n213,n64,n136);
not (n214,n215);
nand (n215,n216,n218);
or (n216,n217,n139);
not (n217,n151);
nand (n218,n219,n142);
not (n219,n220);
nor (n220,n221,n222);
and (n221,n45,n58);
and (n222,n46,n60);
or (n223,n224,n225);
and (n224,n124,n154);
and (n225,n125,n131);
or (n226,n227,n247);
and (n227,n228,n246);
xor (n228,n229,n230);
xor (n229,n171,n182);
or (n230,n231,n245);
and (n231,n232,n244);
xor (n232,n233,n238);
nand (n233,n234,n237);
or (n234,n235,n158);
not (n235,n236);
nand (n237,n160,n157);
nand (n238,n239,n243);
or (n239,n139,n240);
nor (n240,n241,n242);
and (n241,n60,n187);
and (n242,n58,n189);
or (n243,n141,n133);
not (n244,n19);
and (n245,n233,n238);
xor (n246,n18,n123);
and (n247,n229,n230);
or (n248,n249,n391);
and (n249,n250,n315);
xor (n250,n251,n314);
or (n251,n252,n313);
and (n252,n253,n312);
xor (n253,n254,n280);
or (n254,n255,n279);
and (n255,n256,n272);
xor (n256,n257,n265);
nand (n257,n258,n263);
or (n258,n259,n53);
not (n259,n260);
nand (n260,n261,n262);
or (n261,n86,n64);
or (n262,n83,n63);
nand (n263,n264,n67);
not (n264,n54);
nand (n265,n266,n271);
or (n266,n267,n29);
not (n267,n268);
nand (n268,n269,n270);
or (n269,n137,n26);
nand (n270,n26,n137);
nand (n271,n31,n22);
nand (n272,n273,n278);
or (n273,n94,n274);
not (n274,n275);
nor (n275,n276,n277);
and (n276,n156,n87);
and (n277,n157,n84);
or (n278,n88,n98);
and (n279,n257,n265);
or (n280,n281,n311);
and (n281,n282,n304);
xor (n282,n283,n296);
nand (n283,n284,n114);
or (n284,n285,n291);
nand (n285,n286,n290);
or (n286,n287,n288);
not (n288,n289);
nand (n290,n287,n288);
nor (n291,n285,n292);
nor (n292,n293,n295);
and (n293,n294,n114);
not (n294,n287);
and (n295,n287,n113);
nand (n296,n297,n302);
or (n297,n298,n105);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n45,n33);
and (n301,n46,n34);
nand (n302,n303,n111);
not (n303,n116);
nand (n304,n305,n310);
or (n305,n139,n306);
not (n306,n307);
nor (n307,n308,n309);
and (n308,n77,n60);
and (n309,n75,n58);
or (n310,n141,n240);
and (n311,n283,n296);
xor (n312,n50,n103);
and (n313,n254,n280);
xor (n314,n228,n246);
or (n315,n316,n390);
and (n316,n317,n361);
xor (n317,n318,n319);
xor (n318,n232,n244);
or (n319,n320,n360);
and (n320,n321,n335);
xor (n321,n322,n328);
nand (n322,n323,n326);
or (n323,n324,n158);
not (n324,n325);
or (n326,n327,n235);
not (n327,n160);
not (n328,n329);
nor (n329,n330,n334);
and (n330,n291,n331);
nor (n331,n332,n333);
and (n332,n120,n113);
and (n333,n118,n114);
and (n334,n285,n114);
or (n335,n336,n359);
and (n336,n337,n352);
xor (n337,n338,n345);
nand (n338,n339,n344);
or (n339,n340,n105);
not (n340,n341);
nor (n341,n342,n343);
and (n342,n24,n33);
and (n343,n25,n34);
nand (n344,n111,n299);
nand (n345,n346,n351);
or (n346,n347,n139);
not (n347,n348);
nor (n348,n349,n350);
and (n349,n69,n60);
and (n350,n70,n58);
nand (n351,n142,n307);
nand (n352,n353,n354);
or (n353,n259,n54);
nand (n354,n355,n356);
not (n355,n53);
nor (n356,n357,n358);
and (n357,n100,n63);
and (n358,n101,n64);
and (n359,n338,n345);
and (n360,n322,n328);
or (n361,n362,n389);
and (n362,n363,n388);
xor (n363,n364,n387);
or (n364,n365,n386);
and (n365,n366,n381);
xor (n366,n367,n374);
nand (n367,n368,n373);
or (n368,n369,n29);
not (n369,n370);
nor (n370,n371,n372);
and (n371,n189,n26);
and (n372,n187,n27);
nand (n373,n31,n268);
nand (n374,n375,n380);
or (n375,n376,n94);
not (n376,n377);
nor (n377,n378,n379);
and (n378,n235,n87);
and (n379,n236,n84);
nand (n380,n89,n275);
nand (n381,n382,n385);
or (n382,n383,n158);
not (n383,n384);
nand (n385,n160,n325);
and (n386,n367,n374);
xor (n387,n256,n272);
xor (n388,n282,n304);
and (n389,n364,n387);
and (n390,n318,n319);
and (n391,n251,n314);
nand (n392,n14,n248);
nand (n393,n394,n1731);
or (n394,n395,n499);
nor (n395,n396,n498);
or (n396,n397,n497);
and (n397,n398,n401);
xor (n398,n399,n400);
xor (n399,n253,n312);
xor (n400,n317,n361);
or (n401,n402,n496);
and (n402,n403,n465);
xor (n403,n404,n405);
xor (n404,n321,n335);
or (n405,n406,n464);
and (n406,n407,n441);
xor (n407,n329,n408);
or (n408,n409,n440);
and (n409,n410,n433);
xor (n410,n411,n425);
nand (n411,n412,n289);
or (n412,n413,n419);
nand (n413,n414,n418);
or (n414,n415,n417);
not (n415,n416);
nand (n418,n417,n415);
not (n419,n420);
nand (n420,n421,n422);
not (n421,n413);
nand (n422,n423,n424);
or (n423,n415,n289);
nand (n424,n415,n289);
nand (n425,n426,n432);
or (n426,n427,n431);
not (n427,n428);
nand (n428,n429,n430);
or (n429,n46,n113);
nand (n430,n113,n46);
not (n431,n291);
nand (n432,n331,n285);
nand (n433,n434,n439);
or (n434,n435,n29);
not (n435,n436);
nor (n436,n437,n438);
and (n437,n77,n26);
and (n438,n75,n27);
nand (n439,n31,n370);
and (n440,n411,n425);
or (n441,n442,n463);
and (n442,n443,n456);
xor (n443,n444,n449);
nand (n444,n445,n448);
or (n445,n446,n158);
not (n446,n447);
nand (n448,n160,n384);
nand (n449,n450,n455);
or (n450,n451,n139);
not (n451,n452);
nor (n452,n453,n454);
and (n453,n86,n60);
and (n454,n83,n58);
nand (n455,n142,n348);
nand (n456,n457,n458);
or (n457,n340,n110);
or (n458,n105,n459);
not (n459,n460);
nor (n460,n461,n462);
and (n461,n136,n33);
and (n462,n137,n34);
and (n463,n444,n449);
and (n464,n329,n408);
or (n465,n466,n495);
and (n466,n467,n470);
xor (n467,n468,n469);
xor (n468,n366,n381);
xor (n469,n337,n352);
or (n470,n471,n494);
and (n471,n472,n487);
xor (n472,n473,n480);
nand (n473,n474,n479);
or (n474,n475,n53);
not (n475,n476);
nor (n476,n477,n478);
and (n477,n63,n156);
and (n478,n157,n64);
nand (n479,n264,n356);
nand (n480,n481,n486);
or (n481,n482,n94);
not (n482,n483);
nor (n483,n484,n485);
and (n484,n324,n87);
and (n485,n325,n84);
nand (n486,n89,n377);
not (n487,n488);
nor (n488,n489,n493);
and (n489,n419,n490);
nor (n490,n491,n492);
and (n491,n120,n288);
and (n492,n118,n289);
nor (n493,n421,n288);
and (n494,n473,n480);
and (n495,n468,n469);
and (n496,n404,n405);
and (n497,n399,n400);
xor (n498,n250,n315);
not (n499,n500);
nand (n500,n501,n1213);
nor (n501,n502,n1199);
and (n502,n503,n866);
and (n503,n504,n849);
nor (n504,n505,n757);
nor (n505,n506,n679);
xor (n506,n507,n588);
xor (n507,n508,n535);
or (n508,n509,n534);
and (n509,n510,n513);
xor (n510,n511,n512);
xor (n511,n443,n456);
xor (n512,n472,n487);
or (n513,n514,n533);
and (n514,n515,n523);
xor (n515,n516,n488);
nand (n516,n517,n522);
or (n517,n518,n94);
not (n518,n519);
nor (n519,n520,n521);
and (n520,n383,n87);
and (n521,n384,n84);
nand (n522,n89,n483);
nand (n523,n524,n417);
nor (n524,n525,n529);
and (n525,n174,n526);
nand (n526,n527,n528);
or (n527,n75,n33);
nand (n528,n33,n75);
and (n529,n111,n530);
nor (n530,n531,n532);
and (n531,n189,n33);
and (n532,n187,n34);
and (n533,n516,n488);
and (n534,n511,n512);
xor (n535,n536,n587);
xor (n536,n537,n538);
xor (n537,n407,n441);
or (n538,n539,n586);
and (n539,n540,n585);
xor (n540,n541,n562);
or (n541,n542,n561);
and (n542,n543,n555);
xor (n543,n544,n551);
nand (n544,n545,n550);
or (n545,n546,n139);
not (n546,n547);
nand (n547,n548,n549);
or (n548,n101,n60);
nand (n549,n60,n101);
nand (n550,n452,n142);
nand (n551,n552,n554);
or (n552,n553,n105);
not (n553,n530);
nand (n554,n111,n460);
nand (n555,n556,n557);
or (n556,n54,n475);
or (n557,n53,n558);
nor (n558,n559,n560);
and (n559,n236,n63);
and (n560,n64,n235);
and (n561,n544,n551);
or (n562,n563,n584);
and (n563,n564,n577);
xor (n564,n565,n572);
nand (n565,n566,n571);
or (n566,n567,n431);
not (n567,n568);
nor (n568,n569,n570);
and (n569,n24,n113);
and (n570,n25,n114);
nand (n571,n285,n428);
nand (n572,n573,n576);
or (n573,n574,n158);
not (n574,n575);
nand (n576,n160,n447);
nand (n577,n578,n583);
or (n578,n579,n29);
not (n579,n580);
nor (n580,n581,n582);
and (n581,n69,n26);
and (n582,n70,n27);
nand (n583,n31,n436);
and (n584,n565,n572);
xor (n585,n410,n433);
and (n586,n541,n562);
xor (n587,n467,n470);
or (n588,n589,n678);
and (n589,n590,n642);
xor (n590,n591,n592);
xor (n591,n540,n585);
or (n592,n593,n641);
and (n593,n594,n640);
xor (n594,n595,n617);
or (n595,n596,n616);
and (n596,n597,n610);
xor (n597,n598,n605);
nand (n598,n599,n604);
or (n599,n600,n94);
not (n600,n601);
nand (n601,n602,n603);
or (n602,n446,n84);
nand (n603,n84,n446);
nand (n604,n519,n89);
nand (n605,n606,n609);
or (n606,n607,n158);
not (n607,n608);
nand (n609,n160,n575);
nand (n610,n611,n613);
or (n611,n612,n421);
not (n612,n490);
or (n613,n420,n614);
not (n614,n615);
xor (n615,n45,n288);
and (n616,n598,n605);
or (n617,n618,n639);
and (n618,n619,n633);
xor (n619,n620,n627);
nand (n620,n621,n626);
or (n621,n622,n29);
not (n622,n623);
nor (n623,n624,n625);
and (n624,n86,n26);
and (n625,n83,n27);
nand (n626,n31,n580);
nand (n627,n628,n632);
or (n628,n629,n431);
nor (n629,n630,n631);
and (n630,n136,n114);
and (n631,n137,n113);
nand (n632,n568,n285);
nand (n633,n634,n638);
or (n634,n139,n635);
nor (n635,n636,n637);
and (n636,n156,n58);
and (n637,n157,n60);
or (n638,n141,n546);
and (n639,n620,n627);
xor (n640,n543,n555);
and (n641,n595,n617);
or (n642,n643,n677);
and (n643,n644,n647);
xor (n644,n645,n646);
xor (n645,n564,n577);
xor (n646,n515,n523);
and (n647,n648,n671);
or (n648,n649,n670);
and (n649,n650,n665);
xor (n650,n651,n658);
nand (n651,n652,n657);
or (n652,n653,n105);
not (n653,n654);
nor (n654,n655,n656);
and (n655,n69,n33);
and (n656,n70,n34);
nand (n657,n526,n111);
nand (n658,n659,n664);
or (n659,n660,n94);
not (n660,n661);
nand (n661,n662,n663);
or (n662,n575,n87);
nand (n663,n575,n87);
nand (n664,n89,n601);
nand (n665,n666,n669);
or (n666,n667,n158);
not (n667,n668);
nand (n669,n160,n608);
and (n670,n651,n658);
nand (n671,n672,n676);
or (n672,n53,n673);
nor (n673,n674,n675);
and (n674,n63,n325);
and (n675,n64,n324);
or (n676,n54,n558);
and (n677,n645,n646);
and (n678,n591,n592);
or (n679,n680,n756);
and (n680,n681,n684);
xor (n681,n682,n683);
xor (n682,n510,n513);
xor (n683,n590,n642);
or (n684,n685,n755);
and (n685,n686,n719);
xor (n686,n687,n688);
xor (n687,n594,n640);
or (n688,n689,n718);
and (n689,n690,n716);
xor (n690,n691,n715);
or (n691,n692,n714);
and (n692,n693,n708);
xor (n693,n694,n701);
nand (n694,n695,n700);
or (n695,n696,n420);
not (n696,n697);
nor (n697,n698,n699);
and (n698,n24,n288);
and (n699,n25,n289);
nand (n700,n413,n615);
nand (n701,n702,n707);
or (n702,n703,n29);
not (n703,n704);
nor (n704,n705,n706);
and (n705,n100,n26);
and (n706,n101,n27);
nand (n707,n31,n623);
nand (n708,n709,n712);
or (n709,n431,n710);
not (n710,n711);
xor (n711,n189,n113);
or (n712,n629,n713);
not (n713,n285);
and (n714,n694,n701);
xor (n715,n619,n633);
nand (n716,n717,n523);
or (n717,n417,n524);
and (n718,n691,n715);
or (n719,n720,n754);
and (n720,n721,n753);
xor (n721,n722,n723);
xor (n722,n597,n610);
or (n723,n724,n752);
and (n724,n725,n741);
xor (n725,n726,n734);
nand (n726,n727,n732);
or (n727,n728,n139);
not (n728,n729);
nand (n729,n730,n731);
or (n730,n58,n235);
or (n731,n60,n236);
nand (n732,n733,n142);
not (n733,n635);
nand (n734,n735,n740);
or (n735,n736,n53);
not (n736,n737);
nand (n737,n738,n739);
or (n738,n64,n383);
or (n739,n63,n384);
or (n740,n54,n673);
nand (n741,n742,n751);
or (n742,n743,n746);
nand (n743,n744,n417);
not (n744,n745);
not (n746,n747);
nor (n747,n748,n750);
and (n748,n120,n749);
not (n749,n417);
and (n750,n118,n417);
or (n751,n749,n744);
and (n752,n726,n734);
xor (n753,n671,n648);
and (n754,n722,n723);
and (n755,n687,n688);
and (n756,n682,n683);
nor (n757,n758,n759);
xor (n758,n681,n684);
or (n759,n760,n848);
and (n760,n761,n847);
xor (n761,n762,n763);
xor (n762,n644,n647);
or (n763,n764,n846);
and (n764,n765,n845);
xor (n765,n766,n838);
or (n766,n767,n837);
and (n767,n768,n812);
xor (n768,n769,n787);
or (n769,n770,n786);
and (n770,n771,n779);
xor (n771,n772,n773);
and (n772,n160,n668);
nand (n773,n774,n778);
or (n774,n743,n775);
nor (n775,n776,n777);
and (n776,n45,n417);
and (n777,n46,n749);
nand (n778,n747,n745);
nand (n779,n780,n785);
or (n780,n781,n420);
not (n781,n782);
nor (n782,n783,n784);
and (n783,n136,n288);
and (n784,n137,n289);
nand (n785,n413,n697);
and (n786,n772,n773);
or (n787,n788,n811);
and (n788,n789,n804);
xor (n789,n790,n797);
nand (n790,n791,n796);
or (n791,n792,n431);
not (n792,n793);
nor (n793,n794,n795);
and (n794,n77,n113);
and (n795,n75,n114);
nand (n796,n711,n285);
nand (n797,n798,n799);
or (n798,n141,n728);
nand (n799,n800,n140);
not (n800,n801);
nor (n801,n802,n803);
and (n802,n325,n60);
and (n803,n324,n58);
nand (n804,n805,n806);
or (n805,n736,n54);
nand (n806,n807,n355);
not (n807,n808);
nor (n808,n809,n810);
and (n809,n447,n63);
and (n810,n64,n446);
and (n811,n790,n797);
or (n812,n813,n836);
and (n813,n814,n829);
xor (n814,n815,n822);
nand (n815,n816,n821);
or (n816,n817,n94);
not (n817,n818);
nor (n818,n819,n820);
and (n819,n607,n87);
and (n820,n608,n84);
nand (n821,n661,n89);
nand (n822,n823,n828);
or (n823,n824,n105);
not (n824,n825);
nand (n825,n826,n827);
or (n826,n34,n86);
or (n827,n33,n83);
nand (n828,n111,n654);
nand (n829,n830,n835);
or (n830,n29,n831);
not (n831,n832);
nor (n832,n833,n834);
and (n833,n156,n26);
and (n834,n157,n27);
or (n835,n178,n703);
and (n836,n815,n822);
and (n837,n769,n787);
or (n838,n839,n844);
and (n839,n840,n843);
xor (n840,n841,n842);
xor (n841,n650,n665);
xor (n842,n693,n708);
xor (n843,n725,n741);
and (n844,n841,n842);
xor (n845,n690,n716);
and (n846,n766,n838);
xor (n847,n686,n719);
and (n848,n762,n763);
nor (n849,n850,n861);
nor (n850,n851,n852);
xor (n851,n398,n401);
or (n852,n853,n860);
and (n853,n854,n857);
xor (n854,n855,n856);
xor (n855,n363,n388);
xor (n856,n403,n465);
or (n857,n858,n859);
and (n858,n536,n587);
and (n859,n537,n538);
and (n860,n855,n856);
nor (n861,n862,n863);
xor (n862,n854,n857);
or (n863,n864,n865);
and (n864,n507,n588);
and (n865,n508,n535);
nand (n866,n867,n1193);
or (n867,n868,n1175);
not (n868,n869);
nor (n869,n870,n1174);
and (n870,n871,n1112);
nand (n871,n872,n1017);
xor (n872,n873,n1004);
xor (n873,n874,n875);
xor (n874,n840,n843);
or (n875,n876,n1003);
and (n876,n877,n973);
xor (n877,n878,n925);
or (n878,n879,n924);
and (n879,n880,n901);
xor (n880,n881,n887);
nand (n881,n882,n886);
or (n882,n53,n883);
nor (n883,n884,n885);
and (n884,n63,n575);
and (n885,n64,n574);
or (n886,n54,n808);
xor (n887,n888,n894);
nor (n888,n889,n87);
nor (n889,n890,n892);
and (n890,n891,n63);
nand (n891,n668,n91);
and (n892,n667,n893);
not (n893,n91);
nand (n894,n895,n900);
or (n895,n896,n743);
not (n896,n897);
nor (n897,n898,n899);
and (n898,n24,n749);
and (n899,n25,n417);
or (n900,n775,n744);
or (n901,n902,n923);
and (n902,n903,n912);
xor (n903,n904,n905);
and (n904,n89,n668);
nand (n905,n906,n911);
or (n906,n743,n907);
not (n907,n908);
nor (n908,n909,n910);
and (n909,n136,n749);
and (n910,n137,n417);
nand (n911,n897,n745);
nand (n912,n913,n918);
or (n913,n420,n914);
not (n914,n915);
nor (n915,n916,n917);
and (n916,n288,n77);
and (n917,n75,n289);
or (n918,n421,n919);
not (n919,n920);
nor (n920,n921,n922);
and (n921,n189,n288);
and (n922,n187,n289);
and (n923,n904,n905);
and (n924,n881,n887);
xor (n925,n926,n949);
xor (n926,n927,n928);
and (n927,n888,n894);
or (n928,n929,n948);
and (n929,n930,n941);
xor (n930,n931,n934);
nand (n931,n932,n933);
or (n932,n919,n420);
nand (n933,n782,n413);
nand (n934,n935,n940);
or (n935,n936,n94);
not (n936,n937);
nand (n937,n938,n939);
or (n938,n87,n668);
or (n939,n84,n667);
nand (n940,n818,n89);
nand (n941,n942,n943);
or (n942,n824,n110);
or (n943,n105,n944);
not (n944,n945);
nor (n945,n946,n947);
and (n946,n100,n33);
and (n947,n101,n34);
and (n948,n931,n934);
or (n949,n950,n972);
and (n950,n951,n966);
xor (n951,n952,n959);
nand (n952,n953,n958);
or (n953,n954,n29);
not (n954,n955);
nor (n955,n956,n957);
and (n956,n235,n26);
and (n957,n236,n27);
nand (n958,n31,n832);
nand (n959,n960,n965);
or (n960,n961,n431);
not (n961,n962);
nand (n962,n963,n964);
or (n963,n114,n69);
or (n964,n113,n70);
nand (n965,n285,n793);
nand (n966,n967,n971);
or (n967,n139,n968);
nor (n968,n969,n970);
and (n969,n60,n384);
and (n970,n58,n383);
or (n971,n141,n801);
and (n972,n952,n959);
or (n973,n974,n1002);
and (n974,n975,n1001);
xor (n975,n976,n1000);
or (n976,n977,n999);
and (n977,n978,n992);
xor (n978,n979,n986);
nand (n979,n980,n985);
or (n980,n981,n105);
not (n981,n982);
nor (n982,n983,n984);
and (n983,n157,n34);
and (n984,n156,n33);
nand (n985,n111,n945);
nand (n986,n987,n991);
or (n987,n29,n988);
nor (n988,n989,n990);
and (n989,n324,n27);
and (n990,n325,n26);
nand (n991,n31,n955);
nand (n992,n993,n994);
or (n993,n713,n961);
nand (n994,n995,n291);
not (n995,n996);
nor (n996,n997,n998);
and (n997,n113,n83);
and (n998,n114,n86);
and (n999,n979,n986);
xor (n1000,n951,n966);
xor (n1001,n930,n941);
and (n1002,n976,n1000);
and (n1003,n878,n925);
xor (n1004,n1005,n1010);
xor (n1005,n1006,n1009);
or (n1006,n1007,n1008);
and (n1007,n926,n949);
and (n1008,n927,n928);
xor (n1009,n768,n812);
or (n1010,n1011,n1016);
and (n1011,n1012,n1015);
xor (n1012,n1013,n1014);
xor (n1013,n789,n804);
xor (n1014,n771,n779);
xor (n1015,n814,n829);
and (n1016,n1013,n1014);
or (n1017,n1018,n1111);
and (n1018,n1019,n1110);
xor (n1019,n1020,n1021);
xor (n1020,n1012,n1015);
or (n1021,n1022,n1109);
and (n1022,n1023,n1056);
xor (n1023,n1024,n1055);
or (n1024,n1025,n1054);
and (n1025,n1026,n1041);
xor (n1026,n1027,n1034);
nand (n1027,n1028,n1032);
or (n1028,n1029,n139);
nor (n1029,n1030,n1031);
and (n1030,n446,n58);
and (n1031,n447,n60);
nand (n1032,n1033,n142);
not (n1033,n968);
nand (n1034,n1035,n1039);
or (n1035,n53,n1036);
nor (n1036,n1037,n1038);
and (n1037,n63,n608);
and (n1038,n64,n607);
nand (n1039,n1040,n264);
not (n1040,n883);
and (n1041,n1042,n1047);
nor (n1042,n1043,n63);
nor (n1043,n1044,n1046);
and (n1044,n1045,n60);
nand (n1045,n668,n57);
and (n1046,n667,n56);
nand (n1047,n1048,n1053);
or (n1048,n743,n1049);
not (n1049,n1050);
nor (n1050,n1051,n1052);
and (n1051,n189,n749);
and (n1052,n187,n417);
nand (n1053,n908,n745);
and (n1054,n1027,n1034);
xor (n1055,n880,n901);
or (n1056,n1057,n1108);
and (n1057,n1058,n1107);
xor (n1058,n1059,n1084);
or (n1059,n1060,n1083);
and (n1060,n1061,n1076);
xor (n1061,n1062,n1069);
nand (n1062,n1063,n1068);
or (n1063,n1064,n420);
not (n1064,n1065);
nor (n1065,n1066,n1067);
and (n1066,n69,n288);
and (n1067,n70,n289);
nand (n1068,n915,n413);
nand (n1069,n1070,n1075);
or (n1070,n1071,n105);
not (n1071,n1072);
nand (n1072,n1073,n1074);
or (n1073,n34,n235);
or (n1074,n33,n236);
nand (n1075,n111,n982);
nand (n1076,n1077,n1082);
or (n1077,n29,n1078);
not (n1078,n1079);
nor (n1079,n1080,n1081);
and (n1080,n383,n26);
and (n1081,n384,n27);
or (n1082,n178,n988);
and (n1083,n1062,n1069);
or (n1084,n1085,n1106);
and (n1085,n1086,n1100);
xor (n1086,n1087,n1093);
nand (n1087,n1088,n1092);
or (n1088,n431,n1089);
nor (n1089,n1090,n1091);
and (n1090,n101,n113);
and (n1091,n100,n114);
or (n1092,n996,n713);
nand (n1093,n1094,n1099);
or (n1094,n139,n1095);
not (n1095,n1096);
nor (n1096,n1097,n1098);
and (n1097,n574,n60);
and (n1098,n575,n58);
or (n1099,n1029,n141);
nand (n1100,n1101,n1105);
or (n1101,n53,n1102);
nor (n1102,n1103,n1104);
and (n1103,n667,n64);
and (n1104,n668,n63);
or (n1105,n1036,n54);
and (n1106,n1087,n1093);
xor (n1107,n903,n912);
and (n1108,n1059,n1084);
and (n1109,n1024,n1055);
xor (n1110,n877,n973);
and (n1111,n1020,n1021);
nand (n1112,n1113,n1114);
xor (n1113,n1019,n1110);
or (n1114,n1115,n1173);
and (n1115,n1116,n1172);
xor (n1116,n1117,n1118);
xor (n1117,n975,n1001);
or (n1118,n1119,n1171);
and (n1119,n1120,n1123);
xor (n1120,n1121,n1122);
xor (n1121,n978,n992);
xor (n1122,n1026,n1041);
or (n1123,n1124,n1170);
and (n1124,n1125,n1145);
xor (n1125,n1126,n1127);
xor (n1126,n1042,n1047);
or (n1127,n1128,n1144);
and (n1128,n1129,n1138);
xor (n1129,n1130,n1131);
and (n1130,n264,n668);
nand (n1131,n1132,n1137);
or (n1132,n1133,n420);
not (n1133,n1134);
nor (n1134,n1135,n1136);
and (n1135,n86,n288);
and (n1136,n83,n289);
nand (n1137,n413,n1065);
nand (n1138,n1139,n1140);
or (n1139,n1071,n110);
or (n1140,n105,n1141);
nor (n1141,n1142,n1143);
and (n1142,n33,n325);
and (n1143,n34,n324);
and (n1144,n1130,n1131);
or (n1145,n1146,n1169);
and (n1146,n1147,n1162);
xor (n1147,n1148,n1155);
nand (n1148,n1149,n1154);
or (n1149,n1150,n29);
not (n1150,n1151);
nand (n1151,n1152,n1153);
or (n1152,n446,n27);
or (n1153,n26,n447);
nand (n1154,n1079,n31);
nand (n1155,n1156,n1157);
or (n1156,n744,n1049);
nand (n1157,n1158,n1161);
nor (n1158,n1159,n1160);
and (n1159,n77,n749);
and (n1160,n75,n417);
not (n1161,n743);
nand (n1162,n1163,n1168);
or (n1163,n1164,n139);
not (n1164,n1165);
nand (n1165,n1166,n1167);
or (n1166,n58,n607);
or (n1167,n60,n608);
nand (n1168,n1096,n142);
and (n1169,n1148,n1155);
and (n1170,n1126,n1127);
and (n1171,n1121,n1122);
xor (n1172,n1023,n1056);
and (n1173,n1117,n1118);
nor (n1174,n872,n1017);
not (n1175,n1176);
nor (n1176,n1177,n1188);
nor (n1177,n1178,n1179);
xor (n1178,n761,n847);
or (n1179,n1180,n1187);
and (n1180,n1181,n1186);
xor (n1181,n1182,n1183);
xor (n1182,n721,n753);
or (n1183,n1184,n1185);
and (n1184,n1005,n1010);
and (n1185,n1006,n1009);
xor (n1186,n765,n845);
and (n1187,n1182,n1183);
nor (n1188,n1189,n1190);
xor (n1189,n1181,n1186);
or (n1190,n1191,n1192);
and (n1191,n873,n1004);
and (n1192,n874,n875);
nor (n1193,n1194,n1198);
and (n1194,n1195,n1196);
not (n1195,n1177);
not (n1196,n1197);
nand (n1197,n1189,n1190);
and (n1198,n1178,n1179);
nand (n1199,n1200,n1207);
or (n1200,n1201,n1202);
not (n1201,n849);
not (n1202,n1203);
nor (n1203,n1204,n505);
and (n1204,n1205,n1206);
nand (n1205,n679,n506);
nand (n1206,n758,n759);
nor (n1207,n1208,n1212);
and (n1208,n1209,n1210);
not (n1209,n850);
not (n1210,n1211);
nand (n1211,n862,n863);
and (n1212,n851,n852);
nand (n1213,n503,n1214,n1217);
and (n1214,n1176,n1215);
nor (n1215,n1174,n1216);
nor (n1216,n1113,n1114);
nand (n1217,n1218,n1718);
or (n1218,n1219,n1654);
not (n1219,n1220);
nand (n1220,n1221,n1643,n1653);
nand (n1221,n1222,n1449,n1510);
nor (n1222,n1223,n1387);
not (n1223,n1224);
or (n1224,n1225,n1350);
xor (n1225,n1226,n1310);
xor (n1226,n1227,n1257);
xor (n1227,n1228,n1248);
xor (n1228,n1229,n1239);
nand (n1229,n1230,n1235);
or (n1230,n1231,n29);
not (n1231,n1232);
nor (n1232,n1233,n1234);
and (n1233,n607,n26);
and (n1234,n608,n27);
nand (n1235,n31,n1236);
nand (n1236,n1237,n1238);
or (n1237,n27,n574);
or (n1238,n26,n575);
nand (n1239,n1240,n1244);
or (n1240,n1241,n743);
nor (n1241,n1242,n1243);
and (n1242,n749,n83);
and (n1243,n417,n86);
or (n1244,n1245,n744);
nor (n1245,n1246,n1247);
and (n1246,n749,n70);
and (n1247,n417,n69);
nand (n1248,n1249,n1253);
or (n1249,n431,n1250);
nor (n1250,n1251,n1252);
and (n1251,n113,n325);
and (n1252,n114,n324);
or (n1253,n1254,n713);
nor (n1254,n1255,n1256);
and (n1255,n113,n236);
and (n1256,n114,n235);
or (n1257,n1258,n1309);
and (n1258,n1259,n1284);
xor (n1259,n1260,n1266);
nand (n1260,n1261,n1265);
or (n1261,n431,n1262);
nor (n1262,n1263,n1264);
and (n1263,n113,n384);
and (n1264,n114,n383);
or (n1265,n713,n1250);
xor (n1266,n1267,n1273);
and (n1267,n1268,n27);
nand (n1268,n1269,n1270);
or (n1269,n668,n35);
nand (n1270,n1271,n33);
not (n1271,n1272);
and (n1272,n668,n35);
nand (n1273,n1274,n1279);
or (n1274,n1275,n421);
not (n1275,n1276);
nand (n1276,n1277,n1278);
or (n1277,n289,n156);
or (n1278,n288,n157);
nand (n1279,n1280,n419);
not (n1280,n1281);
nor (n1281,n1282,n1283);
and (n1282,n288,n236);
and (n1283,n289,n235);
or (n1284,n1285,n1308);
and (n1285,n1286,n1298);
xor (n1286,n1287,n1288);
and (n1287,n31,n668);
nand (n1288,n1289,n1294);
or (n1289,n744,n1290);
not (n1290,n1291);
nor (n1291,n1292,n1293);
and (n1292,n100,n749);
and (n1293,n101,n417);
or (n1294,n1295,n743);
nor (n1295,n1296,n1297);
and (n1296,n749,n157);
and (n1297,n417,n156);
nand (n1298,n1299,n1303);
or (n1299,n105,n1300);
nor (n1300,n1301,n1302);
and (n1301,n33,n608);
and (n1302,n34,n607);
or (n1303,n110,n1304);
not (n1304,n1305);
nor (n1305,n1306,n1307);
and (n1306,n575,n34);
and (n1307,n574,n33);
and (n1308,n1287,n1288);
and (n1309,n1260,n1266);
xor (n1310,n1311,n1333);
xor (n1311,n1312,n1313);
and (n1312,n1267,n1273);
or (n1313,n1314,n1332);
and (n1314,n1315,n1329);
xor (n1315,n1316,n1322);
nand (n1316,n1317,n1318);
or (n1317,n1304,n105);
nand (n1318,n111,n1319);
nor (n1319,n1320,n1321);
and (n1320,n446,n33);
and (n1321,n447,n34);
nand (n1322,n1323,n1328);
or (n1323,n1324,n29);
not (n1324,n1325);
nand (n1325,n1326,n1327);
or (n1326,n26,n668);
or (n1327,n667,n27);
nand (n1328,n31,n1232);
nand (n1329,n1330,n1331);
or (n1330,n743,n1290);
or (n1331,n1241,n744);
and (n1332,n1316,n1322);
xor (n1333,n1334,n1342);
xor (n1334,n1335,n1336);
and (n1335,n142,n668);
nand (n1336,n1337,n1338);
or (n1337,n1275,n420);
nand (n1338,n413,n1339);
nand (n1339,n1340,n1341);
or (n1340,n289,n100);
or (n1341,n288,n101);
nand (n1342,n1343,n1345);
or (n1343,n1344,n105);
not (n1344,n1319);
nand (n1345,n1346,n111);
not (n1346,n1347);
nor (n1347,n1348,n1349);
and (n1348,n33,n384);
and (n1349,n34,n383);
or (n1350,n1351,n1386);
and (n1351,n1352,n1385);
xor (n1352,n1353,n1354);
xor (n1353,n1315,n1329);
or (n1354,n1355,n1384);
and (n1355,n1356,n1369);
xor (n1356,n1357,n1363);
nand (n1357,n1358,n1362);
or (n1358,n420,n1359);
nor (n1359,n1360,n1361);
and (n1360,n288,n325);
and (n1361,n289,n324);
or (n1362,n421,n1281);
nand (n1363,n1364,n1368);
or (n1364,n431,n1365);
nor (n1365,n1366,n1367);
and (n1366,n113,n447);
and (n1367,n114,n446);
or (n1368,n1262,n713);
and (n1369,n1370,n1377);
nor (n1370,n1371,n33);
nor (n1371,n1372,n1375);
and (n1372,n1373,n113);
not (n1373,n1374);
and (n1374,n668,n108);
and (n1375,n667,n1376);
not (n1376,n108);
nand (n1377,n1378,n1383);
or (n1378,n1379,n743);
not (n1379,n1380);
nor (n1380,n1381,n1382);
and (n1381,n235,n749);
and (n1382,n236,n417);
or (n1383,n1295,n744);
and (n1384,n1357,n1363);
xor (n1385,n1259,n1284);
and (n1386,n1353,n1354);
nand (n1387,n1388,n1443);
not (n1388,n1389);
nor (n1389,n1390,n1418);
xor (n1390,n1391,n1417);
xor (n1391,n1392,n1416);
or (n1392,n1393,n1415);
and (n1393,n1394,n1409);
xor (n1394,n1395,n1403);
nand (n1395,n1396,n1401);
or (n1396,n1397,n105);
not (n1397,n1398);
nand (n1398,n1399,n1400);
or (n1399,n33,n668);
or (n1400,n34,n667);
nand (n1401,n1402,n111);
not (n1402,n1300);
nand (n1403,n1404,n1408);
or (n1404,n420,n1405);
nor (n1405,n1406,n1407);
and (n1406,n288,n384);
and (n1407,n289,n383);
or (n1408,n1359,n421);
nand (n1409,n1410,n1414);
or (n1410,n431,n1411);
nor (n1411,n1412,n1413);
and (n1412,n113,n575);
and (n1413,n114,n574);
or (n1414,n1365,n713);
and (n1415,n1395,n1403);
xor (n1416,n1286,n1298);
xor (n1417,n1356,n1369);
or (n1418,n1419,n1442);
and (n1419,n1420,n1441);
xor (n1420,n1421,n1422);
xor (n1421,n1370,n1377);
or (n1422,n1423,n1440);
and (n1423,n1424,n1433);
xor (n1424,n1425,n1426);
and (n1425,n111,n668);
nand (n1426,n1427,n1432);
or (n1427,n743,n1428);
not (n1428,n1429);
nor (n1429,n1430,n1431);
and (n1430,n325,n417);
and (n1431,n324,n749);
nand (n1432,n1380,n745);
nand (n1433,n1434,n1439);
or (n1434,n420,n1435);
not (n1435,n1436);
nor (n1436,n1437,n1438);
and (n1437,n446,n288);
and (n1438,n447,n289);
or (n1439,n421,n1405);
and (n1440,n1425,n1426);
xor (n1441,n1394,n1409);
and (n1442,n1421,n1422);
not (n1443,n1444);
nor (n1444,n1445,n1446);
xor (n1445,n1352,n1385);
or (n1446,n1447,n1448);
and (n1447,n1391,n1417);
and (n1448,n1392,n1416);
nand (n1449,n1450,n1506);
not (n1450,n1451);
xor (n1451,n1452,n1503);
xor (n1452,n1453,n1483);
xor (n1453,n1454,n1468);
xor (n1454,n1455,n1462);
nand (n1455,n1456,n1457);
or (n1456,n1164,n141);
nand (n1457,n1458,n140);
not (n1458,n1459);
nor (n1459,n1460,n1461);
and (n1460,n667,n58);
and (n1461,n60,n668);
nand (n1462,n1463,n1464);
or (n1463,n431,n1254);
or (n1464,n713,n1465);
nor (n1465,n1466,n1467);
and (n1466,n113,n157);
and (n1467,n114,n156);
nand (n1468,n1469,n1482);
or (n1469,n1470,n1477);
not (n1470,n1471);
nand (n1471,n1472,n58);
nand (n1472,n1473,n1474);
or (n1473,n668,n145);
nand (n1474,n1475,n26);
not (n1475,n1476);
and (n1476,n668,n145);
not (n1477,n1478);
nand (n1478,n1479,n1481);
or (n1479,n1480,n420);
not (n1480,n1339);
nand (n1481,n413,n1134);
or (n1482,n1478,n1471);
xor (n1483,n1484,n1491);
xor (n1484,n1485,n1488);
or (n1485,n1486,n1487);
and (n1486,n1334,n1342);
and (n1487,n1335,n1336);
or (n1488,n1489,n1490);
and (n1489,n1228,n1248);
and (n1490,n1229,n1239);
xor (n1491,n1492,n1499);
xor (n1492,n1493,n1496);
nand (n1493,n1494,n1495);
or (n1494,n105,n1347);
or (n1495,n1141,n110);
nand (n1496,n1497,n1498);
or (n1497,n1150,n178);
nand (n1498,n30,n1236);
nand (n1499,n1500,n1501);
or (n1500,n1245,n743);
or (n1501,n1502,n744);
not (n1502,n1158);
or (n1503,n1504,n1505);
and (n1504,n1311,n1333);
and (n1505,n1312,n1313);
not (n1506,n1507);
or (n1507,n1508,n1509);
and (n1508,n1226,n1310);
and (n1509,n1227,n1257);
or (n1510,n1511,n1642);
and (n1511,n1512,n1539);
xor (n1512,n1513,n1538);
or (n1513,n1514,n1537);
and (n1514,n1515,n1536);
xor (n1515,n1516,n1523);
nand (n1516,n1517,n1522);
or (n1517,n431,n1518);
not (n1518,n1519);
nor (n1519,n1520,n1521);
and (n1520,n608,n114);
and (n1521,n607,n113);
or (n1522,n1411,n713);
and (n1523,n1524,n1530);
nor (n1524,n1525,n113);
nor (n1525,n1526,n1529);
and (n1526,n1527,n288);
not (n1527,n1528);
and (n1528,n668,n287);
and (n1529,n667,n294);
nand (n1530,n1531,n1532);
or (n1531,n744,n1428);
nand (n1532,n1533,n1161);
nand (n1533,n1534,n1535);
or (n1534,n384,n749);
nand (n1535,n749,n384);
xor (n1536,n1424,n1433);
and (n1537,n1516,n1523);
xor (n1538,n1420,n1441);
or (n1539,n1540,n1641);
and (n1540,n1541,n1560);
xor (n1541,n1542,n1559);
or (n1542,n1543,n1558);
and (n1543,n1544,n1557);
xor (n1544,n1545,n1550);
nand (n1545,n1546,n1549);
or (n1546,n1547,n420);
not (n1547,n1548);
xor (n1548,n574,n288);
nand (n1549,n413,n1436);
nand (n1550,n1551,n1556);
or (n1551,n1552,n431);
not (n1552,n1553);
nand (n1553,n1554,n1555);
or (n1554,n113,n668);
or (n1555,n667,n114);
nand (n1556,n1519,n285);
xor (n1557,n1524,n1530);
and (n1558,n1545,n1550);
xor (n1559,n1515,n1536);
or (n1560,n1561,n1640);
and (n1561,n1562,n1584);
xor (n1562,n1563,n1583);
or (n1563,n1564,n1582);
and (n1564,n1565,n1574);
xor (n1565,n1566,n1567);
and (n1566,n285,n668);
nand (n1567,n1568,n1573);
or (n1568,n1569,n420);
not (n1569,n1570);
nor (n1570,n1571,n1572);
and (n1571,n607,n288);
and (n1572,n608,n289);
nand (n1573,n413,n1548);
nand (n1574,n1575,n1580);
or (n1575,n743,n1576);
not (n1576,n1577);
nand (n1577,n1578,n1579);
or (n1578,n447,n749);
nand (n1579,n749,n447);
or (n1580,n1581,n744);
not (n1581,n1533);
and (n1582,n1566,n1567);
xor (n1583,n1544,n1557);
nand (n1584,n1585,n1639);
or (n1585,n1586,n1601);
nor (n1586,n1587,n1588);
xor (n1587,n1565,n1574);
nor (n1588,n1589,n1596);
not (n1589,n1590);
nand (n1590,n1591,n1595);
or (n1591,n743,n1592);
nor (n1592,n1593,n1594);
and (n1593,n574,n417);
and (n1594,n575,n749);
nand (n1595,n1577,n745);
nand (n1596,n1597,n289);
nand (n1597,n1598,n1600);
or (n1598,n1599,n417);
and (n1599,n668,n416);
or (n1600,n668,n416);
nor (n1601,n1602,n1638);
and (n1602,n1603,n1614);
nand (n1603,n1604,n1608);
nor (n1604,n1605,n1606);
and (n1605,n1596,n1590);
and (n1606,n1607,n1589);
not (n1607,n1596);
nor (n1608,n1609,n1613);
and (n1609,n419,n1610);
nand (n1610,n1611,n1612);
or (n1611,n288,n668);
or (n1612,n667,n289);
and (n1613,n413,n1570);
nand (n1614,n1615,n1637);
or (n1615,n1616,n1631);
not (n1616,n1617);
nor (n1617,n1618,n1629);
not (n1618,n1619);
nand (n1619,n1620,n1625);
or (n1620,n744,n1621);
not (n1621,n1622);
nor (n1622,n1623,n1624);
and (n1623,n607,n749);
and (n1624,n608,n417);
nand (n1625,n1626,n1161);
nor (n1626,n1627,n1628);
and (n1627,n667,n749);
and (n1628,n668,n417);
nand (n1629,n1630,n417);
nand (n1630,n668,n745);
not (n1631,n1632);
nand (n1632,n1633,n1636);
nor (n1633,n1634,n1635);
nor (n1634,n1621,n743);
nor (n1635,n1592,n744);
nand (n1636,n668,n413);
or (n1637,n1633,n1636);
nor (n1638,n1608,n1604);
nand (n1639,n1587,n1588);
and (n1640,n1563,n1583);
and (n1641,n1542,n1559);
and (n1642,n1513,n1538);
nand (n1643,n1644,n1449);
or (n1644,n1645,n1647);
not (n1645,n1646);
nand (n1646,n1225,n1350);
not (n1647,n1648);
nand (n1648,n1224,n1649);
nand (n1649,n1650,n1652);
or (n1650,n1444,n1651);
nand (n1651,n1390,n1418);
nand (n1652,n1445,n1446);
nand (n1653,n1451,n1507);
not (n1654,n1655);
nor (n1655,n1656,n1681);
nor (n1656,n1657,n1658);
xor (n1657,n1116,n1172);
or (n1658,n1659,n1680);
and (n1659,n1660,n1663);
xor (n1660,n1661,n1662);
xor (n1661,n1058,n1107);
xor (n1662,n1120,n1123);
or (n1663,n1664,n1679);
and (n1664,n1665,n1668);
xor (n1665,n1666,n1667);
xor (n1666,n1086,n1100);
xor (n1667,n1061,n1076);
or (n1668,n1669,n1678);
and (n1669,n1670,n1675);
xor (n1670,n1671,n1674);
nand (n1671,n1672,n1673);
or (n1672,n431,n1465);
or (n1673,n1089,n713);
nor (n1674,n1477,n1471);
or (n1675,n1676,n1677);
and (n1676,n1492,n1499);
and (n1677,n1493,n1496);
and (n1678,n1671,n1674);
and (n1679,n1666,n1667);
and (n1680,n1661,n1662);
nand (n1681,n1682,n1711);
nor (n1682,n1683,n1706);
nor (n1683,n1684,n1697);
xor (n1684,n1685,n1696);
xor (n1685,n1686,n1687);
xor (n1686,n1125,n1145);
or (n1687,n1688,n1695);
and (n1688,n1689,n1692);
xor (n1689,n1690,n1691);
xor (n1690,n1147,n1162);
xor (n1691,n1129,n1138);
or (n1692,n1693,n1694);
and (n1693,n1454,n1468);
and (n1694,n1455,n1462);
and (n1695,n1690,n1691);
xor (n1696,n1665,n1668);
or (n1697,n1698,n1705);
and (n1698,n1699,n1704);
xor (n1699,n1700,n1701);
xor (n1700,n1670,n1675);
or (n1701,n1702,n1703);
and (n1702,n1484,n1491);
and (n1703,n1485,n1488);
xor (n1704,n1689,n1692);
and (n1705,n1700,n1701);
nor (n1706,n1707,n1710);
or (n1707,n1708,n1709);
and (n1708,n1452,n1503);
and (n1709,n1453,n1483);
xor (n1710,n1699,n1704);
nand (n1711,n1712,n1714);
not (n1712,n1713);
xor (n1713,n1660,n1663);
not (n1714,n1715);
or (n1715,n1716,n1717);
and (n1716,n1685,n1696);
and (n1717,n1686,n1687);
nor (n1718,n1719,n1730);
and (n1719,n1720,n1729);
nand (n1720,n1721,n1728);
or (n1721,n1722,n1723);
not (n1722,n1711);
not (n1723,n1724);
nand (n1724,n1725,n1727);
or (n1725,n1683,n1726);
nand (n1726,n1707,n1710);
nand (n1727,n1684,n1697);
nand (n1728,n1713,n1715);
not (n1729,n1656);
and (n1730,n1657,n1658);
nand (n1731,n498,n396);
nand (n1732,n393,n11);
not (n1733,n1734);
nand (n1734,n1735,n6);
not (n1735,n7);
wire s0n1736,s1n1736,notn1736;
or (n1736,s0n1736,s1n1736);
not(notn1736,n7);
and (s0n1736,notn1736,n1737);
and (s1n1736,n7,1'b0);
wire s0n1737,s1n1737,notn1737;
or (n1737,s0n1737,s1n1737);
not(notn1737,n6);
and (s0n1737,notn1737,n3);
and (s1n1737,n6,n1738);
xor (n1738,n1739,n3005);
xor (n1739,n1740,n3004);
xor (n1740,n1741,n2953);
xor (n1741,n1742,n130);
xor (n1742,n1743,n2890);
xor (n1743,n1744,n2889);
xor (n1744,n1745,n2823);
xor (n1745,n1746,n2822);
xor (n1746,n1747,n2747);
xor (n1747,n1748,n2746);
xor (n1748,n1749,n2670);
xor (n1749,n1750,n153);
xor (n1750,n1751,n2584);
xor (n1751,n1752,n2583);
xor (n1752,n1753,n2500);
xor (n1753,n1754,n2499);
or (n1754,n1755,n2405);
and (n1755,n1756,n2404);
or (n1756,n1757,n2318);
and (n1757,n1758,n2317);
or (n1758,n1759,n2223);
and (n1759,n1760,n2222);
or (n1760,n1761,n2130);
and (n1761,n1762,n333);
or (n1762,n1763,n2036);
and (n1763,n1764,n2035);
or (n1764,n1765,n1948);
and (n1765,n1766,n492);
or (n1766,n1767,n1854);
and (n1767,n1768,n1853);
and (n1768,n750,n1769);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
and (n1771,n118,n745);
and (n1772,n46,n417);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1778);
and (n1776,n1777,n899);
and (n1777,n46,n745);
and (n1778,n1779,n1780);
xor (n1779,n1777,n899);
or (n1780,n1781,n1783);
and (n1781,n1782,n910);
and (n1782,n25,n745);
and (n1783,n1784,n1785);
xor (n1784,n1782,n910);
or (n1785,n1786,n1788);
and (n1786,n1787,n1052);
and (n1787,n137,n745);
and (n1788,n1789,n1790);
xor (n1789,n1787,n1052);
or (n1790,n1791,n1793);
and (n1791,n1792,n1160);
and (n1792,n187,n745);
and (n1793,n1794,n1795);
xor (n1794,n1792,n1160);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
and (n1797,n75,n745);
and (n1798,n70,n417);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
and (n1803,n70,n745);
and (n1804,n83,n417);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1810);
and (n1808,n1809,n1293);
and (n1809,n83,n745);
and (n1810,n1811,n1812);
xor (n1811,n1809,n1293);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
and (n1814,n101,n745);
and (n1815,n157,n417);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1821);
and (n1819,n1820,n1382);
and (n1820,n157,n745);
and (n1821,n1822,n1823);
xor (n1822,n1820,n1382);
or (n1823,n1824,n1826);
and (n1824,n1825,n1430);
and (n1825,n236,n745);
and (n1826,n1827,n1828);
xor (n1827,n1825,n1430);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
and (n1830,n325,n745);
and (n1831,n384,n417);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1838);
and (n1835,n1836,n1837);
and (n1836,n384,n745);
and (n1837,n447,n417);
and (n1838,n1839,n1840);
xor (n1839,n1836,n1837);
or (n1840,n1841,n1844);
and (n1841,n1842,n1843);
and (n1842,n447,n745);
and (n1843,n575,n417);
and (n1844,n1845,n1846);
xor (n1845,n1842,n1843);
or (n1846,n1847,n1849);
and (n1847,n1848,n1624);
and (n1848,n575,n745);
and (n1849,n1850,n1851);
xor (n1850,n1848,n1624);
and (n1851,n1852,n1628);
and (n1852,n608,n745);
and (n1853,n118,n416);
and (n1854,n1855,n1856);
xor (n1855,n1768,n1853);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n750,n1769);
and (n1859,n46,n416);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1774,n1775);
and (n1865,n25,n416);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
or (n1868,n1869,n1872);
and (n1869,n1870,n1871);
xor (n1870,n1779,n1780);
and (n1871,n137,n416);
and (n1872,n1873,n1874);
xor (n1873,n1870,n1871);
or (n1874,n1875,n1878);
and (n1875,n1876,n1877);
xor (n1876,n1784,n1785);
and (n1877,n187,n416);
and (n1878,n1879,n1880);
xor (n1879,n1876,n1877);
or (n1880,n1881,n1884);
and (n1881,n1882,n1883);
xor (n1882,n1789,n1790);
and (n1883,n75,n416);
and (n1884,n1885,n1886);
xor (n1885,n1882,n1883);
or (n1886,n1887,n1890);
and (n1887,n1888,n1889);
xor (n1888,n1794,n1795);
and (n1889,n70,n416);
and (n1890,n1891,n1892);
xor (n1891,n1888,n1889);
or (n1892,n1893,n1896);
and (n1893,n1894,n1895);
xor (n1894,n1800,n1801);
and (n1895,n83,n416);
and (n1896,n1897,n1898);
xor (n1897,n1894,n1895);
or (n1898,n1899,n1902);
and (n1899,n1900,n1901);
xor (n1900,n1806,n1807);
and (n1901,n101,n416);
and (n1902,n1903,n1904);
xor (n1903,n1900,n1901);
or (n1904,n1905,n1908);
and (n1905,n1906,n1907);
xor (n1906,n1811,n1812);
and (n1907,n157,n416);
and (n1908,n1909,n1910);
xor (n1909,n1906,n1907);
or (n1910,n1911,n1914);
and (n1911,n1912,n1913);
xor (n1912,n1817,n1818);
and (n1913,n236,n416);
and (n1914,n1915,n1916);
xor (n1915,n1912,n1913);
or (n1916,n1917,n1920);
and (n1917,n1918,n1919);
xor (n1918,n1822,n1823);
and (n1919,n325,n416);
and (n1920,n1921,n1922);
xor (n1921,n1918,n1919);
or (n1922,n1923,n1926);
and (n1923,n1924,n1925);
xor (n1924,n1827,n1828);
and (n1925,n384,n416);
and (n1926,n1927,n1928);
xor (n1927,n1924,n1925);
or (n1928,n1929,n1932);
and (n1929,n1930,n1931);
xor (n1930,n1833,n1834);
and (n1931,n447,n416);
and (n1932,n1933,n1934);
xor (n1933,n1930,n1931);
or (n1934,n1935,n1938);
and (n1935,n1936,n1937);
xor (n1936,n1839,n1840);
and (n1937,n575,n416);
and (n1938,n1939,n1940);
xor (n1939,n1936,n1937);
or (n1940,n1941,n1944);
and (n1941,n1942,n1943);
xor (n1942,n1845,n1846);
and (n1943,n608,n416);
and (n1944,n1945,n1946);
xor (n1945,n1942,n1943);
and (n1946,n1947,n1599);
xor (n1947,n1850,n1851);
and (n1948,n1949,n1950);
xor (n1949,n1766,n492);
or (n1950,n1951,n1954);
and (n1951,n1952,n1953);
xor (n1952,n1855,n1856);
and (n1953,n46,n289);
and (n1954,n1955,n1956);
xor (n1955,n1952,n1953);
or (n1956,n1957,n1959);
and (n1957,n1958,n699);
xor (n1958,n1861,n1862);
and (n1959,n1960,n1961);
xor (n1960,n1958,n699);
or (n1961,n1962,n1964);
and (n1962,n1963,n784);
xor (n1963,n1867,n1868);
and (n1964,n1965,n1966);
xor (n1965,n1963,n784);
or (n1966,n1967,n1969);
and (n1967,n1968,n922);
xor (n1968,n1873,n1874);
and (n1969,n1970,n1971);
xor (n1970,n1968,n922);
or (n1971,n1972,n1974);
and (n1972,n1973,n917);
xor (n1973,n1879,n1880);
and (n1974,n1975,n1976);
xor (n1975,n1973,n917);
or (n1976,n1977,n1979);
and (n1977,n1978,n1067);
xor (n1978,n1885,n1886);
and (n1979,n1980,n1981);
xor (n1980,n1978,n1067);
or (n1981,n1982,n1984);
and (n1982,n1983,n1136);
xor (n1983,n1891,n1892);
and (n1984,n1985,n1986);
xor (n1985,n1983,n1136);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1897,n1898);
and (n1989,n101,n289);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1996);
and (n1993,n1994,n1995);
xor (n1994,n1903,n1904);
and (n1995,n157,n289);
and (n1996,n1997,n1998);
xor (n1997,n1994,n1995);
or (n1998,n1999,n2002);
and (n1999,n2000,n2001);
xor (n2000,n1909,n1910);
and (n2001,n236,n289);
and (n2002,n2003,n2004);
xor (n2003,n2000,n2001);
or (n2004,n2005,n2008);
and (n2005,n2006,n2007);
xor (n2006,n1915,n1916);
and (n2007,n325,n289);
and (n2008,n2009,n2010);
xor (n2009,n2006,n2007);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1921,n1922);
and (n2013,n384,n289);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
or (n2016,n2017,n2019);
and (n2017,n2018,n1438);
xor (n2018,n1927,n1928);
and (n2019,n2020,n2021);
xor (n2020,n2018,n1438);
or (n2021,n2022,n2025);
and (n2022,n2023,n2024);
xor (n2023,n1933,n1934);
and (n2024,n575,n289);
and (n2025,n2026,n2027);
xor (n2026,n2023,n2024);
or (n2027,n2028,n2030);
and (n2028,n2029,n1572);
xor (n2029,n1939,n1940);
and (n2030,n2031,n2032);
xor (n2031,n2029,n1572);
and (n2032,n2033,n2034);
xor (n2033,n1945,n1946);
and (n2034,n668,n289);
and (n2035,n118,n287);
and (n2036,n2037,n2038);
xor (n2037,n1764,n2035);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
xor (n2040,n1949,n1950);
and (n2041,n46,n287);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
or (n2044,n2045,n2048);
and (n2045,n2046,n2047);
xor (n2046,n1955,n1956);
and (n2047,n25,n287);
and (n2048,n2049,n2050);
xor (n2049,n2046,n2047);
or (n2050,n2051,n2054);
and (n2051,n2052,n2053);
xor (n2052,n1960,n1961);
and (n2053,n137,n287);
and (n2054,n2055,n2056);
xor (n2055,n2052,n2053);
or (n2056,n2057,n2060);
and (n2057,n2058,n2059);
xor (n2058,n1965,n1966);
and (n2059,n187,n287);
and (n2060,n2061,n2062);
xor (n2061,n2058,n2059);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
xor (n2064,n1970,n1971);
and (n2065,n75,n287);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n1975,n1976);
and (n2071,n70,n287);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2078);
and (n2075,n2076,n2077);
xor (n2076,n1980,n1981);
and (n2077,n83,n287);
and (n2078,n2079,n2080);
xor (n2079,n2076,n2077);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n1985,n1986);
and (n2083,n101,n287);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n1991,n1992);
and (n2089,n157,n287);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n1997,n1998);
and (n2095,n236,n287);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2003,n2004);
and (n2101,n325,n287);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2009,n2010);
and (n2107,n384,n287);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2015,n2016);
and (n2113,n447,n287);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2020,n2021);
and (n2119,n575,n287);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n2026,n2027);
and (n2125,n608,n287);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
and (n2128,n2129,n1528);
xor (n2129,n2031,n2032);
and (n2130,n2131,n2132);
xor (n2131,n1762,n333);
or (n2132,n2133,n2136);
and (n2133,n2134,n2135);
xor (n2134,n2037,n2038);
and (n2135,n46,n114);
and (n2136,n2137,n2138);
xor (n2137,n2134,n2135);
or (n2138,n2139,n2141);
and (n2139,n2140,n570);
xor (n2140,n2043,n2044);
and (n2141,n2142,n2143);
xor (n2142,n2140,n570);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2049,n2050);
and (n2146,n137,n114);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2055,n2056);
and (n2152,n187,n114);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2158);
and (n2156,n2157,n795);
xor (n2157,n2061,n2062);
and (n2158,n2159,n2160);
xor (n2159,n2157,n795);
or (n2160,n2161,n2164);
and (n2161,n2162,n2163);
xor (n2162,n2067,n2068);
and (n2163,n70,n114);
and (n2164,n2165,n2166);
xor (n2165,n2162,n2163);
or (n2166,n2167,n2170);
and (n2167,n2168,n2169);
xor (n2168,n2073,n2074);
and (n2169,n83,n114);
and (n2170,n2171,n2172);
xor (n2171,n2168,n2169);
or (n2172,n2173,n2176);
and (n2173,n2174,n2175);
xor (n2174,n2079,n2080);
and (n2175,n101,n114);
and (n2176,n2177,n2178);
xor (n2177,n2174,n2175);
or (n2178,n2179,n2182);
and (n2179,n2180,n2181);
xor (n2180,n2085,n2086);
and (n2181,n157,n114);
and (n2182,n2183,n2184);
xor (n2183,n2180,n2181);
or (n2184,n2185,n2188);
and (n2185,n2186,n2187);
xor (n2186,n2091,n2092);
and (n2187,n236,n114);
and (n2188,n2189,n2190);
xor (n2189,n2186,n2187);
or (n2190,n2191,n2194);
and (n2191,n2192,n2193);
xor (n2192,n2097,n2098);
and (n2193,n325,n114);
and (n2194,n2195,n2196);
xor (n2195,n2192,n2193);
or (n2196,n2197,n2200);
and (n2197,n2198,n2199);
xor (n2198,n2103,n2104);
and (n2199,n384,n114);
and (n2200,n2201,n2202);
xor (n2201,n2198,n2199);
or (n2202,n2203,n2206);
and (n2203,n2204,n2205);
xor (n2204,n2109,n2110);
and (n2205,n447,n114);
and (n2206,n2207,n2208);
xor (n2207,n2204,n2205);
or (n2208,n2209,n2212);
and (n2209,n2210,n2211);
xor (n2210,n2115,n2116);
and (n2211,n575,n114);
and (n2212,n2213,n2214);
xor (n2213,n2210,n2211);
or (n2214,n2215,n2217);
and (n2215,n2216,n1520);
xor (n2216,n2121,n2122);
and (n2217,n2218,n2219);
xor (n2218,n2216,n1520);
and (n2219,n2220,n2221);
xor (n2220,n2127,n2128);
and (n2221,n668,n114);
and (n2222,n118,n108);
and (n2223,n2224,n2225);
xor (n2224,n1760,n2222);
or (n2225,n2226,n2229);
and (n2226,n2227,n2228);
xor (n2227,n2131,n2132);
and (n2228,n46,n108);
and (n2229,n2230,n2231);
xor (n2230,n2227,n2228);
or (n2231,n2232,n2235);
and (n2232,n2233,n2234);
xor (n2233,n2137,n2138);
and (n2234,n25,n108);
and (n2235,n2236,n2237);
xor (n2236,n2233,n2234);
or (n2237,n2238,n2241);
and (n2238,n2239,n2240);
xor (n2239,n2142,n2143);
and (n2240,n137,n108);
and (n2241,n2242,n2243);
xor (n2242,n2239,n2240);
or (n2243,n2244,n2247);
and (n2244,n2245,n2246);
xor (n2245,n2148,n2149);
and (n2246,n187,n108);
and (n2247,n2248,n2249);
xor (n2248,n2245,n2246);
or (n2249,n2250,n2253);
and (n2250,n2251,n2252);
xor (n2251,n2154,n2155);
and (n2252,n75,n108);
and (n2253,n2254,n2255);
xor (n2254,n2251,n2252);
or (n2255,n2256,n2259);
and (n2256,n2257,n2258);
xor (n2257,n2159,n2160);
and (n2258,n70,n108);
and (n2259,n2260,n2261);
xor (n2260,n2257,n2258);
or (n2261,n2262,n2265);
and (n2262,n2263,n2264);
xor (n2263,n2165,n2166);
and (n2264,n83,n108);
and (n2265,n2266,n2267);
xor (n2266,n2263,n2264);
or (n2267,n2268,n2271);
and (n2268,n2269,n2270);
xor (n2269,n2171,n2172);
and (n2270,n101,n108);
and (n2271,n2272,n2273);
xor (n2272,n2269,n2270);
or (n2273,n2274,n2277);
and (n2274,n2275,n2276);
xor (n2275,n2177,n2178);
and (n2276,n157,n108);
and (n2277,n2278,n2279);
xor (n2278,n2275,n2276);
or (n2279,n2280,n2283);
and (n2280,n2281,n2282);
xor (n2281,n2183,n2184);
and (n2282,n236,n108);
and (n2283,n2284,n2285);
xor (n2284,n2281,n2282);
or (n2285,n2286,n2289);
and (n2286,n2287,n2288);
xor (n2287,n2189,n2190);
and (n2288,n325,n108);
and (n2289,n2290,n2291);
xor (n2290,n2287,n2288);
or (n2291,n2292,n2295);
and (n2292,n2293,n2294);
xor (n2293,n2195,n2196);
and (n2294,n384,n108);
and (n2295,n2296,n2297);
xor (n2296,n2293,n2294);
or (n2297,n2298,n2301);
and (n2298,n2299,n2300);
xor (n2299,n2201,n2202);
and (n2300,n447,n108);
and (n2301,n2302,n2303);
xor (n2302,n2299,n2300);
or (n2303,n2304,n2307);
and (n2304,n2305,n2306);
xor (n2305,n2207,n2208);
and (n2306,n575,n108);
and (n2307,n2308,n2309);
xor (n2308,n2305,n2306);
or (n2309,n2310,n2313);
and (n2310,n2311,n2312);
xor (n2311,n2213,n2214);
and (n2312,n608,n108);
and (n2313,n2314,n2315);
xor (n2314,n2311,n2312);
and (n2315,n2316,n1374);
xor (n2316,n2218,n2219);
and (n2317,n118,n34);
and (n2318,n2319,n2320);
xor (n2319,n1758,n2317);
or (n2320,n2321,n2323);
and (n2321,n2322,n301);
xor (n2322,n2224,n2225);
and (n2323,n2324,n2325);
xor (n2324,n2322,n301);
or (n2325,n2326,n2328);
and (n2326,n2327,n343);
xor (n2327,n2230,n2231);
and (n2328,n2329,n2330);
xor (n2329,n2327,n343);
or (n2330,n2331,n2333);
and (n2331,n2332,n462);
xor (n2332,n2236,n2237);
and (n2333,n2334,n2335);
xor (n2334,n2332,n462);
or (n2335,n2336,n2338);
and (n2336,n2337,n532);
xor (n2337,n2242,n2243);
and (n2338,n2339,n2340);
xor (n2339,n2337,n532);
or (n2340,n2341,n2344);
and (n2341,n2342,n2343);
xor (n2342,n2248,n2249);
and (n2343,n75,n34);
and (n2344,n2345,n2346);
xor (n2345,n2342,n2343);
or (n2346,n2347,n2349);
and (n2347,n2348,n656);
xor (n2348,n2254,n2255);
and (n2349,n2350,n2351);
xor (n2350,n2348,n656);
or (n2351,n2352,n2355);
and (n2352,n2353,n2354);
xor (n2353,n2260,n2261);
and (n2354,n83,n34);
and (n2355,n2356,n2357);
xor (n2356,n2353,n2354);
or (n2357,n2358,n2360);
and (n2358,n2359,n947);
xor (n2359,n2266,n2267);
and (n2360,n2361,n2362);
xor (n2361,n2359,n947);
or (n2362,n2363,n2365);
and (n2363,n2364,n983);
xor (n2364,n2272,n2273);
and (n2365,n2366,n2367);
xor (n2366,n2364,n983);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2278,n2279);
and (n2370,n236,n34);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2284,n2285);
and (n2376,n325,n34);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2290,n2291);
and (n2382,n384,n34);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2388);
and (n2386,n2387,n1321);
xor (n2387,n2296,n2297);
and (n2388,n2389,n2390);
xor (n2389,n2387,n1321);
or (n2390,n2391,n2393);
and (n2391,n2392,n1306);
xor (n2392,n2302,n2303);
and (n2393,n2394,n2395);
xor (n2394,n2392,n1306);
or (n2395,n2396,n2399);
and (n2396,n2397,n2398);
xor (n2397,n2308,n2309);
and (n2398,n608,n34);
and (n2399,n2400,n2401);
xor (n2400,n2397,n2398);
and (n2401,n2402,n2403);
xor (n2402,n2314,n2315);
and (n2403,n668,n34);
and (n2404,n118,n35);
and (n2405,n2406,n2407);
xor (n2406,n1756,n2404);
or (n2407,n2408,n2411);
and (n2408,n2409,n2410);
xor (n2409,n2319,n2320);
and (n2410,n46,n35);
and (n2411,n2412,n2413);
xor (n2412,n2409,n2410);
or (n2413,n2414,n2417);
and (n2414,n2415,n2416);
xor (n2415,n2324,n2325);
and (n2416,n25,n35);
and (n2417,n2418,n2419);
xor (n2418,n2415,n2416);
or (n2419,n2420,n2423);
and (n2420,n2421,n2422);
xor (n2421,n2329,n2330);
and (n2422,n137,n35);
and (n2423,n2424,n2425);
xor (n2424,n2421,n2422);
or (n2425,n2426,n2429);
and (n2426,n2427,n2428);
xor (n2427,n2334,n2335);
and (n2428,n187,n35);
and (n2429,n2430,n2431);
xor (n2430,n2427,n2428);
or (n2431,n2432,n2435);
and (n2432,n2433,n2434);
xor (n2433,n2339,n2340);
and (n2434,n75,n35);
and (n2435,n2436,n2437);
xor (n2436,n2433,n2434);
or (n2437,n2438,n2441);
and (n2438,n2439,n2440);
xor (n2439,n2345,n2346);
and (n2440,n70,n35);
and (n2441,n2442,n2443);
xor (n2442,n2439,n2440);
or (n2443,n2444,n2447);
and (n2444,n2445,n2446);
xor (n2445,n2350,n2351);
and (n2446,n83,n35);
and (n2447,n2448,n2449);
xor (n2448,n2445,n2446);
or (n2449,n2450,n2453);
and (n2450,n2451,n2452);
xor (n2451,n2356,n2357);
and (n2452,n101,n35);
and (n2453,n2454,n2455);
xor (n2454,n2451,n2452);
or (n2455,n2456,n2459);
and (n2456,n2457,n2458);
xor (n2457,n2361,n2362);
and (n2458,n157,n35);
and (n2459,n2460,n2461);
xor (n2460,n2457,n2458);
or (n2461,n2462,n2465);
and (n2462,n2463,n2464);
xor (n2463,n2366,n2367);
and (n2464,n236,n35);
and (n2465,n2466,n2467);
xor (n2466,n2463,n2464);
or (n2467,n2468,n2471);
and (n2468,n2469,n2470);
xor (n2469,n2372,n2373);
and (n2470,n325,n35);
and (n2471,n2472,n2473);
xor (n2472,n2469,n2470);
or (n2473,n2474,n2477);
and (n2474,n2475,n2476);
xor (n2475,n2378,n2379);
and (n2476,n384,n35);
and (n2477,n2478,n2479);
xor (n2478,n2475,n2476);
or (n2479,n2480,n2483);
and (n2480,n2481,n2482);
xor (n2481,n2384,n2385);
and (n2482,n447,n35);
and (n2483,n2484,n2485);
xor (n2484,n2481,n2482);
or (n2485,n2486,n2489);
and (n2486,n2487,n2488);
xor (n2487,n2389,n2390);
and (n2488,n575,n35);
and (n2489,n2490,n2491);
xor (n2490,n2487,n2488);
or (n2491,n2492,n2495);
and (n2492,n2493,n2494);
xor (n2493,n2394,n2395);
and (n2494,n608,n35);
and (n2495,n2496,n2497);
xor (n2496,n2493,n2494);
and (n2497,n2498,n1272);
xor (n2498,n2400,n2401);
and (n2499,n118,n27);
or (n2500,n2501,n2504);
and (n2501,n2502,n2503);
xor (n2502,n2406,n2407);
and (n2503,n46,n27);
and (n2504,n2505,n2506);
xor (n2505,n2502,n2503);
or (n2506,n2507,n2509);
and (n2507,n2508,n28);
xor (n2508,n2412,n2413);
and (n2509,n2510,n2511);
xor (n2510,n2508,n28);
or (n2511,n2512,n2515);
and (n2512,n2513,n2514);
xor (n2513,n2418,n2419);
and (n2514,n137,n27);
and (n2515,n2516,n2517);
xor (n2516,n2513,n2514);
or (n2517,n2518,n2520);
and (n2518,n2519,n372);
xor (n2519,n2424,n2425);
and (n2520,n2521,n2522);
xor (n2521,n2519,n372);
or (n2522,n2523,n2525);
and (n2523,n2524,n438);
xor (n2524,n2430,n2431);
and (n2525,n2526,n2527);
xor (n2526,n2524,n438);
or (n2527,n2528,n2530);
and (n2528,n2529,n582);
xor (n2529,n2436,n2437);
and (n2530,n2531,n2532);
xor (n2531,n2529,n582);
or (n2532,n2533,n2535);
and (n2533,n2534,n625);
xor (n2534,n2442,n2443);
and (n2535,n2536,n2537);
xor (n2536,n2534,n625);
or (n2537,n2538,n2540);
and (n2538,n2539,n706);
xor (n2539,n2448,n2449);
and (n2540,n2541,n2542);
xor (n2541,n2539,n706);
or (n2542,n2543,n2545);
and (n2543,n2544,n834);
xor (n2544,n2454,n2455);
and (n2545,n2546,n2547);
xor (n2546,n2544,n834);
or (n2547,n2548,n2550);
and (n2548,n2549,n957);
xor (n2549,n2460,n2461);
and (n2550,n2551,n2552);
xor (n2551,n2549,n957);
or (n2552,n2553,n2556);
and (n2553,n2554,n2555);
xor (n2554,n2466,n2467);
and (n2555,n325,n27);
and (n2556,n2557,n2558);
xor (n2557,n2554,n2555);
or (n2558,n2559,n2561);
and (n2559,n2560,n1081);
xor (n2560,n2472,n2473);
and (n2561,n2562,n2563);
xor (n2562,n2560,n1081);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2478,n2479);
and (n2566,n447,n27);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2484,n2485);
and (n2572,n575,n27);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
or (n2575,n2576,n2578);
and (n2576,n2577,n1234);
xor (n2577,n2490,n2491);
and (n2578,n2579,n2580);
xor (n2579,n2577,n1234);
and (n2580,n2581,n2582);
xor (n2581,n2496,n2497);
and (n2582,n668,n27);
and (n2583,n46,n145);
or (n2584,n2585,n2588);
and (n2585,n2586,n2587);
xor (n2586,n2505,n2506);
and (n2587,n25,n145);
and (n2588,n2589,n2590);
xor (n2589,n2586,n2587);
or (n2590,n2591,n2594);
and (n2591,n2592,n2593);
xor (n2592,n2510,n2511);
and (n2593,n137,n145);
and (n2594,n2595,n2596);
xor (n2595,n2592,n2593);
or (n2596,n2597,n2600);
and (n2597,n2598,n2599);
xor (n2598,n2516,n2517);
and (n2599,n187,n145);
and (n2600,n2601,n2602);
xor (n2601,n2598,n2599);
or (n2602,n2603,n2606);
and (n2603,n2604,n2605);
xor (n2604,n2521,n2522);
and (n2605,n75,n145);
and (n2606,n2607,n2608);
xor (n2607,n2604,n2605);
or (n2608,n2609,n2612);
and (n2609,n2610,n2611);
xor (n2610,n2526,n2527);
and (n2611,n70,n145);
and (n2612,n2613,n2614);
xor (n2613,n2610,n2611);
or (n2614,n2615,n2618);
and (n2615,n2616,n2617);
xor (n2616,n2531,n2532);
and (n2617,n83,n145);
and (n2618,n2619,n2620);
xor (n2619,n2616,n2617);
or (n2620,n2621,n2624);
and (n2621,n2622,n2623);
xor (n2622,n2536,n2537);
and (n2623,n101,n145);
and (n2624,n2625,n2626);
xor (n2625,n2622,n2623);
or (n2626,n2627,n2630);
and (n2627,n2628,n2629);
xor (n2628,n2541,n2542);
and (n2629,n157,n145);
and (n2630,n2631,n2632);
xor (n2631,n2628,n2629);
or (n2632,n2633,n2636);
and (n2633,n2634,n2635);
xor (n2634,n2546,n2547);
and (n2635,n236,n145);
and (n2636,n2637,n2638);
xor (n2637,n2634,n2635);
or (n2638,n2639,n2642);
and (n2639,n2640,n2641);
xor (n2640,n2551,n2552);
and (n2641,n325,n145);
and (n2642,n2643,n2644);
xor (n2643,n2640,n2641);
or (n2644,n2645,n2648);
and (n2645,n2646,n2647);
xor (n2646,n2557,n2558);
and (n2647,n384,n145);
and (n2648,n2649,n2650);
xor (n2649,n2646,n2647);
or (n2650,n2651,n2654);
and (n2651,n2652,n2653);
xor (n2652,n2562,n2563);
and (n2653,n447,n145);
and (n2654,n2655,n2656);
xor (n2655,n2652,n2653);
or (n2656,n2657,n2660);
and (n2657,n2658,n2659);
xor (n2658,n2568,n2569);
and (n2659,n575,n145);
and (n2660,n2661,n2662);
xor (n2661,n2658,n2659);
or (n2662,n2663,n2666);
and (n2663,n2664,n2665);
xor (n2664,n2574,n2575);
and (n2665,n608,n145);
and (n2666,n2667,n2668);
xor (n2667,n2664,n2665);
and (n2668,n2669,n1476);
xor (n2669,n2579,n2580);
or (n2670,n2671,n2673);
and (n2671,n2672,n138);
xor (n2672,n2589,n2590);
and (n2673,n2674,n2675);
xor (n2674,n2672,n138);
or (n2675,n2676,n2679);
and (n2676,n2677,n2678);
xor (n2677,n2595,n2596);
and (n2678,n187,n58);
and (n2679,n2680,n2681);
xor (n2680,n2677,n2678);
or (n2681,n2682,n2684);
and (n2682,n2683,n309);
xor (n2683,n2601,n2602);
and (n2684,n2685,n2686);
xor (n2685,n2683,n309);
or (n2686,n2687,n2689);
and (n2687,n2688,n350);
xor (n2688,n2607,n2608);
and (n2689,n2690,n2691);
xor (n2690,n2688,n350);
or (n2691,n2692,n2694);
and (n2692,n2693,n454);
xor (n2693,n2613,n2614);
and (n2694,n2695,n2696);
xor (n2695,n2693,n454);
or (n2696,n2697,n2700);
and (n2697,n2698,n2699);
xor (n2698,n2619,n2620);
and (n2699,n101,n58);
and (n2700,n2701,n2702);
xor (n2701,n2698,n2699);
or (n2702,n2703,n2706);
and (n2703,n2704,n2705);
xor (n2704,n2625,n2626);
and (n2705,n157,n58);
and (n2706,n2707,n2708);
xor (n2707,n2704,n2705);
or (n2708,n2709,n2712);
and (n2709,n2710,n2711);
xor (n2710,n2631,n2632);
and (n2711,n236,n58);
and (n2712,n2713,n2714);
xor (n2713,n2710,n2711);
or (n2714,n2715,n2718);
and (n2715,n2716,n2717);
xor (n2716,n2637,n2638);
and (n2717,n325,n58);
and (n2718,n2719,n2720);
xor (n2719,n2716,n2717);
or (n2720,n2721,n2724);
and (n2721,n2722,n2723);
xor (n2722,n2643,n2644);
and (n2723,n384,n58);
and (n2724,n2725,n2726);
xor (n2725,n2722,n2723);
or (n2726,n2727,n2730);
and (n2727,n2728,n2729);
xor (n2728,n2649,n2650);
and (n2729,n447,n58);
and (n2730,n2731,n2732);
xor (n2731,n2728,n2729);
or (n2732,n2733,n2735);
and (n2733,n2734,n1098);
xor (n2734,n2655,n2656);
and (n2735,n2736,n2737);
xor (n2736,n2734,n1098);
or (n2737,n2738,n2741);
and (n2738,n2739,n2740);
xor (n2739,n2661,n2662);
and (n2740,n608,n58);
and (n2741,n2742,n2743);
xor (n2742,n2739,n2740);
and (n2743,n2744,n2745);
xor (n2744,n2667,n2668);
and (n2745,n668,n58);
and (n2746,n137,n57);
or (n2747,n2748,n2751);
and (n2748,n2749,n2750);
xor (n2749,n2674,n2675);
and (n2750,n187,n57);
and (n2751,n2752,n2753);
xor (n2752,n2749,n2750);
or (n2753,n2754,n2757);
and (n2754,n2755,n2756);
xor (n2755,n2680,n2681);
and (n2756,n75,n57);
and (n2757,n2758,n2759);
xor (n2758,n2755,n2756);
or (n2759,n2760,n2763);
and (n2760,n2761,n2762);
xor (n2761,n2685,n2686);
and (n2762,n70,n57);
and (n2763,n2764,n2765);
xor (n2764,n2761,n2762);
or (n2765,n2766,n2769);
and (n2766,n2767,n2768);
xor (n2767,n2690,n2691);
and (n2768,n83,n57);
and (n2769,n2770,n2771);
xor (n2770,n2767,n2768);
or (n2771,n2772,n2775);
and (n2772,n2773,n2774);
xor (n2773,n2695,n2696);
and (n2774,n101,n57);
and (n2775,n2776,n2777);
xor (n2776,n2773,n2774);
or (n2777,n2778,n2781);
and (n2778,n2779,n2780);
xor (n2779,n2701,n2702);
and (n2780,n157,n57);
and (n2781,n2782,n2783);
xor (n2782,n2779,n2780);
or (n2783,n2784,n2787);
and (n2784,n2785,n2786);
xor (n2785,n2707,n2708);
and (n2786,n236,n57);
and (n2787,n2788,n2789);
xor (n2788,n2785,n2786);
or (n2789,n2790,n2793);
and (n2790,n2791,n2792);
xor (n2791,n2713,n2714);
and (n2792,n325,n57);
and (n2793,n2794,n2795);
xor (n2794,n2791,n2792);
or (n2795,n2796,n2799);
and (n2796,n2797,n2798);
xor (n2797,n2719,n2720);
and (n2798,n384,n57);
and (n2799,n2800,n2801);
xor (n2800,n2797,n2798);
or (n2801,n2802,n2805);
and (n2802,n2803,n2804);
xor (n2803,n2725,n2726);
and (n2804,n447,n57);
and (n2805,n2806,n2807);
xor (n2806,n2803,n2804);
or (n2807,n2808,n2811);
and (n2808,n2809,n2810);
xor (n2809,n2731,n2732);
and (n2810,n575,n57);
and (n2811,n2812,n2813);
xor (n2812,n2809,n2810);
or (n2813,n2814,n2817);
and (n2814,n2815,n2816);
xor (n2815,n2736,n2737);
and (n2816,n608,n57);
and (n2817,n2818,n2819);
xor (n2818,n2815,n2816);
and (n2819,n2820,n2821);
xor (n2820,n2742,n2743);
not (n2821,n1045);
and (n2822,n187,n64);
or (n2823,n2824,n2827);
and (n2824,n2825,n2826);
xor (n2825,n2752,n2753);
and (n2826,n75,n64);
and (n2827,n2828,n2829);
xor (n2828,n2825,n2826);
or (n2829,n2830,n2832);
and (n2830,n2831,n71);
xor (n2831,n2758,n2759);
and (n2832,n2833,n2834);
xor (n2833,n2831,n71);
or (n2834,n2835,n2838);
and (n2835,n2836,n2837);
xor (n2836,n2764,n2765);
and (n2837,n83,n64);
and (n2838,n2839,n2840);
xor (n2839,n2836,n2837);
or (n2840,n2841,n2843);
and (n2841,n2842,n358);
xor (n2842,n2770,n2771);
and (n2843,n2844,n2845);
xor (n2844,n2842,n358);
or (n2845,n2846,n2848);
and (n2846,n2847,n478);
xor (n2847,n2776,n2777);
and (n2848,n2849,n2850);
xor (n2849,n2847,n478);
or (n2850,n2851,n2854);
and (n2851,n2852,n2853);
xor (n2852,n2782,n2783);
and (n2853,n236,n64);
and (n2854,n2855,n2856);
xor (n2855,n2852,n2853);
or (n2856,n2857,n2860);
and (n2857,n2858,n2859);
xor (n2858,n2788,n2789);
and (n2859,n325,n64);
and (n2860,n2861,n2862);
xor (n2861,n2858,n2859);
or (n2862,n2863,n2866);
and (n2863,n2864,n2865);
xor (n2864,n2794,n2795);
and (n2865,n384,n64);
and (n2866,n2867,n2868);
xor (n2867,n2864,n2865);
or (n2868,n2869,n2872);
and (n2869,n2870,n2871);
xor (n2870,n2800,n2801);
and (n2871,n447,n64);
and (n2872,n2873,n2874);
xor (n2873,n2870,n2871);
or (n2874,n2875,n2878);
and (n2875,n2876,n2877);
xor (n2876,n2806,n2807);
and (n2877,n575,n64);
and (n2878,n2879,n2880);
xor (n2879,n2876,n2877);
or (n2880,n2881,n2884);
and (n2881,n2882,n2883);
xor (n2882,n2812,n2813);
and (n2883,n608,n64);
and (n2884,n2885,n2886);
xor (n2885,n2882,n2883);
and (n2886,n2887,n2888);
xor (n2887,n2818,n2819);
and (n2888,n668,n64);
and (n2889,n75,n91);
or (n2890,n2891,n2894);
and (n2891,n2892,n2893);
xor (n2892,n2828,n2829);
and (n2893,n70,n91);
and (n2894,n2895,n2896);
xor (n2895,n2892,n2893);
or (n2896,n2897,n2900);
and (n2897,n2898,n2899);
xor (n2898,n2833,n2834);
and (n2899,n83,n91);
and (n2900,n2901,n2902);
xor (n2901,n2898,n2899);
or (n2902,n2903,n2906);
and (n2903,n2904,n2905);
xor (n2904,n2839,n2840);
and (n2905,n101,n91);
and (n2906,n2907,n2908);
xor (n2907,n2904,n2905);
or (n2908,n2909,n2912);
and (n2909,n2910,n2911);
xor (n2910,n2844,n2845);
and (n2911,n157,n91);
and (n2912,n2913,n2914);
xor (n2913,n2910,n2911);
or (n2914,n2915,n2918);
and (n2915,n2916,n2917);
xor (n2916,n2849,n2850);
and (n2917,n236,n91);
and (n2918,n2919,n2920);
xor (n2919,n2916,n2917);
or (n2920,n2921,n2924);
and (n2921,n2922,n2923);
xor (n2922,n2855,n2856);
and (n2923,n325,n91);
and (n2924,n2925,n2926);
xor (n2925,n2922,n2923);
or (n2926,n2927,n2930);
and (n2927,n2928,n2929);
xor (n2928,n2861,n2862);
and (n2929,n384,n91);
and (n2930,n2931,n2932);
xor (n2931,n2928,n2929);
or (n2932,n2933,n2936);
and (n2933,n2934,n2935);
xor (n2934,n2867,n2868);
and (n2935,n447,n91);
and (n2936,n2937,n2938);
xor (n2937,n2934,n2935);
or (n2938,n2939,n2942);
and (n2939,n2940,n2941);
xor (n2940,n2873,n2874);
and (n2941,n575,n91);
and (n2942,n2943,n2944);
xor (n2943,n2940,n2941);
or (n2944,n2945,n2948);
and (n2945,n2946,n2947);
xor (n2946,n2879,n2880);
and (n2947,n608,n91);
and (n2948,n2949,n2950);
xor (n2949,n2946,n2947);
and (n2950,n2951,n2952);
xor (n2951,n2885,n2886);
not (n2952,n891);
or (n2953,n2954,n2956);
and (n2954,n2955,n82);
xor (n2955,n2895,n2896);
and (n2956,n2957,n2958);
xor (n2957,n2955,n82);
or (n2958,n2959,n2962);
and (n2959,n2960,n2961);
xor (n2960,n2901,n2902);
and (n2961,n101,n84);
and (n2962,n2963,n2964);
xor (n2963,n2960,n2961);
or (n2964,n2965,n2967);
and (n2965,n2966,n277);
xor (n2966,n2907,n2908);
and (n2967,n2968,n2969);
xor (n2968,n2966,n277);
or (n2969,n2970,n2972);
and (n2970,n2971,n379);
xor (n2971,n2913,n2914);
and (n2972,n2973,n2974);
xor (n2973,n2971,n379);
or (n2974,n2975,n2977);
and (n2975,n2976,n485);
xor (n2976,n2919,n2920);
and (n2977,n2978,n2979);
xor (n2978,n2976,n485);
or (n2979,n2980,n2982);
and (n2980,n2981,n521);
xor (n2981,n2925,n2926);
and (n2982,n2983,n2984);
xor (n2983,n2981,n521);
or (n2984,n2985,n2988);
and (n2985,n2986,n2987);
xor (n2986,n2931,n2932);
and (n2987,n447,n84);
and (n2988,n2989,n2990);
xor (n2989,n2986,n2987);
or (n2990,n2991,n2994);
and (n2991,n2992,n2993);
xor (n2992,n2937,n2938);
and (n2993,n575,n84);
and (n2994,n2995,n2996);
xor (n2995,n2992,n2993);
or (n2996,n2997,n2999);
and (n2997,n2998,n820);
xor (n2998,n2943,n2944);
and (n2999,n3000,n3001);
xor (n3000,n2998,n820);
and (n3001,n3002,n3003);
xor (n3002,n2949,n2950);
and (n3003,n668,n84);
and (n3004,n83,n162);
or (n3005,n3006,n3009);
and (n3006,n3007,n3008);
xor (n3007,n2957,n2958);
and (n3008,n101,n162);
and (n3009,n3010,n3011);
xor (n3010,n3007,n3008);
or (n3011,n3012,n3015);
and (n3012,n3013,n3014);
xor (n3013,n2963,n2964);
and (n3014,n157,n162);
and (n3015,n3016,n3017);
xor (n3016,n3013,n3014);
or (n3017,n3018,n3021);
and (n3018,n3019,n3020);
xor (n3019,n2968,n2969);
and (n3020,n236,n162);
and (n3021,n3022,n3023);
xor (n3022,n3019,n3020);
or (n3023,n3024,n3027);
and (n3024,n3025,n3026);
xor (n3025,n2973,n2974);
and (n3026,n325,n162);
and (n3027,n3028,n3029);
xor (n3028,n3025,n3026);
or (n3029,n3030,n3033);
and (n3030,n3031,n3032);
xor (n3031,n2978,n2979);
and (n3032,n384,n162);
and (n3033,n3034,n3035);
xor (n3034,n3031,n3032);
or (n3035,n3036,n3039);
and (n3036,n3037,n3038);
xor (n3037,n2983,n2984);
and (n3038,n447,n162);
and (n3039,n3040,n3041);
xor (n3040,n3037,n3038);
or (n3041,n3042,n3045);
and (n3042,n3043,n3044);
xor (n3043,n2989,n2990);
and (n3044,n575,n162);
and (n3045,n3046,n3047);
xor (n3046,n3043,n3044);
or (n3047,n3048,n3051);
and (n3048,n3049,n3050);
xor (n3049,n2995,n2996);
and (n3050,n608,n162);
and (n3051,n3052,n3053);
xor (n3052,n3049,n3050);
and (n3053,n3054,n3055);
xor (n3054,n3000,n3001);
and (n3055,n668,n162);
endmodule
