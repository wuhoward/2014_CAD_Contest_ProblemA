module top (out,n17,n18,n22,n31,n36,n40,n46,n56,n57
        ,n61,n65,n74,n81,n87,n103,n130,n131,n203,n226
        ,n232,n242,n244,n250,n262,n310,n334,n391,n412,n413
        ,n443,n715,n748,n808,n885);
output out;
input n17;
input n18;
input n22;
input n31;
input n36;
input n40;
input n46;
input n56;
input n57;
input n61;
input n65;
input n74;
input n81;
input n87;
input n103;
input n130;
input n131;
input n203;
input n226;
input n232;
input n242;
input n244;
input n250;
input n262;
input n310;
input n334;
input n391;
input n412;
input n413;
input n443;
input n715;
input n748;
input n808;
input n885;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n243;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
xor (out,n0,n1893);
nor (n0,n1,n1890);
and (n1,n2,n181);
nor (n2,n3,n180);
not (n3,n4);
nand (n4,n5,n155);
or (n5,n6,n154);
and (n6,n7,n118);
xor (n7,n8,n66);
xor (n8,n9,n49);
xor (n9,n10,n25);
nand (n10,n11,n22);
or (n11,n12,n14);
and (n12,n13,n20);
not (n13,n14);
nand (n14,n15,n19);
or (n15,n16,n18);
not (n16,n17);
nand (n19,n18,n16);
nand (n20,n21,n23);
nand (n21,n22,n16);
nand (n23,n17,n24);
not (n24,n22);
nand (n25,n26,n43);
or (n26,n27,n38);
nand (n27,n28,n33);
nor (n28,n29,n32);
and (n29,n30,n22);
not (n30,n31);
and (n32,n31,n24);
nor (n33,n34,n37);
and (n34,n30,n35);
not (n35,n36);
and (n37,n31,n36);
nor (n38,n39,n41);
and (n39,n35,n40);
and (n41,n36,n42);
not (n42,n40);
or (n43,n28,n44);
nor (n44,n45,n47);
and (n45,n35,n46);
and (n47,n36,n48);
not (n48,n46);
nand (n49,n50,n62);
or (n50,n51,n60);
not (n51,n52);
nor (n52,n53,n59);
nand (n53,n54,n58);
or (n54,n55,n57);
not (n55,n56);
nand (n58,n57,n55);
not (n59,n57);
not (n60,n61);
or (n62,n63,n64);
not (n63,n53);
not (n64,n65);
xor (n66,n67,n97);
xor (n67,n68,n90);
nand (n68,n69,n84);
or (n69,n70,n79);
nand (n70,n71,n76);
not (n71,n72);
nand (n72,n73,n75);
or (n73,n35,n74);
nand (n75,n74,n35);
nand (n76,n77,n78);
or (n77,n74,n55);
nand (n78,n55,n74);
nor (n79,n80,n82);
and (n80,n55,n81);
and (n82,n56,n83);
not (n83,n81);
or (n84,n71,n85);
nor (n85,n86,n88);
and (n86,n55,n87);
and (n88,n56,n89);
not (n89,n87);
nand (n90,n91,n96);
or (n91,n92,n93);
not (n92,n12);
nor (n93,n94,n95);
and (n94,n24,n46);
and (n95,n22,n48);
or (n96,n13,n24);
or (n97,n98,n117);
and (n98,n99,n111);
xor (n99,n100,n105);
nand (n100,n101,n104);
or (n101,n102,n51);
not (n102,n103);
nand (n104,n53,n61);
nand (n105,n106,n110);
or (n106,n27,n107);
nor (n107,n108,n109);
and (n108,n35,n87);
and (n109,n36,n89);
or (n110,n28,n38);
nand (n111,n112,n116);
or (n112,n70,n113);
nor (n113,n114,n115);
and (n114,n55,n65);
and (n115,n56,n64);
or (n116,n71,n79);
and (n117,n100,n105);
or (n118,n119,n153);
and (n119,n120,n152);
xor (n120,n121,n122);
not (n121,n90);
or (n122,n123,n151);
and (n123,n124,n145);
xor (n124,n125,n139);
nand (n125,n126,n18);
or (n126,n127,n133);
nand (n127,n128,n132);
or (n128,n129,n131);
not (n129,n130);
nand (n132,n129,n131);
nor (n133,n127,n134);
nor (n134,n135,n137);
and (n135,n136,n131);
not (n136,n18);
and (n137,n18,n138);
not (n138,n131);
nand (n139,n140,n144);
or (n140,n92,n141);
nor (n141,n142,n143);
and (n142,n42,n22);
and (n143,n40,n24);
or (n144,n13,n93);
nand (n145,n146,n150);
or (n146,n70,n147);
nor (n147,n148,n149);
and (n148,n55,n61);
and (n149,n56,n60);
or (n150,n71,n113);
and (n151,n125,n139);
xor (n152,n99,n111);
and (n153,n121,n122);
and (n154,n8,n66);
xor (n155,n156,n177);
xor (n156,n157,n160);
or (n157,n158,n159);
and (n158,n9,n49);
and (n159,n10,n25);
xor (n160,n161,n171);
xor (n161,n162,n168);
nand (n162,n163,n164);
or (n163,n70,n85);
or (n164,n71,n165);
nor (n165,n166,n167);
and (n166,n55,n40);
and (n167,n56,n42);
nand (n168,n169,n170);
or (n169,n51,n64);
or (n170,n63,n83);
nor (n171,n172,n175);
and (n172,n173,n174);
not (n173,n27);
not (n174,n44);
and (n175,n176,n36);
not (n176,n28);
or (n177,n178,n179);
and (n178,n67,n97);
and (n179,n68,n90);
nor (n180,n5,n155);
nand (n181,n182,n1871);
or (n182,n183,n639);
not (n183,n184);
nor (n184,n185,n634);
nand (n185,n186,n621);
and (n186,n187,n593);
nor (n187,n188,n547);
nor (n188,n189,n494);
or (n189,n190,n493);
and (n190,n191,n397);
xor (n191,n192,n303);
xor (n192,n193,n284);
xor (n193,n194,n235);
or (n194,n195,n234);
and (n195,n196,n220);
xor (n196,n197,n209);
nand (n197,n198,n205);
or (n198,n199,n27);
not (n199,n200);
nand (n200,n201,n204);
or (n201,n202,n36);
not (n202,n203);
or (n204,n203,n35);
nand (n205,n176,n206);
nor (n206,n207,n208);
and (n207,n35,n102);
and (n208,n103,n36);
nand (n209,n210,n216);
or (n210,n211,n215);
not (n211,n212);
nand (n212,n213,n214);
or (n213,n81,n136);
nand (n214,n136,n81);
not (n215,n133);
nand (n216,n127,n217);
nor (n217,n218,n219);
and (n218,n89,n136);
and (n219,n87,n18);
nand (n220,n221,n228);
or (n221,n70,n222);
not (n222,n223);
nor (n223,n224,n227);
and (n224,n225,n55);
not (n225,n226);
and (n227,n226,n56);
or (n228,n71,n229);
nor (n229,n230,n233);
and (n230,n231,n56);
not (n231,n232);
and (n233,n232,n55);
and (n234,n197,n209);
or (n235,n236,n283);
and (n236,n237,n273);
xor (n237,n238,n253);
nand (n238,n239,n250);
or (n239,n240,n246);
nand (n240,n241,n245);
or (n241,n242,n243);
not (n243,n244);
nand (n245,n242,n243);
nor (n246,n240,n247);
nor (n247,n248,n251);
and (n248,n249,n250);
not (n249,n242);
and (n251,n242,n252);
not (n252,n250);
nand (n253,n254,n268);
or (n254,n255,n259);
not (n255,n256);
nor (n256,n257,n258);
and (n257,n42,n129);
and (n258,n40,n130);
nand (n259,n260,n264);
nand (n260,n261,n263);
or (n261,n262,n129);
nand (n263,n129,n262);
not (n264,n265);
nand (n265,n266,n267);
or (n266,n252,n262);
nand (n267,n262,n252);
nand (n268,n269,n265);
not (n269,n270);
nor (n270,n271,n272);
and (n271,n129,n46);
and (n272,n130,n48);
nand (n273,n274,n279);
or (n274,n92,n275);
not (n275,n276);
nor (n276,n277,n278);
and (n277,n60,n24);
and (n278,n61,n22);
or (n279,n13,n280);
nor (n280,n281,n282);
and (n281,n24,n65);
and (n282,n22,n64);
and (n283,n238,n253);
xor (n284,n285,n300);
xor (n285,n286,n293);
nand (n286,n287,n289);
or (n287,n27,n288);
not (n288,n206);
or (n289,n290,n28);
nor (n290,n291,n292);
and (n291,n61,n35);
and (n292,n36,n60);
nand (n293,n294,n299);
or (n294,n295,n71);
not (n295,n296);
nor (n296,n297,n298);
and (n297,n203,n56);
and (n298,n202,n55);
or (n299,n70,n229);
nand (n300,n301,n302);
or (n301,n259,n270);
or (n302,n264,n129);
xor (n303,n304,n368);
xor (n304,n305,n328);
xor (n305,n306,n319);
xor (n306,n307,n312);
nand (n307,n308,n311);
or (n308,n309,n51);
not (n309,n310);
nand (n311,n53,n226);
nand (n312,n313,n314);
or (n313,n92,n280);
or (n314,n13,n315);
not (n315,n316);
nor (n316,n317,n318);
and (n317,n83,n24);
and (n318,n81,n22);
not (n319,n320);
nand (n320,n321,n323);
or (n321,n322,n215);
not (n322,n217);
nand (n323,n324,n127);
not (n324,n325);
nor (n325,n326,n327);
and (n326,n42,n18);
and (n327,n40,n136);
or (n328,n329,n367);
and (n329,n330,n343);
xor (n330,n331,n336);
nand (n331,n332,n335);
or (n332,n333,n51);
not (n333,n334);
or (n335,n63,n309);
not (n336,n337);
nor (n337,n338,n342);
and (n338,n246,n339);
nor (n339,n340,n341);
and (n340,n48,n252);
and (n341,n46,n250);
and (n342,n240,n250);
or (n343,n344,n366);
and (n344,n345,n360);
xor (n345,n346,n353);
nand (n346,n347,n352);
or (n347,n348,n259);
not (n348,n349);
nor (n349,n350,n351);
and (n350,n89,n129);
and (n351,n87,n130);
nand (n352,n265,n256);
nand (n353,n354,n359);
or (n354,n355,n92);
not (n355,n356);
nor (n356,n357,n358);
and (n357,n102,n24);
and (n358,n103,n22);
nand (n359,n14,n276);
nand (n360,n361,n362);
or (n361,n199,n28);
nand (n362,n173,n363);
nor (n363,n364,n365);
and (n364,n231,n35);
and (n365,n232,n36);
and (n366,n346,n353);
and (n367,n331,n336);
or (n368,n369,n396);
and (n369,n370,n395);
xor (n370,n371,n394);
or (n371,n372,n393);
and (n372,n373,n388);
xor (n373,n374,n381);
nand (n374,n375,n380);
or (n375,n376,n215);
not (n376,n377);
nor (n377,n378,n379);
and (n378,n64,n136);
and (n379,n65,n18);
nand (n380,n127,n212);
nand (n381,n382,n387);
or (n382,n383,n70);
not (n383,n384);
nor (n384,n385,n386);
and (n385,n309,n55);
and (n386,n310,n56);
nand (n387,n72,n223);
nand (n388,n389,n392);
or (n389,n390,n51);
not (n390,n391);
nand (n392,n53,n334);
and (n393,n374,n381);
xor (n394,n196,n220);
xor (n395,n237,n273);
and (n396,n371,n394);
or (n397,n398,n492);
and (n398,n399,n461);
xor (n399,n400,n401);
xor (n400,n330,n343);
or (n401,n402,n460);
and (n402,n403,n437);
xor (n403,n337,n404);
or (n404,n405,n436);
and (n405,n406,n429);
xor (n406,n407,n421);
nand (n407,n408,n244);
or (n408,n409,n415);
nand (n409,n410,n414);
or (n410,n411,n413);
not (n411,n412);
nand (n414,n413,n411);
not (n415,n416);
nand (n416,n417,n418);
not (n417,n409);
nand (n418,n419,n420);
or (n419,n411,n244);
nand (n420,n411,n244);
nand (n421,n422,n428);
or (n422,n423,n427);
not (n423,n424);
nand (n424,n425,n426);
or (n425,n40,n252);
nand (n426,n252,n40);
not (n427,n246);
nand (n428,n339,n240);
nand (n429,n430,n435);
or (n430,n431,n215);
not (n431,n432);
nor (n432,n433,n434);
and (n433,n60,n136);
and (n434,n61,n18);
nand (n435,n127,n377);
and (n436,n407,n421);
or (n437,n438,n459);
and (n438,n439,n452);
xor (n439,n440,n445);
nand (n440,n441,n444);
or (n441,n442,n51);
not (n442,n443);
nand (n444,n53,n391);
nand (n445,n446,n451);
or (n446,n447,n92);
not (n447,n448);
nor (n448,n449,n450);
and (n449,n202,n24);
and (n450,n203,n22);
nand (n451,n14,n356);
nand (n452,n453,n454);
or (n453,n348,n264);
or (n454,n259,n455);
not (n455,n456);
nor (n456,n457,n458);
and (n457,n83,n129);
and (n458,n81,n130);
and (n459,n440,n445);
and (n460,n337,n404);
or (n461,n462,n491);
and (n462,n463,n466);
xor (n463,n464,n465);
xor (n464,n373,n388);
xor (n465,n345,n360);
or (n466,n467,n490);
and (n467,n468,n483);
xor (n468,n469,n476);
nand (n469,n470,n475);
or (n470,n471,n27);
not (n471,n472);
nor (n472,n473,n474);
and (n473,n35,n225);
and (n474,n226,n36);
nand (n475,n176,n363);
nand (n476,n477,n482);
or (n477,n478,n70);
not (n478,n479);
nor (n479,n480,n481);
and (n480,n333,n55);
and (n481,n334,n56);
nand (n482,n72,n384);
not (n483,n484);
nor (n484,n485,n489);
and (n485,n415,n486);
nor (n486,n487,n488);
and (n487,n48,n243);
and (n488,n46,n244);
nor (n489,n417,n243);
and (n490,n469,n476);
and (n491,n464,n465);
and (n492,n400,n401);
and (n493,n192,n303);
xor (n494,n495,n544);
xor (n495,n496,n499);
or (n496,n497,n498);
and (n497,n193,n284);
and (n498,n194,n235);
xor (n499,n500,n522);
xor (n500,n501,n519);
xor (n501,n502,n513);
xor (n502,n503,n506);
nand (n503,n504,n130);
or (n504,n265,n505);
not (n505,n259);
nand (n506,n507,n508);
or (n507,n215,n325);
or (n508,n509,n510);
not (n509,n127);
nor (n510,n511,n512);
and (n511,n136,n46);
and (n512,n18,n48);
nand (n513,n514,n515);
or (n514,n27,n290);
or (n515,n28,n516);
nor (n516,n517,n518);
and (n517,n35,n65);
and (n518,n36,n64);
or (n519,n520,n521);
and (n520,n306,n319);
and (n521,n307,n312);
xor (n522,n523,n527);
xor (n523,n320,n524);
or (n524,n525,n526);
and (n525,n285,n300);
and (n526,n286,n293);
xor (n527,n528,n541);
xor (n528,n529,n535);
nand (n529,n530,n531);
or (n530,n295,n70);
nand (n531,n72,n532);
nor (n532,n533,n534);
and (n533,n102,n55);
and (n534,n103,n56);
nand (n535,n536,n537);
or (n536,n315,n92);
nand (n537,n14,n538);
nor (n538,n539,n540);
and (n539,n89,n24);
and (n540,n87,n22);
nand (n541,n542,n543);
or (n542,n225,n51);
nand (n543,n53,n232);
or (n544,n545,n546);
and (n545,n304,n368);
and (n546,n305,n328);
nor (n547,n548,n590);
xor (n548,n549,n587);
xor (n549,n550,n553);
or (n550,n551,n552);
and (n551,n523,n527);
and (n552,n320,n524);
xor (n553,n554,n570);
xor (n554,n555,n558);
or (n555,n556,n557);
and (n556,n502,n513);
and (n557,n503,n506);
xor (n558,n559,n567);
xor (n559,n560,n564);
nand (n560,n561,n563);
or (n561,n70,n562);
not (n562,n532);
or (n563,n71,n147);
nand (n564,n565,n566);
or (n565,n231,n51);
nand (n566,n53,n203);
nand (n567,n568,n569);
or (n568,n215,n510);
or (n569,n509,n136);
xor (n570,n571,n584);
xor (n571,n572,n578);
nand (n572,n573,n574);
or (n573,n27,n516);
or (n574,n28,n575);
nor (n575,n576,n577);
and (n576,n35,n81);
and (n577,n36,n83);
not (n578,n579);
nand (n579,n580,n582);
or (n580,n581,n92);
not (n581,n538);
nand (n582,n583,n14);
not (n583,n141);
or (n584,n585,n586);
and (n585,n528,n541);
and (n586,n529,n535);
or (n587,n588,n589);
and (n588,n500,n522);
and (n589,n501,n519);
or (n590,n591,n592);
and (n591,n495,n544);
and (n592,n496,n499);
nand (n593,n594,n617);
not (n594,n595);
xor (n595,n596,n614);
xor (n596,n597,n600);
or (n597,n598,n599);
and (n598,n571,n584);
and (n599,n572,n578);
xor (n600,n601,n606);
xor (n601,n602,n605);
or (n602,n603,n604);
and (n603,n559,n567);
and (n604,n560,n564);
xor (n605,n124,n145);
xor (n606,n607,n579);
xor (n607,n608,n611);
nand (n608,n609,n610);
or (n609,n51,n202);
or (n610,n63,n102);
nand (n611,n612,n613);
or (n612,n27,n575);
or (n613,n107,n28);
or (n614,n615,n616);
and (n615,n554,n570);
and (n616,n555,n558);
not (n617,n618);
or (n618,n619,n620);
and (n619,n549,n587);
and (n620,n550,n553);
or (n621,n622,n625);
or (n622,n623,n624);
and (n623,n596,n614);
and (n624,n597,n600);
xor (n625,n626,n631);
xor (n626,n627,n630);
or (n627,n628,n629);
and (n628,n607,n579);
and (n629,n608,n611);
xor (n630,n120,n152);
or (n631,n632,n633);
and (n632,n601,n606);
and (n633,n602,n605);
nor (n634,n635,n638);
or (n635,n636,n637);
and (n636,n626,n631);
and (n637,n627,n630);
xor (n638,n7,n118);
not (n639,n640);
nand (n640,n641,n1353);
nor (n641,n642,n1339);
and (n642,n643,n1006);
and (n643,n644,n989);
nor (n644,n645,n897);
nor (n645,n646,n819);
xor (n646,n647,n728);
xor (n647,n648,n675);
or (n648,n649,n674);
and (n649,n650,n653);
xor (n650,n651,n652);
xor (n651,n439,n452);
xor (n652,n468,n483);
or (n653,n654,n673);
and (n654,n655,n663);
xor (n655,n656,n484);
nand (n656,n657,n662);
or (n657,n658,n70);
not (n658,n659);
nor (n659,n660,n661);
and (n660,n390,n55);
and (n661,n391,n56);
nand (n662,n72,n479);
nand (n663,n664,n413);
nor (n664,n665,n669);
and (n665,n505,n666);
nand (n666,n667,n668);
or (n667,n61,n129);
nand (n668,n129,n61);
and (n669,n265,n670);
nor (n670,n671,n672);
and (n671,n64,n129);
and (n672,n65,n130);
and (n673,n656,n484);
and (n674,n651,n652);
xor (n675,n676,n727);
xor (n676,n677,n678);
xor (n677,n403,n437);
or (n678,n679,n726);
and (n679,n680,n725);
xor (n680,n681,n702);
or (n681,n682,n701);
and (n682,n683,n695);
xor (n683,n684,n691);
nand (n684,n685,n690);
or (n685,n686,n92);
not (n686,n687);
nand (n687,n688,n689);
or (n688,n232,n24);
nand (n689,n24,n232);
nand (n690,n448,n14);
nand (n691,n692,n694);
or (n692,n693,n259);
not (n693,n670);
nand (n694,n265,n456);
nand (n695,n696,n697);
or (n696,n28,n471);
or (n697,n27,n698);
nor (n698,n699,n700);
and (n699,n310,n35);
and (n700,n36,n309);
and (n701,n684,n691);
or (n702,n703,n724);
and (n703,n704,n717);
xor (n704,n705,n712);
nand (n705,n706,n711);
or (n706,n707,n427);
not (n707,n708);
nor (n708,n709,n710);
and (n709,n89,n252);
and (n710,n87,n250);
nand (n711,n240,n424);
nand (n712,n713,n716);
or (n713,n714,n51);
not (n714,n715);
nand (n716,n53,n443);
nand (n717,n718,n723);
or (n718,n719,n215);
not (n719,n720);
nor (n720,n721,n722);
and (n721,n102,n136);
and (n722,n103,n18);
nand (n723,n127,n432);
and (n724,n705,n712);
xor (n725,n406,n429);
and (n726,n681,n702);
xor (n727,n463,n466);
or (n728,n729,n818);
and (n729,n730,n782);
xor (n730,n731,n732);
xor (n731,n680,n725);
or (n732,n733,n781);
and (n733,n734,n780);
xor (n734,n735,n757);
or (n735,n736,n756);
and (n736,n737,n750);
xor (n737,n738,n745);
nand (n738,n739,n744);
or (n739,n740,n70);
not (n740,n741);
nand (n741,n742,n743);
or (n742,n442,n56);
nand (n743,n56,n442);
nand (n744,n659,n72);
nand (n745,n746,n749);
or (n746,n747,n51);
not (n747,n748);
nand (n749,n53,n715);
nand (n750,n751,n753);
or (n751,n752,n417);
not (n752,n486);
or (n753,n416,n754);
not (n754,n755);
xor (n755,n42,n243);
and (n756,n738,n745);
or (n757,n758,n779);
and (n758,n759,n773);
xor (n759,n760,n767);
nand (n760,n761,n766);
or (n761,n762,n215);
not (n762,n763);
nor (n763,n764,n765);
and (n764,n202,n136);
and (n765,n203,n18);
nand (n766,n127,n720);
nand (n767,n768,n772);
or (n768,n769,n427);
nor (n769,n770,n771);
and (n770,n83,n250);
and (n771,n81,n252);
nand (n772,n708,n240);
nand (n773,n774,n778);
or (n774,n92,n775);
nor (n775,n776,n777);
and (n776,n225,n22);
and (n777,n226,n24);
or (n778,n13,n686);
and (n779,n760,n767);
xor (n780,n683,n695);
and (n781,n735,n757);
or (n782,n783,n817);
and (n783,n784,n787);
xor (n784,n785,n786);
xor (n785,n704,n717);
xor (n786,n655,n663);
and (n787,n788,n811);
or (n788,n789,n810);
and (n789,n790,n805);
xor (n790,n791,n798);
nand (n791,n792,n797);
or (n792,n793,n259);
not (n793,n794);
nor (n794,n795,n796);
and (n795,n102,n129);
and (n796,n103,n130);
nand (n797,n666,n265);
nand (n798,n799,n804);
or (n799,n800,n70);
not (n800,n801);
nand (n801,n802,n803);
or (n802,n715,n55);
nand (n803,n715,n55);
nand (n804,n72,n741);
nand (n805,n806,n809);
or (n806,n807,n51);
not (n807,n808);
nand (n809,n53,n748);
and (n810,n791,n798);
nand (n811,n812,n816);
or (n812,n27,n813);
nor (n813,n814,n815);
and (n814,n35,n334);
and (n815,n36,n333);
or (n816,n28,n698);
and (n817,n785,n786);
and (n818,n731,n732);
or (n819,n820,n896);
and (n820,n821,n824);
xor (n821,n822,n823);
xor (n822,n650,n653);
xor (n823,n730,n782);
or (n824,n825,n895);
and (n825,n826,n859);
xor (n826,n827,n828);
xor (n827,n734,n780);
or (n828,n829,n858);
and (n829,n830,n856);
xor (n830,n831,n855);
or (n831,n832,n854);
and (n832,n833,n848);
xor (n833,n834,n841);
nand (n834,n835,n840);
or (n835,n836,n416);
not (n836,n837);
nor (n837,n838,n839);
and (n838,n89,n243);
and (n839,n87,n244);
nand (n840,n409,n755);
nand (n841,n842,n847);
or (n842,n843,n215);
not (n843,n844);
nor (n844,n845,n846);
and (n845,n231,n136);
and (n846,n232,n18);
nand (n847,n127,n763);
nand (n848,n849,n852);
or (n849,n427,n850);
not (n850,n851);
xor (n851,n64,n252);
or (n852,n769,n853);
not (n853,n240);
and (n854,n834,n841);
xor (n855,n759,n773);
nand (n856,n857,n663);
or (n857,n413,n664);
and (n858,n831,n855);
or (n859,n860,n894);
and (n860,n861,n893);
xor (n861,n862,n863);
xor (n862,n737,n750);
or (n863,n864,n892);
and (n864,n865,n881);
xor (n865,n866,n874);
nand (n866,n867,n872);
or (n867,n868,n92);
not (n868,n869);
nand (n869,n870,n871);
or (n870,n22,n309);
or (n871,n24,n310);
nand (n872,n873,n14);
not (n873,n775);
nand (n874,n875,n880);
or (n875,n876,n27);
not (n876,n877);
nand (n877,n878,n879);
or (n878,n36,n390);
or (n879,n35,n391);
or (n880,n28,n813);
nand (n881,n882,n891);
or (n882,n883,n886);
nand (n883,n884,n413);
not (n884,n885);
not (n886,n887);
nor (n887,n888,n890);
and (n888,n48,n889);
not (n889,n413);
and (n890,n46,n413);
or (n891,n889,n884);
and (n892,n866,n874);
xor (n893,n811,n788);
and (n894,n862,n863);
and (n895,n827,n828);
and (n896,n822,n823);
nor (n897,n898,n899);
xor (n898,n821,n824);
or (n899,n900,n988);
and (n900,n901,n987);
xor (n901,n902,n903);
xor (n902,n784,n787);
or (n903,n904,n986);
and (n904,n905,n985);
xor (n905,n906,n978);
or (n906,n907,n977);
and (n907,n908,n952);
xor (n908,n909,n927);
or (n909,n910,n926);
and (n910,n911,n919);
xor (n911,n912,n913);
and (n912,n53,n808);
nand (n913,n914,n918);
or (n914,n883,n915);
nor (n915,n916,n917);
and (n916,n42,n413);
and (n917,n40,n889);
nand (n918,n887,n885);
nand (n919,n920,n925);
or (n920,n921,n416);
not (n921,n922);
nor (n922,n923,n924);
and (n923,n83,n243);
and (n924,n81,n244);
nand (n925,n409,n837);
and (n926,n912,n913);
or (n927,n928,n951);
and (n928,n929,n944);
xor (n929,n930,n937);
nand (n930,n931,n936);
or (n931,n932,n427);
not (n932,n933);
nor (n933,n934,n935);
and (n934,n60,n252);
and (n935,n61,n250);
nand (n936,n851,n240);
nand (n937,n938,n939);
or (n938,n13,n868);
nand (n939,n940,n12);
not (n940,n941);
nor (n941,n942,n943);
and (n942,n334,n24);
and (n943,n333,n22);
nand (n944,n945,n946);
or (n945,n876,n28);
nand (n946,n947,n173);
not (n947,n948);
nor (n948,n949,n950);
and (n949,n443,n35);
and (n950,n36,n442);
and (n951,n930,n937);
or (n952,n953,n976);
and (n953,n954,n969);
xor (n954,n955,n962);
nand (n955,n956,n961);
or (n956,n957,n70);
not (n957,n958);
nor (n958,n959,n960);
and (n959,n747,n55);
and (n960,n748,n56);
nand (n961,n801,n72);
nand (n962,n963,n968);
or (n963,n964,n259);
not (n964,n965);
nand (n965,n966,n967);
or (n966,n130,n202);
or (n967,n129,n203);
nand (n968,n265,n794);
nand (n969,n970,n975);
or (n970,n215,n971);
not (n971,n972);
nor (n972,n973,n974);
and (n973,n225,n136);
and (n974,n226,n18);
or (n975,n509,n843);
and (n976,n955,n962);
and (n977,n909,n927);
or (n978,n979,n984);
and (n979,n980,n983);
xor (n980,n981,n982);
xor (n981,n790,n805);
xor (n982,n833,n848);
xor (n983,n865,n881);
and (n984,n981,n982);
xor (n985,n830,n856);
and (n986,n906,n978);
xor (n987,n826,n859);
and (n988,n902,n903);
nor (n989,n990,n1001);
nor (n990,n991,n992);
xor (n991,n191,n397);
or (n992,n993,n1000);
and (n993,n994,n997);
xor (n994,n995,n996);
xor (n995,n370,n395);
xor (n996,n399,n461);
or (n997,n998,n999);
and (n998,n676,n727);
and (n999,n677,n678);
and (n1000,n995,n996);
nor (n1001,n1002,n1003);
xor (n1002,n994,n997);
or (n1003,n1004,n1005);
and (n1004,n647,n728);
and (n1005,n648,n675);
nand (n1006,n1007,n1333);
or (n1007,n1008,n1315);
not (n1008,n1009);
nor (n1009,n1010,n1314);
and (n1010,n1011,n1252);
nand (n1011,n1012,n1157);
xor (n1012,n1013,n1144);
xor (n1013,n1014,n1015);
xor (n1014,n980,n983);
or (n1015,n1016,n1143);
and (n1016,n1017,n1113);
xor (n1017,n1018,n1065);
or (n1018,n1019,n1064);
and (n1019,n1020,n1041);
xor (n1020,n1021,n1027);
nand (n1021,n1022,n1026);
or (n1022,n27,n1023);
nor (n1023,n1024,n1025);
and (n1024,n35,n715);
and (n1025,n36,n714);
or (n1026,n28,n948);
xor (n1027,n1028,n1034);
nor (n1028,n1029,n55);
nor (n1029,n1030,n1032);
and (n1030,n1031,n35);
nand (n1031,n808,n74);
and (n1032,n807,n1033);
not (n1033,n74);
nand (n1034,n1035,n1040);
or (n1035,n1036,n883);
not (n1036,n1037);
nor (n1037,n1038,n1039);
and (n1038,n89,n889);
and (n1039,n87,n413);
or (n1040,n915,n884);
or (n1041,n1042,n1063);
and (n1042,n1043,n1052);
xor (n1043,n1044,n1045);
and (n1044,n72,n808);
nand (n1045,n1046,n1051);
or (n1046,n883,n1047);
not (n1047,n1048);
nor (n1048,n1049,n1050);
and (n1049,n83,n889);
and (n1050,n81,n413);
nand (n1051,n1037,n885);
nand (n1052,n1053,n1058);
or (n1053,n416,n1054);
not (n1054,n1055);
nor (n1055,n1056,n1057);
and (n1056,n243,n60);
and (n1057,n61,n244);
or (n1058,n417,n1059);
not (n1059,n1060);
nor (n1060,n1061,n1062);
and (n1061,n64,n243);
and (n1062,n65,n244);
and (n1063,n1044,n1045);
and (n1064,n1021,n1027);
xor (n1065,n1066,n1089);
xor (n1066,n1067,n1068);
and (n1067,n1028,n1034);
or (n1068,n1069,n1088);
and (n1069,n1070,n1081);
xor (n1070,n1071,n1074);
nand (n1071,n1072,n1073);
or (n1072,n1059,n416);
nand (n1073,n922,n409);
nand (n1074,n1075,n1080);
or (n1075,n1076,n70);
not (n1076,n1077);
nand (n1077,n1078,n1079);
or (n1078,n55,n808);
or (n1079,n56,n807);
nand (n1080,n958,n72);
nand (n1081,n1082,n1083);
or (n1082,n964,n264);
or (n1083,n259,n1084);
not (n1084,n1085);
nor (n1085,n1086,n1087);
and (n1086,n231,n129);
and (n1087,n232,n130);
and (n1088,n1071,n1074);
or (n1089,n1090,n1112);
and (n1090,n1091,n1106);
xor (n1091,n1092,n1099);
nand (n1092,n1093,n1098);
or (n1093,n1094,n215);
not (n1094,n1095);
nor (n1095,n1096,n1097);
and (n1096,n309,n136);
and (n1097,n310,n18);
nand (n1098,n127,n972);
nand (n1099,n1100,n1105);
or (n1100,n1101,n427);
not (n1101,n1102);
nand (n1102,n1103,n1104);
or (n1103,n250,n102);
or (n1104,n252,n103);
nand (n1105,n240,n933);
nand (n1106,n1107,n1111);
or (n1107,n92,n1108);
nor (n1108,n1109,n1110);
and (n1109,n24,n391);
and (n1110,n22,n390);
or (n1111,n13,n941);
and (n1112,n1092,n1099);
or (n1113,n1114,n1142);
and (n1114,n1115,n1141);
xor (n1115,n1116,n1140);
or (n1116,n1117,n1139);
and (n1117,n1118,n1132);
xor (n1118,n1119,n1126);
nand (n1119,n1120,n1125);
or (n1120,n1121,n259);
not (n1121,n1122);
nor (n1122,n1123,n1124);
and (n1123,n226,n130);
and (n1124,n225,n129);
nand (n1125,n265,n1085);
nand (n1126,n1127,n1131);
or (n1127,n215,n1128);
nor (n1128,n1129,n1130);
and (n1129,n333,n18);
and (n1130,n334,n136);
nand (n1131,n127,n1095);
nand (n1132,n1133,n1134);
or (n1133,n853,n1101);
nand (n1134,n1135,n246);
not (n1135,n1136);
nor (n1136,n1137,n1138);
and (n1137,n252,n203);
and (n1138,n250,n202);
and (n1139,n1119,n1126);
xor (n1140,n1091,n1106);
xor (n1141,n1070,n1081);
and (n1142,n1116,n1140);
and (n1143,n1018,n1065);
xor (n1144,n1145,n1150);
xor (n1145,n1146,n1149);
or (n1146,n1147,n1148);
and (n1147,n1066,n1089);
and (n1148,n1067,n1068);
xor (n1149,n908,n952);
or (n1150,n1151,n1156);
and (n1151,n1152,n1155);
xor (n1152,n1153,n1154);
xor (n1153,n929,n944);
xor (n1154,n911,n919);
xor (n1155,n954,n969);
and (n1156,n1153,n1154);
or (n1157,n1158,n1251);
and (n1158,n1159,n1250);
xor (n1159,n1160,n1161);
xor (n1160,n1152,n1155);
or (n1161,n1162,n1249);
and (n1162,n1163,n1196);
xor (n1163,n1164,n1195);
or (n1164,n1165,n1194);
and (n1165,n1166,n1181);
xor (n1166,n1167,n1174);
nand (n1167,n1168,n1172);
or (n1168,n1169,n92);
nor (n1169,n1170,n1171);
and (n1170,n442,n22);
and (n1171,n443,n24);
nand (n1172,n1173,n14);
not (n1173,n1108);
nand (n1174,n1175,n1179);
or (n1175,n27,n1176);
nor (n1176,n1177,n1178);
and (n1177,n35,n748);
and (n1178,n36,n747);
nand (n1179,n1180,n176);
not (n1180,n1023);
and (n1181,n1182,n1187);
nor (n1182,n1183,n35);
nor (n1183,n1184,n1186);
and (n1184,n1185,n24);
nand (n1185,n808,n31);
and (n1186,n807,n30);
nand (n1187,n1188,n1193);
or (n1188,n883,n1189);
not (n1189,n1190);
nor (n1190,n1191,n1192);
and (n1191,n64,n889);
and (n1192,n65,n413);
nand (n1193,n1048,n885);
and (n1194,n1167,n1174);
xor (n1195,n1020,n1041);
or (n1196,n1197,n1248);
and (n1197,n1198,n1247);
xor (n1198,n1199,n1224);
or (n1199,n1200,n1223);
and (n1200,n1201,n1216);
xor (n1201,n1202,n1209);
nand (n1202,n1203,n1208);
or (n1203,n1204,n416);
not (n1204,n1205);
nor (n1205,n1206,n1207);
and (n1206,n102,n243);
and (n1207,n103,n244);
nand (n1208,n1055,n409);
nand (n1209,n1210,n1215);
or (n1210,n1211,n259);
not (n1211,n1212);
nand (n1212,n1213,n1214);
or (n1213,n130,n309);
or (n1214,n129,n310);
nand (n1215,n265,n1122);
nand (n1216,n1217,n1222);
or (n1217,n215,n1218);
not (n1218,n1219);
nor (n1219,n1220,n1221);
and (n1220,n390,n136);
and (n1221,n391,n18);
or (n1222,n509,n1128);
and (n1223,n1202,n1209);
or (n1224,n1225,n1246);
and (n1225,n1226,n1240);
xor (n1226,n1227,n1233);
nand (n1227,n1228,n1232);
or (n1228,n427,n1229);
nor (n1229,n1230,n1231);
and (n1230,n232,n252);
and (n1231,n231,n250);
or (n1232,n1136,n853);
nand (n1233,n1234,n1239);
or (n1234,n92,n1235);
not (n1235,n1236);
nor (n1236,n1237,n1238);
and (n1237,n714,n24);
and (n1238,n715,n22);
or (n1239,n1169,n13);
nand (n1240,n1241,n1245);
or (n1241,n27,n1242);
nor (n1242,n1243,n1244);
and (n1243,n807,n36);
and (n1244,n808,n35);
or (n1245,n1176,n28);
and (n1246,n1227,n1233);
xor (n1247,n1043,n1052);
and (n1248,n1199,n1224);
and (n1249,n1164,n1195);
xor (n1250,n1017,n1113);
and (n1251,n1160,n1161);
nand (n1252,n1253,n1254);
xor (n1253,n1159,n1250);
or (n1254,n1255,n1313);
and (n1255,n1256,n1312);
xor (n1256,n1257,n1258);
xor (n1257,n1115,n1141);
or (n1258,n1259,n1311);
and (n1259,n1260,n1263);
xor (n1260,n1261,n1262);
xor (n1261,n1118,n1132);
xor (n1262,n1166,n1181);
or (n1263,n1264,n1310);
and (n1264,n1265,n1285);
xor (n1265,n1266,n1267);
xor (n1266,n1182,n1187);
or (n1267,n1268,n1284);
and (n1268,n1269,n1278);
xor (n1269,n1270,n1271);
and (n1270,n176,n808);
nand (n1271,n1272,n1277);
or (n1272,n1273,n416);
not (n1273,n1274);
nor (n1274,n1275,n1276);
and (n1275,n202,n243);
and (n1276,n203,n244);
nand (n1277,n409,n1205);
nand (n1278,n1279,n1280);
or (n1279,n1211,n264);
or (n1280,n259,n1281);
nor (n1281,n1282,n1283);
and (n1282,n129,n334);
and (n1283,n130,n333);
and (n1284,n1270,n1271);
or (n1285,n1286,n1309);
and (n1286,n1287,n1302);
xor (n1287,n1288,n1295);
nand (n1288,n1289,n1294);
or (n1289,n1290,n215);
not (n1290,n1291);
nand (n1291,n1292,n1293);
or (n1292,n442,n18);
or (n1293,n136,n443);
nand (n1294,n1219,n127);
nand (n1295,n1296,n1297);
or (n1296,n884,n1189);
nand (n1297,n1298,n1301);
nor (n1298,n1299,n1300);
and (n1299,n60,n889);
and (n1300,n61,n413);
not (n1301,n883);
nand (n1302,n1303,n1308);
or (n1303,n1304,n92);
not (n1304,n1305);
nand (n1305,n1306,n1307);
or (n1306,n22,n747);
or (n1307,n24,n748);
nand (n1308,n1236,n14);
and (n1309,n1288,n1295);
and (n1310,n1266,n1267);
and (n1311,n1261,n1262);
xor (n1312,n1163,n1196);
and (n1313,n1257,n1258);
nor (n1314,n1012,n1157);
not (n1315,n1316);
nor (n1316,n1317,n1328);
nor (n1317,n1318,n1319);
xor (n1318,n901,n987);
or (n1319,n1320,n1327);
and (n1320,n1321,n1326);
xor (n1321,n1322,n1323);
xor (n1322,n861,n893);
or (n1323,n1324,n1325);
and (n1324,n1145,n1150);
and (n1325,n1146,n1149);
xor (n1326,n905,n985);
and (n1327,n1322,n1323);
nor (n1328,n1329,n1330);
xor (n1329,n1321,n1326);
or (n1330,n1331,n1332);
and (n1331,n1013,n1144);
and (n1332,n1014,n1015);
nor (n1333,n1334,n1338);
and (n1334,n1335,n1336);
not (n1335,n1317);
not (n1336,n1337);
nand (n1337,n1329,n1330);
and (n1338,n1318,n1319);
nand (n1339,n1340,n1347);
or (n1340,n1341,n1342);
not (n1341,n989);
not (n1342,n1343);
nor (n1343,n1344,n645);
and (n1344,n1345,n1346);
nand (n1345,n819,n646);
nand (n1346,n898,n899);
nor (n1347,n1348,n1352);
and (n1348,n1349,n1350);
not (n1349,n990);
not (n1350,n1351);
nand (n1351,n1002,n1003);
and (n1352,n991,n992);
nand (n1353,n643,n1354,n1357);
and (n1354,n1316,n1355);
nor (n1355,n1314,n1356);
nor (n1356,n1253,n1254);
nand (n1357,n1358,n1858);
or (n1358,n1359,n1794);
not (n1359,n1360);
nand (n1360,n1361,n1783,n1793);
nand (n1361,n1362,n1589,n1650);
nor (n1362,n1363,n1527);
not (n1363,n1364);
or (n1364,n1365,n1490);
xor (n1365,n1366,n1450);
xor (n1366,n1367,n1397);
xor (n1367,n1368,n1388);
xor (n1368,n1369,n1379);
nand (n1369,n1370,n1375);
or (n1370,n1371,n215);
not (n1371,n1372);
nor (n1372,n1373,n1374);
and (n1373,n747,n136);
and (n1374,n748,n18);
nand (n1375,n127,n1376);
nand (n1376,n1377,n1378);
or (n1377,n18,n714);
or (n1378,n136,n715);
nand (n1379,n1380,n1384);
or (n1380,n1381,n883);
nor (n1381,n1382,n1383);
and (n1382,n889,n203);
and (n1383,n413,n202);
or (n1384,n1385,n884);
nor (n1385,n1386,n1387);
and (n1386,n889,n103);
and (n1387,n413,n102);
nand (n1388,n1389,n1393);
or (n1389,n427,n1390);
nor (n1390,n1391,n1392);
and (n1391,n252,n334);
and (n1392,n250,n333);
or (n1393,n1394,n853);
nor (n1394,n1395,n1396);
and (n1395,n252,n310);
and (n1396,n250,n309);
or (n1397,n1398,n1449);
and (n1398,n1399,n1424);
xor (n1399,n1400,n1406);
nand (n1400,n1401,n1405);
or (n1401,n427,n1402);
nor (n1402,n1403,n1404);
and (n1403,n252,n391);
and (n1404,n250,n390);
or (n1405,n853,n1390);
xor (n1406,n1407,n1413);
and (n1407,n1408,n18);
nand (n1408,n1409,n1410);
or (n1409,n808,n131);
nand (n1410,n1411,n129);
not (n1411,n1412);
and (n1412,n808,n131);
nand (n1413,n1414,n1419);
or (n1414,n1415,n417);
not (n1415,n1416);
nand (n1416,n1417,n1418);
or (n1417,n244,n225);
or (n1418,n243,n226);
nand (n1419,n1420,n415);
not (n1420,n1421);
nor (n1421,n1422,n1423);
and (n1422,n243,n310);
and (n1423,n244,n309);
or (n1424,n1425,n1448);
and (n1425,n1426,n1438);
xor (n1426,n1427,n1428);
and (n1427,n127,n808);
nand (n1428,n1429,n1434);
or (n1429,n884,n1430);
not (n1430,n1431);
nor (n1431,n1432,n1433);
and (n1432,n231,n889);
and (n1433,n232,n413);
or (n1434,n1435,n883);
nor (n1435,n1436,n1437);
and (n1436,n889,n226);
and (n1437,n413,n225);
nand (n1438,n1439,n1443);
or (n1439,n259,n1440);
nor (n1440,n1441,n1442);
and (n1441,n129,n748);
and (n1442,n130,n747);
or (n1443,n264,n1444);
not (n1444,n1445);
nor (n1445,n1446,n1447);
and (n1446,n715,n130);
and (n1447,n714,n129);
and (n1448,n1427,n1428);
and (n1449,n1400,n1406);
xor (n1450,n1451,n1473);
xor (n1451,n1452,n1453);
and (n1452,n1407,n1413);
or (n1453,n1454,n1472);
and (n1454,n1455,n1469);
xor (n1455,n1456,n1462);
nand (n1456,n1457,n1458);
or (n1457,n1444,n259);
nand (n1458,n265,n1459);
nor (n1459,n1460,n1461);
and (n1460,n442,n129);
and (n1461,n443,n130);
nand (n1462,n1463,n1468);
or (n1463,n1464,n215);
not (n1464,n1465);
nand (n1465,n1466,n1467);
or (n1466,n136,n808);
or (n1467,n807,n18);
nand (n1468,n127,n1372);
nand (n1469,n1470,n1471);
or (n1470,n883,n1430);
or (n1471,n1381,n884);
and (n1472,n1456,n1462);
xor (n1473,n1474,n1482);
xor (n1474,n1475,n1476);
and (n1475,n14,n808);
nand (n1476,n1477,n1478);
or (n1477,n1415,n416);
nand (n1478,n409,n1479);
nand (n1479,n1480,n1481);
or (n1480,n244,n231);
or (n1481,n243,n232);
nand (n1482,n1483,n1485);
or (n1483,n1484,n259);
not (n1484,n1459);
nand (n1485,n1486,n265);
not (n1486,n1487);
nor (n1487,n1488,n1489);
and (n1488,n129,n391);
and (n1489,n130,n390);
or (n1490,n1491,n1526);
and (n1491,n1492,n1525);
xor (n1492,n1493,n1494);
xor (n1493,n1455,n1469);
or (n1494,n1495,n1524);
and (n1495,n1496,n1509);
xor (n1496,n1497,n1503);
nand (n1497,n1498,n1502);
or (n1498,n416,n1499);
nor (n1499,n1500,n1501);
and (n1500,n243,n334);
and (n1501,n244,n333);
or (n1502,n417,n1421);
nand (n1503,n1504,n1508);
or (n1504,n427,n1505);
nor (n1505,n1506,n1507);
and (n1506,n252,n443);
and (n1507,n250,n442);
or (n1508,n1402,n853);
and (n1509,n1510,n1517);
nor (n1510,n1511,n129);
nor (n1511,n1512,n1515);
and (n1512,n1513,n252);
not (n1513,n1514);
and (n1514,n808,n262);
and (n1515,n807,n1516);
not (n1516,n262);
nand (n1517,n1518,n1523);
or (n1518,n1519,n883);
not (n1519,n1520);
nor (n1520,n1521,n1522);
and (n1521,n309,n889);
and (n1522,n310,n413);
or (n1523,n1435,n884);
and (n1524,n1497,n1503);
xor (n1525,n1399,n1424);
and (n1526,n1493,n1494);
nand (n1527,n1528,n1583);
not (n1528,n1529);
nor (n1529,n1530,n1558);
xor (n1530,n1531,n1557);
xor (n1531,n1532,n1556);
or (n1532,n1533,n1555);
and (n1533,n1534,n1549);
xor (n1534,n1535,n1543);
nand (n1535,n1536,n1541);
or (n1536,n1537,n259);
not (n1537,n1538);
nand (n1538,n1539,n1540);
or (n1539,n129,n808);
or (n1540,n130,n807);
nand (n1541,n1542,n265);
not (n1542,n1440);
nand (n1543,n1544,n1548);
or (n1544,n416,n1545);
nor (n1545,n1546,n1547);
and (n1546,n243,n391);
and (n1547,n244,n390);
or (n1548,n1499,n417);
nand (n1549,n1550,n1554);
or (n1550,n427,n1551);
nor (n1551,n1552,n1553);
and (n1552,n252,n715);
and (n1553,n250,n714);
or (n1554,n1505,n853);
and (n1555,n1535,n1543);
xor (n1556,n1426,n1438);
xor (n1557,n1496,n1509);
or (n1558,n1559,n1582);
and (n1559,n1560,n1581);
xor (n1560,n1561,n1562);
xor (n1561,n1510,n1517);
or (n1562,n1563,n1580);
and (n1563,n1564,n1573);
xor (n1564,n1565,n1566);
and (n1565,n265,n808);
nand (n1566,n1567,n1572);
or (n1567,n883,n1568);
not (n1568,n1569);
nor (n1569,n1570,n1571);
and (n1570,n334,n413);
and (n1571,n333,n889);
nand (n1572,n1520,n885);
nand (n1573,n1574,n1579);
or (n1574,n416,n1575);
not (n1575,n1576);
nor (n1576,n1577,n1578);
and (n1577,n442,n243);
and (n1578,n443,n244);
or (n1579,n417,n1545);
and (n1580,n1565,n1566);
xor (n1581,n1534,n1549);
and (n1582,n1561,n1562);
not (n1583,n1584);
nor (n1584,n1585,n1586);
xor (n1585,n1492,n1525);
or (n1586,n1587,n1588);
and (n1587,n1531,n1557);
and (n1588,n1532,n1556);
nand (n1589,n1590,n1646);
not (n1590,n1591);
xor (n1591,n1592,n1643);
xor (n1592,n1593,n1623);
xor (n1593,n1594,n1608);
xor (n1594,n1595,n1602);
nand (n1595,n1596,n1597);
or (n1596,n1304,n13);
nand (n1597,n1598,n12);
not (n1598,n1599);
nor (n1599,n1600,n1601);
and (n1600,n807,n22);
and (n1601,n24,n808);
nand (n1602,n1603,n1604);
or (n1603,n427,n1394);
or (n1604,n853,n1605);
nor (n1605,n1606,n1607);
and (n1606,n252,n226);
and (n1607,n250,n225);
nand (n1608,n1609,n1622);
or (n1609,n1610,n1617);
not (n1610,n1611);
nand (n1611,n1612,n22);
nand (n1612,n1613,n1614);
or (n1613,n808,n17);
nand (n1614,n1615,n136);
not (n1615,n1616);
and (n1616,n808,n17);
not (n1617,n1618);
nand (n1618,n1619,n1621);
or (n1619,n1620,n416);
not (n1620,n1479);
nand (n1621,n409,n1274);
or (n1622,n1618,n1611);
xor (n1623,n1624,n1631);
xor (n1624,n1625,n1628);
or (n1625,n1626,n1627);
and (n1626,n1474,n1482);
and (n1627,n1475,n1476);
or (n1628,n1629,n1630);
and (n1629,n1368,n1388);
and (n1630,n1369,n1379);
xor (n1631,n1632,n1639);
xor (n1632,n1633,n1636);
nand (n1633,n1634,n1635);
or (n1634,n259,n1487);
or (n1635,n1281,n264);
nand (n1636,n1637,n1638);
or (n1637,n1290,n509);
nand (n1638,n133,n1376);
nand (n1639,n1640,n1641);
or (n1640,n1385,n883);
or (n1641,n1642,n884);
not (n1642,n1298);
or (n1643,n1644,n1645);
and (n1644,n1451,n1473);
and (n1645,n1452,n1453);
not (n1646,n1647);
or (n1647,n1648,n1649);
and (n1648,n1366,n1450);
and (n1649,n1367,n1397);
or (n1650,n1651,n1782);
and (n1651,n1652,n1679);
xor (n1652,n1653,n1678);
or (n1653,n1654,n1677);
and (n1654,n1655,n1676);
xor (n1655,n1656,n1663);
nand (n1656,n1657,n1662);
or (n1657,n427,n1658);
not (n1658,n1659);
nor (n1659,n1660,n1661);
and (n1660,n748,n250);
and (n1661,n747,n252);
or (n1662,n1551,n853);
and (n1663,n1664,n1670);
nor (n1664,n1665,n252);
nor (n1665,n1666,n1669);
and (n1666,n1667,n243);
not (n1667,n1668);
and (n1668,n808,n242);
and (n1669,n807,n249);
nand (n1670,n1671,n1672);
or (n1671,n884,n1568);
nand (n1672,n1673,n1301);
nand (n1673,n1674,n1675);
or (n1674,n391,n889);
nand (n1675,n889,n391);
xor (n1676,n1564,n1573);
and (n1677,n1656,n1663);
xor (n1678,n1560,n1581);
or (n1679,n1680,n1781);
and (n1680,n1681,n1700);
xor (n1681,n1682,n1699);
or (n1682,n1683,n1698);
and (n1683,n1684,n1697);
xor (n1684,n1685,n1690);
nand (n1685,n1686,n1689);
or (n1686,n1687,n416);
not (n1687,n1688);
xor (n1688,n714,n243);
nand (n1689,n409,n1576);
nand (n1690,n1691,n1696);
or (n1691,n1692,n427);
not (n1692,n1693);
nand (n1693,n1694,n1695);
or (n1694,n252,n808);
or (n1695,n807,n250);
nand (n1696,n1659,n240);
xor (n1697,n1664,n1670);
and (n1698,n1685,n1690);
xor (n1699,n1655,n1676);
or (n1700,n1701,n1780);
and (n1701,n1702,n1724);
xor (n1702,n1703,n1723);
or (n1703,n1704,n1722);
and (n1704,n1705,n1714);
xor (n1705,n1706,n1707);
and (n1706,n240,n808);
nand (n1707,n1708,n1713);
or (n1708,n1709,n416);
not (n1709,n1710);
nor (n1710,n1711,n1712);
and (n1711,n747,n243);
and (n1712,n748,n244);
nand (n1713,n409,n1688);
nand (n1714,n1715,n1720);
or (n1715,n883,n1716);
not (n1716,n1717);
nand (n1717,n1718,n1719);
or (n1718,n443,n889);
nand (n1719,n889,n443);
or (n1720,n1721,n884);
not (n1721,n1673);
and (n1722,n1706,n1707);
xor (n1723,n1684,n1697);
nand (n1724,n1725,n1779);
or (n1725,n1726,n1741);
nor (n1726,n1727,n1728);
xor (n1727,n1705,n1714);
nor (n1728,n1729,n1736);
not (n1729,n1730);
nand (n1730,n1731,n1735);
or (n1731,n883,n1732);
nor (n1732,n1733,n1734);
and (n1733,n714,n413);
and (n1734,n715,n889);
nand (n1735,n1717,n885);
nand (n1736,n1737,n244);
nand (n1737,n1738,n1740);
or (n1738,n1739,n413);
and (n1739,n808,n412);
or (n1740,n808,n412);
nor (n1741,n1742,n1778);
and (n1742,n1743,n1754);
nand (n1743,n1744,n1748);
nor (n1744,n1745,n1746);
and (n1745,n1736,n1730);
and (n1746,n1747,n1729);
not (n1747,n1736);
nor (n1748,n1749,n1753);
and (n1749,n415,n1750);
nand (n1750,n1751,n1752);
or (n1751,n243,n808);
or (n1752,n807,n244);
and (n1753,n409,n1710);
nand (n1754,n1755,n1777);
or (n1755,n1756,n1771);
not (n1756,n1757);
nor (n1757,n1758,n1769);
not (n1758,n1759);
nand (n1759,n1760,n1765);
or (n1760,n884,n1761);
not (n1761,n1762);
nor (n1762,n1763,n1764);
and (n1763,n747,n889);
and (n1764,n748,n413);
nand (n1765,n1766,n1301);
nor (n1766,n1767,n1768);
and (n1767,n807,n889);
and (n1768,n808,n413);
nand (n1769,n1770,n413);
nand (n1770,n808,n885);
not (n1771,n1772);
nand (n1772,n1773,n1776);
nor (n1773,n1774,n1775);
nor (n1774,n1761,n883);
nor (n1775,n1732,n884);
nand (n1776,n808,n409);
or (n1777,n1773,n1776);
nor (n1778,n1748,n1744);
nand (n1779,n1727,n1728);
and (n1780,n1703,n1723);
and (n1781,n1682,n1699);
and (n1782,n1653,n1678);
nand (n1783,n1784,n1589);
or (n1784,n1785,n1787);
not (n1785,n1786);
nand (n1786,n1365,n1490);
not (n1787,n1788);
nand (n1788,n1364,n1789);
nand (n1789,n1790,n1792);
or (n1790,n1584,n1791);
nand (n1791,n1530,n1558);
nand (n1792,n1585,n1586);
nand (n1793,n1591,n1647);
not (n1794,n1795);
nor (n1795,n1796,n1821);
nor (n1796,n1797,n1798);
xor (n1797,n1256,n1312);
or (n1798,n1799,n1820);
and (n1799,n1800,n1803);
xor (n1800,n1801,n1802);
xor (n1801,n1198,n1247);
xor (n1802,n1260,n1263);
or (n1803,n1804,n1819);
and (n1804,n1805,n1808);
xor (n1805,n1806,n1807);
xor (n1806,n1226,n1240);
xor (n1807,n1201,n1216);
or (n1808,n1809,n1818);
and (n1809,n1810,n1815);
xor (n1810,n1811,n1814);
nand (n1811,n1812,n1813);
or (n1812,n427,n1605);
or (n1813,n1229,n853);
nor (n1814,n1617,n1611);
or (n1815,n1816,n1817);
and (n1816,n1632,n1639);
and (n1817,n1633,n1636);
and (n1818,n1811,n1814);
and (n1819,n1806,n1807);
and (n1820,n1801,n1802);
nand (n1821,n1822,n1851);
nor (n1822,n1823,n1846);
nor (n1823,n1824,n1837);
xor (n1824,n1825,n1836);
xor (n1825,n1826,n1827);
xor (n1826,n1265,n1285);
or (n1827,n1828,n1835);
and (n1828,n1829,n1832);
xor (n1829,n1830,n1831);
xor (n1830,n1287,n1302);
xor (n1831,n1269,n1278);
or (n1832,n1833,n1834);
and (n1833,n1594,n1608);
and (n1834,n1595,n1602);
and (n1835,n1830,n1831);
xor (n1836,n1805,n1808);
or (n1837,n1838,n1845);
and (n1838,n1839,n1844);
xor (n1839,n1840,n1841);
xor (n1840,n1810,n1815);
or (n1841,n1842,n1843);
and (n1842,n1624,n1631);
and (n1843,n1625,n1628);
xor (n1844,n1829,n1832);
and (n1845,n1840,n1841);
nor (n1846,n1847,n1850);
or (n1847,n1848,n1849);
and (n1848,n1592,n1643);
and (n1849,n1593,n1623);
xor (n1850,n1839,n1844);
nand (n1851,n1852,n1854);
not (n1852,n1853);
xor (n1853,n1800,n1803);
not (n1854,n1855);
or (n1855,n1856,n1857);
and (n1856,n1825,n1836);
and (n1857,n1826,n1827);
nor (n1858,n1859,n1870);
and (n1859,n1860,n1869);
nand (n1860,n1861,n1868);
or (n1861,n1862,n1863);
not (n1862,n1851);
not (n1863,n1864);
nand (n1864,n1865,n1867);
or (n1865,n1823,n1866);
nand (n1866,n1847,n1850);
nand (n1867,n1824,n1837);
nand (n1868,n1853,n1855);
not (n1869,n1796);
and (n1870,n1797,n1798);
nor (n1871,n1872,n1888);
and (n1872,n1873,n1887);
nand (n1873,n1874,n1886);
or (n1874,n1875,n1876);
not (n1875,n621);
not (n1876,n1877);
nand (n1877,n1878,n1885);
or (n1878,n1879,n1880);
not (n1879,n593);
not (n1880,n1881);
nand (n1881,n1882,n1884);
or (n1882,n1883,n547);
nand (n1883,n494,n189);
nand (n1884,n548,n590);
nand (n1885,n618,n595);
nand (n1886,n622,n625);
not (n1887,n634);
not (n1888,n1889);
nand (n1889,n635,n638);
and (n1890,n1891,n1892);
not (n1891,n2);
not (n1892,n181);
xor (n1893,n1894,n3276);
xor (n1894,n1895,n3275);
xor (n1895,n1896,n3201);
xor (n1896,n1897,n3200);
xor (n1897,n1898,n3113);
xor (n1898,n1899,n3112);
xor (n1899,n1900,n3022);
xor (n1900,n1901,n3021);
or (n1901,n1902,n2926);
and (n1902,n1903,n2925);
or (n1903,n1904,n2836);
and (n1904,n1905,n2835);
or (n1905,n1906,n2741);
and (n1906,n1907,n2740);
or (n1907,n1908,n2655);
and (n1908,n1909,n2654);
or (n1909,n1910,n2560);
and (n1910,n1911,n2559);
or (n1911,n1912,n2473);
and (n1912,n1913,n2472);
or (n1913,n1914,n2378);
and (n1914,n1915,n2377);
or (n1915,n1916,n2285);
and (n1916,n1917,n341);
or (n1917,n1918,n2191);
and (n1918,n1919,n2190);
or (n1919,n1920,n2103);
and (n1920,n1921,n488);
or (n1921,n1922,n2009);
and (n1922,n1923,n2008);
and (n1923,n890,n1924);
or (n1924,n1925,n1928);
and (n1925,n1926,n1927);
and (n1926,n46,n885);
and (n1927,n40,n413);
and (n1928,n1929,n1930);
xor (n1929,n1926,n1927);
or (n1930,n1931,n1933);
and (n1931,n1932,n1039);
and (n1932,n40,n885);
and (n1933,n1934,n1935);
xor (n1934,n1932,n1039);
or (n1935,n1936,n1938);
and (n1936,n1937,n1050);
and (n1937,n87,n885);
and (n1938,n1939,n1940);
xor (n1939,n1937,n1050);
or (n1940,n1941,n1943);
and (n1941,n1942,n1192);
and (n1942,n81,n885);
and (n1943,n1944,n1945);
xor (n1944,n1942,n1192);
or (n1945,n1946,n1948);
and (n1946,n1947,n1300);
and (n1947,n65,n885);
and (n1948,n1949,n1950);
xor (n1949,n1947,n1300);
or (n1950,n1951,n1954);
and (n1951,n1952,n1953);
and (n1952,n61,n885);
and (n1953,n103,n413);
and (n1954,n1955,n1956);
xor (n1955,n1952,n1953);
or (n1956,n1957,n1960);
and (n1957,n1958,n1959);
and (n1958,n103,n885);
and (n1959,n203,n413);
and (n1960,n1961,n1962);
xor (n1961,n1958,n1959);
or (n1962,n1963,n1965);
and (n1963,n1964,n1433);
and (n1964,n203,n885);
and (n1965,n1966,n1967);
xor (n1966,n1964,n1433);
or (n1967,n1968,n1971);
and (n1968,n1969,n1970);
and (n1969,n232,n885);
and (n1970,n226,n413);
and (n1971,n1972,n1973);
xor (n1972,n1969,n1970);
or (n1973,n1974,n1976);
and (n1974,n1975,n1522);
and (n1975,n226,n885);
and (n1976,n1977,n1978);
xor (n1977,n1975,n1522);
or (n1978,n1979,n1981);
and (n1979,n1980,n1570);
and (n1980,n310,n885);
and (n1981,n1982,n1983);
xor (n1982,n1980,n1570);
or (n1983,n1984,n1987);
and (n1984,n1985,n1986);
and (n1985,n334,n885);
and (n1986,n391,n413);
and (n1987,n1988,n1989);
xor (n1988,n1985,n1986);
or (n1989,n1990,n1993);
and (n1990,n1991,n1992);
and (n1991,n391,n885);
and (n1992,n443,n413);
and (n1993,n1994,n1995);
xor (n1994,n1991,n1992);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
and (n1997,n443,n885);
and (n1998,n715,n413);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2004);
and (n2002,n2003,n1764);
and (n2003,n715,n885);
and (n2004,n2005,n2006);
xor (n2005,n2003,n1764);
and (n2006,n2007,n1768);
and (n2007,n748,n885);
and (n2008,n46,n412);
and (n2009,n2010,n2011);
xor (n2010,n1923,n2008);
or (n2011,n2012,n2015);
and (n2012,n2013,n2014);
xor (n2013,n890,n1924);
and (n2014,n40,n412);
and (n2015,n2016,n2017);
xor (n2016,n2013,n2014);
or (n2017,n2018,n2021);
and (n2018,n2019,n2020);
xor (n2019,n1929,n1930);
and (n2020,n87,n412);
and (n2021,n2022,n2023);
xor (n2022,n2019,n2020);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
xor (n2025,n1934,n1935);
and (n2026,n81,n412);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1939,n1940);
and (n2032,n65,n412);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1944,n1945);
and (n2038,n61,n412);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
or (n2041,n2042,n2045);
and (n2042,n2043,n2044);
xor (n2043,n1949,n1950);
and (n2044,n103,n412);
and (n2045,n2046,n2047);
xor (n2046,n2043,n2044);
or (n2047,n2048,n2051);
and (n2048,n2049,n2050);
xor (n2049,n1955,n1956);
and (n2050,n203,n412);
and (n2051,n2052,n2053);
xor (n2052,n2049,n2050);
or (n2053,n2054,n2057);
and (n2054,n2055,n2056);
xor (n2055,n1961,n1962);
and (n2056,n232,n412);
and (n2057,n2058,n2059);
xor (n2058,n2055,n2056);
or (n2059,n2060,n2063);
and (n2060,n2061,n2062);
xor (n2061,n1966,n1967);
and (n2062,n226,n412);
and (n2063,n2064,n2065);
xor (n2064,n2061,n2062);
or (n2065,n2066,n2069);
and (n2066,n2067,n2068);
xor (n2067,n1972,n1973);
and (n2068,n310,n412);
and (n2069,n2070,n2071);
xor (n2070,n2067,n2068);
or (n2071,n2072,n2075);
and (n2072,n2073,n2074);
xor (n2073,n1977,n1978);
and (n2074,n334,n412);
and (n2075,n2076,n2077);
xor (n2076,n2073,n2074);
or (n2077,n2078,n2081);
and (n2078,n2079,n2080);
xor (n2079,n1982,n1983);
and (n2080,n391,n412);
and (n2081,n2082,n2083);
xor (n2082,n2079,n2080);
or (n2083,n2084,n2087);
and (n2084,n2085,n2086);
xor (n2085,n1988,n1989);
and (n2086,n443,n412);
and (n2087,n2088,n2089);
xor (n2088,n2085,n2086);
or (n2089,n2090,n2093);
and (n2090,n2091,n2092);
xor (n2091,n1994,n1995);
and (n2092,n715,n412);
and (n2093,n2094,n2095);
xor (n2094,n2091,n2092);
or (n2095,n2096,n2099);
and (n2096,n2097,n2098);
xor (n2097,n2000,n2001);
and (n2098,n748,n412);
and (n2099,n2100,n2101);
xor (n2100,n2097,n2098);
and (n2101,n2102,n1739);
xor (n2102,n2005,n2006);
and (n2103,n2104,n2105);
xor (n2104,n1921,n488);
or (n2105,n2106,n2109);
and (n2106,n2107,n2108);
xor (n2107,n2010,n2011);
and (n2108,n40,n244);
and (n2109,n2110,n2111);
xor (n2110,n2107,n2108);
or (n2111,n2112,n2114);
and (n2112,n2113,n839);
xor (n2113,n2016,n2017);
and (n2114,n2115,n2116);
xor (n2115,n2113,n839);
or (n2116,n2117,n2119);
and (n2117,n2118,n924);
xor (n2118,n2022,n2023);
and (n2119,n2120,n2121);
xor (n2120,n2118,n924);
or (n2121,n2122,n2124);
and (n2122,n2123,n1062);
xor (n2123,n2028,n2029);
and (n2124,n2125,n2126);
xor (n2125,n2123,n1062);
or (n2126,n2127,n2129);
and (n2127,n2128,n1057);
xor (n2128,n2034,n2035);
and (n2129,n2130,n2131);
xor (n2130,n2128,n1057);
or (n2131,n2132,n2134);
and (n2132,n2133,n1207);
xor (n2133,n2040,n2041);
and (n2134,n2135,n2136);
xor (n2135,n2133,n1207);
or (n2136,n2137,n2139);
and (n2137,n2138,n1276);
xor (n2138,n2046,n2047);
and (n2139,n2140,n2141);
xor (n2140,n2138,n1276);
or (n2141,n2142,n2145);
and (n2142,n2143,n2144);
xor (n2143,n2052,n2053);
and (n2144,n232,n244);
and (n2145,n2146,n2147);
xor (n2146,n2143,n2144);
or (n2147,n2148,n2151);
and (n2148,n2149,n2150);
xor (n2149,n2058,n2059);
and (n2150,n226,n244);
and (n2151,n2152,n2153);
xor (n2152,n2149,n2150);
or (n2153,n2154,n2157);
and (n2154,n2155,n2156);
xor (n2155,n2064,n2065);
and (n2156,n310,n244);
and (n2157,n2158,n2159);
xor (n2158,n2155,n2156);
or (n2159,n2160,n2163);
and (n2160,n2161,n2162);
xor (n2161,n2070,n2071);
and (n2162,n334,n244);
and (n2163,n2164,n2165);
xor (n2164,n2161,n2162);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2076,n2077);
and (n2168,n391,n244);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2174);
and (n2172,n2173,n1578);
xor (n2173,n2082,n2083);
and (n2174,n2175,n2176);
xor (n2175,n2173,n1578);
or (n2176,n2177,n2180);
and (n2177,n2178,n2179);
xor (n2178,n2088,n2089);
and (n2179,n715,n244);
and (n2180,n2181,n2182);
xor (n2181,n2178,n2179);
or (n2182,n2183,n2185);
and (n2183,n2184,n1712);
xor (n2184,n2094,n2095);
and (n2185,n2186,n2187);
xor (n2186,n2184,n1712);
and (n2187,n2188,n2189);
xor (n2188,n2100,n2101);
and (n2189,n808,n244);
and (n2190,n46,n242);
and (n2191,n2192,n2193);
xor (n2192,n1919,n2190);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
xor (n2195,n2104,n2105);
and (n2196,n40,n242);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2110,n2111);
and (n2202,n87,n242);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
xor (n2207,n2115,n2116);
and (n2208,n81,n242);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2215);
and (n2212,n2213,n2214);
xor (n2213,n2120,n2121);
and (n2214,n65,n242);
and (n2215,n2216,n2217);
xor (n2216,n2213,n2214);
or (n2217,n2218,n2221);
and (n2218,n2219,n2220);
xor (n2219,n2125,n2126);
and (n2220,n61,n242);
and (n2221,n2222,n2223);
xor (n2222,n2219,n2220);
or (n2223,n2224,n2227);
and (n2224,n2225,n2226);
xor (n2225,n2130,n2131);
and (n2226,n103,n242);
and (n2227,n2228,n2229);
xor (n2228,n2225,n2226);
or (n2229,n2230,n2233);
and (n2230,n2231,n2232);
xor (n2231,n2135,n2136);
and (n2232,n203,n242);
and (n2233,n2234,n2235);
xor (n2234,n2231,n2232);
or (n2235,n2236,n2239);
and (n2236,n2237,n2238);
xor (n2237,n2140,n2141);
and (n2238,n232,n242);
and (n2239,n2240,n2241);
xor (n2240,n2237,n2238);
or (n2241,n2242,n2245);
and (n2242,n2243,n2244);
xor (n2243,n2146,n2147);
and (n2244,n226,n242);
and (n2245,n2246,n2247);
xor (n2246,n2243,n2244);
or (n2247,n2248,n2251);
and (n2248,n2249,n2250);
xor (n2249,n2152,n2153);
and (n2250,n310,n242);
and (n2251,n2252,n2253);
xor (n2252,n2249,n2250);
or (n2253,n2254,n2257);
and (n2254,n2255,n2256);
xor (n2255,n2158,n2159);
and (n2256,n334,n242);
and (n2257,n2258,n2259);
xor (n2258,n2255,n2256);
or (n2259,n2260,n2263);
and (n2260,n2261,n2262);
xor (n2261,n2164,n2165);
and (n2262,n391,n242);
and (n2263,n2264,n2265);
xor (n2264,n2261,n2262);
or (n2265,n2266,n2269);
and (n2266,n2267,n2268);
xor (n2267,n2170,n2171);
and (n2268,n443,n242);
and (n2269,n2270,n2271);
xor (n2270,n2267,n2268);
or (n2271,n2272,n2275);
and (n2272,n2273,n2274);
xor (n2273,n2175,n2176);
and (n2274,n715,n242);
and (n2275,n2276,n2277);
xor (n2276,n2273,n2274);
or (n2277,n2278,n2281);
and (n2278,n2279,n2280);
xor (n2279,n2181,n2182);
and (n2280,n748,n242);
and (n2281,n2282,n2283);
xor (n2282,n2279,n2280);
and (n2283,n2284,n1668);
xor (n2284,n2186,n2187);
and (n2285,n2286,n2287);
xor (n2286,n1917,n341);
or (n2287,n2288,n2291);
and (n2288,n2289,n2290);
xor (n2289,n2192,n2193);
and (n2290,n40,n250);
and (n2291,n2292,n2293);
xor (n2292,n2289,n2290);
or (n2293,n2294,n2296);
and (n2294,n2295,n710);
xor (n2295,n2198,n2199);
and (n2296,n2297,n2298);
xor (n2297,n2295,n710);
or (n2298,n2299,n2302);
and (n2299,n2300,n2301);
xor (n2300,n2204,n2205);
and (n2301,n81,n250);
and (n2302,n2303,n2304);
xor (n2303,n2300,n2301);
or (n2304,n2305,n2308);
and (n2305,n2306,n2307);
xor (n2306,n2210,n2211);
and (n2307,n65,n250);
and (n2308,n2309,n2310);
xor (n2309,n2306,n2307);
or (n2310,n2311,n2313);
and (n2311,n2312,n935);
xor (n2312,n2216,n2217);
and (n2313,n2314,n2315);
xor (n2314,n2312,n935);
or (n2315,n2316,n2319);
and (n2316,n2317,n2318);
xor (n2317,n2222,n2223);
and (n2318,n103,n250);
and (n2319,n2320,n2321);
xor (n2320,n2317,n2318);
or (n2321,n2322,n2325);
and (n2322,n2323,n2324);
xor (n2323,n2228,n2229);
and (n2324,n203,n250);
and (n2325,n2326,n2327);
xor (n2326,n2323,n2324);
or (n2327,n2328,n2331);
and (n2328,n2329,n2330);
xor (n2329,n2234,n2235);
and (n2330,n232,n250);
and (n2331,n2332,n2333);
xor (n2332,n2329,n2330);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2240,n2241);
and (n2336,n226,n250);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
or (n2339,n2340,n2343);
and (n2340,n2341,n2342);
xor (n2341,n2246,n2247);
and (n2342,n310,n250);
and (n2343,n2344,n2345);
xor (n2344,n2341,n2342);
or (n2345,n2346,n2349);
and (n2346,n2347,n2348);
xor (n2347,n2252,n2253);
and (n2348,n334,n250);
and (n2349,n2350,n2351);
xor (n2350,n2347,n2348);
or (n2351,n2352,n2355);
and (n2352,n2353,n2354);
xor (n2353,n2258,n2259);
and (n2354,n391,n250);
and (n2355,n2356,n2357);
xor (n2356,n2353,n2354);
or (n2357,n2358,n2361);
and (n2358,n2359,n2360);
xor (n2359,n2264,n2265);
and (n2360,n443,n250);
and (n2361,n2362,n2363);
xor (n2362,n2359,n2360);
or (n2363,n2364,n2367);
and (n2364,n2365,n2366);
xor (n2365,n2270,n2271);
and (n2366,n715,n250);
and (n2367,n2368,n2369);
xor (n2368,n2365,n2366);
or (n2369,n2370,n2372);
and (n2370,n2371,n1660);
xor (n2371,n2276,n2277);
and (n2372,n2373,n2374);
xor (n2373,n2371,n1660);
and (n2374,n2375,n2376);
xor (n2375,n2282,n2283);
and (n2376,n808,n250);
and (n2377,n46,n262);
and (n2378,n2379,n2380);
xor (n2379,n1915,n2377);
or (n2380,n2381,n2384);
and (n2381,n2382,n2383);
xor (n2382,n2286,n2287);
and (n2383,n40,n262);
and (n2384,n2385,n2386);
xor (n2385,n2382,n2383);
or (n2386,n2387,n2390);
and (n2387,n2388,n2389);
xor (n2388,n2292,n2293);
and (n2389,n87,n262);
and (n2390,n2391,n2392);
xor (n2391,n2388,n2389);
or (n2392,n2393,n2396);
and (n2393,n2394,n2395);
xor (n2394,n2297,n2298);
and (n2395,n81,n262);
and (n2396,n2397,n2398);
xor (n2397,n2394,n2395);
or (n2398,n2399,n2402);
and (n2399,n2400,n2401);
xor (n2400,n2303,n2304);
and (n2401,n65,n262);
and (n2402,n2403,n2404);
xor (n2403,n2400,n2401);
or (n2404,n2405,n2408);
and (n2405,n2406,n2407);
xor (n2406,n2309,n2310);
and (n2407,n61,n262);
and (n2408,n2409,n2410);
xor (n2409,n2406,n2407);
or (n2410,n2411,n2414);
and (n2411,n2412,n2413);
xor (n2412,n2314,n2315);
and (n2413,n103,n262);
and (n2414,n2415,n2416);
xor (n2415,n2412,n2413);
or (n2416,n2417,n2420);
and (n2417,n2418,n2419);
xor (n2418,n2320,n2321);
and (n2419,n203,n262);
and (n2420,n2421,n2422);
xor (n2421,n2418,n2419);
or (n2422,n2423,n2426);
and (n2423,n2424,n2425);
xor (n2424,n2326,n2327);
and (n2425,n232,n262);
and (n2426,n2427,n2428);
xor (n2427,n2424,n2425);
or (n2428,n2429,n2432);
and (n2429,n2430,n2431);
xor (n2430,n2332,n2333);
and (n2431,n226,n262);
and (n2432,n2433,n2434);
xor (n2433,n2430,n2431);
or (n2434,n2435,n2438);
and (n2435,n2436,n2437);
xor (n2436,n2338,n2339);
and (n2437,n310,n262);
and (n2438,n2439,n2440);
xor (n2439,n2436,n2437);
or (n2440,n2441,n2444);
and (n2441,n2442,n2443);
xor (n2442,n2344,n2345);
and (n2443,n334,n262);
and (n2444,n2445,n2446);
xor (n2445,n2442,n2443);
or (n2446,n2447,n2450);
and (n2447,n2448,n2449);
xor (n2448,n2350,n2351);
and (n2449,n391,n262);
and (n2450,n2451,n2452);
xor (n2451,n2448,n2449);
or (n2452,n2453,n2456);
and (n2453,n2454,n2455);
xor (n2454,n2356,n2357);
and (n2455,n443,n262);
and (n2456,n2457,n2458);
xor (n2457,n2454,n2455);
or (n2458,n2459,n2462);
and (n2459,n2460,n2461);
xor (n2460,n2362,n2363);
and (n2461,n715,n262);
and (n2462,n2463,n2464);
xor (n2463,n2460,n2461);
or (n2464,n2465,n2468);
and (n2465,n2466,n2467);
xor (n2466,n2368,n2369);
and (n2467,n748,n262);
and (n2468,n2469,n2470);
xor (n2469,n2466,n2467);
and (n2470,n2471,n1514);
xor (n2471,n2373,n2374);
and (n2472,n46,n130);
and (n2473,n2474,n2475);
xor (n2474,n1913,n2472);
or (n2475,n2476,n2478);
and (n2476,n2477,n258);
xor (n2477,n2379,n2380);
and (n2478,n2479,n2480);
xor (n2479,n2477,n258);
or (n2480,n2481,n2483);
and (n2481,n2482,n351);
xor (n2482,n2385,n2386);
and (n2483,n2484,n2485);
xor (n2484,n2482,n351);
or (n2485,n2486,n2488);
and (n2486,n2487,n458);
xor (n2487,n2391,n2392);
and (n2488,n2489,n2490);
xor (n2489,n2487,n458);
or (n2490,n2491,n2493);
and (n2491,n2492,n672);
xor (n2492,n2397,n2398);
and (n2493,n2494,n2495);
xor (n2494,n2492,n672);
or (n2495,n2496,n2499);
and (n2496,n2497,n2498);
xor (n2497,n2403,n2404);
and (n2498,n61,n130);
and (n2499,n2500,n2501);
xor (n2500,n2497,n2498);
or (n2501,n2502,n2504);
and (n2502,n2503,n796);
xor (n2503,n2409,n2410);
and (n2504,n2505,n2506);
xor (n2505,n2503,n796);
or (n2506,n2507,n2510);
and (n2507,n2508,n2509);
xor (n2508,n2415,n2416);
and (n2509,n203,n130);
and (n2510,n2511,n2512);
xor (n2511,n2508,n2509);
or (n2512,n2513,n2515);
and (n2513,n2514,n1087);
xor (n2514,n2421,n2422);
and (n2515,n2516,n2517);
xor (n2516,n2514,n1087);
or (n2517,n2518,n2520);
and (n2518,n2519,n1123);
xor (n2519,n2427,n2428);
and (n2520,n2521,n2522);
xor (n2521,n2519,n1123);
or (n2522,n2523,n2526);
and (n2523,n2524,n2525);
xor (n2524,n2433,n2434);
and (n2525,n310,n130);
and (n2526,n2527,n2528);
xor (n2527,n2524,n2525);
or (n2528,n2529,n2532);
and (n2529,n2530,n2531);
xor (n2530,n2439,n2440);
and (n2531,n334,n130);
and (n2532,n2533,n2534);
xor (n2533,n2530,n2531);
or (n2534,n2535,n2538);
and (n2535,n2536,n2537);
xor (n2536,n2445,n2446);
and (n2537,n391,n130);
and (n2538,n2539,n2540);
xor (n2539,n2536,n2537);
or (n2540,n2541,n2543);
and (n2541,n2542,n1461);
xor (n2542,n2451,n2452);
and (n2543,n2544,n2545);
xor (n2544,n2542,n1461);
or (n2545,n2546,n2548);
and (n2546,n2547,n1446);
xor (n2547,n2457,n2458);
and (n2548,n2549,n2550);
xor (n2549,n2547,n1446);
or (n2550,n2551,n2554);
and (n2551,n2552,n2553);
xor (n2552,n2463,n2464);
and (n2553,n748,n130);
and (n2554,n2555,n2556);
xor (n2555,n2552,n2553);
and (n2556,n2557,n2558);
xor (n2557,n2469,n2470);
and (n2558,n808,n130);
and (n2559,n46,n131);
and (n2560,n2561,n2562);
xor (n2561,n1911,n2559);
or (n2562,n2563,n2566);
and (n2563,n2564,n2565);
xor (n2564,n2474,n2475);
and (n2565,n40,n131);
and (n2566,n2567,n2568);
xor (n2567,n2564,n2565);
or (n2568,n2569,n2572);
and (n2569,n2570,n2571);
xor (n2570,n2479,n2480);
and (n2571,n87,n131);
and (n2572,n2573,n2574);
xor (n2573,n2570,n2571);
or (n2574,n2575,n2578);
and (n2575,n2576,n2577);
xor (n2576,n2484,n2485);
and (n2577,n81,n131);
and (n2578,n2579,n2580);
xor (n2579,n2576,n2577);
or (n2580,n2581,n2584);
and (n2581,n2582,n2583);
xor (n2582,n2489,n2490);
and (n2583,n65,n131);
and (n2584,n2585,n2586);
xor (n2585,n2582,n2583);
or (n2586,n2587,n2590);
and (n2587,n2588,n2589);
xor (n2588,n2494,n2495);
and (n2589,n61,n131);
and (n2590,n2591,n2592);
xor (n2591,n2588,n2589);
or (n2592,n2593,n2596);
and (n2593,n2594,n2595);
xor (n2594,n2500,n2501);
and (n2595,n103,n131);
and (n2596,n2597,n2598);
xor (n2597,n2594,n2595);
or (n2598,n2599,n2602);
and (n2599,n2600,n2601);
xor (n2600,n2505,n2506);
and (n2601,n203,n131);
and (n2602,n2603,n2604);
xor (n2603,n2600,n2601);
or (n2604,n2605,n2608);
and (n2605,n2606,n2607);
xor (n2606,n2511,n2512);
and (n2607,n232,n131);
and (n2608,n2609,n2610);
xor (n2609,n2606,n2607);
or (n2610,n2611,n2614);
and (n2611,n2612,n2613);
xor (n2612,n2516,n2517);
and (n2613,n226,n131);
and (n2614,n2615,n2616);
xor (n2615,n2612,n2613);
or (n2616,n2617,n2620);
and (n2617,n2618,n2619);
xor (n2618,n2521,n2522);
and (n2619,n310,n131);
and (n2620,n2621,n2622);
xor (n2621,n2618,n2619);
or (n2622,n2623,n2626);
and (n2623,n2624,n2625);
xor (n2624,n2527,n2528);
and (n2625,n334,n131);
and (n2626,n2627,n2628);
xor (n2627,n2624,n2625);
or (n2628,n2629,n2632);
and (n2629,n2630,n2631);
xor (n2630,n2533,n2534);
and (n2631,n391,n131);
and (n2632,n2633,n2634);
xor (n2633,n2630,n2631);
or (n2634,n2635,n2638);
and (n2635,n2636,n2637);
xor (n2636,n2539,n2540);
and (n2637,n443,n131);
and (n2638,n2639,n2640);
xor (n2639,n2636,n2637);
or (n2640,n2641,n2644);
and (n2641,n2642,n2643);
xor (n2642,n2544,n2545);
and (n2643,n715,n131);
and (n2644,n2645,n2646);
xor (n2645,n2642,n2643);
or (n2646,n2647,n2650);
and (n2647,n2648,n2649);
xor (n2648,n2549,n2550);
and (n2649,n748,n131);
and (n2650,n2651,n2652);
xor (n2651,n2648,n2649);
and (n2652,n2653,n1412);
xor (n2653,n2555,n2556);
and (n2654,n46,n18);
and (n2655,n2656,n2657);
xor (n2656,n1909,n2654);
or (n2657,n2658,n2661);
and (n2658,n2659,n2660);
xor (n2659,n2561,n2562);
and (n2660,n40,n18);
and (n2661,n2662,n2663);
xor (n2662,n2659,n2660);
or (n2663,n2664,n2666);
and (n2664,n2665,n219);
xor (n2665,n2567,n2568);
and (n2666,n2667,n2668);
xor (n2667,n2665,n219);
or (n2668,n2669,n2672);
and (n2669,n2670,n2671);
xor (n2670,n2573,n2574);
and (n2671,n81,n18);
and (n2672,n2673,n2674);
xor (n2673,n2670,n2671);
or (n2674,n2675,n2677);
and (n2675,n2676,n379);
xor (n2676,n2579,n2580);
and (n2677,n2678,n2679);
xor (n2678,n2676,n379);
or (n2679,n2680,n2682);
and (n2680,n2681,n434);
xor (n2681,n2585,n2586);
and (n2682,n2683,n2684);
xor (n2683,n2681,n434);
or (n2684,n2685,n2687);
and (n2685,n2686,n722);
xor (n2686,n2591,n2592);
and (n2687,n2688,n2689);
xor (n2688,n2686,n722);
or (n2689,n2690,n2692);
and (n2690,n2691,n765);
xor (n2691,n2597,n2598);
and (n2692,n2693,n2694);
xor (n2693,n2691,n765);
or (n2694,n2695,n2697);
and (n2695,n2696,n846);
xor (n2696,n2603,n2604);
and (n2697,n2698,n2699);
xor (n2698,n2696,n846);
or (n2699,n2700,n2702);
and (n2700,n2701,n974);
xor (n2701,n2609,n2610);
and (n2702,n2703,n2704);
xor (n2703,n2701,n974);
or (n2704,n2705,n2707);
and (n2705,n2706,n1097);
xor (n2706,n2615,n2616);
and (n2707,n2708,n2709);
xor (n2708,n2706,n1097);
or (n2709,n2710,n2713);
and (n2710,n2711,n2712);
xor (n2711,n2621,n2622);
and (n2712,n334,n18);
and (n2713,n2714,n2715);
xor (n2714,n2711,n2712);
or (n2715,n2716,n2718);
and (n2716,n2717,n1221);
xor (n2717,n2627,n2628);
and (n2718,n2719,n2720);
xor (n2719,n2717,n1221);
or (n2720,n2721,n2724);
and (n2721,n2722,n2723);
xor (n2722,n2633,n2634);
and (n2723,n443,n18);
and (n2724,n2725,n2726);
xor (n2725,n2722,n2723);
or (n2726,n2727,n2730);
and (n2727,n2728,n2729);
xor (n2728,n2639,n2640);
and (n2729,n715,n18);
and (n2730,n2731,n2732);
xor (n2731,n2728,n2729);
or (n2732,n2733,n2735);
and (n2733,n2734,n1374);
xor (n2734,n2645,n2646);
and (n2735,n2736,n2737);
xor (n2736,n2734,n1374);
and (n2737,n2738,n2739);
xor (n2738,n2651,n2652);
and (n2739,n808,n18);
and (n2740,n46,n17);
and (n2741,n2742,n2743);
xor (n2742,n1907,n2740);
or (n2743,n2744,n2747);
and (n2744,n2745,n2746);
xor (n2745,n2656,n2657);
and (n2746,n40,n17);
and (n2747,n2748,n2749);
xor (n2748,n2745,n2746);
or (n2749,n2750,n2753);
and (n2750,n2751,n2752);
xor (n2751,n2662,n2663);
and (n2752,n87,n17);
and (n2753,n2754,n2755);
xor (n2754,n2751,n2752);
or (n2755,n2756,n2759);
and (n2756,n2757,n2758);
xor (n2757,n2667,n2668);
and (n2758,n81,n17);
and (n2759,n2760,n2761);
xor (n2760,n2757,n2758);
or (n2761,n2762,n2765);
and (n2762,n2763,n2764);
xor (n2763,n2673,n2674);
and (n2764,n65,n17);
and (n2765,n2766,n2767);
xor (n2766,n2763,n2764);
or (n2767,n2768,n2771);
and (n2768,n2769,n2770);
xor (n2769,n2678,n2679);
and (n2770,n61,n17);
and (n2771,n2772,n2773);
xor (n2772,n2769,n2770);
or (n2773,n2774,n2777);
and (n2774,n2775,n2776);
xor (n2775,n2683,n2684);
and (n2776,n103,n17);
and (n2777,n2778,n2779);
xor (n2778,n2775,n2776);
or (n2779,n2780,n2783);
and (n2780,n2781,n2782);
xor (n2781,n2688,n2689);
and (n2782,n203,n17);
and (n2783,n2784,n2785);
xor (n2784,n2781,n2782);
or (n2785,n2786,n2789);
and (n2786,n2787,n2788);
xor (n2787,n2693,n2694);
and (n2788,n232,n17);
and (n2789,n2790,n2791);
xor (n2790,n2787,n2788);
or (n2791,n2792,n2795);
and (n2792,n2793,n2794);
xor (n2793,n2698,n2699);
and (n2794,n226,n17);
and (n2795,n2796,n2797);
xor (n2796,n2793,n2794);
or (n2797,n2798,n2801);
and (n2798,n2799,n2800);
xor (n2799,n2703,n2704);
and (n2800,n310,n17);
and (n2801,n2802,n2803);
xor (n2802,n2799,n2800);
or (n2803,n2804,n2807);
and (n2804,n2805,n2806);
xor (n2805,n2708,n2709);
and (n2806,n334,n17);
and (n2807,n2808,n2809);
xor (n2808,n2805,n2806);
or (n2809,n2810,n2813);
and (n2810,n2811,n2812);
xor (n2811,n2714,n2715);
and (n2812,n391,n17);
and (n2813,n2814,n2815);
xor (n2814,n2811,n2812);
or (n2815,n2816,n2819);
and (n2816,n2817,n2818);
xor (n2817,n2719,n2720);
and (n2818,n443,n17);
and (n2819,n2820,n2821);
xor (n2820,n2817,n2818);
or (n2821,n2822,n2825);
and (n2822,n2823,n2824);
xor (n2823,n2725,n2726);
and (n2824,n715,n17);
and (n2825,n2826,n2827);
xor (n2826,n2823,n2824);
or (n2827,n2828,n2831);
and (n2828,n2829,n2830);
xor (n2829,n2731,n2732);
and (n2830,n748,n17);
and (n2831,n2832,n2833);
xor (n2832,n2829,n2830);
and (n2833,n2834,n1616);
xor (n2834,n2736,n2737);
and (n2835,n46,n22);
and (n2836,n2837,n2838);
xor (n2837,n1905,n2835);
or (n2838,n2839,n2842);
and (n2839,n2840,n2841);
xor (n2840,n2742,n2743);
and (n2841,n40,n22);
and (n2842,n2843,n2844);
xor (n2843,n2840,n2841);
or (n2844,n2845,n2847);
and (n2845,n2846,n540);
xor (n2846,n2748,n2749);
and (n2847,n2848,n2849);
xor (n2848,n2846,n540);
or (n2849,n2850,n2852);
and (n2850,n2851,n318);
xor (n2851,n2754,n2755);
and (n2852,n2853,n2854);
xor (n2853,n2851,n318);
or (n2854,n2855,n2858);
and (n2855,n2856,n2857);
xor (n2856,n2760,n2761);
and (n2857,n65,n22);
and (n2858,n2859,n2860);
xor (n2859,n2856,n2857);
or (n2860,n2861,n2863);
and (n2861,n2862,n278);
xor (n2862,n2766,n2767);
and (n2863,n2864,n2865);
xor (n2864,n2862,n278);
or (n2865,n2866,n2868);
and (n2866,n2867,n358);
xor (n2867,n2772,n2773);
and (n2868,n2869,n2870);
xor (n2869,n2867,n358);
or (n2870,n2871,n2873);
and (n2871,n2872,n450);
xor (n2872,n2778,n2779);
and (n2873,n2874,n2875);
xor (n2874,n2872,n450);
or (n2875,n2876,n2879);
and (n2876,n2877,n2878);
xor (n2877,n2784,n2785);
and (n2878,n232,n22);
and (n2879,n2880,n2881);
xor (n2880,n2877,n2878);
or (n2881,n2882,n2885);
and (n2882,n2883,n2884);
xor (n2883,n2790,n2791);
and (n2884,n226,n22);
and (n2885,n2886,n2887);
xor (n2886,n2883,n2884);
or (n2887,n2888,n2891);
and (n2888,n2889,n2890);
xor (n2889,n2796,n2797);
and (n2890,n310,n22);
and (n2891,n2892,n2893);
xor (n2892,n2889,n2890);
or (n2893,n2894,n2897);
and (n2894,n2895,n2896);
xor (n2895,n2802,n2803);
and (n2896,n334,n22);
and (n2897,n2898,n2899);
xor (n2898,n2895,n2896);
or (n2899,n2900,n2903);
and (n2900,n2901,n2902);
xor (n2901,n2808,n2809);
and (n2902,n391,n22);
and (n2903,n2904,n2905);
xor (n2904,n2901,n2902);
or (n2905,n2906,n2909);
and (n2906,n2907,n2908);
xor (n2907,n2814,n2815);
and (n2908,n443,n22);
and (n2909,n2910,n2911);
xor (n2910,n2907,n2908);
or (n2911,n2912,n2914);
and (n2912,n2913,n1238);
xor (n2913,n2820,n2821);
and (n2914,n2915,n2916);
xor (n2915,n2913,n1238);
or (n2916,n2917,n2920);
and (n2917,n2918,n2919);
xor (n2918,n2826,n2827);
and (n2919,n748,n22);
and (n2920,n2921,n2922);
xor (n2921,n2918,n2919);
and (n2922,n2923,n2924);
xor (n2923,n2832,n2833);
and (n2924,n808,n22);
and (n2925,n46,n31);
and (n2926,n2927,n2928);
xor (n2927,n1903,n2925);
or (n2928,n2929,n2932);
and (n2929,n2930,n2931);
xor (n2930,n2837,n2838);
and (n2931,n40,n31);
and (n2932,n2933,n2934);
xor (n2933,n2930,n2931);
or (n2934,n2935,n2938);
and (n2935,n2936,n2937);
xor (n2936,n2843,n2844);
and (n2937,n87,n31);
and (n2938,n2939,n2940);
xor (n2939,n2936,n2937);
or (n2940,n2941,n2944);
and (n2941,n2942,n2943);
xor (n2942,n2848,n2849);
and (n2943,n81,n31);
and (n2944,n2945,n2946);
xor (n2945,n2942,n2943);
or (n2946,n2947,n2950);
and (n2947,n2948,n2949);
xor (n2948,n2853,n2854);
and (n2949,n65,n31);
and (n2950,n2951,n2952);
xor (n2951,n2948,n2949);
or (n2952,n2953,n2956);
and (n2953,n2954,n2955);
xor (n2954,n2859,n2860);
and (n2955,n61,n31);
and (n2956,n2957,n2958);
xor (n2957,n2954,n2955);
or (n2958,n2959,n2962);
and (n2959,n2960,n2961);
xor (n2960,n2864,n2865);
and (n2961,n103,n31);
and (n2962,n2963,n2964);
xor (n2963,n2960,n2961);
or (n2964,n2965,n2968);
and (n2965,n2966,n2967);
xor (n2966,n2869,n2870);
and (n2967,n203,n31);
and (n2968,n2969,n2970);
xor (n2969,n2966,n2967);
or (n2970,n2971,n2974);
and (n2971,n2972,n2973);
xor (n2972,n2874,n2875);
and (n2973,n232,n31);
and (n2974,n2975,n2976);
xor (n2975,n2972,n2973);
or (n2976,n2977,n2980);
and (n2977,n2978,n2979);
xor (n2978,n2880,n2881);
and (n2979,n226,n31);
and (n2980,n2981,n2982);
xor (n2981,n2978,n2979);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
xor (n2984,n2886,n2887);
and (n2985,n310,n31);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
or (n2988,n2989,n2992);
and (n2989,n2990,n2991);
xor (n2990,n2892,n2893);
and (n2991,n334,n31);
and (n2992,n2993,n2994);
xor (n2993,n2990,n2991);
or (n2994,n2995,n2998);
and (n2995,n2996,n2997);
xor (n2996,n2898,n2899);
and (n2997,n391,n31);
and (n2998,n2999,n3000);
xor (n2999,n2996,n2997);
or (n3000,n3001,n3004);
and (n3001,n3002,n3003);
xor (n3002,n2904,n2905);
and (n3003,n443,n31);
and (n3004,n3005,n3006);
xor (n3005,n3002,n3003);
or (n3006,n3007,n3010);
and (n3007,n3008,n3009);
xor (n3008,n2910,n2911);
and (n3009,n715,n31);
and (n3010,n3011,n3012);
xor (n3011,n3008,n3009);
or (n3012,n3013,n3016);
and (n3013,n3014,n3015);
xor (n3014,n2915,n2916);
and (n3015,n748,n31);
and (n3016,n3017,n3018);
xor (n3017,n3014,n3015);
and (n3018,n3019,n3020);
xor (n3019,n2921,n2922);
not (n3020,n1185);
and (n3021,n46,n36);
or (n3022,n3023,n3026);
and (n3023,n3024,n3025);
xor (n3024,n2927,n2928);
and (n3025,n40,n36);
and (n3026,n3027,n3028);
xor (n3027,n3024,n3025);
or (n3028,n3029,n3032);
and (n3029,n3030,n3031);
xor (n3030,n2933,n2934);
and (n3031,n87,n36);
and (n3032,n3033,n3034);
xor (n3033,n3030,n3031);
or (n3034,n3035,n3038);
and (n3035,n3036,n3037);
xor (n3036,n2939,n2940);
and (n3037,n81,n36);
and (n3038,n3039,n3040);
xor (n3039,n3036,n3037);
or (n3040,n3041,n3044);
and (n3041,n3042,n3043);
xor (n3042,n2945,n2946);
and (n3043,n65,n36);
and (n3044,n3045,n3046);
xor (n3045,n3042,n3043);
or (n3046,n3047,n3050);
and (n3047,n3048,n3049);
xor (n3048,n2951,n2952);
and (n3049,n61,n36);
and (n3050,n3051,n3052);
xor (n3051,n3048,n3049);
or (n3052,n3053,n3055);
and (n3053,n3054,n208);
xor (n3054,n2957,n2958);
and (n3055,n3056,n3057);
xor (n3056,n3054,n208);
or (n3057,n3058,n3061);
and (n3058,n3059,n3060);
xor (n3059,n2963,n2964);
and (n3060,n203,n36);
and (n3061,n3062,n3063);
xor (n3062,n3059,n3060);
or (n3063,n3064,n3066);
and (n3064,n3065,n365);
xor (n3065,n2969,n2970);
and (n3066,n3067,n3068);
xor (n3067,n3065,n365);
or (n3068,n3069,n3071);
and (n3069,n3070,n474);
xor (n3070,n2975,n2976);
and (n3071,n3072,n3073);
xor (n3072,n3070,n474);
or (n3073,n3074,n3077);
and (n3074,n3075,n3076);
xor (n3075,n2981,n2982);
and (n3076,n310,n36);
and (n3077,n3078,n3079);
xor (n3078,n3075,n3076);
or (n3079,n3080,n3083);
and (n3080,n3081,n3082);
xor (n3081,n2987,n2988);
and (n3082,n334,n36);
and (n3083,n3084,n3085);
xor (n3084,n3081,n3082);
or (n3085,n3086,n3089);
and (n3086,n3087,n3088);
xor (n3087,n2993,n2994);
and (n3088,n391,n36);
and (n3089,n3090,n3091);
xor (n3090,n3087,n3088);
or (n3091,n3092,n3095);
and (n3092,n3093,n3094);
xor (n3093,n2999,n3000);
and (n3094,n443,n36);
and (n3095,n3096,n3097);
xor (n3096,n3093,n3094);
or (n3097,n3098,n3101);
and (n3098,n3099,n3100);
xor (n3099,n3005,n3006);
and (n3100,n715,n36);
and (n3101,n3102,n3103);
xor (n3102,n3099,n3100);
or (n3103,n3104,n3107);
and (n3104,n3105,n3106);
xor (n3105,n3011,n3012);
and (n3106,n748,n36);
and (n3107,n3108,n3109);
xor (n3108,n3105,n3106);
and (n3109,n3110,n3111);
xor (n3110,n3017,n3018);
and (n3111,n808,n36);
and (n3112,n40,n74);
or (n3113,n3114,n3117);
and (n3114,n3115,n3116);
xor (n3115,n3027,n3028);
and (n3116,n87,n74);
and (n3117,n3118,n3119);
xor (n3118,n3115,n3116);
or (n3119,n3120,n3123);
and (n3120,n3121,n3122);
xor (n3121,n3033,n3034);
and (n3122,n81,n74);
and (n3123,n3124,n3125);
xor (n3124,n3121,n3122);
or (n3125,n3126,n3129);
and (n3126,n3127,n3128);
xor (n3127,n3039,n3040);
and (n3128,n65,n74);
and (n3129,n3130,n3131);
xor (n3130,n3127,n3128);
or (n3131,n3132,n3135);
and (n3132,n3133,n3134);
xor (n3133,n3045,n3046);
and (n3134,n61,n74);
and (n3135,n3136,n3137);
xor (n3136,n3133,n3134);
or (n3137,n3138,n3141);
and (n3138,n3139,n3140);
xor (n3139,n3051,n3052);
and (n3140,n103,n74);
and (n3141,n3142,n3143);
xor (n3142,n3139,n3140);
or (n3143,n3144,n3147);
and (n3144,n3145,n3146);
xor (n3145,n3056,n3057);
and (n3146,n203,n74);
and (n3147,n3148,n3149);
xor (n3148,n3145,n3146);
or (n3149,n3150,n3153);
and (n3150,n3151,n3152);
xor (n3151,n3062,n3063);
and (n3152,n232,n74);
and (n3153,n3154,n3155);
xor (n3154,n3151,n3152);
or (n3155,n3156,n3159);
and (n3156,n3157,n3158);
xor (n3157,n3067,n3068);
and (n3158,n226,n74);
and (n3159,n3160,n3161);
xor (n3160,n3157,n3158);
or (n3161,n3162,n3165);
and (n3162,n3163,n3164);
xor (n3163,n3072,n3073);
and (n3164,n310,n74);
and (n3165,n3166,n3167);
xor (n3166,n3163,n3164);
or (n3167,n3168,n3171);
and (n3168,n3169,n3170);
xor (n3169,n3078,n3079);
and (n3170,n334,n74);
and (n3171,n3172,n3173);
xor (n3172,n3169,n3170);
or (n3173,n3174,n3177);
and (n3174,n3175,n3176);
xor (n3175,n3084,n3085);
and (n3176,n391,n74);
and (n3177,n3178,n3179);
xor (n3178,n3175,n3176);
or (n3179,n3180,n3183);
and (n3180,n3181,n3182);
xor (n3181,n3090,n3091);
and (n3182,n443,n74);
and (n3183,n3184,n3185);
xor (n3184,n3181,n3182);
or (n3185,n3186,n3189);
and (n3186,n3187,n3188);
xor (n3187,n3096,n3097);
and (n3188,n715,n74);
and (n3189,n3190,n3191);
xor (n3190,n3187,n3188);
or (n3191,n3192,n3195);
and (n3192,n3193,n3194);
xor (n3193,n3102,n3103);
and (n3194,n748,n74);
and (n3195,n3196,n3197);
xor (n3196,n3193,n3194);
and (n3197,n3198,n3199);
xor (n3198,n3108,n3109);
not (n3199,n1031);
and (n3200,n87,n56);
or (n3201,n3202,n3205);
and (n3202,n3203,n3204);
xor (n3203,n3118,n3119);
and (n3204,n81,n56);
and (n3205,n3206,n3207);
xor (n3206,n3203,n3204);
or (n3207,n3208,n3211);
and (n3208,n3209,n3210);
xor (n3209,n3124,n3125);
and (n3210,n65,n56);
and (n3211,n3212,n3213);
xor (n3212,n3209,n3210);
or (n3213,n3214,n3217);
and (n3214,n3215,n3216);
xor (n3215,n3130,n3131);
and (n3216,n61,n56);
and (n3217,n3218,n3219);
xor (n3218,n3215,n3216);
or (n3219,n3220,n3222);
and (n3220,n3221,n534);
xor (n3221,n3136,n3137);
and (n3222,n3223,n3224);
xor (n3223,n3221,n534);
or (n3224,n3225,n3227);
and (n3225,n3226,n297);
xor (n3226,n3142,n3143);
and (n3227,n3228,n3229);
xor (n3228,n3226,n297);
or (n3229,n3230,n3233);
and (n3230,n3231,n3232);
xor (n3231,n3148,n3149);
and (n3232,n232,n56);
and (n3233,n3234,n3235);
xor (n3234,n3231,n3232);
or (n3235,n3236,n3238);
and (n3236,n3237,n227);
xor (n3237,n3154,n3155);
and (n3238,n3239,n3240);
xor (n3239,n3237,n227);
or (n3240,n3241,n3243);
and (n3241,n3242,n386);
xor (n3242,n3160,n3161);
and (n3243,n3244,n3245);
xor (n3244,n3242,n386);
or (n3245,n3246,n3248);
and (n3246,n3247,n481);
xor (n3247,n3166,n3167);
and (n3248,n3249,n3250);
xor (n3249,n3247,n481);
or (n3250,n3251,n3253);
and (n3251,n3252,n661);
xor (n3252,n3172,n3173);
and (n3253,n3254,n3255);
xor (n3254,n3252,n661);
or (n3255,n3256,n3259);
and (n3256,n3257,n3258);
xor (n3257,n3178,n3179);
and (n3258,n443,n56);
and (n3259,n3260,n3261);
xor (n3260,n3257,n3258);
or (n3261,n3262,n3265);
and (n3262,n3263,n3264);
xor (n3263,n3184,n3185);
and (n3264,n715,n56);
and (n3265,n3266,n3267);
xor (n3266,n3263,n3264);
or (n3267,n3268,n3270);
and (n3268,n3269,n960);
xor (n3269,n3190,n3191);
and (n3270,n3271,n3272);
xor (n3271,n3269,n960);
and (n3272,n3273,n3274);
xor (n3273,n3196,n3197);
and (n3274,n808,n56);
and (n3275,n81,n57);
or (n3276,n3277,n3280);
and (n3277,n3278,n3279);
xor (n3278,n3206,n3207);
and (n3279,n65,n57);
and (n3280,n3281,n3282);
xor (n3281,n3278,n3279);
or (n3282,n3283,n3286);
and (n3283,n3284,n3285);
xor (n3284,n3212,n3213);
and (n3285,n61,n57);
and (n3286,n3287,n3288);
xor (n3287,n3284,n3285);
or (n3288,n3289,n3292);
and (n3289,n3290,n3291);
xor (n3290,n3218,n3219);
and (n3291,n103,n57);
and (n3292,n3293,n3294);
xor (n3293,n3290,n3291);
or (n3294,n3295,n3298);
and (n3295,n3296,n3297);
xor (n3296,n3223,n3224);
and (n3297,n203,n57);
and (n3298,n3299,n3300);
xor (n3299,n3296,n3297);
or (n3300,n3301,n3304);
and (n3301,n3302,n3303);
xor (n3302,n3228,n3229);
and (n3303,n232,n57);
and (n3304,n3305,n3306);
xor (n3305,n3302,n3303);
or (n3306,n3307,n3310);
and (n3307,n3308,n3309);
xor (n3308,n3234,n3235);
and (n3309,n226,n57);
and (n3310,n3311,n3312);
xor (n3311,n3308,n3309);
or (n3312,n3313,n3316);
and (n3313,n3314,n3315);
xor (n3314,n3239,n3240);
and (n3315,n310,n57);
and (n3316,n3317,n3318);
xor (n3317,n3314,n3315);
or (n3318,n3319,n3322);
and (n3319,n3320,n3321);
xor (n3320,n3244,n3245);
and (n3321,n334,n57);
and (n3322,n3323,n3324);
xor (n3323,n3320,n3321);
or (n3324,n3325,n3328);
and (n3325,n3326,n3327);
xor (n3326,n3249,n3250);
and (n3327,n391,n57);
and (n3328,n3329,n3330);
xor (n3329,n3326,n3327);
or (n3330,n3331,n3334);
and (n3331,n3332,n3333);
xor (n3332,n3254,n3255);
and (n3333,n443,n57);
and (n3334,n3335,n3336);
xor (n3335,n3332,n3333);
or (n3336,n3337,n3340);
and (n3337,n3338,n3339);
xor (n3338,n3260,n3261);
and (n3339,n715,n57);
and (n3340,n3341,n3342);
xor (n3341,n3338,n3339);
or (n3342,n3343,n3346);
and (n3343,n3344,n3345);
xor (n3344,n3266,n3267);
and (n3345,n748,n57);
and (n3346,n3347,n3348);
xor (n3347,n3344,n3345);
and (n3348,n3349,n3350);
xor (n3349,n3271,n3272);
and (n3350,n808,n57);
endmodule
