module top (out,n19,n20,n25,n29,n36,n46,n48,n53,n59
        ,n65,n73,n79,n83,n89,n98,n99,n103,n107,n109
        ,n113,n120,n127,n136,n142,n152,n160,n166,n174,n180
        ,n184,n190,n199,n207,n214);
output out;
input n19;
input n20;
input n25;
input n29;
input n36;
input n46;
input n48;
input n53;
input n59;
input n65;
input n73;
input n79;
input n83;
input n89;
input n98;
input n99;
input n103;
input n107;
input n109;
input n113;
input n120;
input n127;
input n136;
input n142;
input n152;
input n160;
input n166;
input n174;
input n180;
input n184;
input n190;
input n199;
input n207;
input n214;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n108;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
xor (out,n0,n1012);
nand (n0,n1,n1011);
or (n1,n2,n488);
not (n2,n3);
nand (n3,n4,n487);
not (n4,n5);
nor (n5,n6,n428);
xor (n6,n7,n362);
xor (n7,n8,n217);
xor (n8,n9,n145);
xor (n9,n10,n92);
xor (n10,n11,n68);
xor (n11,n12,n39);
nand (n12,n13,n32);
or (n13,n14,n27);
not (n14,n15);
nor (n15,n16,n22);
nand (n16,n17,n21);
or (n17,n18,n20);
not (n18,n19);
nand (n21,n20,n18);
nor (n22,n23,n26);
and (n23,n24,n19);
not (n24,n25);
and (n26,n25,n18);
nor (n27,n28,n30);
and (n28,n24,n29);
and (n30,n25,n31);
not (n31,n29);
or (n32,n33,n34);
not (n33,n16);
nor (n34,n35,n37);
and (n35,n24,n36);
and (n37,n25,n38);
not (n38,n36);
nand (n39,n40,n62);
or (n40,n41,n57);
not (n41,n42);
nor (n42,n43,n50);
not (n43,n44);
nand (n44,n45,n49);
or (n45,n46,n47);
not (n47,n48);
nand (n49,n47,n46);
not (n50,n51);
nor (n51,n52,n55);
and (n52,n53,n54);
not (n54,n46);
and (n55,n56,n46);
not (n56,n53);
nor (n57,n58,n60);
and (n58,n47,n59);
and (n60,n48,n61);
not (n61,n59);
or (n62,n51,n63);
nor (n63,n64,n66);
and (n64,n47,n65);
and (n66,n48,n67);
not (n67,n65);
nand (n68,n69,n86);
or (n69,n70,n81);
nand (n70,n71,n76);
nor (n71,n72,n74);
and (n72,n47,n73);
and (n74,n48,n75);
not (n75,n73);
nand (n76,n77,n80);
or (n77,n73,n78);
not (n78,n79);
nand (n80,n78,n73);
nor (n81,n82,n84);
and (n82,n78,n83);
and (n84,n79,n85);
not (n85,n83);
or (n86,n71,n87);
nor (n87,n88,n90);
and (n88,n78,n89);
and (n90,n79,n91);
not (n91,n89);
xor (n92,n93,n122);
xor (n93,n94,n104);
nor (n94,n95,n102);
nor (n95,n96,n100);
and (n96,n97,n99);
not (n97,n98);
and (n100,n98,n101);
not (n101,n99);
not (n102,n103);
nand (n104,n105,n116);
or (n105,n106,n110);
nand (n106,n107,n108);
not (n108,n109);
nor (n110,n111,n114);
and (n111,n112,n113);
not (n112,n107);
and (n114,n107,n115);
not (n115,n113);
or (n116,n117,n108);
nor (n117,n118,n121);
and (n118,n119,n107);
not (n119,n120);
and (n121,n120,n112);
nand (n122,n123,n139);
or (n123,n124,n134);
nand (n124,n125,n130);
nor (n125,n126,n128);
and (n126,n112,n127);
and (n128,n107,n129);
not (n129,n127);
nand (n130,n131,n133);
or (n131,n127,n132);
not (n132,n20);
nand (n133,n132,n127);
nor (n134,n135,n137);
and (n135,n132,n136);
and (n137,n20,n138);
not (n138,n136);
or (n139,n125,n140);
nor (n140,n141,n143);
and (n141,n132,n142);
and (n143,n20,n144);
not (n144,n142);
xor (n145,n146,n193);
xor (n146,n147,n169);
nand (n147,n148,n163);
or (n148,n149,n158);
nand (n149,n150,n155);
nor (n150,n151,n153);
and (n151,n78,n152);
and (n153,n79,n154);
not (n154,n152);
nand (n155,n156,n157);
or (n156,n152,n97);
nand (n157,n97,n152);
nor (n158,n159,n161);
and (n159,n97,n160);
and (n161,n98,n162);
not (n162,n160);
or (n163,n150,n164);
nor (n164,n165,n167);
and (n165,n97,n166);
and (n167,n98,n168);
not (n168,n166);
nand (n169,n170,n187);
or (n170,n171,n182);
nand (n171,n172,n177);
nor (n172,n173,n175);
and (n173,n24,n174);
and (n175,n25,n176);
not (n176,n174);
nand (n177,n178,n181);
or (n178,n174,n179);
not (n179,n180);
nand (n181,n179,n174);
nor (n182,n183,n185);
and (n183,n179,n184);
and (n185,n180,n186);
not (n186,n184);
or (n187,n172,n188);
nor (n188,n189,n191);
and (n189,n179,n190);
and (n191,n180,n192);
not (n192,n190);
nand (n193,n194,n210);
or (n194,n195,n205);
not (n195,n196);
nor (n196,n197,n201);
nand (n197,n198,n200);
or (n198,n199,n179);
nand (n200,n199,n179);
nor (n201,n202,n203);
and (n202,n56,n199);
and (n203,n53,n204);
not (n204,n199);
nor (n205,n206,n208);
and (n206,n56,n207);
and (n208,n53,n209);
not (n209,n207);
or (n210,n211,n212);
not (n211,n197);
nor (n212,n213,n215);
and (n213,n56,n214);
and (n215,n53,n216);
not (n216,n214);
or (n217,n218,n361);
and (n218,n219,n293);
xor (n219,n220,n258);
or (n220,n221,n257);
and (n221,n222,n241);
xor (n222,n223,n232);
nand (n223,n224,n228);
or (n224,n41,n225);
nor (n225,n226,n227);
and (n226,n47,n83);
and (n227,n48,n85);
or (n228,n51,n229);
nor (n229,n230,n231);
and (n230,n47,n89);
and (n231,n48,n91);
nand (n232,n233,n237);
or (n233,n70,n234);
nor (n234,n235,n236);
and (n235,n78,n160);
and (n236,n79,n162);
or (n237,n71,n238);
nor (n238,n239,n240);
and (n239,n78,n166);
and (n240,n79,n168);
and (n241,n242,n248);
nor (n242,n243,n78);
nor (n243,n244,n247);
and (n244,n245,n47);
not (n245,n246);
and (n246,n103,n73);
and (n247,n102,n75);
nand (n248,n249,n253);
or (n249,n106,n250);
nor (n250,n251,n252);
and (n251,n112,n36);
and (n252,n107,n38);
or (n253,n254,n108);
nor (n254,n255,n256);
and (n255,n138,n107);
and (n256,n136,n112);
and (n257,n223,n232);
xor (n258,n259,n276);
xor (n259,n260,n263);
nand (n260,n261,n262);
or (n261,n70,n238);
or (n262,n71,n81);
xor (n263,n264,n270);
nor (n264,n265,n97);
nor (n265,n266,n269);
and (n266,n267,n78);
not (n267,n268);
and (n268,n103,n152);
and (n269,n102,n154);
nand (n270,n271,n275);
or (n271,n106,n272);
nor (n272,n273,n274);
and (n273,n112,n142);
and (n274,n107,n144);
or (n275,n110,n108);
or (n276,n277,n292);
and (n277,n278,n283);
xor (n278,n279,n280);
nor (n279,n150,n102);
nand (n280,n281,n282);
or (n281,n106,n254);
or (n282,n272,n108);
nand (n283,n284,n288);
or (n284,n124,n285);
nor (n285,n286,n287);
and (n286,n31,n20);
and (n287,n29,n132);
or (n288,n125,n289);
nor (n289,n290,n291);
and (n290,n132,n36);
and (n291,n20,n38);
and (n292,n279,n280);
or (n293,n294,n360);
and (n294,n295,n359);
xor (n295,n296,n332);
or (n296,n297,n331);
and (n297,n298,n320);
xor (n298,n299,n308);
nand (n299,n300,n305);
or (n300,n301,n124);
not (n301,n302);
nor (n302,n303,n304);
and (n303,n190,n20);
and (n304,n192,n132);
nand (n305,n306,n307);
not (n306,n285);
not (n307,n125);
nand (n308,n309,n314);
or (n309,n310,n171);
not (n310,n311);
nand (n311,n312,n313);
or (n312,n180,n67);
or (n313,n179,n65);
nand (n314,n315,n319);
not (n315,n316);
nor (n316,n317,n318);
and (n317,n179,n207);
and (n318,n180,n209);
not (n319,n172);
nand (n320,n321,n326);
or (n321,n322,n195);
not (n322,n323);
nor (n323,n324,n325);
and (n324,n89,n53);
and (n325,n91,n56);
nand (n326,n327,n197);
not (n327,n328);
nor (n328,n329,n330);
and (n329,n56,n59);
and (n330,n53,n61);
and (n331,n299,n308);
or (n332,n333,n358);
and (n333,n334,n352);
xor (n334,n335,n345);
nand (n335,n336,n340);
or (n336,n337,n14);
nor (n337,n338,n339);
and (n338,n216,n25);
and (n339,n214,n24);
nand (n340,n341,n16);
not (n341,n342);
nor (n342,n343,n344);
and (n343,n24,n184);
and (n344,n25,n186);
nand (n345,n346,n350);
or (n346,n347,n41);
nor (n347,n348,n349);
and (n348,n47,n166);
and (n349,n48,n168);
nand (n350,n351,n50);
not (n351,n225);
nand (n352,n353,n357);
or (n353,n70,n354);
nor (n354,n355,n356);
and (n355,n102,n79);
and (n356,n103,n78);
or (n357,n71,n234);
and (n358,n335,n345);
xor (n359,n278,n283);
and (n360,n296,n332);
and (n361,n220,n258);
xor (n362,n363,n409);
xor (n363,n364,n367);
or (n364,n365,n366);
and (n365,n259,n276);
and (n366,n260,n263);
xor (n367,n368,n390);
xor (n368,n369,n370);
and (n369,n264,n270);
or (n370,n371,n389);
and (n371,n372,n383);
xor (n372,n373,n377);
nand (n373,n374,n375);
or (n374,n289,n124);
nand (n375,n376,n307);
not (n376,n134);
nand (n377,n378,n382);
or (n378,n149,n379);
nor (n379,n380,n381);
and (n380,n102,n98);
and (n381,n103,n97);
or (n382,n150,n158);
nand (n383,n384,n388);
or (n384,n171,n385);
nor (n385,n386,n387);
and (n386,n179,n214);
and (n387,n180,n216);
or (n388,n172,n182);
and (n389,n373,n377);
or (n390,n391,n408);
and (n391,n392,n405);
xor (n392,n393,n399);
nand (n393,n394,n398);
or (n394,n195,n395);
nor (n395,n396,n397);
and (n396,n56,n65);
and (n397,n53,n67);
or (n398,n211,n205);
nand (n399,n400,n404);
or (n400,n14,n401);
nor (n401,n402,n403);
and (n402,n24,n190);
and (n403,n25,n192);
or (n404,n33,n27);
nand (n405,n406,n407);
or (n406,n41,n229);
or (n407,n51,n57);
and (n408,n393,n399);
or (n409,n410,n427);
and (n410,n411,n426);
xor (n411,n412,n425);
or (n412,n413,n424);
and (n413,n414,n421);
xor (n414,n415,n418);
nand (n415,n416,n417);
or (n416,n171,n316);
or (n417,n172,n385);
nand (n418,n419,n420);
or (n419,n195,n328);
or (n420,n211,n395);
nand (n421,n422,n423);
or (n422,n14,n342);
or (n423,n33,n401);
and (n424,n415,n418);
xor (n425,n392,n405);
xor (n426,n372,n383);
and (n427,n412,n425);
or (n428,n429,n486);
and (n429,n430,n485);
xor (n430,n431,n432);
xor (n431,n411,n426);
or (n432,n433,n484);
and (n433,n434,n437);
xor (n434,n435,n436);
xor (n435,n414,n421);
xor (n436,n222,n241);
or (n437,n438,n483);
and (n438,n439,n460);
xor (n439,n440,n441);
xor (n440,n242,n248);
or (n441,n442,n459);
and (n442,n443,n452);
xor (n443,n444,n445);
nor (n444,n71,n102);
nand (n445,n446,n451);
or (n446,n447,n124);
not (n447,n448);
nand (n448,n449,n450);
or (n449,n20,n186);
or (n450,n132,n184);
nand (n451,n307,n302);
nand (n452,n453,n458);
or (n453,n171,n454);
not (n454,n455);
nor (n455,n456,n457);
and (n456,n61,n179);
and (n457,n59,n180);
or (n458,n172,n310);
and (n459,n444,n445);
or (n460,n461,n482);
and (n461,n462,n476);
xor (n462,n463,n470);
nand (n463,n464,n469);
or (n464,n465,n195);
not (n465,n466);
nor (n466,n467,n468);
and (n467,n85,n56);
and (n468,n83,n53);
nand (n469,n197,n323);
nand (n470,n471,n475);
or (n471,n106,n472);
nor (n472,n473,n474);
and (n473,n112,n29);
and (n474,n107,n31);
or (n475,n250,n108);
nand (n476,n477,n481);
or (n477,n41,n478);
nor (n478,n479,n480);
and (n479,n47,n160);
and (n480,n48,n162);
or (n481,n51,n347);
and (n482,n463,n470);
and (n483,n440,n441);
and (n484,n435,n436);
xor (n485,n219,n293);
and (n486,n431,n432);
nand (n487,n6,n428);
not (n488,n489);
or (n489,n490,n1010);
and (n490,n491,n552);
xor (n491,n492,n551);
or (n492,n493,n550);
and (n493,n494,n497);
xor (n494,n495,n496);
xor (n495,n295,n359);
xor (n496,n434,n437);
or (n497,n498,n549);
and (n498,n499,n502);
xor (n499,n500,n501);
xor (n500,n334,n352);
xor (n501,n298,n320);
or (n502,n503,n548);
and (n503,n504,n526);
xor (n504,n505,n511);
nand (n505,n506,n510);
or (n506,n14,n507);
nor (n507,n508,n509);
and (n508,n24,n207);
and (n509,n25,n209);
or (n510,n33,n337);
nor (n511,n512,n520);
not (n512,n513);
nand (n513,n514,n519);
or (n514,n515,n124);
not (n515,n516);
nand (n516,n517,n518);
or (n517,n20,n216);
or (n518,n132,n214);
nand (n519,n307,n448);
nand (n520,n521,n48);
nand (n521,n522,n523);
or (n522,n103,n46);
nand (n523,n524,n56);
not (n524,n525);
and (n525,n103,n46);
or (n526,n527,n547);
and (n527,n528,n541);
xor (n528,n529,n535);
nand (n529,n530,n531);
or (n530,n454,n172);
or (n531,n171,n532);
nor (n532,n533,n534);
and (n533,n179,n89);
and (n534,n180,n91);
nand (n535,n536,n540);
or (n536,n195,n537);
or (n537,n538,n539);
and (n538,n166,n53);
and (n539,n168,n56);
nand (n540,n197,n466);
nand (n541,n542,n546);
or (n542,n106,n543);
nor (n543,n544,n545);
and (n544,n112,n190);
and (n545,n107,n192);
or (n546,n472,n108);
and (n547,n529,n535);
and (n548,n505,n511);
and (n549,n500,n501);
and (n550,n495,n496);
xor (n551,n430,n485);
or (n552,n553,n1009);
and (n553,n554,n588);
xor (n554,n555,n587);
or (n555,n556,n586);
and (n556,n557,n585);
xor (n557,n558,n559);
xor (n558,n439,n460);
or (n559,n560,n584);
and (n560,n561,n564);
xor (n561,n562,n563);
xor (n562,n462,n476);
xor (n563,n443,n452);
or (n564,n565,n583);
and (n565,n566,n579);
xor (n566,n567,n573);
nand (n567,n568,n572);
or (n568,n41,n569);
nor (n569,n570,n571);
and (n570,n102,n48);
and (n571,n47,n103);
or (n572,n51,n478);
nand (n573,n574,n578);
or (n574,n14,n575);
nor (n575,n576,n577);
and (n576,n24,n65);
and (n577,n25,n67);
or (n578,n33,n507);
nand (n579,n580,n582);
or (n580,n581,n512);
not (n581,n520);
or (n582,n513,n520);
and (n583,n567,n573);
and (n584,n562,n563);
xor (n585,n499,n502);
and (n586,n558,n559);
xor (n587,n494,n497);
nand (n588,n589,n1003);
nand (n589,n590,n986);
nand (n590,n591,n985);
or (n591,n592,n723);
not (n592,n593);
nand (n593,n594,n685);
not (n594,n595);
xor (n595,n596,n643);
xor (n596,n597,n598);
xor (n597,n566,n579);
xor (n598,n599,n642);
xor (n599,n600,n618);
or (n600,n601,n617);
and (n601,n602,n611);
xor (n602,n603,n604);
nor (n603,n51,n102);
nand (n604,n605,n610);
or (n605,n606,n124);
not (n606,n607);
nand (n607,n608,n609);
or (n608,n20,n209);
or (n609,n132,n207);
nand (n610,n307,n516);
nand (n611,n612,n616);
or (n612,n171,n613);
nor (n613,n614,n615);
and (n614,n179,n83);
and (n615,n180,n85);
or (n616,n172,n532);
and (n617,n603,n604);
or (n618,n619,n641);
and (n619,n620,n635);
xor (n620,n621,n629);
nand (n621,n622,n627);
or (n622,n623,n195);
not (n623,n624);
nand (n624,n625,n626);
or (n625,n53,n162);
or (n626,n56,n160);
nand (n627,n628,n197);
not (n628,n537);
nand (n629,n630,n634);
or (n630,n106,n631);
nor (n631,n632,n633);
and (n632,n112,n184);
and (n633,n107,n186);
or (n634,n543,n108);
nand (n635,n636,n640);
or (n636,n14,n637);
nor (n637,n638,n639);
and (n638,n24,n59);
and (n639,n25,n61);
or (n640,n33,n575);
and (n641,n621,n629);
xor (n642,n528,n541);
or (n643,n644,n684);
and (n644,n645,n683);
xor (n645,n646,n660);
and (n646,n647,n653);
and (n647,n648,n53);
nand (n648,n649,n650);
or (n649,n103,n199);
nand (n650,n651,n179);
not (n651,n652);
and (n652,n103,n199);
nand (n653,n654,n659);
or (n654,n655,n124);
not (n655,n656);
nor (n656,n657,n658);
and (n657,n65,n20);
and (n658,n67,n132);
nand (n659,n307,n607);
or (n660,n661,n682);
and (n661,n662,n676);
xor (n662,n663,n670);
nand (n663,n664,n668);
or (n664,n665,n171);
nor (n665,n666,n667);
and (n666,n166,n179);
and (n667,n168,n180);
nand (n668,n669,n319);
not (n669,n613);
nand (n670,n671,n672);
or (n671,n623,n211);
nand (n672,n196,n673);
nand (n673,n674,n675);
or (n674,n103,n56);
or (n675,n102,n53);
nand (n676,n677,n681);
or (n677,n106,n678);
nor (n678,n679,n680);
and (n679,n112,n214);
and (n680,n107,n216);
or (n681,n631,n108);
and (n682,n663,n670);
xor (n683,n602,n611);
and (n684,n646,n660);
not (n685,n686);
or (n686,n687,n722);
and (n687,n688,n721);
xor (n688,n689,n690);
xor (n689,n620,n635);
or (n690,n691,n720);
and (n691,n692,n700);
xor (n692,n693,n699);
nand (n693,n694,n698);
or (n694,n14,n695);
nor (n695,n696,n697);
and (n696,n24,n89);
and (n697,n25,n91);
or (n698,n33,n637);
xor (n699,n647,n653);
or (n700,n701,n719);
and (n701,n702,n712);
xor (n702,n703,n704);
and (n703,n197,n103);
nand (n704,n705,n706);
or (n705,n678,n108);
nand (n706,n707,n711);
not (n707,n708);
nor (n708,n709,n710);
and (n709,n112,n207);
and (n710,n107,n209);
not (n711,n106);
nand (n712,n713,n718);
or (n713,n714,n171);
not (n714,n715);
nor (n715,n716,n717);
and (n716,n160,n180);
and (n717,n162,n179);
or (n718,n172,n665);
and (n719,n703,n704);
and (n720,n693,n699);
xor (n721,n645,n683);
and (n722,n689,n690);
not (n723,n724);
nand (n724,n725,n984);
or (n725,n726,n769);
not (n726,n727);
nand (n727,n728,n730);
not (n728,n729);
xor (n729,n688,n721);
not (n730,n731);
or (n731,n732,n768);
and (n732,n733,n767);
xor (n733,n734,n735);
xor (n734,n662,n676);
or (n735,n736,n766);
and (n736,n737,n753);
xor (n737,n738,n745);
nand (n738,n739,n744);
or (n739,n740,n124);
not (n740,n741);
nor (n741,n742,n743);
and (n742,n59,n20);
and (n743,n61,n132);
nand (n744,n307,n656);
nand (n745,n746,n751);
or (n746,n747,n14);
not (n747,n748);
nand (n748,n749,n750);
or (n749,n25,n85);
or (n750,n24,n83);
nand (n751,n752,n16);
not (n752,n695);
and (n753,n754,n760);
nor (n754,n755,n179);
nor (n755,n756,n759);
and (n756,n757,n24);
not (n757,n758);
and (n758,n103,n174);
and (n759,n102,n176);
nand (n760,n761,n765);
or (n761,n106,n762);
nor (n762,n763,n764);
and (n763,n65,n112);
and (n764,n67,n107);
or (n765,n708,n108);
and (n766,n738,n745);
xor (n767,n692,n700);
and (n768,n734,n735);
not (n769,n770);
nand (n770,n771,n980,n983);
nand (n771,n772,n960,n973);
nand (n772,n773,n959);
or (n773,n774,n849);
not (n774,n775);
nand (n775,n776,n823);
not (n776,n777);
xor (n777,n778,n803);
xor (n778,n779,n780);
xor (n779,n754,n760);
or (n780,n781,n802);
and (n781,n782,n792);
xor (n782,n783,n784);
and (n783,n319,n103);
nand (n784,n785,n790);
or (n785,n106,n786);
not (n786,n787);
nor (n787,n788,n789);
and (n788,n61,n112);
and (n789,n59,n107);
nand (n790,n791,n109);
not (n791,n762);
nand (n792,n793,n798);
or (n793,n794,n124);
not (n794,n795);
nor (n795,n796,n797);
and (n796,n85,n132);
and (n797,n83,n20);
nand (n798,n307,n799);
nor (n799,n800,n801);
and (n800,n89,n20);
and (n801,n91,n132);
and (n802,n783,n784);
xor (n803,n804,n816);
xor (n804,n805,n812);
nand (n805,n806,n811);
or (n806,n807,n171);
not (n807,n808);
nand (n808,n809,n810);
or (n809,n179,n103);
or (n810,n102,n180);
nand (n811,n319,n715);
nand (n812,n813,n815);
or (n813,n814,n124);
not (n814,n799);
nand (n815,n307,n741);
nand (n816,n817,n822);
or (n817,n818,n14);
not (n818,n819);
nand (n819,n820,n821);
or (n820,n25,n168);
or (n821,n24,n166);
nand (n822,n16,n748);
not (n823,n824);
or (n824,n825,n848);
and (n825,n826,n847);
xor (n826,n827,n834);
nand (n827,n828,n833);
or (n828,n829,n14);
not (n829,n830);
nor (n830,n831,n832);
and (n831,n160,n25);
and (n832,n162,n24);
nand (n833,n16,n819);
and (n834,n835,n840);
and (n835,n836,n25);
nand (n836,n837,n839);
or (n837,n838,n20);
and (n838,n103,n19);
or (n839,n103,n19);
nand (n840,n841,n842);
or (n841,n108,n786);
nand (n842,n843,n711);
not (n843,n844);
nor (n844,n845,n846);
and (n845,n89,n112);
and (n846,n91,n107);
xor (n847,n782,n792);
and (n848,n827,n834);
not (n849,n850);
nand (n850,n851,n958);
or (n851,n852,n876);
not (n852,n853);
nand (n853,n854,n856);
not (n854,n855);
xor (n855,n826,n847);
not (n856,n857);
or (n857,n858,n875);
and (n858,n859,n874);
xor (n859,n860,n867);
nand (n860,n861,n866);
or (n861,n862,n124);
not (n862,n863);
nor (n863,n864,n865);
and (n864,n168,n132);
and (n865,n166,n20);
nand (n866,n307,n795);
nand (n867,n868,n873);
or (n868,n869,n14);
not (n869,n870);
nand (n870,n871,n872);
or (n871,n103,n24);
or (n872,n25,n102);
nand (n873,n16,n830);
xor (n874,n835,n840);
and (n875,n860,n867);
not (n876,n877);
nand (n877,n878,n957);
or (n878,n879,n903);
not (n879,n880);
nand (n880,n881,n883);
not (n881,n882);
xor (n882,n859,n874);
not (n883,n884);
or (n884,n885,n902);
and (n885,n886,n895);
xor (n886,n887,n888);
and (n887,n16,n103);
nand (n888,n889,n894);
or (n889,n890,n124);
not (n890,n891);
nor (n891,n892,n893);
and (n892,n160,n20);
and (n893,n162,n132);
nand (n894,n307,n863);
nand (n895,n896,n901);
or (n896,n106,n897);
not (n897,n898);
nor (n898,n899,n900);
and (n899,n85,n112);
and (n900,n83,n107);
or (n901,n844,n108);
and (n902,n887,n888);
not (n903,n904);
nand (n904,n905,n956);
or (n905,n906,n921);
nor (n906,n907,n908);
xor (n907,n886,n895);
and (n908,n909,n915);
nor (n909,n910,n132);
and (n910,n911,n914);
nand (n911,n912,n112);
not (n912,n913);
and (n913,n103,n127);
nand (n914,n102,n129);
nand (n915,n916,n917);
or (n916,n108,n897);
nand (n917,n918,n711);
nand (n918,n919,n920);
or (n919,n166,n112);
nand (n920,n112,n166);
not (n921,n922);
or (n922,n923,n955);
and (n923,n924,n933);
xor (n924,n925,n932);
nand (n925,n926,n931);
or (n926,n927,n124);
not (n927,n928);
nand (n928,n929,n930);
or (n929,n132,n103);
or (n930,n20,n102);
nand (n931,n307,n891);
xor (n932,n909,n915);
nand (n933,n934,n954);
or (n934,n935,n944);
nor (n935,n936,n943);
nand (n936,n937,n939);
or (n937,n108,n938);
not (n938,n918);
nand (n939,n940,n711);
nand (n940,n941,n942);
or (n941,n160,n112);
nand (n942,n112,n160);
and (n943,n307,n103);
nand (n944,n945,n952);
nand (n945,n946,n948);
or (n946,n108,n947);
not (n947,n940);
nand (n948,n949,n711);
nor (n949,n950,n951);
and (n950,n102,n112);
and (n951,n103,n107);
nor (n952,n953,n112);
nor (n953,n102,n108);
nand (n954,n936,n943);
and (n955,n925,n932);
nand (n956,n907,n908);
nand (n957,n882,n884);
nand (n958,n855,n857);
nand (n959,n824,n777);
nand (n960,n961,n963);
not (n961,n962);
xor (n962,n733,n767);
not (n963,n964);
or (n964,n965,n972);
and (n965,n966,n971);
xor (n966,n967,n970);
or (n967,n968,n969);
and (n968,n804,n816);
and (n969,n805,n812);
xor (n970,n702,n712);
xor (n971,n737,n753);
and (n972,n967,n970);
nand (n973,n974,n976);
not (n974,n975);
xor (n975,n966,n971);
not (n976,n977);
or (n977,n978,n979);
and (n978,n778,n803);
and (n979,n779,n780);
nand (n980,n960,n981);
not (n981,n982);
nand (n982,n975,n977);
nand (n983,n962,n964);
or (n984,n728,n730);
nand (n985,n595,n686);
nor (n986,n987,n998);
nor (n987,n988,n989);
xor (n988,n557,n585);
or (n989,n990,n997);
and (n990,n991,n996);
xor (n991,n992,n993);
xor (n992,n504,n526);
or (n993,n994,n995);
and (n994,n599,n642);
and (n995,n600,n618);
xor (n996,n561,n564);
and (n997,n992,n993);
nor (n998,n999,n1000);
xor (n999,n991,n996);
or (n1000,n1001,n1002);
and (n1001,n596,n643);
and (n1002,n597,n598);
nor (n1003,n1004,n1008);
and (n1004,n1005,n1006);
not (n1005,n987);
not (n1006,n1007);
nand (n1007,n999,n1000);
and (n1008,n988,n989);
and (n1009,n555,n587);
and (n1010,n492,n551);
or (n1011,n489,n3);
xor (n1012,n1013,n1711);
xor (n1013,n1014,n1708);
xor (n1014,n1015,n1707);
xor (n1015,n1016,n1699);
xor (n1016,n1017,n1698);
xor (n1017,n1018,n1683);
xor (n1018,n1019,n1682);
xor (n1019,n1020,n1662);
xor (n1020,n1021,n1661);
xor (n1021,n1022,n1634);
xor (n1022,n1023,n1633);
xor (n1023,n1024,n1601);
xor (n1024,n1025,n1600);
xor (n1025,n1026,n1564);
xor (n1026,n1027,n1563);
xor (n1027,n1028,n1519);
xor (n1028,n1029,n1518);
xor (n1029,n1030,n1469);
xor (n1030,n1031,n1468);
xor (n1031,n1032,n1412);
xor (n1032,n1033,n1411);
xor (n1033,n1034,n1349);
xor (n1034,n1035,n1348);
xor (n1035,n1036,n1280);
xor (n1036,n1037,n1279);
xor (n1037,n1038,n1211);
xor (n1038,n1039,n1210);
xor (n1039,n1040,n1130);
xor (n1040,n1041,n1129);
xor (n1041,n1042,n1045);
xor (n1042,n1043,n1044);
and (n1043,n120,n109);
and (n1044,n113,n107);
or (n1045,n1046,n1049);
and (n1046,n1047,n1048);
and (n1047,n113,n109);
and (n1048,n142,n107);
and (n1049,n1050,n1051);
xor (n1050,n1047,n1048);
or (n1051,n1052,n1055);
and (n1052,n1053,n1054);
and (n1053,n142,n109);
and (n1054,n136,n107);
and (n1055,n1056,n1057);
xor (n1056,n1053,n1054);
or (n1057,n1058,n1061);
and (n1058,n1059,n1060);
and (n1059,n136,n109);
and (n1060,n36,n107);
and (n1061,n1062,n1063);
xor (n1062,n1059,n1060);
or (n1063,n1064,n1067);
and (n1064,n1065,n1066);
and (n1065,n36,n109);
and (n1066,n29,n107);
and (n1067,n1068,n1069);
xor (n1068,n1065,n1066);
or (n1069,n1070,n1073);
and (n1070,n1071,n1072);
and (n1071,n29,n109);
and (n1072,n190,n107);
and (n1073,n1074,n1075);
xor (n1074,n1071,n1072);
or (n1075,n1076,n1079);
and (n1076,n1077,n1078);
and (n1077,n190,n109);
and (n1078,n184,n107);
and (n1079,n1080,n1081);
xor (n1080,n1077,n1078);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
and (n1083,n184,n109);
and (n1084,n214,n107);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
and (n1089,n214,n109);
and (n1090,n207,n107);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
and (n1095,n207,n109);
and (n1096,n65,n107);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
or (n1099,n1100,n1102);
and (n1100,n1101,n789);
and (n1101,n65,n109);
and (n1102,n1103,n1104);
xor (n1103,n1101,n789);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
and (n1106,n59,n109);
and (n1107,n89,n107);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1113);
and (n1111,n1112,n900);
and (n1112,n89,n109);
and (n1113,n1114,n1115);
xor (n1114,n1112,n900);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n83,n109);
and (n1118,n166,n107);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n166,n109);
and (n1124,n160,n107);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
and (n1127,n1128,n951);
and (n1128,n160,n109);
and (n1129,n142,n127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1050,n1051);
and (n1133,n136,n127);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1056,n1057);
and (n1139,n36,n127);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1062,n1063);
and (n1145,n29,n127);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1068,n1069);
and (n1151,n190,n127);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1074,n1075);
and (n1157,n184,n127);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1080,n1081);
and (n1163,n214,n127);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1086,n1087);
and (n1169,n207,n127);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
or (n1172,n1173,n1176);
and (n1173,n1174,n1175);
xor (n1174,n1092,n1093);
and (n1175,n65,n127);
and (n1176,n1177,n1178);
xor (n1177,n1174,n1175);
or (n1178,n1179,n1182);
and (n1179,n1180,n1181);
xor (n1180,n1098,n1099);
and (n1181,n59,n127);
and (n1182,n1183,n1184);
xor (n1183,n1180,n1181);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1103,n1104);
and (n1187,n89,n127);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1109,n1110);
and (n1193,n83,n127);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
or (n1196,n1197,n1200);
and (n1197,n1198,n1199);
xor (n1198,n1114,n1115);
and (n1199,n166,n127);
and (n1200,n1201,n1202);
xor (n1201,n1198,n1199);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
xor (n1204,n1120,n1121);
and (n1205,n160,n127);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
and (n1208,n1209,n913);
xor (n1209,n1126,n1127);
and (n1210,n136,n20);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1135,n1136);
and (n1214,n36,n20);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1141,n1142);
and (n1220,n29,n20);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
or (n1223,n1224,n1226);
and (n1224,n1225,n303);
xor (n1225,n1147,n1148);
and (n1226,n1227,n1228);
xor (n1227,n1225,n303);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1153,n1154);
and (n1231,n184,n20);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1159,n1160);
and (n1237,n214,n20);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1165,n1166);
and (n1243,n207,n20);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1249);
and (n1247,n1248,n657);
xor (n1248,n1171,n1172);
and (n1249,n1250,n1251);
xor (n1250,n1248,n657);
or (n1251,n1252,n1254);
and (n1252,n1253,n742);
xor (n1253,n1177,n1178);
and (n1254,n1255,n1256);
xor (n1255,n1253,n742);
or (n1256,n1257,n1259);
and (n1257,n1258,n800);
xor (n1258,n1183,n1184);
and (n1259,n1260,n1261);
xor (n1260,n1258,n800);
or (n1261,n1262,n1264);
and (n1262,n1263,n797);
xor (n1263,n1189,n1190);
and (n1264,n1265,n1266);
xor (n1265,n1263,n797);
or (n1266,n1267,n1269);
and (n1267,n1268,n865);
xor (n1268,n1195,n1196);
and (n1269,n1270,n1271);
xor (n1270,n1268,n865);
or (n1271,n1272,n1274);
and (n1272,n1273,n892);
xor (n1273,n1201,n1202);
and (n1274,n1275,n1276);
xor (n1275,n1273,n892);
and (n1276,n1277,n1278);
xor (n1277,n1207,n1208);
and (n1278,n103,n20);
and (n1279,n36,n19);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1216,n1217);
and (n1283,n29,n19);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1222,n1223);
and (n1289,n190,n19);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1227,n1228);
and (n1295,n184,n19);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1233,n1234);
and (n1301,n214,n19);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1239,n1240);
and (n1307,n207,n19);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1245,n1246);
and (n1313,n65,n19);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1250,n1251);
and (n1319,n59,n19);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1255,n1256);
and (n1325,n89,n19);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1260,n1261);
and (n1331,n83,n19);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1265,n1266);
and (n1337,n166,n19);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1270,n1271);
and (n1343,n160,n19);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
and (n1346,n1347,n838);
xor (n1347,n1275,n1276);
and (n1348,n29,n25);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1285,n1286);
and (n1352,n190,n25);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
or (n1355,n1356,n1359);
and (n1356,n1357,n1358);
xor (n1357,n1291,n1292);
and (n1358,n184,n25);
and (n1359,n1360,n1361);
xor (n1360,n1357,n1358);
or (n1361,n1362,n1365);
and (n1362,n1363,n1364);
xor (n1363,n1297,n1298);
and (n1364,n214,n25);
and (n1365,n1366,n1367);
xor (n1366,n1363,n1364);
or (n1367,n1368,n1371);
and (n1368,n1369,n1370);
xor (n1369,n1303,n1304);
and (n1370,n207,n25);
and (n1371,n1372,n1373);
xor (n1372,n1369,n1370);
or (n1373,n1374,n1377);
and (n1374,n1375,n1376);
xor (n1375,n1309,n1310);
and (n1376,n65,n25);
and (n1377,n1378,n1379);
xor (n1378,n1375,n1376);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1315,n1316);
and (n1382,n59,n25);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
or (n1385,n1386,n1389);
and (n1386,n1387,n1388);
xor (n1387,n1321,n1322);
and (n1388,n89,n25);
and (n1389,n1390,n1391);
xor (n1390,n1387,n1388);
or (n1391,n1392,n1395);
and (n1392,n1393,n1394);
xor (n1393,n1327,n1328);
and (n1394,n83,n25);
and (n1395,n1396,n1397);
xor (n1396,n1393,n1394);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1333,n1334);
and (n1400,n166,n25);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
or (n1403,n1404,n1406);
and (n1404,n1405,n831);
xor (n1405,n1339,n1340);
and (n1406,n1407,n1408);
xor (n1407,n1405,n831);
and (n1408,n1409,n1410);
xor (n1409,n1345,n1346);
and (n1410,n103,n25);
and (n1411,n190,n174);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1354,n1355);
and (n1415,n184,n174);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1360,n1361);
and (n1421,n214,n174);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1366,n1367);
and (n1427,n207,n174);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1372,n1373);
and (n1433,n65,n174);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1378,n1379);
and (n1439,n59,n174);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1384,n1385);
and (n1445,n89,n174);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1390,n1391);
and (n1451,n83,n174);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1396,n1397);
and (n1457,n166,n174);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1402,n1403);
and (n1463,n160,n174);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
and (n1466,n1467,n758);
xor (n1467,n1407,n1408);
and (n1468,n184,n180);
or (n1469,n1470,n1473);
and (n1470,n1471,n1472);
xor (n1471,n1417,n1418);
and (n1472,n214,n180);
and (n1473,n1474,n1475);
xor (n1474,n1471,n1472);
or (n1475,n1476,n1479);
and (n1476,n1477,n1478);
xor (n1477,n1423,n1424);
and (n1478,n207,n180);
and (n1479,n1480,n1481);
xor (n1480,n1477,n1478);
or (n1481,n1482,n1485);
and (n1482,n1483,n1484);
xor (n1483,n1429,n1430);
and (n1484,n65,n180);
and (n1485,n1486,n1487);
xor (n1486,n1483,n1484);
or (n1487,n1488,n1490);
and (n1488,n1489,n457);
xor (n1489,n1435,n1436);
and (n1490,n1491,n1492);
xor (n1491,n1489,n457);
or (n1492,n1493,n1496);
and (n1493,n1494,n1495);
xor (n1494,n1441,n1442);
and (n1495,n89,n180);
and (n1496,n1497,n1498);
xor (n1497,n1494,n1495);
or (n1498,n1499,n1502);
and (n1499,n1500,n1501);
xor (n1500,n1447,n1448);
and (n1501,n83,n180);
and (n1502,n1503,n1504);
xor (n1503,n1500,n1501);
or (n1504,n1505,n1508);
and (n1505,n1506,n1507);
xor (n1506,n1453,n1454);
and (n1507,n166,n180);
and (n1508,n1509,n1510);
xor (n1509,n1506,n1507);
or (n1510,n1511,n1513);
and (n1511,n1512,n716);
xor (n1512,n1459,n1460);
and (n1513,n1514,n1515);
xor (n1514,n1512,n716);
and (n1515,n1516,n1517);
xor (n1516,n1465,n1466);
and (n1517,n103,n180);
and (n1518,n214,n199);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1474,n1475);
and (n1522,n207,n199);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1480,n1481);
and (n1528,n65,n199);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1486,n1487);
and (n1534,n59,n199);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1491,n1492);
and (n1540,n89,n199);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1497,n1498);
and (n1546,n83,n199);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1503,n1504);
and (n1552,n166,n199);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1509,n1510);
and (n1558,n160,n199);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
and (n1561,n1562,n652);
xor (n1562,n1514,n1515);
and (n1563,n207,n53);
or (n1564,n1565,n1568);
and (n1565,n1566,n1567);
xor (n1566,n1524,n1525);
and (n1567,n65,n53);
and (n1568,n1569,n1570);
xor (n1569,n1566,n1567);
or (n1570,n1571,n1574);
and (n1571,n1572,n1573);
xor (n1572,n1530,n1531);
and (n1573,n59,n53);
and (n1574,n1575,n1576);
xor (n1575,n1572,n1573);
or (n1576,n1577,n1579);
and (n1577,n1578,n324);
xor (n1578,n1536,n1537);
and (n1579,n1580,n1581);
xor (n1580,n1578,n324);
or (n1581,n1582,n1584);
and (n1582,n1583,n468);
xor (n1583,n1542,n1543);
and (n1584,n1585,n1586);
xor (n1585,n1583,n468);
or (n1586,n1587,n1589);
and (n1587,n1588,n538);
xor (n1588,n1548,n1549);
and (n1589,n1590,n1591);
xor (n1590,n1588,n538);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1554,n1555);
and (n1594,n160,n53);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
and (n1597,n1598,n1599);
xor (n1598,n1560,n1561);
and (n1599,n103,n53);
and (n1600,n65,n46);
or (n1601,n1602,n1605);
and (n1602,n1603,n1604);
xor (n1603,n1569,n1570);
and (n1604,n59,n46);
and (n1605,n1606,n1607);
xor (n1606,n1603,n1604);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1575,n1576);
and (n1610,n89,n46);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1580,n1581);
and (n1616,n83,n46);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1585,n1586);
and (n1622,n166,n46);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1590,n1591);
and (n1628,n160,n46);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
and (n1631,n1632,n525);
xor (n1632,n1596,n1597);
and (n1633,n59,n48);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1606,n1607);
and (n1637,n89,n48);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1612,n1613);
and (n1643,n83,n48);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1618,n1619);
and (n1649,n166,n48);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1624,n1625);
and (n1655,n160,n48);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
and (n1658,n1659,n1660);
xor (n1659,n1630,n1631);
and (n1660,n103,n48);
and (n1661,n89,n73);
or (n1662,n1663,n1666);
and (n1663,n1664,n1665);
xor (n1664,n1639,n1640);
and (n1665,n83,n73);
and (n1666,n1667,n1668);
xor (n1667,n1664,n1665);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1645,n1646);
and (n1671,n166,n73);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1651,n1652);
and (n1677,n160,n73);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
and (n1680,n1681,n246);
xor (n1681,n1657,n1658);
and (n1682,n83,n79);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1667,n1668);
and (n1686,n166,n79);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
or (n1689,n1690,n1693);
and (n1690,n1691,n1692);
xor (n1691,n1673,n1674);
and (n1692,n160,n79);
and (n1693,n1694,n1695);
xor (n1694,n1691,n1692);
and (n1695,n1696,n1697);
xor (n1696,n1679,n1680);
and (n1697,n103,n79);
and (n1698,n166,n152);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1688,n1689);
and (n1702,n160,n152);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
and (n1705,n1706,n268);
xor (n1706,n1694,n1695);
and (n1707,n160,n98);
and (n1708,n1709,n1710);
xor (n1709,n1704,n1705);
and (n1710,n103,n98);
and (n1711,n103,n99);
endmodule
