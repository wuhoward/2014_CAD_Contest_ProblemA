module top (out,n23,n24,n26,n27,n32,n39,n46,n53,n60
        ,n67,n74,n81,n88,n94,n96,n149,n196,n237,n272
        ,n301,n324,n341,n352,n357,n380,n381,n383,n384,n389
        ,n396,n403,n410,n417,n424,n431,n438,n445,n451,n453
        ,n506,n553,n594,n629,n658,n681,n698,n709,n714,n715);
output out;
input n23;
input n24;
input n26;
input n27;
input n32;
input n39;
input n46;
input n53;
input n60;
input n67;
input n74;
input n81;
input n88;
input n94;
input n96;
input n149;
input n196;
input n237;
input n272;
input n301;
input n324;
input n341;
input n352;
input n357;
input n380;
input n381;
input n383;
input n384;
input n389;
input n396;
input n403;
input n410;
input n417;
input n424;
input n431;
input n438;
input n445;
input n451;
input n453;
input n506;
input n553;
input n594;
input n629;
input n658;
input n681;
input n698;
input n709;
input n714;
input n715;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n353;
wire n354;
wire n355;
wire n356;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n382;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n452;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n710;
wire n711;
wire n712;
wire n713;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
xor (out,n0,n716);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n715);
and (s0n0,notn0,n1);
and (s1n0,n715,n358);
xor (n1,n2,n356);
xor (n2,n3,n353);
xor (n3,n4,n351);
xor (n4,n5,n342);
xor (n5,n6,n340);
xor (n6,n7,n325);
xor (n7,n8,n323);
xor (n8,n9,n302);
xor (n9,n10,n300);
xor (n10,n11,n273);
xor (n11,n12,n271);
xor (n12,n13,n238);
xor (n13,n14,n236);
xor (n14,n15,n197);
xor (n15,n16,n195);
xor (n16,n17,n150);
xor (n17,n18,n148);
xor (n18,n19,n97);
xor (n19,n20,n95);
xor (n20,n21,n28);
xor (n21,n22,n25);
and (n22,n23,n24);
and (n25,n26,n27);
or (n28,n29,n33);
and (n29,n30,n31);
and (n30,n26,n24);
and (n31,n32,n27);
and (n33,n34,n35);
xor (n34,n30,n31);
or (n35,n36,n40);
and (n36,n37,n38);
and (n37,n32,n24);
and (n38,n39,n27);
and (n40,n41,n42);
xor (n41,n37,n38);
or (n42,n43,n47);
and (n43,n44,n45);
and (n44,n39,n24);
and (n45,n46,n27);
and (n47,n48,n49);
xor (n48,n44,n45);
or (n49,n50,n54);
and (n50,n51,n52);
and (n51,n46,n24);
and (n52,n53,n27);
and (n54,n55,n56);
xor (n55,n51,n52);
or (n56,n57,n61);
and (n57,n58,n59);
and (n58,n53,n24);
and (n59,n60,n27);
and (n61,n62,n63);
xor (n62,n58,n59);
or (n63,n64,n68);
and (n64,n65,n66);
and (n65,n60,n24);
and (n66,n67,n27);
and (n68,n69,n70);
xor (n69,n65,n66);
or (n70,n71,n75);
and (n71,n72,n73);
and (n72,n67,n24);
and (n73,n74,n27);
and (n75,n76,n77);
xor (n76,n72,n73);
or (n77,n78,n82);
and (n78,n79,n80);
and (n79,n74,n24);
and (n80,n81,n27);
and (n82,n83,n84);
xor (n83,n79,n80);
or (n84,n85,n89);
and (n85,n86,n87);
and (n86,n81,n24);
and (n87,n88,n27);
and (n89,n90,n91);
xor (n90,n86,n87);
and (n91,n92,n93);
and (n92,n88,n24);
and (n93,n94,n27);
and (n95,n32,n96);
or (n97,n98,n101);
and (n98,n99,n100);
xor (n99,n34,n35);
and (n100,n39,n96);
and (n101,n102,n103);
xor (n102,n99,n100);
or (n103,n104,n107);
and (n104,n105,n106);
xor (n105,n41,n42);
and (n106,n46,n96);
and (n107,n108,n109);
xor (n108,n105,n106);
or (n109,n110,n113);
and (n110,n111,n112);
xor (n111,n48,n49);
and (n112,n53,n96);
and (n113,n114,n115);
xor (n114,n111,n112);
or (n115,n116,n119);
and (n116,n117,n118);
xor (n117,n55,n56);
and (n118,n60,n96);
and (n119,n120,n121);
xor (n120,n117,n118);
or (n121,n122,n125);
and (n122,n123,n124);
xor (n123,n62,n63);
and (n124,n67,n96);
and (n125,n126,n127);
xor (n126,n123,n124);
or (n127,n128,n131);
and (n128,n129,n130);
xor (n129,n69,n70);
and (n130,n74,n96);
and (n131,n132,n133);
xor (n132,n129,n130);
or (n133,n134,n137);
and (n134,n135,n136);
xor (n135,n76,n77);
and (n136,n81,n96);
and (n137,n138,n139);
xor (n138,n135,n136);
or (n139,n140,n143);
and (n140,n141,n142);
xor (n141,n83,n84);
and (n142,n88,n96);
and (n143,n144,n145);
xor (n144,n141,n142);
and (n145,n146,n147);
xor (n146,n90,n91);
and (n147,n94,n96);
and (n148,n39,n149);
or (n150,n151,n154);
and (n151,n152,n153);
xor (n152,n102,n103);
and (n153,n46,n149);
and (n154,n155,n156);
xor (n155,n152,n153);
or (n156,n157,n160);
and (n157,n158,n159);
xor (n158,n108,n109);
and (n159,n53,n149);
and (n160,n161,n162);
xor (n161,n158,n159);
or (n162,n163,n166);
and (n163,n164,n165);
xor (n164,n114,n115);
and (n165,n60,n149);
and (n166,n167,n168);
xor (n167,n164,n165);
or (n168,n169,n172);
and (n169,n170,n171);
xor (n170,n120,n121);
and (n171,n67,n149);
and (n172,n173,n174);
xor (n173,n170,n171);
or (n174,n175,n178);
and (n175,n176,n177);
xor (n176,n126,n127);
and (n177,n74,n149);
and (n178,n179,n180);
xor (n179,n176,n177);
or (n180,n181,n184);
and (n181,n182,n183);
xor (n182,n132,n133);
and (n183,n81,n149);
and (n184,n185,n186);
xor (n185,n182,n183);
or (n186,n187,n190);
and (n187,n188,n189);
xor (n188,n138,n139);
and (n189,n88,n149);
and (n190,n191,n192);
xor (n191,n188,n189);
and (n192,n193,n194);
xor (n193,n144,n145);
and (n194,n94,n149);
and (n195,n46,n196);
or (n197,n198,n201);
and (n198,n199,n200);
xor (n199,n155,n156);
and (n200,n53,n196);
and (n201,n202,n203);
xor (n202,n199,n200);
or (n203,n204,n207);
and (n204,n205,n206);
xor (n205,n161,n162);
and (n206,n60,n196);
and (n207,n208,n209);
xor (n208,n205,n206);
or (n209,n210,n213);
and (n210,n211,n212);
xor (n211,n167,n168);
and (n212,n67,n196);
and (n213,n214,n215);
xor (n214,n211,n212);
or (n215,n216,n219);
and (n216,n217,n218);
xor (n217,n173,n174);
and (n218,n74,n196);
and (n219,n220,n221);
xor (n220,n217,n218);
or (n221,n222,n225);
and (n222,n223,n224);
xor (n223,n179,n180);
and (n224,n81,n196);
and (n225,n226,n227);
xor (n226,n223,n224);
or (n227,n228,n231);
and (n228,n229,n230);
xor (n229,n185,n186);
and (n230,n88,n196);
and (n231,n232,n233);
xor (n232,n229,n230);
and (n233,n234,n235);
xor (n234,n191,n192);
and (n235,n94,n196);
and (n236,n53,n237);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n202,n203);
and (n241,n60,n237);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n208,n209);
and (n247,n67,n237);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n214,n215);
and (n253,n74,n237);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n220,n221);
and (n259,n81,n237);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n226,n227);
and (n265,n88,n237);
and (n266,n267,n268);
xor (n267,n264,n265);
and (n268,n269,n270);
xor (n269,n232,n233);
and (n270,n94,n237);
and (n271,n60,n272);
or (n273,n274,n277);
and (n274,n275,n276);
xor (n275,n243,n244);
and (n276,n67,n272);
and (n277,n278,n279);
xor (n278,n275,n276);
or (n279,n280,n283);
and (n280,n281,n282);
xor (n281,n249,n250);
and (n282,n74,n272);
and (n283,n284,n285);
xor (n284,n281,n282);
or (n285,n286,n289);
and (n286,n287,n288);
xor (n287,n255,n256);
and (n288,n81,n272);
and (n289,n290,n291);
xor (n290,n287,n288);
or (n291,n292,n295);
and (n292,n293,n294);
xor (n293,n261,n262);
and (n294,n88,n272);
and (n295,n296,n297);
xor (n296,n293,n294);
and (n297,n298,n299);
xor (n298,n267,n268);
and (n299,n94,n272);
and (n300,n67,n301);
or (n302,n303,n306);
and (n303,n304,n305);
xor (n304,n278,n279);
and (n305,n74,n301);
and (n306,n307,n308);
xor (n307,n304,n305);
or (n308,n309,n312);
and (n309,n310,n311);
xor (n310,n284,n285);
and (n311,n81,n301);
and (n312,n313,n314);
xor (n313,n310,n311);
or (n314,n315,n318);
and (n315,n316,n317);
xor (n316,n290,n291);
and (n317,n88,n301);
and (n318,n319,n320);
xor (n319,n316,n317);
and (n320,n321,n322);
xor (n321,n296,n297);
and (n322,n94,n301);
and (n323,n74,n324);
or (n325,n326,n329);
and (n326,n327,n328);
xor (n327,n307,n308);
and (n328,n81,n324);
and (n329,n330,n331);
xor (n330,n327,n328);
or (n331,n332,n335);
and (n332,n333,n334);
xor (n333,n313,n314);
and (n334,n88,n324);
and (n335,n336,n337);
xor (n336,n333,n334);
and (n337,n338,n339);
xor (n338,n319,n320);
and (n339,n94,n324);
and (n340,n81,n341);
or (n342,n343,n346);
and (n343,n344,n345);
xor (n344,n330,n331);
and (n345,n88,n341);
and (n346,n347,n348);
xor (n347,n344,n345);
and (n348,n349,n350);
xor (n349,n336,n337);
and (n350,n94,n341);
and (n351,n88,n352);
and (n353,n354,n355);
xor (n354,n347,n348);
and (n355,n94,n352);
and (n356,n94,n357);
xor (n358,n359,n713);
xor (n359,n360,n710);
xor (n360,n361,n708);
xor (n361,n362,n699);
xor (n362,n363,n697);
xor (n363,n364,n682);
xor (n364,n365,n680);
xor (n365,n366,n659);
xor (n366,n367,n657);
xor (n367,n368,n630);
xor (n368,n369,n628);
xor (n369,n370,n595);
xor (n370,n371,n593);
xor (n371,n372,n554);
xor (n372,n373,n552);
xor (n373,n374,n507);
xor (n374,n375,n505);
xor (n375,n376,n454);
xor (n376,n377,n452);
xor (n377,n378,n385);
xor (n378,n379,n382);
and (n379,n380,n381);
and (n382,n383,n384);
or (n385,n386,n390);
and (n386,n387,n388);
and (n387,n383,n381);
and (n388,n389,n384);
and (n390,n391,n392);
xor (n391,n387,n388);
or (n392,n393,n397);
and (n393,n394,n395);
and (n394,n389,n381);
and (n395,n396,n384);
and (n397,n398,n399);
xor (n398,n394,n395);
or (n399,n400,n404);
and (n400,n401,n402);
and (n401,n396,n381);
and (n402,n403,n384);
and (n404,n405,n406);
xor (n405,n401,n402);
or (n406,n407,n411);
and (n407,n408,n409);
and (n408,n403,n381);
and (n409,n410,n384);
and (n411,n412,n413);
xor (n412,n408,n409);
or (n413,n414,n418);
and (n414,n415,n416);
and (n415,n410,n381);
and (n416,n417,n384);
and (n418,n419,n420);
xor (n419,n415,n416);
or (n420,n421,n425);
and (n421,n422,n423);
and (n422,n417,n381);
and (n423,n424,n384);
and (n425,n426,n427);
xor (n426,n422,n423);
or (n427,n428,n432);
and (n428,n429,n430);
and (n429,n424,n381);
and (n430,n431,n384);
and (n432,n433,n434);
xor (n433,n429,n430);
or (n434,n435,n439);
and (n435,n436,n437);
and (n436,n431,n381);
and (n437,n438,n384);
and (n439,n440,n441);
xor (n440,n436,n437);
or (n441,n442,n446);
and (n442,n443,n444);
and (n443,n438,n381);
and (n444,n445,n384);
and (n446,n447,n448);
xor (n447,n443,n444);
and (n448,n449,n450);
and (n449,n445,n381);
and (n450,n451,n384);
and (n452,n389,n453);
or (n454,n455,n458);
and (n455,n456,n457);
xor (n456,n391,n392);
and (n457,n396,n453);
and (n458,n459,n460);
xor (n459,n456,n457);
or (n460,n461,n464);
and (n461,n462,n463);
xor (n462,n398,n399);
and (n463,n403,n453);
and (n464,n465,n466);
xor (n465,n462,n463);
or (n466,n467,n470);
and (n467,n468,n469);
xor (n468,n405,n406);
and (n469,n410,n453);
and (n470,n471,n472);
xor (n471,n468,n469);
or (n472,n473,n476);
and (n473,n474,n475);
xor (n474,n412,n413);
and (n475,n417,n453);
and (n476,n477,n478);
xor (n477,n474,n475);
or (n478,n479,n482);
and (n479,n480,n481);
xor (n480,n419,n420);
and (n481,n424,n453);
and (n482,n483,n484);
xor (n483,n480,n481);
or (n484,n485,n488);
and (n485,n486,n487);
xor (n486,n426,n427);
and (n487,n431,n453);
and (n488,n489,n490);
xor (n489,n486,n487);
or (n490,n491,n494);
and (n491,n492,n493);
xor (n492,n433,n434);
and (n493,n438,n453);
and (n494,n495,n496);
xor (n495,n492,n493);
or (n496,n497,n500);
and (n497,n498,n499);
xor (n498,n440,n441);
and (n499,n445,n453);
and (n500,n501,n502);
xor (n501,n498,n499);
and (n502,n503,n504);
xor (n503,n447,n448);
and (n504,n451,n453);
and (n505,n396,n506);
or (n507,n508,n511);
and (n508,n509,n510);
xor (n509,n459,n460);
and (n510,n403,n506);
and (n511,n512,n513);
xor (n512,n509,n510);
or (n513,n514,n517);
and (n514,n515,n516);
xor (n515,n465,n466);
and (n516,n410,n506);
and (n517,n518,n519);
xor (n518,n515,n516);
or (n519,n520,n523);
and (n520,n521,n522);
xor (n521,n471,n472);
and (n522,n417,n506);
and (n523,n524,n525);
xor (n524,n521,n522);
or (n525,n526,n529);
and (n526,n527,n528);
xor (n527,n477,n478);
and (n528,n424,n506);
and (n529,n530,n531);
xor (n530,n527,n528);
or (n531,n532,n535);
and (n532,n533,n534);
xor (n533,n483,n484);
and (n534,n431,n506);
and (n535,n536,n537);
xor (n536,n533,n534);
or (n537,n538,n541);
and (n538,n539,n540);
xor (n539,n489,n490);
and (n540,n438,n506);
and (n541,n542,n543);
xor (n542,n539,n540);
or (n543,n544,n547);
and (n544,n545,n546);
xor (n545,n495,n496);
and (n546,n445,n506);
and (n547,n548,n549);
xor (n548,n545,n546);
and (n549,n550,n551);
xor (n550,n501,n502);
and (n551,n451,n506);
and (n552,n403,n553);
or (n554,n555,n558);
and (n555,n556,n557);
xor (n556,n512,n513);
and (n557,n410,n553);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
xor (n562,n518,n519);
and (n563,n417,n553);
and (n564,n565,n566);
xor (n565,n562,n563);
or (n566,n567,n570);
and (n567,n568,n569);
xor (n568,n524,n525);
and (n569,n424,n553);
and (n570,n571,n572);
xor (n571,n568,n569);
or (n572,n573,n576);
and (n573,n574,n575);
xor (n574,n530,n531);
and (n575,n431,n553);
and (n576,n577,n578);
xor (n577,n574,n575);
or (n578,n579,n582);
and (n579,n580,n581);
xor (n580,n536,n537);
and (n581,n438,n553);
and (n582,n583,n584);
xor (n583,n580,n581);
or (n584,n585,n588);
and (n585,n586,n587);
xor (n586,n542,n543);
and (n587,n445,n553);
and (n588,n589,n590);
xor (n589,n586,n587);
and (n590,n591,n592);
xor (n591,n548,n549);
and (n592,n451,n553);
and (n593,n410,n594);
or (n595,n596,n599);
and (n596,n597,n598);
xor (n597,n559,n560);
and (n598,n417,n594);
and (n599,n600,n601);
xor (n600,n597,n598);
or (n601,n602,n605);
and (n602,n603,n604);
xor (n603,n565,n566);
and (n604,n424,n594);
and (n605,n606,n607);
xor (n606,n603,n604);
or (n607,n608,n611);
and (n608,n609,n610);
xor (n609,n571,n572);
and (n610,n431,n594);
and (n611,n612,n613);
xor (n612,n609,n610);
or (n613,n614,n617);
and (n614,n615,n616);
xor (n615,n577,n578);
and (n616,n438,n594);
and (n617,n618,n619);
xor (n618,n615,n616);
or (n619,n620,n623);
and (n620,n621,n622);
xor (n621,n583,n584);
and (n622,n445,n594);
and (n623,n624,n625);
xor (n624,n621,n622);
and (n625,n626,n627);
xor (n626,n589,n590);
and (n627,n451,n594);
and (n628,n417,n629);
or (n630,n631,n634);
and (n631,n632,n633);
xor (n632,n600,n601);
and (n633,n424,n629);
and (n634,n635,n636);
xor (n635,n632,n633);
or (n636,n637,n640);
and (n637,n638,n639);
xor (n638,n606,n607);
and (n639,n431,n629);
and (n640,n641,n642);
xor (n641,n638,n639);
or (n642,n643,n646);
and (n643,n644,n645);
xor (n644,n612,n613);
and (n645,n438,n629);
and (n646,n647,n648);
xor (n647,n644,n645);
or (n648,n649,n652);
and (n649,n650,n651);
xor (n650,n618,n619);
and (n651,n445,n629);
and (n652,n653,n654);
xor (n653,n650,n651);
and (n654,n655,n656);
xor (n655,n624,n625);
and (n656,n451,n629);
and (n657,n424,n658);
or (n659,n660,n663);
and (n660,n661,n662);
xor (n661,n635,n636);
and (n662,n431,n658);
and (n663,n664,n665);
xor (n664,n661,n662);
or (n665,n666,n669);
and (n666,n667,n668);
xor (n667,n641,n642);
and (n668,n438,n658);
and (n669,n670,n671);
xor (n670,n667,n668);
or (n671,n672,n675);
and (n672,n673,n674);
xor (n673,n647,n648);
and (n674,n445,n658);
and (n675,n676,n677);
xor (n676,n673,n674);
and (n677,n678,n679);
xor (n678,n653,n654);
and (n679,n451,n658);
and (n680,n431,n681);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n664,n665);
and (n685,n438,n681);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n670,n671);
and (n691,n445,n681);
and (n692,n693,n694);
xor (n693,n690,n691);
and (n694,n695,n696);
xor (n695,n676,n677);
and (n696,n451,n681);
and (n697,n438,n698);
or (n699,n700,n703);
and (n700,n701,n702);
xor (n701,n687,n688);
and (n702,n445,n698);
and (n703,n704,n705);
xor (n704,n701,n702);
and (n705,n706,n707);
xor (n706,n693,n694);
and (n707,n451,n698);
and (n708,n445,n709);
and (n710,n711,n712);
xor (n711,n704,n705);
and (n712,n451,n709);
and (n713,n451,n714);
xor (n716,n717,n1071);
xor (n717,n718,n1068);
xor (n718,n719,n1066);
xor (n719,n720,n1057);
xor (n720,n721,n1055);
xor (n721,n722,n1040);
xor (n722,n723,n1038);
xor (n723,n724,n1017);
xor (n724,n725,n1015);
xor (n725,n726,n988);
xor (n726,n727,n986);
xor (n727,n728,n953);
xor (n728,n729,n951);
xor (n729,n730,n912);
xor (n730,n731,n910);
xor (n731,n732,n865);
xor (n732,n733,n863);
xor (n733,n734,n812);
xor (n734,n735,n810);
xor (n735,n736,n743);
xor (n736,n737,n740);
and (n737,n738,n739);
wire s0n738,s1n738,notn738;
or (n738,s0n738,s1n738);
not(notn738,n715);
and (s0n738,notn738,n23);
and (s1n738,n715,n380);
wire s0n739,s1n739,notn739;
or (n739,s0n739,s1n739);
not(notn739,n715);
and (s0n739,notn739,n24);
and (s1n739,n715,n381);
and (n740,n741,n742);
wire s0n741,s1n741,notn741;
or (n741,s0n741,s1n741);
not(notn741,n715);
and (s0n741,notn741,n26);
and (s1n741,n715,n383);
wire s0n742,s1n742,notn742;
or (n742,s0n742,s1n742);
not(notn742,n715);
and (s0n742,notn742,n27);
and (s1n742,n715,n384);
or (n743,n744,n748);
and (n744,n745,n746);
and (n745,n741,n739);
and (n746,n747,n742);
wire s0n747,s1n747,notn747;
or (n747,s0n747,s1n747);
not(notn747,n715);
and (s0n747,notn747,n32);
and (s1n747,n715,n389);
and (n748,n749,n750);
xor (n749,n745,n746);
or (n750,n751,n755);
and (n751,n752,n753);
and (n752,n747,n739);
and (n753,n754,n742);
wire s0n754,s1n754,notn754;
or (n754,s0n754,s1n754);
not(notn754,n715);
and (s0n754,notn754,n39);
and (s1n754,n715,n396);
and (n755,n756,n757);
xor (n756,n752,n753);
or (n757,n758,n762);
and (n758,n759,n760);
and (n759,n754,n739);
and (n760,n761,n742);
wire s0n761,s1n761,notn761;
or (n761,s0n761,s1n761);
not(notn761,n715);
and (s0n761,notn761,n46);
and (s1n761,n715,n403);
and (n762,n763,n764);
xor (n763,n759,n760);
or (n764,n765,n769);
and (n765,n766,n767);
and (n766,n761,n739);
and (n767,n768,n742);
wire s0n768,s1n768,notn768;
or (n768,s0n768,s1n768);
not(notn768,n715);
and (s0n768,notn768,n53);
and (s1n768,n715,n410);
and (n769,n770,n771);
xor (n770,n766,n767);
or (n771,n772,n776);
and (n772,n773,n774);
and (n773,n768,n739);
and (n774,n775,n742);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n715);
and (s0n775,notn775,n60);
and (s1n775,n715,n417);
and (n776,n777,n778);
xor (n777,n773,n774);
or (n778,n779,n783);
and (n779,n780,n781);
and (n780,n775,n739);
and (n781,n782,n742);
wire s0n782,s1n782,notn782;
or (n782,s0n782,s1n782);
not(notn782,n715);
and (s0n782,notn782,n67);
and (s1n782,n715,n424);
and (n783,n784,n785);
xor (n784,n780,n781);
or (n785,n786,n790);
and (n786,n787,n788);
and (n787,n782,n739);
and (n788,n789,n742);
wire s0n789,s1n789,notn789;
or (n789,s0n789,s1n789);
not(notn789,n715);
and (s0n789,notn789,n74);
and (s1n789,n715,n431);
and (n790,n791,n792);
xor (n791,n787,n788);
or (n792,n793,n797);
and (n793,n794,n795);
and (n794,n789,n739);
and (n795,n796,n742);
wire s0n796,s1n796,notn796;
or (n796,s0n796,s1n796);
not(notn796,n715);
and (s0n796,notn796,n81);
and (s1n796,n715,n438);
and (n797,n798,n799);
xor (n798,n794,n795);
or (n799,n800,n804);
and (n800,n801,n802);
and (n801,n796,n739);
and (n802,n803,n742);
wire s0n803,s1n803,notn803;
or (n803,s0n803,s1n803);
not(notn803,n715);
and (s0n803,notn803,n88);
and (s1n803,n715,n445);
and (n804,n805,n806);
xor (n805,n801,n802);
and (n806,n807,n808);
and (n807,n803,n739);
and (n808,n809,n742);
wire s0n809,s1n809,notn809;
or (n809,s0n809,s1n809);
not(notn809,n715);
and (s0n809,notn809,n94);
and (s1n809,n715,n451);
and (n810,n747,n811);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n715);
and (s0n811,notn811,n96);
and (s1n811,n715,n453);
or (n812,n813,n816);
and (n813,n814,n815);
xor (n814,n749,n750);
and (n815,n754,n811);
and (n816,n817,n818);
xor (n817,n814,n815);
or (n818,n819,n822);
and (n819,n820,n821);
xor (n820,n756,n757);
and (n821,n761,n811);
and (n822,n823,n824);
xor (n823,n820,n821);
or (n824,n825,n828);
and (n825,n826,n827);
xor (n826,n763,n764);
and (n827,n768,n811);
and (n828,n829,n830);
xor (n829,n826,n827);
or (n830,n831,n834);
and (n831,n832,n833);
xor (n832,n770,n771);
and (n833,n775,n811);
and (n834,n835,n836);
xor (n835,n832,n833);
or (n836,n837,n840);
and (n837,n838,n839);
xor (n838,n777,n778);
and (n839,n782,n811);
and (n840,n841,n842);
xor (n841,n838,n839);
or (n842,n843,n846);
and (n843,n844,n845);
xor (n844,n784,n785);
and (n845,n789,n811);
and (n846,n847,n848);
xor (n847,n844,n845);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n791,n792);
and (n851,n796,n811);
and (n852,n853,n854);
xor (n853,n850,n851);
or (n854,n855,n858);
and (n855,n856,n857);
xor (n856,n798,n799);
and (n857,n803,n811);
and (n858,n859,n860);
xor (n859,n856,n857);
and (n860,n861,n862);
xor (n861,n805,n806);
and (n862,n809,n811);
and (n863,n754,n864);
wire s0n864,s1n864,notn864;
or (n864,s0n864,s1n864);
not(notn864,n715);
and (s0n864,notn864,n149);
and (s1n864,n715,n506);
or (n865,n866,n869);
and (n866,n867,n868);
xor (n867,n817,n818);
and (n868,n761,n864);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n875);
and (n872,n873,n874);
xor (n873,n823,n824);
and (n874,n768,n864);
and (n875,n876,n877);
xor (n876,n873,n874);
or (n877,n878,n881);
and (n878,n879,n880);
xor (n879,n829,n830);
and (n880,n775,n864);
and (n881,n882,n883);
xor (n882,n879,n880);
or (n883,n884,n887);
and (n884,n885,n886);
xor (n885,n835,n836);
and (n886,n782,n864);
and (n887,n888,n889);
xor (n888,n885,n886);
or (n889,n890,n893);
and (n890,n891,n892);
xor (n891,n841,n842);
and (n892,n789,n864);
and (n893,n894,n895);
xor (n894,n891,n892);
or (n895,n896,n899);
and (n896,n897,n898);
xor (n897,n847,n848);
and (n898,n796,n864);
and (n899,n900,n901);
xor (n900,n897,n898);
or (n901,n902,n905);
and (n902,n903,n904);
xor (n903,n853,n854);
and (n904,n803,n864);
and (n905,n906,n907);
xor (n906,n903,n904);
and (n907,n908,n909);
xor (n908,n859,n860);
and (n909,n809,n864);
and (n910,n761,n911);
wire s0n911,s1n911,notn911;
or (n911,s0n911,s1n911);
not(notn911,n715);
and (s0n911,notn911,n196);
and (s1n911,n715,n553);
or (n912,n913,n916);
and (n913,n914,n915);
xor (n914,n870,n871);
and (n915,n768,n911);
and (n916,n917,n918);
xor (n917,n914,n915);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n876,n877);
and (n921,n775,n911);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n882,n883);
and (n927,n782,n911);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n888,n889);
and (n933,n789,n911);
and (n934,n935,n936);
xor (n935,n932,n933);
or (n936,n937,n940);
and (n937,n938,n939);
xor (n938,n894,n895);
and (n939,n796,n911);
and (n940,n941,n942);
xor (n941,n938,n939);
or (n942,n943,n946);
and (n943,n944,n945);
xor (n944,n900,n901);
and (n945,n803,n911);
and (n946,n947,n948);
xor (n947,n944,n945);
and (n948,n949,n950);
xor (n949,n906,n907);
and (n950,n809,n911);
and (n951,n768,n952);
wire s0n952,s1n952,notn952;
or (n952,s0n952,s1n952);
not(notn952,n715);
and (s0n952,notn952,n237);
and (s1n952,n715,n594);
or (n953,n954,n957);
and (n954,n955,n956);
xor (n955,n917,n918);
and (n956,n775,n952);
and (n957,n958,n959);
xor (n958,n955,n956);
or (n959,n960,n963);
and (n960,n961,n962);
xor (n961,n923,n924);
and (n962,n782,n952);
and (n963,n964,n965);
xor (n964,n961,n962);
or (n965,n966,n969);
and (n966,n967,n968);
xor (n967,n929,n930);
and (n968,n789,n952);
and (n969,n970,n971);
xor (n970,n967,n968);
or (n971,n972,n975);
and (n972,n973,n974);
xor (n973,n935,n936);
and (n974,n796,n952);
and (n975,n976,n977);
xor (n976,n973,n974);
or (n977,n978,n981);
and (n978,n979,n980);
xor (n979,n941,n942);
and (n980,n803,n952);
and (n981,n982,n983);
xor (n982,n979,n980);
and (n983,n984,n985);
xor (n984,n947,n948);
and (n985,n809,n952);
and (n986,n775,n987);
wire s0n987,s1n987,notn987;
or (n987,s0n987,s1n987);
not(notn987,n715);
and (s0n987,notn987,n272);
and (s1n987,n715,n629);
or (n988,n989,n992);
and (n989,n990,n991);
xor (n990,n958,n959);
and (n991,n782,n987);
and (n992,n993,n994);
xor (n993,n990,n991);
or (n994,n995,n998);
and (n995,n996,n997);
xor (n996,n964,n965);
and (n997,n789,n987);
and (n998,n999,n1000);
xor (n999,n996,n997);
or (n1000,n1001,n1004);
and (n1001,n1002,n1003);
xor (n1002,n970,n971);
and (n1003,n796,n987);
and (n1004,n1005,n1006);
xor (n1005,n1002,n1003);
or (n1006,n1007,n1010);
and (n1007,n1008,n1009);
xor (n1008,n976,n977);
and (n1009,n803,n987);
and (n1010,n1011,n1012);
xor (n1011,n1008,n1009);
and (n1012,n1013,n1014);
xor (n1013,n982,n983);
and (n1014,n809,n987);
and (n1015,n782,n1016);
wire s0n1016,s1n1016,notn1016;
or (n1016,s0n1016,s1n1016);
not(notn1016,n715);
and (s0n1016,notn1016,n301);
and (s1n1016,n715,n658);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
xor (n1019,n993,n994);
and (n1020,n789,n1016);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
or (n1023,n1024,n1027);
and (n1024,n1025,n1026);
xor (n1025,n999,n1000);
and (n1026,n796,n1016);
and (n1027,n1028,n1029);
xor (n1028,n1025,n1026);
or (n1029,n1030,n1033);
and (n1030,n1031,n1032);
xor (n1031,n1005,n1006);
and (n1032,n803,n1016);
and (n1033,n1034,n1035);
xor (n1034,n1031,n1032);
and (n1035,n1036,n1037);
xor (n1036,n1011,n1012);
and (n1037,n809,n1016);
and (n1038,n789,n1039);
wire s0n1039,s1n1039,notn1039;
or (n1039,s0n1039,s1n1039);
not(notn1039,n715);
and (s0n1039,notn1039,n324);
and (s1n1039,n715,n681);
or (n1040,n1041,n1044);
and (n1041,n1042,n1043);
xor (n1042,n1022,n1023);
and (n1043,n796,n1039);
and (n1044,n1045,n1046);
xor (n1045,n1042,n1043);
or (n1046,n1047,n1050);
and (n1047,n1048,n1049);
xor (n1048,n1028,n1029);
and (n1049,n803,n1039);
and (n1050,n1051,n1052);
xor (n1051,n1048,n1049);
and (n1052,n1053,n1054);
xor (n1053,n1034,n1035);
and (n1054,n809,n1039);
and (n1055,n796,n1056);
wire s0n1056,s1n1056,notn1056;
or (n1056,s0n1056,s1n1056);
not(notn1056,n715);
and (s0n1056,notn1056,n341);
and (s1n1056,n715,n698);
or (n1057,n1058,n1061);
and (n1058,n1059,n1060);
xor (n1059,n1045,n1046);
and (n1060,n803,n1056);
and (n1061,n1062,n1063);
xor (n1062,n1059,n1060);
and (n1063,n1064,n1065);
xor (n1064,n1051,n1052);
and (n1065,n809,n1056);
and (n1066,n803,n1067);
wire s0n1067,s1n1067,notn1067;
or (n1067,s0n1067,s1n1067);
not(notn1067,n715);
and (s0n1067,notn1067,n352);
and (s1n1067,n715,n709);
and (n1068,n1069,n1070);
xor (n1069,n1062,n1063);
and (n1070,n809,n1067);
and (n1071,n809,n1072);
wire s0n1072,s1n1072,notn1072;
or (n1072,s0n1072,s1n1072);
not(notn1072,n715);
and (s0n1072,notn1072,n357);
and (s1n1072,n715,n714);
endmodule
