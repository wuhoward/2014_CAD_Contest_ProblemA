module top (out,n12,n14,n15,n17,n20,n24,n26,n28,n31
        ,n35,n37,n39,n42,n48,n50,n52,n55,n59,n61
        ,n63,n66,n71,n73,n74,n88,n102,n103,n175,n184
        ,n185,n221,n293,n323,n324,n469,n473,n475,n501,n502
        ,n609,n626,n627,n794,n798,n800,n811,n823,n837);
output out;
input n12;
input n14;
input n15;
input n17;
input n20;
input n24;
input n26;
input n28;
input n31;
input n35;
input n37;
input n39;
input n42;
input n48;
input n50;
input n52;
input n55;
input n59;
input n61;
input n63;
input n66;
input n71;
input n73;
input n74;
input n88;
input n102;
input n103;
input n175;
input n184;
input n185;
input n221;
input n293;
input n323;
input n324;
input n469;
input n473;
input n475;
input n501;
input n502;
input n609;
input n626;
input n627;
input n794;
input n798;
input n800;
input n811;
input n823;
input n837;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n16;
wire n18;
wire n19;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n36;
wire n38;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n51;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n60;
wire n62;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n470;
wire n471;
wire n472;
wire n474;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n795;
wire n796;
wire n797;
wire n799;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
xor (out,n0,n2797);
xnor (n0,n1,n2739);
nand (n1,n2,n366);
nand (n2,n3,n243);
xor (n3,n4,n200);
xor (n4,n5,n91);
xor (n5,n6,n78);
xor (n6,n7,n43);
xor (n7,n8,n32);
xor (n8,n9,n21);
xor (n9,n10,n20);
or (n10,n11,n16);
and (n11,n12,n13);
xor (n13,n14,n15);
and (n16,n17,n18);
nor (n18,n13,n19);
xnor (n19,n20,n14);
xor (n21,n22,n31);
or (n22,n23,n27);
and (n23,n24,n25);
xor (n25,n26,n20);
and (n27,n28,n29);
nor (n29,n25,n30);
xnor (n30,n31,n26);
xor (n32,n33,n42);
or (n33,n34,n38);
and (n34,n35,n36);
xor (n36,n37,n31);
and (n38,n39,n40);
nor (n40,n36,n41);
xnor (n41,n42,n37);
xor (n43,n44,n67);
xor (n44,n45,n56);
xor (n45,n46,n55);
or (n46,n47,n51);
and (n47,n48,n49);
xor (n49,n50,n42);
and (n51,n52,n53);
nor (n53,n49,n54);
xnor (n54,n55,n50);
xor (n56,n57,n66);
or (n57,n58,n62);
and (n58,n59,n60);
xor (n60,n61,n55);
and (n62,n63,n64);
nor (n64,n60,n65);
xnor (n65,n66,n61);
not (n67,n68);
xor (n68,n69,n15);
or (n69,n70,n75);
and (n70,n71,n72);
xor (n72,n73,n74);
and (n75,n71,n76);
nor (n76,n72,n77);
xnor (n77,n15,n73);
nand (n78,n79,n89,n90);
nand (n79,n80,n84);
xor (n80,n81,n55);
or (n81,n82,n83);
and (n82,n52,n49);
and (n83,n59,n53);
xor (n84,n85,n66);
or (n85,n86,n87);
and (n86,n63,n60);
and (n87,n88,n64);
nand (n89,n66,n84);
nand (n90,n80,n66);
xor (n91,n92,n162);
xor (n92,n93,n128);
xor (n93,n94,n116);
xor (n94,n66,n95);
nand (n95,n96,n110,n115);
nand (n96,n97,n107);
not (n97,n98);
xor (n98,n99,n74);
or (n99,n100,n104);
and (n100,n71,n101);
xor (n101,n102,n103);
and (n104,n71,n105);
nor (n105,n101,n106);
xnor (n106,n74,n102);
xor (n107,n108,n15);
or (n108,n70,n109);
and (n109,n12,n76);
nand (n110,n111,n107);
xor (n111,n112,n31);
or (n112,n113,n114);
and (n113,n28,n25);
and (n114,n35,n29);
nand (n115,n97,n111);
nand (n116,n117,n122,n127);
nand (n117,n118,n98);
xor (n118,n119,n20);
or (n119,n120,n121);
and (n120,n17,n13);
and (n121,n24,n18);
nand (n122,n123,n98);
xor (n123,n124,n42);
or (n124,n125,n126);
and (n125,n39,n36);
and (n126,n48,n40);
nand (n127,n118,n123);
nand (n128,n129,n148,n161);
nand (n129,n130,n132);
xor (n130,n131,n111);
xor (n131,n97,n107);
nand (n132,n133,n142,n147);
nand (n133,n134,n138);
xor (n134,n135,n15);
or (n135,n136,n137);
and (n136,n12,n72);
and (n137,n17,n76);
xor (n138,n139,n31);
or (n139,n140,n141);
and (n140,n35,n25);
and (n141,n39,n29);
nand (n142,n143,n138);
xor (n143,n144,n20);
or (n144,n145,n146);
and (n145,n24,n13);
and (n146,n28,n18);
nand (n147,n134,n143);
nand (n148,n149,n132);
nand (n149,n150,n155,n160);
nand (n150,n97,n151);
xor (n151,n152,n42);
or (n152,n153,n154);
and (n153,n48,n36);
and (n154,n52,n40);
nand (n155,n156,n151);
xor (n156,n157,n55);
or (n157,n158,n159);
and (n158,n59,n49);
and (n159,n63,n53);
nand (n160,n97,n156);
nand (n161,n130,n149);
nand (n162,n163,n168,n199);
nand (n163,n164,n166);
xor (n164,n165,n66);
xor (n165,n80,n84);
xor (n166,n167,n123);
xor (n167,n118,n98);
nand (n168,n169,n166);
nand (n169,n170,n176,n198);
nand (n170,n171,n66);
xor (n171,n172,n66);
or (n172,n173,n174);
and (n173,n88,n60);
and (n174,n175,n64);
nand (n176,n177,n66);
nand (n177,n178,n192,n197);
nand (n178,n179,n189);
not (n179,n180);
xor (n180,n181,n103);
or (n181,n182,n186);
and (n182,n71,n183);
xor (n183,n184,n185);
and (n186,n71,n187);
nor (n187,n183,n188);
xnor (n188,n103,n184);
xor (n189,n190,n74);
or (n190,n100,n191);
and (n191,n12,n105);
nand (n192,n193,n189);
xor (n193,n194,n15);
or (n194,n195,n196);
and (n195,n17,n72);
and (n196,n24,n76);
nand (n197,n179,n193);
nand (n198,n171,n177);
nand (n199,n164,n169);
nand (n200,n201,n239,n242);
nand (n201,n202,n237);
nand (n202,n203,n223,n236);
nand (n203,n204,n206);
xor (n204,n205,n143);
xor (n205,n134,n138);
nand (n206,n207,n216,n222);
nand (n207,n208,n212);
xor (n208,n209,n20);
or (n209,n210,n211);
and (n210,n28,n13);
and (n211,n35,n18);
xor (n212,n213,n31);
or (n213,n214,n215);
and (n214,n39,n25);
and (n215,n48,n29);
nand (n216,n217,n212);
xor (n217,n218,n66);
or (n218,n219,n220);
and (n219,n175,n60);
and (n220,n221,n64);
nand (n222,n208,n217);
nand (n223,n224,n206);
nand (n224,n225,n230,n235);
nand (n225,n180,n226);
xor (n226,n227,n42);
or (n227,n228,n229);
and (n228,n52,n36);
and (n229,n59,n40);
nand (n230,n231,n226);
xor (n231,n232,n55);
or (n232,n233,n234);
and (n233,n63,n49);
and (n234,n88,n53);
nand (n235,n180,n231);
nand (n236,n204,n224);
xor (n237,n238,n149);
xor (n238,n130,n132);
nand (n239,n240,n237);
xor (n240,n241,n169);
xor (n241,n164,n166);
nand (n242,n202,n240);
nand (n243,n244,n276,n365);
nand (n244,n245,n274);
nand (n245,n246,n250,n273);
nand (n246,n247,n249);
xor (n247,n248,n156);
xor (n248,n97,n151);
xor (n249,n172,n177);
nand (n250,n251,n249);
nand (n251,n252,n255,n272);
nand (n252,n66,n253);
xor (n253,n254,n193);
xor (n254,n179,n189);
nand (n255,n256,n253);
nand (n256,n257,n266,n271);
nand (n257,n258,n262);
xor (n258,n259,n74);
or (n259,n260,n261);
and (n260,n12,n101);
and (n261,n17,n105);
xor (n262,n263,n15);
or (n263,n264,n265);
and (n264,n24,n72);
and (n265,n28,n76);
nand (n266,n267,n262);
xor (n267,n268,n20);
or (n268,n269,n270);
and (n269,n35,n13);
and (n270,n39,n18);
nand (n271,n258,n267);
nand (n272,n66,n256);
nand (n273,n247,n251);
xor (n274,n275,n240);
xor (n275,n202,n237);
nand (n276,n277,n274);
nand (n277,n278,n302,n364);
nand (n278,n279,n281);
xor (n279,n280,n224);
xor (n280,n204,n206);
nand (n281,n282,n298,n301);
nand (n282,n283,n296);
nand (n283,n284,n294,n295);
nand (n284,n285,n289);
xor (n285,n286,n31);
or (n286,n287,n288);
and (n287,n48,n25);
and (n288,n52,n29);
xor (n289,n290,n66);
or (n290,n291,n292);
and (n291,n221,n60);
and (n292,n293,n64);
nand (n294,n179,n289);
nand (n295,n285,n179);
xor (n296,n297,n217);
xor (n297,n208,n212);
nand (n298,n299,n296);
xor (n299,n300,n231);
xor (n300,n180,n226);
nand (n301,n283,n299);
nand (n302,n303,n281);
nand (n303,n304,n360,n363);
nand (n304,n305,n338);
nand (n305,n306,n315,n337);
nand (n306,n307,n311);
xor (n307,n308,n42);
or (n308,n309,n310);
and (n309,n59,n36);
and (n310,n63,n40);
xor (n311,n312,n55);
or (n312,n313,n314);
and (n313,n88,n49);
and (n314,n175,n53);
nand (n315,n316,n311);
nand (n316,n317,n331,n336);
nand (n317,n318,n328);
not (n318,n319);
xor (n319,n320,n185);
or (n320,n321,n325);
and (n321,n71,n322);
xor (n322,n323,n324);
and (n325,n71,n326);
nor (n326,n322,n327);
xnor (n327,n185,n323);
xor (n328,n329,n103);
or (n329,n182,n330);
and (n330,n12,n187);
nand (n331,n332,n328);
xor (n332,n333,n15);
or (n333,n334,n335);
and (n334,n28,n72);
and (n335,n35,n76);
nand (n336,n318,n332);
nand (n337,n307,n316);
nand (n338,n339,n342,n359);
nand (n339,n66,n340);
xor (n340,n341,n267);
xor (n341,n258,n262);
nand (n342,n343,n340);
nand (n343,n344,n353,n358);
nand (n344,n345,n349);
xor (n345,n346,n74);
or (n346,n347,n348);
and (n347,n17,n101);
and (n348,n24,n105);
xor (n349,n350,n20);
or (n350,n351,n352);
and (n351,n39,n13);
and (n352,n48,n18);
nand (n353,n354,n349);
xor (n354,n355,n31);
or (n355,n356,n357);
and (n356,n52,n25);
and (n357,n59,n29);
nand (n358,n345,n354);
nand (n359,n66,n343);
nand (n360,n361,n338);
xor (n361,n362,n256);
xor (n362,n66,n253);
nand (n363,n305,n361);
nand (n364,n279,n303);
nand (n365,n245,n277);
nand (n366,n367,n2737);
nand (n367,n368,n775);
nor (n368,n369,n769);
nor (n369,n370,n745);
nor (n370,n371,n743);
nor (n371,n372,n718);
nand (n372,n373,n680);
nand (n373,n374,n596,n679);
nand (n374,n375,n459);
xor (n375,n376,n449);
xor (n376,n377,n399);
xor (n377,n378,n383);
xor (n378,n379,n66);
xor (n379,n380,n42);
or (n380,n381,n382);
and (n381,n63,n36);
and (n382,n88,n40);
nand (n383,n384,n393,n398);
nand (n384,n385,n389);
xor (n385,n386,n15);
or (n386,n387,n388);
and (n387,n35,n72);
and (n388,n39,n76);
xor (n389,n390,n103);
or (n390,n391,n392);
and (n391,n12,n183);
and (n392,n17,n187);
nand (n393,n394,n389);
xor (n394,n395,n74);
or (n395,n396,n397);
and (n396,n24,n101);
and (n397,n28,n105);
nand (n398,n385,n394);
nand (n399,n400,n431,n448);
nand (n400,n401,n417);
nand (n401,n402,n411,n416);
nand (n402,n403,n407);
xor (n403,n404,n15);
or (n404,n405,n406);
and (n405,n39,n72);
and (n406,n48,n76);
xor (n407,n408,n103);
or (n408,n409,n410);
and (n409,n17,n183);
and (n410,n24,n187);
nand (n411,n412,n407);
xor (n412,n413,n20);
or (n413,n414,n415);
and (n414,n52,n13);
and (n415,n59,n18);
nand (n416,n403,n412);
xor (n417,n418,n427);
xor (n418,n419,n423);
xor (n419,n420,n20);
or (n420,n421,n422);
and (n421,n48,n13);
and (n422,n52,n18);
xor (n423,n424,n31);
or (n424,n425,n426);
and (n425,n59,n25);
and (n426,n63,n29);
xor (n427,n428,n55);
or (n428,n429,n430);
and (n429,n221,n49);
and (n430,n293,n53);
nand (n431,n432,n417);
nand (n432,n433,n442,n447);
nand (n433,n434,n438);
xor (n434,n435,n185);
or (n435,n436,n437);
and (n436,n12,n322);
and (n437,n17,n326);
xor (n438,n439,n31);
or (n439,n440,n441);
and (n440,n63,n25);
and (n441,n88,n29);
nand (n442,n443,n438);
xor (n443,n444,n42);
or (n444,n445,n446);
and (n445,n175,n36);
and (n446,n221,n40);
nand (n447,n434,n443);
nand (n448,n401,n432);
xor (n449,n450,n455);
xor (n450,n451,n453);
xor (n451,n452,n332);
xor (n452,n318,n328);
xor (n453,n454,n354);
xor (n454,n345,n349);
nand (n455,n456,n457,n458);
nand (n456,n419,n423);
nand (n457,n427,n423);
nand (n458,n419,n427);
xor (n459,n460,n535);
xor (n460,n461,n515);
nand (n461,n462,n488,n514);
nand (n462,n463,n478);
nand (n463,n464,n476,n477);
nand (n464,n465,n470);
xor (n465,n466,n55);
or (n466,n467,n468);
and (n467,n293,n49);
and (n468,n469,n53);
xor (n470,n471,n66);
or (n471,n472,n474);
and (n472,n473,n60);
and (n474,n475,n64);
nand (n476,n66,n470);
nand (n477,n465,n66);
xor (n478,n479,n484);
xor (n479,n480,n318);
xor (n480,n481,n66);
or (n481,n482,n483);
and (n482,n469,n60);
and (n483,n473,n64);
xor (n484,n485,n42);
or (n485,n486,n487);
and (n486,n88,n36);
and (n487,n175,n40);
nand (n488,n489,n478);
xor (n489,n490,n512);
xor (n490,n66,n491);
nand (n491,n492,n506,n511);
nand (n492,n493,n496);
xor (n493,n494,n185);
or (n494,n321,n495);
and (n495,n12,n326);
not (n496,n497);
xor (n497,n498,n324);
or (n498,n499,n503);
and (n499,n71,n500);
xor (n500,n501,n502);
and (n503,n71,n504);
nor (n504,n500,n505);
xnor (n505,n324,n501);
nand (n506,n507,n496);
xor (n507,n508,n74);
or (n508,n509,n510);
and (n509,n28,n101);
and (n510,n35,n105);
nand (n511,n493,n507);
xor (n512,n513,n394);
xor (n513,n385,n389);
nand (n514,n463,n489);
xor (n515,n516,n531);
xor (n516,n517,n521);
nand (n517,n518,n519,n520);
nand (n518,n480,n318);
nand (n519,n484,n318);
nand (n520,n480,n484);
xor (n521,n522,n319);
xor (n522,n523,n527);
xor (n523,n524,n55);
or (n524,n525,n526);
and (n525,n175,n49);
and (n526,n221,n53);
xor (n527,n528,n66);
or (n528,n529,n530);
and (n529,n293,n60);
and (n530,n469,n64);
nand (n531,n532,n533,n534);
nand (n532,n66,n491);
nand (n533,n512,n491);
nand (n534,n66,n512);
nand (n535,n536,n592,n595);
nand (n536,n537,n557);
nand (n537,n538,n553,n556);
nand (n538,n539,n551);
nand (n539,n540,n545,n550);
nand (n540,n497,n541);
xor (n541,n542,n74);
or (n542,n543,n544);
and (n543,n35,n101);
and (n544,n39,n105);
nand (n545,n546,n541);
xor (n546,n547,n15);
or (n547,n548,n549);
and (n548,n48,n72);
and (n549,n52,n76);
nand (n550,n497,n546);
xor (n551,n552,n412);
xor (n552,n403,n407);
nand (n553,n554,n551);
xor (n554,n555,n507);
xor (n555,n493,n496);
nand (n556,n539,n554);
nand (n557,n558,n588,n591);
nand (n558,n559,n572);
nand (n559,n560,n566,n571);
nand (n560,n561,n565);
xor (n561,n562,n103);
or (n562,n563,n564);
and (n563,n24,n183);
and (n564,n28,n187);
not (n565,n434);
nand (n566,n567,n565);
xor (n567,n568,n20);
or (n568,n569,n570);
and (n569,n59,n13);
and (n570,n63,n18);
nand (n571,n561,n567);
nand (n572,n573,n582,n587);
nand (n573,n574,n578);
xor (n574,n575,n31);
or (n575,n576,n577);
and (n576,n88,n25);
and (n577,n175,n29);
xor (n578,n579,n42);
or (n579,n580,n581);
and (n580,n221,n36);
and (n581,n293,n40);
nand (n582,n583,n578);
xor (n583,n584,n55);
or (n584,n585,n586);
and (n585,n469,n49);
and (n586,n473,n53);
nand (n587,n574,n583);
nand (n588,n589,n572);
xor (n589,n590,n443);
xor (n590,n434,n438);
nand (n591,n559,n589);
nand (n592,n593,n557);
xor (n593,n594,n432);
xor (n594,n401,n417);
nand (n595,n537,n593);
nand (n596,n597,n459);
nand (n597,n598,n675,n678);
nand (n598,n599,n601);
xor (n599,n600,n489);
xor (n600,n463,n478);
nand (n601,n602,n635,n674);
nand (n602,n603,n633);
nand (n603,n604,n610,n632);
nand (n604,n605,n66);
xor (n605,n606,n66);
or (n606,n607,n608);
and (n607,n475,n60);
and (n608,n609,n64);
nand (n610,n611,n66);
nand (n611,n612,n620,n631);
nand (n612,n613,n616);
xor (n613,n614,n324);
or (n614,n499,n615);
and (n615,n12,n504);
xor (n616,n617,n185);
or (n617,n618,n619);
and (n618,n17,n322);
and (n619,n24,n326);
nand (n620,n621,n616);
not (n621,n622);
xor (n622,n623,n502);
or (n623,n624,n628);
and (n624,n71,n625);
xor (n625,n626,n627);
and (n628,n71,n629);
nor (n629,n625,n630);
xnor (n630,n502,n626);
nand (n631,n613,n621);
nand (n632,n605,n611);
xor (n633,n634,n66);
xor (n634,n465,n470);
nand (n635,n636,n633);
nand (n636,n637,n656,n673);
nand (n637,n638,n654);
nand (n638,n639,n648,n653);
nand (n639,n640,n644);
xor (n640,n641,n103);
or (n641,n642,n643);
and (n642,n28,n183);
and (n643,n35,n187);
xor (n644,n645,n74);
or (n645,n646,n647);
and (n646,n39,n101);
and (n647,n48,n105);
nand (n648,n649,n644);
xor (n649,n650,n15);
or (n650,n651,n652);
and (n651,n52,n72);
and (n652,n59,n76);
nand (n653,n640,n649);
xor (n654,n655,n546);
xor (n655,n497,n541);
nand (n656,n657,n654);
nand (n657,n658,n667,n672);
nand (n658,n659,n663);
xor (n659,n660,n31);
or (n660,n661,n662);
and (n661,n175,n25);
and (n662,n221,n29);
xor (n663,n664,n324);
or (n664,n665,n666);
and (n665,n12,n500);
and (n666,n17,n504);
nand (n667,n668,n663);
xor (n668,n669,n20);
or (n669,n670,n671);
and (n670,n63,n13);
and (n671,n88,n18);
nand (n672,n659,n668);
nand (n673,n638,n657);
nand (n674,n603,n636);
nand (n675,n676,n601);
xor (n676,n677,n593);
xor (n677,n537,n557);
nand (n678,n599,n676);
nand (n679,n375,n597);
xor (n680,n681,n714);
xor (n681,n682,n686);
nand (n682,n683,n684,n685);
nand (n683,n377,n399);
nand (n684,n449,n399);
nand (n685,n377,n449);
xor (n686,n687,n702);
xor (n687,n688,n692);
nand (n688,n689,n690,n691);
nand (n689,n517,n521);
nand (n690,n531,n521);
nand (n691,n517,n531);
xor (n692,n693,n700);
xor (n693,n694,n698);
nand (n694,n695,n696,n697);
nand (n695,n523,n527);
nand (n696,n319,n527);
nand (n697,n523,n319);
xor (n698,n699,n316);
xor (n699,n307,n311);
xor (n700,n701,n179);
xor (n701,n285,n289);
xor (n702,n703,n710);
xor (n703,n704,n708);
nand (n704,n705,n706,n707);
nand (n705,n379,n66);
nand (n706,n383,n66);
nand (n707,n379,n383);
xor (n708,n709,n343);
xor (n709,n66,n340);
nand (n710,n711,n712,n713);
nand (n711,n451,n453);
nand (n712,n455,n453);
nand (n713,n451,n455);
nand (n714,n715,n716,n717);
nand (n715,n461,n515);
nand (n716,n535,n515);
nand (n717,n461,n535);
nor (n718,n719,n723);
nand (n719,n720,n721,n722);
nand (n720,n682,n686);
nand (n721,n714,n686);
nand (n722,n682,n714);
xor (n723,n724,n739);
xor (n724,n725,n727);
xor (n725,n726,n361);
xor (n726,n305,n338);
xor (n727,n728,n735);
xor (n728,n729,n731);
xor (n729,n730,n299);
xor (n730,n283,n296);
nand (n731,n732,n733,n734);
nand (n732,n694,n698);
nand (n733,n700,n698);
nand (n734,n694,n700);
nand (n735,n736,n737,n738);
nand (n736,n704,n708);
nand (n737,n710,n708);
nand (n738,n704,n710);
nand (n739,n740,n741,n742);
nand (n740,n688,n692);
nand (n741,n702,n692);
nand (n742,n688,n702);
not (n743,n744);
nand (n744,n719,n723);
not (n745,n746);
nor (n746,n747,n762);
nor (n747,n748,n752);
nand (n748,n749,n750,n751);
nand (n749,n725,n727);
nand (n750,n739,n727);
nand (n751,n725,n739);
xor (n752,n753,n758);
xor (n753,n754,n756);
xor (n754,n755,n251);
xor (n755,n247,n249);
xor (n756,n757,n303);
xor (n757,n279,n281);
nand (n758,n759,n760,n761);
nand (n759,n729,n731);
nand (n760,n735,n731);
nand (n761,n729,n735);
nor (n762,n763,n767);
nand (n763,n764,n765,n766);
nand (n764,n754,n756);
nand (n765,n758,n756);
nand (n766,n754,n758);
xor (n767,n768,n277);
xor (n768,n245,n274);
not (n769,n770);
nor (n770,n771,n773);
nor (n771,n772,n762);
nand (n772,n748,n752);
not (n773,n774);
nand (n774,n763,n767);
nand (n775,n776,n2733);
nand (n776,n777,n2307);
nor (n777,n778,n2275);
nor (n778,n779,n1748);
nor (n779,n780,n1733);
nor (n780,n781,n1454);
nand (n781,n782,n1237);
nor (n782,n783,n1136);
nor (n783,n784,n1046);
nand (n784,n785,n961,n1045);
nand (n785,n786,n863);
xor (n786,n787,n839);
xor (n787,n788,n813);
xor (n788,n789,n801);
xor (n789,n790,n795);
xor (n790,n791,n20);
or (n791,n792,n793);
and (n792,n609,n13);
and (n793,n794,n18);
xor (n795,n796,n31);
or (n796,n797,n799);
and (n797,n798,n25);
and (n799,n800,n29);
xor (n801,n802,n806);
xor (n802,n803,n502);
or (n803,n804,n805);
and (n804,n39,n625);
and (n805,n48,n629);
xnor (n806,n807,n627);
nor (n807,n808,n812);
and (n808,n35,n809);
and (n809,n810,n627);
not (n810,n811);
and (n812,n28,n811);
nand (n813,n814,n824,n838);
nand (n814,n815,n819);
xor (n815,n816,n20);
or (n816,n817,n818);
and (n817,n794,n13);
and (n818,n798,n18);
xor (n819,n820,n31);
or (n820,n821,n822);
and (n821,n800,n25);
and (n822,n823,n29);
nand (n824,n825,n819);
xor (n825,n826,n835);
xor (n826,n827,n831);
xor (n827,n828,n502);
or (n828,n829,n830);
and (n829,n48,n625);
and (n830,n52,n629);
xor (n831,n832,n185);
or (n832,n833,n834);
and (n833,n88,n322);
and (n834,n175,n326);
xnor (n835,n836,n42);
nand (n836,n837,n36);
nand (n838,n815,n825);
xor (n839,n840,n849);
xor (n840,n841,n845);
xor (n841,n842,n42);
or (n842,n843,n844);
and (n843,n823,n36);
and (n844,n837,n40);
nand (n845,n846,n847,n848);
nand (n846,n827,n831);
nand (n847,n835,n831);
nand (n848,n827,n835);
xor (n849,n850,n859);
xor (n850,n851,n855);
xor (n851,n852,n185);
or (n852,n853,n854);
and (n853,n63,n322);
and (n854,n88,n326);
xor (n855,n856,n324);
or (n856,n857,n858);
and (n857,n52,n500);
and (n858,n59,n504);
xor (n859,n860,n103);
or (n860,n861,n862);
and (n861,n175,n183);
and (n862,n221,n187);
nand (n863,n864,n918,n960);
nand (n864,n865,n867);
xor (n865,n866,n825);
xor (n866,n815,n819);
xor (n867,n868,n907);
xor (n868,n869,n885);
nand (n869,n870,n879,n884);
nand (n870,n871,n875);
xor (n871,n872,n185);
or (n872,n873,n874);
and (n873,n175,n322);
and (n874,n221,n326);
xor (n875,n876,n324);
or (n876,n877,n878);
and (n877,n63,n500);
and (n878,n88,n504);
nand (n879,n880,n875);
xor (n880,n881,n103);
or (n881,n882,n883);
and (n882,n293,n183);
and (n883,n469,n187);
nand (n884,n871,n880);
nand (n885,n886,n901,n906);
nand (n886,n887,n896);
xor (n887,n888,n892);
xnor (n888,n889,n627);
nor (n889,n890,n891);
and (n890,n48,n809);
and (n891,n39,n811);
xor (n892,n893,n502);
or (n893,n894,n895);
and (n894,n52,n625);
and (n895,n59,n629);
and (n896,n897,n31);
xnor (n897,n898,n627);
nor (n898,n899,n900);
and (n899,n52,n809);
and (n900,n48,n811);
nand (n901,n902,n896);
xor (n902,n903,n74);
or (n903,n904,n905);
and (n904,n473,n101);
and (n905,n475,n105);
nand (n906,n887,n902);
xor (n907,n908,n914);
xor (n908,n909,n913);
xor (n909,n910,n74);
or (n910,n911,n912);
and (n911,n469,n101);
and (n912,n473,n105);
and (n913,n888,n892);
xor (n914,n915,n15);
or (n915,n916,n917);
and (n916,n475,n72);
and (n917,n609,n76);
nand (n918,n919,n867);
nand (n919,n920,n944,n959);
nand (n920,n921,n942);
nand (n921,n922,n936,n941);
nand (n922,n923,n932);
and (n923,n924,n928);
xnor (n924,n925,n627);
nor (n925,n926,n927);
and (n926,n59,n809);
and (n927,n52,n811);
xor (n928,n929,n502);
or (n929,n930,n931);
and (n930,n63,n625);
and (n931,n88,n629);
xor (n932,n933,n74);
or (n933,n934,n935);
and (n934,n475,n101);
and (n935,n609,n105);
nand (n936,n937,n932);
xor (n937,n938,n15);
or (n938,n939,n940);
and (n939,n794,n72);
and (n940,n798,n76);
nand (n941,n923,n937);
xor (n942,n943,n902);
xor (n943,n887,n896);
nand (n944,n945,n942);
xor (n945,n946,n955);
xor (n946,n947,n951);
xor (n947,n948,n15);
or (n948,n949,n950);
and (n949,n609,n72);
and (n950,n794,n76);
xor (n951,n952,n20);
or (n952,n953,n954);
and (n953,n798,n13);
and (n954,n800,n18);
xor (n955,n956,n31);
or (n956,n957,n958);
and (n957,n823,n25);
and (n958,n837,n29);
nand (n959,n921,n945);
nand (n960,n865,n919);
nand (n961,n962,n863);
xor (n962,n963,n1002);
xor (n963,n964,n968);
nand (n964,n965,n966,n967);
nand (n965,n869,n885);
nand (n966,n907,n885);
nand (n967,n869,n907);
xor (n968,n969,n991);
xor (n969,n970,n987);
nand (n970,n971,n981,n986);
nand (n971,n972,n976);
xor (n972,n973,n324);
or (n973,n974,n975);
and (n974,n59,n500);
and (n975,n63,n504);
xor (n976,n977,n42);
xnor (n977,n978,n627);
nor (n978,n979,n980);
and (n979,n39,n809);
and (n980,n35,n811);
nand (n981,n982,n976);
xor (n982,n983,n103);
or (n983,n984,n985);
and (n984,n221,n183);
and (n985,n293,n187);
nand (n986,n972,n982);
nand (n987,n988,n989,n990);
nand (n988,n909,n913);
nand (n989,n914,n913);
nand (n990,n909,n914);
xor (n991,n992,n998);
xor (n992,n993,n994);
and (n993,n977,n42);
xor (n994,n995,n74);
or (n995,n996,n997);
and (n996,n293,n101);
and (n997,n469,n105);
xor (n998,n999,n15);
or (n999,n1000,n1001);
and (n1000,n473,n72);
and (n1001,n475,n76);
nand (n1002,n1003,n1010,n1044);
nand (n1003,n1004,n1008);
nand (n1004,n1005,n1006,n1007);
nand (n1005,n947,n951);
nand (n1006,n955,n951);
nand (n1007,n947,n955);
xor (n1008,n1009,n982);
xor (n1009,n972,n976);
nand (n1010,n1011,n1008);
nand (n1011,n1012,n1029,n1043);
nand (n1012,n1013,n1027);
nand (n1013,n1014,n1023,n1026);
nand (n1014,n1015,n1019);
xor (n1015,n1016,n502);
or (n1016,n1017,n1018);
and (n1017,n59,n625);
and (n1018,n63,n629);
xor (n1019,n1020,n185);
or (n1020,n1021,n1022);
and (n1021,n221,n322);
and (n1022,n293,n326);
nand (n1023,n1024,n1019);
xnor (n1024,n1025,n31);
nand (n1025,n837,n25);
nand (n1026,n1015,n1024);
xor (n1027,n1028,n880);
xor (n1028,n871,n875);
nand (n1029,n1030,n1027);
nand (n1030,n1031,n1037,n1042);
nand (n1031,n1032,n1036);
xor (n1032,n1033,n324);
or (n1033,n1034,n1035);
and (n1034,n88,n500);
and (n1035,n175,n504);
xor (n1036,n897,n31);
nand (n1037,n1038,n1036);
xor (n1038,n1039,n103);
or (n1039,n1040,n1041);
and (n1040,n469,n183);
and (n1041,n473,n187);
nand (n1042,n1032,n1038);
nand (n1043,n1013,n1030);
nand (n1044,n1004,n1011);
nand (n1045,n786,n962);
xor (n1046,n1047,n1132);
xor (n1047,n1048,n1069);
xor (n1048,n1049,n1065);
xor (n1049,n1050,n1061);
xor (n1050,n1051,n1057);
xor (n1051,n1052,n1056);
xor (n1052,n1053,n31);
or (n1053,n1054,n1055);
and (n1054,n794,n25);
and (n1055,n798,n29);
and (n1056,n802,n806);
xor (n1057,n1058,n42);
or (n1058,n1059,n1060);
and (n1059,n800,n36);
and (n1060,n823,n40);
nand (n1061,n1062,n1063,n1064);
nand (n1062,n841,n845);
nand (n1063,n849,n845);
nand (n1064,n841,n849);
nand (n1065,n1066,n1067,n1068);
nand (n1066,n970,n987);
nand (n1067,n991,n987);
nand (n1068,n970,n991);
xor (n1069,n1070,n1128);
xor (n1070,n1071,n1095);
xor (n1071,n1072,n1091);
xor (n1072,n1073,n1077);
nand (n1073,n1074,n1075,n1076);
nand (n1074,n993,n994);
nand (n1075,n998,n994);
nand (n1076,n993,n998);
xor (n1077,n1078,n1087);
xor (n1078,n1079,n1083);
xnor (n1079,n1080,n627);
nor (n1080,n1081,n1082);
and (n1081,n28,n809);
and (n1082,n24,n811);
xor (n1083,n1084,n185);
or (n1084,n1085,n1086);
and (n1085,n59,n322);
and (n1086,n63,n326);
xor (n1087,n1088,n324);
or (n1088,n1089,n1090);
and (n1089,n48,n500);
and (n1090,n52,n504);
nand (n1091,n1092,n1093,n1094);
nand (n1092,n851,n855);
nand (n1093,n859,n855);
nand (n1094,n851,n859);
xor (n1095,n1096,n1114);
xor (n1096,n1097,n1101);
nand (n1097,n1098,n1099,n1100);
nand (n1098,n790,n795);
nand (n1099,n801,n795);
nand (n1100,n790,n801);
xor (n1101,n1102,n1112);
xor (n1102,n1103,n1107);
xor (n1103,n1104,n103);
or (n1104,n1105,n1106);
and (n1105,n88,n183);
and (n1106,n175,n187);
xor (n1107,n55,n1108);
xor (n1108,n1109,n502);
or (n1109,n1110,n1111);
and (n1110,n35,n625);
and (n1111,n39,n629);
xnor (n1112,n1113,n55);
nand (n1113,n837,n49);
xor (n1114,n1115,n1124);
xor (n1115,n1116,n1120);
xor (n1116,n1117,n74);
or (n1117,n1118,n1119);
and (n1118,n221,n101);
and (n1119,n293,n105);
xor (n1120,n1121,n15);
or (n1121,n1122,n1123);
and (n1122,n469,n72);
and (n1123,n473,n76);
xor (n1124,n1125,n20);
or (n1125,n1126,n1127);
and (n1126,n475,n13);
and (n1127,n609,n18);
nand (n1128,n1129,n1130,n1131);
nand (n1129,n788,n813);
nand (n1130,n839,n813);
nand (n1131,n788,n839);
nand (n1132,n1133,n1134,n1135);
nand (n1133,n964,n968);
nand (n1134,n1002,n968);
nand (n1135,n964,n1002);
nor (n1136,n1137,n1141);
nand (n1137,n1138,n1139,n1140);
nand (n1138,n1048,n1069);
nand (n1139,n1132,n1069);
nand (n1140,n1048,n1132);
xor (n1141,n1142,n1151);
xor (n1142,n1143,n1147);
nand (n1143,n1144,n1145,n1146);
nand (n1144,n1050,n1061);
nand (n1145,n1065,n1061);
nand (n1146,n1050,n1065);
nand (n1147,n1148,n1149,n1150);
nand (n1148,n1071,n1095);
nand (n1149,n1128,n1095);
nand (n1150,n1071,n1128);
xor (n1151,n1152,n1213);
xor (n1152,n1153,n1184);
xor (n1153,n1154,n1173);
xor (n1154,n1155,n1169);
xor (n1155,n1156,n1165);
xor (n1156,n1157,n1161);
xor (n1157,n1158,n185);
or (n1158,n1159,n1160);
and (n1159,n52,n322);
and (n1160,n59,n326);
xor (n1161,n1162,n324);
or (n1162,n1163,n1164);
and (n1163,n39,n500);
and (n1164,n48,n504);
xor (n1165,n1166,n103);
or (n1166,n1167,n1168);
and (n1167,n63,n183);
and (n1168,n88,n187);
nand (n1169,n1170,n1171,n1172);
nand (n1170,n1103,n1107);
nand (n1171,n1112,n1107);
nand (n1172,n1103,n1112);
xor (n1173,n1174,n1180);
xor (n1174,n1175,n1179);
xor (n1175,n1176,n74);
or (n1176,n1177,n1178);
and (n1177,n175,n101);
and (n1178,n221,n105);
and (n1179,n55,n1108);
xor (n1180,n1181,n15);
or (n1181,n1182,n1183);
and (n1182,n293,n72);
and (n1183,n469,n76);
xor (n1184,n1185,n1209);
xor (n1185,n1186,n1190);
nand (n1186,n1187,n1188,n1189);
nand (n1187,n1116,n1120);
nand (n1188,n1124,n1120);
nand (n1189,n1116,n1124);
xor (n1190,n1191,n1200);
xor (n1191,n1192,n1196);
xor (n1192,n1193,n20);
or (n1193,n1194,n1195);
and (n1194,n473,n13);
and (n1195,n475,n18);
xor (n1196,n1197,n31);
or (n1197,n1198,n1199);
and (n1198,n609,n25);
and (n1199,n794,n29);
xor (n1200,n1201,n1205);
xnor (n1201,n1202,n627);
nor (n1202,n1203,n1204);
and (n1203,n24,n809);
and (n1204,n17,n811);
xor (n1205,n1206,n502);
or (n1206,n1207,n1208);
and (n1207,n28,n625);
and (n1208,n35,n629);
nand (n1209,n1210,n1211,n1212);
nand (n1210,n1052,n1056);
nand (n1211,n1057,n1056);
nand (n1212,n1052,n1057);
xor (n1213,n1214,n1233);
xor (n1214,n1215,n1229);
xor (n1215,n1216,n1225);
xor (n1216,n1217,n1221);
xor (n1217,n1218,n42);
or (n1218,n1219,n1220);
and (n1219,n798,n36);
and (n1220,n800,n40);
xor (n1221,n1222,n55);
or (n1222,n1223,n1224);
and (n1223,n823,n49);
and (n1224,n837,n53);
nand (n1225,n1226,n1227,n1228);
nand (n1226,n1079,n1083);
nand (n1227,n1087,n1083);
nand (n1228,n1079,n1087);
nand (n1229,n1230,n1231,n1232);
nand (n1230,n1073,n1077);
nand (n1231,n1091,n1077);
nand (n1232,n1073,n1091);
nand (n1233,n1234,n1235,n1236);
nand (n1234,n1097,n1101);
nand (n1235,n1114,n1101);
nand (n1236,n1097,n1114);
nor (n1237,n1238,n1343);
nor (n1238,n1239,n1243);
nand (n1239,n1240,n1241,n1242);
nand (n1240,n1143,n1147);
nand (n1241,n1151,n1147);
nand (n1242,n1143,n1151);
xor (n1243,n1244,n1339);
xor (n1244,n1245,n1279);
xor (n1245,n1246,n1275);
xor (n1246,n1247,n1251);
nand (n1247,n1248,n1249,n1250);
nand (n1248,n1155,n1169);
nand (n1249,n1173,n1169);
nand (n1250,n1155,n1173);
xor (n1251,n1252,n1261);
xor (n1252,n1253,n1257);
xor (n1253,n1254,n55);
or (n1254,n1255,n1256);
and (n1255,n800,n49);
and (n1256,n823,n53);
nand (n1257,n1258,n1259,n1260);
nand (n1258,n1175,n1179);
nand (n1259,n1180,n1179);
nand (n1260,n1175,n1180);
xor (n1261,n1262,n1271);
xor (n1262,n1263,n1267);
xor (n1263,n1264,n185);
or (n1264,n1265,n1266);
and (n1265,n48,n322);
and (n1266,n52,n326);
xnor (n1267,n1268,n627);
nor (n1268,n1269,n1270);
and (n1269,n17,n809);
and (n1270,n12,n811);
xor (n1271,n1272,n324);
or (n1272,n1273,n1274);
and (n1273,n35,n500);
and (n1274,n39,n504);
nand (n1275,n1276,n1277,n1278);
nand (n1276,n1186,n1190);
nand (n1277,n1209,n1190);
nand (n1278,n1186,n1209);
xor (n1279,n1280,n1335);
xor (n1280,n1281,n1303);
xor (n1281,n1282,n1291);
xor (n1282,n1283,n1287);
nand (n1283,n1284,n1285,n1286);
nand (n1284,n1157,n1161);
nand (n1285,n1165,n1161);
nand (n1286,n1157,n1165);
nand (n1287,n1288,n1289,n1290);
nand (n1288,n1192,n1196);
nand (n1289,n1200,n1196);
nand (n1290,n1192,n1200);
xor (n1291,n1292,n1299);
xor (n1292,n1293,n1297);
xor (n1293,n1294,n103);
or (n1294,n1295,n1296);
and (n1295,n59,n183);
and (n1296,n63,n187);
xnor (n1297,n1298,n66);
nand (n1298,n837,n60);
xor (n1299,n1300,n74);
or (n1300,n1301,n1302);
and (n1301,n88,n101);
and (n1302,n175,n105);
xor (n1303,n1304,n1323);
xor (n1304,n1305,n1309);
nand (n1305,n1306,n1307,n1308);
nand (n1306,n1217,n1221);
nand (n1307,n1225,n1221);
nand (n1308,n1217,n1225);
xor (n1309,n1310,n1319);
xor (n1310,n1311,n1315);
xor (n1311,n1312,n15);
or (n1312,n1313,n1314);
and (n1313,n221,n72);
and (n1314,n293,n76);
xor (n1315,n1316,n20);
or (n1316,n1317,n1318);
and (n1317,n469,n13);
and (n1318,n473,n18);
xor (n1319,n1320,n31);
or (n1320,n1321,n1322);
and (n1321,n475,n25);
and (n1322,n609,n29);
xor (n1323,n1324,n1331);
xor (n1324,n1325,n1330);
xor (n1325,n66,n1326);
xor (n1326,n1327,n502);
or (n1327,n1328,n1329);
and (n1328,n24,n625);
and (n1329,n28,n629);
and (n1330,n1201,n1205);
xor (n1331,n1332,n42);
or (n1332,n1333,n1334);
and (n1333,n794,n36);
and (n1334,n798,n40);
nand (n1335,n1336,n1337,n1338);
nand (n1336,n1215,n1229);
nand (n1337,n1233,n1229);
nand (n1338,n1215,n1233);
nand (n1339,n1340,n1341,n1342);
nand (n1340,n1153,n1184);
nand (n1341,n1213,n1184);
nand (n1342,n1153,n1213);
nor (n1343,n1344,n1348);
nand (n1344,n1345,n1346,n1347);
nand (n1345,n1245,n1279);
nand (n1346,n1339,n1279);
nand (n1347,n1245,n1339);
xor (n1348,n1349,n1358);
xor (n1349,n1350,n1354);
nand (n1350,n1351,n1352,n1353);
nand (n1351,n1247,n1251);
nand (n1352,n1275,n1251);
nand (n1353,n1247,n1275);
nand (n1354,n1355,n1356,n1357);
nand (n1355,n1281,n1303);
nand (n1356,n1335,n1303);
nand (n1357,n1281,n1335);
xor (n1358,n1359,n1420);
xor (n1359,n1360,n1384);
xor (n1360,n1361,n1380);
xor (n1361,n1362,n1366);
nand (n1362,n1363,n1364,n1365);
nand (n1363,n1311,n1315);
nand (n1364,n1319,n1315);
nand (n1365,n1311,n1319);
xor (n1366,n1367,n1376);
xor (n1367,n1368,n1372);
xor (n1368,n1369,n74);
or (n1369,n1370,n1371);
and (n1370,n63,n101);
and (n1371,n88,n105);
xor (n1372,n1373,n15);
or (n1373,n1374,n1375);
and (n1374,n175,n72);
and (n1375,n221,n76);
xor (n1376,n1377,n20);
or (n1377,n1378,n1379);
and (n1378,n293,n13);
and (n1379,n469,n18);
nand (n1380,n1381,n1382,n1383);
nand (n1381,n1325,n1330);
nand (n1382,n1331,n1330);
nand (n1383,n1325,n1331);
xor (n1384,n1385,n1406);
xor (n1385,n1386,n1402);
xor (n1386,n1387,n1401);
xor (n1387,n1388,n1392);
xor (n1388,n1389,n31);
or (n1389,n1390,n1391);
and (n1390,n473,n25);
and (n1391,n475,n29);
xor (n1392,n1393,n1397);
xnor (n1393,n1394,n627);
nor (n1394,n1395,n1396);
and (n1395,n12,n809);
and (n1396,n71,n811);
xor (n1397,n1398,n502);
or (n1398,n1399,n1400);
and (n1399,n17,n625);
and (n1400,n24,n629);
and (n1401,n66,n1326);
nand (n1402,n1403,n1404,n1405);
nand (n1403,n1253,n1257);
nand (n1404,n1261,n1257);
nand (n1405,n1253,n1261);
xor (n1406,n1407,n1416);
xor (n1407,n1408,n1412);
xor (n1408,n1409,n42);
or (n1409,n1410,n1411);
and (n1410,n609,n36);
and (n1411,n794,n40);
xor (n1412,n1413,n66);
or (n1413,n1414,n1415);
and (n1414,n823,n60);
and (n1415,n837,n64);
xor (n1416,n1417,n55);
or (n1417,n1418,n1419);
and (n1418,n798,n49);
and (n1419,n800,n53);
xor (n1420,n1421,n1450);
xor (n1421,n1422,n1446);
xor (n1422,n1423,n1442);
xor (n1423,n1424,n1428);
nand (n1424,n1425,n1426,n1427);
nand (n1425,n1263,n1267);
nand (n1426,n1271,n1267);
nand (n1427,n1263,n1271);
xor (n1428,n1429,n1438);
xor (n1429,n1430,n1434);
xor (n1430,n1431,n185);
or (n1431,n1432,n1433);
and (n1432,n39,n322);
and (n1433,n48,n326);
xor (n1434,n1435,n324);
or (n1435,n1436,n1437);
and (n1436,n28,n500);
and (n1437,n35,n504);
xor (n1438,n1439,n103);
or (n1439,n1440,n1441);
and (n1440,n52,n183);
and (n1441,n59,n187);
nand (n1442,n1443,n1444,n1445);
nand (n1443,n1293,n1297);
nand (n1444,n1299,n1297);
nand (n1445,n1293,n1299);
nand (n1446,n1447,n1448,n1449);
nand (n1447,n1283,n1287);
nand (n1448,n1291,n1287);
nand (n1449,n1283,n1291);
nand (n1450,n1451,n1452,n1453);
nand (n1451,n1305,n1309);
nand (n1452,n1323,n1309);
nand (n1453,n1305,n1323);
nor (n1454,n1455,n1727);
nor (n1455,n1456,n1703);
nor (n1456,n1457,n1701);
nor (n1457,n1458,n1676);
nand (n1458,n1459,n1638);
nand (n1459,n1460,n1585,n1637);
nand (n1460,n1461,n1512);
xor (n1461,n1462,n1499);
xor (n1462,n1463,n1484);
nand (n1463,n1464,n1478,n1483);
nand (n1464,n1465,n1474);
and (n1465,n1466,n1470);
xnor (n1466,n1467,n627);
nor (n1467,n1468,n1469);
and (n1468,n88,n809);
and (n1469,n63,n811);
xor (n1470,n1471,n502);
or (n1471,n1472,n1473);
and (n1472,n175,n625);
and (n1473,n221,n629);
xor (n1474,n1475,n74);
or (n1475,n1476,n1477);
and (n1476,n794,n101);
and (n1477,n798,n105);
nand (n1478,n1479,n1474);
xor (n1479,n1480,n15);
or (n1480,n1481,n1482);
and (n1481,n800,n72);
and (n1482,n823,n76);
nand (n1483,n1465,n1479);
xor (n1484,n1485,n1494);
xor (n1485,n1486,n1490);
xor (n1486,n1487,n185);
or (n1487,n1488,n1489);
and (n1488,n293,n322);
and (n1489,n469,n326);
xor (n1490,n1491,n324);
or (n1491,n1492,n1493);
and (n1492,n175,n500);
and (n1493,n221,n504);
and (n1494,n1495,n20);
xnor (n1495,n1496,n627);
nor (n1496,n1497,n1498);
and (n1497,n63,n809);
and (n1498,n59,n811);
nand (n1499,n1500,n1506,n1511);
nand (n1500,n1501,n1505);
xor (n1501,n1502,n324);
or (n1502,n1503,n1504);
and (n1503,n221,n500);
and (n1504,n293,n504);
xor (n1505,n1495,n20);
nand (n1506,n1507,n1505);
xor (n1507,n1508,n103);
or (n1508,n1509,n1510);
and (n1509,n475,n183);
and (n1510,n609,n187);
nand (n1511,n1501,n1507);
xor (n1512,n1513,n1549);
xor (n1513,n1514,n1525);
xor (n1514,n1515,n1521);
xor (n1515,n1516,n1520);
xor (n1516,n1517,n103);
or (n1517,n1518,n1519);
and (n1518,n473,n183);
and (n1519,n475,n187);
xor (n1520,n924,n928);
xor (n1521,n1522,n74);
or (n1522,n1523,n1524);
and (n1523,n609,n101);
and (n1524,n794,n105);
xor (n1525,n1526,n1535);
xor (n1526,n1527,n1531);
xor (n1527,n1528,n15);
or (n1528,n1529,n1530);
and (n1529,n798,n72);
and (n1530,n800,n76);
xor (n1531,n1532,n20);
or (n1532,n1533,n1534);
and (n1533,n823,n13);
and (n1534,n837,n18);
nand (n1535,n1536,n1543,n1548);
nand (n1536,n1537,n1541);
xor (n1537,n1538,n502);
or (n1538,n1539,n1540);
and (n1539,n88,n625);
and (n1540,n175,n629);
xnor (n1541,n1542,n20);
nand (n1542,n837,n13);
nand (n1543,n1544,n1541);
xor (n1544,n1545,n185);
or (n1545,n1546,n1547);
and (n1546,n469,n322);
and (n1547,n473,n326);
nand (n1548,n1537,n1544);
nand (n1549,n1550,n1570,n1584);
nand (n1550,n1551,n1553);
xor (n1551,n1552,n1544);
xor (n1552,n1537,n1541);
nand (n1553,n1554,n1563,n1569);
nand (n1554,n1555,n1559);
xor (n1555,n1556,n185);
or (n1556,n1557,n1558);
and (n1557,n473,n322);
and (n1558,n475,n326);
xor (n1559,n1560,n324);
or (n1560,n1561,n1562);
and (n1561,n293,n500);
and (n1562,n469,n504);
nand (n1563,n1564,n1559);
and (n1564,n1565,n15);
xnor (n1565,n1566,n627);
nor (n1566,n1567,n1568);
and (n1567,n175,n809);
and (n1568,n88,n811);
nand (n1569,n1555,n1564);
nand (n1570,n1571,n1553);
nand (n1571,n1572,n1578,n1583);
nand (n1572,n1573,n1577);
xor (n1573,n1574,n103);
or (n1574,n1575,n1576);
and (n1575,n609,n183);
and (n1576,n794,n187);
xor (n1577,n1466,n1470);
nand (n1578,n1579,n1577);
xor (n1579,n1580,n74);
or (n1580,n1581,n1582);
and (n1581,n798,n101);
and (n1582,n800,n105);
nand (n1583,n1573,n1579);
nand (n1584,n1551,n1571);
nand (n1585,n1586,n1512);
nand (n1586,n1587,n1592,n1636);
nand (n1587,n1588,n1590);
xor (n1588,n1589,n1479);
xor (n1589,n1465,n1474);
xor (n1590,n1591,n1507);
xor (n1591,n1501,n1505);
nand (n1592,n1593,n1590);
nand (n1593,n1594,n1613,n1635);
nand (n1594,n1595,n1599);
xor (n1595,n1596,n15);
or (n1596,n1597,n1598);
and (n1597,n823,n72);
and (n1598,n837,n76);
nand (n1599,n1600,n1607,n1612);
nand (n1600,n1601,n1605);
xor (n1601,n1602,n502);
or (n1602,n1603,n1604);
and (n1603,n221,n625);
and (n1604,n293,n629);
xnor (n1605,n1606,n15);
nand (n1606,n837,n72);
nand (n1607,n1608,n1605);
xor (n1608,n1609,n185);
or (n1609,n1610,n1611);
and (n1610,n475,n322);
and (n1611,n609,n326);
nand (n1612,n1601,n1608);
nand (n1613,n1614,n1599);
nand (n1614,n1615,n1629,n1634);
nand (n1615,n1616,n1620);
xor (n1616,n1617,n324);
or (n1617,n1618,n1619);
and (n1618,n469,n500);
and (n1619,n473,n504);
and (n1620,n1621,n1625);
xnor (n1621,n1622,n627);
nor (n1622,n1623,n1624);
and (n1623,n221,n809);
and (n1624,n175,n811);
xor (n1625,n1626,n502);
or (n1626,n1627,n1628);
and (n1627,n293,n625);
and (n1628,n469,n629);
nand (n1629,n1630,n1620);
xor (n1630,n1631,n103);
or (n1631,n1632,n1633);
and (n1632,n794,n183);
and (n1633,n798,n187);
nand (n1634,n1616,n1630);
nand (n1635,n1595,n1614);
nand (n1636,n1588,n1593);
nand (n1637,n1461,n1586);
xor (n1638,n1639,n1654);
xor (n1639,n1640,n1650);
xor (n1640,n1641,n1648);
xor (n1641,n1642,n1646);
nand (n1642,n1643,n1644,n1645);
nand (n1643,n1486,n1490);
nand (n1644,n1494,n1490);
nand (n1645,n1486,n1494);
xor (n1646,n1647,n937);
xor (n1647,n923,n932);
xor (n1648,n1649,n1038);
xor (n1649,n1032,n1036);
nand (n1650,n1651,n1652,n1653);
nand (n1651,n1514,n1525);
nand (n1652,n1549,n1525);
nand (n1653,n1514,n1549);
xor (n1654,n1655,n1664);
xor (n1655,n1656,n1660);
nand (n1656,n1657,n1658,n1659);
nand (n1657,n1527,n1531);
nand (n1658,n1535,n1531);
nand (n1659,n1527,n1535);
nand (n1660,n1661,n1662,n1663);
nand (n1661,n1463,n1484);
nand (n1662,n1499,n1484);
nand (n1663,n1463,n1499);
xor (n1664,n1665,n1674);
xor (n1665,n1666,n1670);
xor (n1666,n1667,n20);
or (n1667,n1668,n1669);
and (n1668,n800,n13);
and (n1669,n823,n18);
nand (n1670,n1671,n1672,n1673);
nand (n1671,n1516,n1520);
nand (n1672,n1521,n1520);
nand (n1673,n1516,n1521);
xor (n1674,n1675,n1024);
xor (n1675,n1015,n1019);
nor (n1676,n1677,n1681);
nand (n1677,n1678,n1679,n1680);
nand (n1678,n1640,n1650);
nand (n1679,n1654,n1650);
nand (n1680,n1640,n1654);
xor (n1681,n1682,n1689);
xor (n1682,n1683,n1685);
xor (n1683,n1684,n945);
xor (n1684,n921,n942);
nand (n1685,n1686,n1687,n1688);
nand (n1686,n1656,n1660);
nand (n1687,n1664,n1660);
nand (n1688,n1656,n1664);
xor (n1689,n1690,n1699);
xor (n1690,n1691,n1695);
nand (n1691,n1692,n1693,n1694);
nand (n1692,n1666,n1670);
nand (n1693,n1674,n1670);
nand (n1694,n1666,n1674);
nand (n1695,n1696,n1697,n1698);
nand (n1696,n1642,n1646);
nand (n1697,n1648,n1646);
nand (n1698,n1642,n1648);
xor (n1699,n1700,n1030);
xor (n1700,n1013,n1027);
not (n1701,n1702);
nand (n1702,n1677,n1681);
not (n1703,n1704);
nor (n1704,n1705,n1720);
nor (n1705,n1706,n1710);
nand (n1706,n1707,n1708,n1709);
nand (n1707,n1683,n1685);
nand (n1708,n1689,n1685);
nand (n1709,n1683,n1689);
xor (n1710,n1711,n1718);
xor (n1711,n1712,n1714);
xor (n1712,n1713,n1011);
xor (n1713,n1004,n1008);
nand (n1714,n1715,n1716,n1717);
nand (n1715,n1691,n1695);
nand (n1716,n1699,n1695);
nand (n1717,n1691,n1699);
xor (n1718,n1719,n919);
xor (n1719,n865,n867);
nor (n1720,n1721,n1725);
nand (n1721,n1722,n1723,n1724);
nand (n1722,n1712,n1714);
nand (n1723,n1718,n1714);
nand (n1724,n1712,n1718);
xor (n1725,n1726,n962);
xor (n1726,n786,n863);
not (n1727,n1728);
nor (n1728,n1729,n1731);
nor (n1729,n1730,n1720);
nand (n1730,n1706,n1710);
not (n1731,n1732);
nand (n1732,n1721,n1725);
not (n1733,n1734);
nor (n1734,n1735,n1742);
nor (n1735,n1736,n1741);
nor (n1736,n1737,n1739);
nor (n1737,n1738,n1136);
nand (n1738,n784,n1046);
not (n1739,n1740);
nand (n1740,n1137,n1141);
not (n1741,n1237);
not (n1742,n1743);
nor (n1743,n1744,n1746);
nor (n1744,n1745,n1343);
nand (n1745,n1239,n1243);
not (n1746,n1747);
nand (n1747,n1344,n1348);
not (n1748,n1749);
nor (n1749,n1750,n2165);
nand (n1750,n1751,n1978);
nor (n1751,n1752,n1864);
nor (n1752,n1753,n1757);
nand (n1753,n1754,n1755,n1756);
nand (n1754,n1350,n1354);
nand (n1755,n1358,n1354);
nand (n1756,n1350,n1358);
xor (n1757,n1758,n1860);
xor (n1758,n1759,n1792);
xor (n1759,n1760,n1788);
xor (n1760,n1761,n1784);
xor (n1761,n1762,n1780);
xor (n1762,n1763,n1776);
xor (n1763,n1764,n1773);
xor (n1764,n1765,n1769);
xor (n1765,n1766,n502);
or (n1766,n1767,n1768);
and (n1767,n12,n625);
and (n1768,n17,n629);
xor (n1769,n1770,n324);
or (n1770,n1771,n1772);
and (n1771,n24,n500);
and (n1772,n28,n504);
xnor (n1773,n1774,n627);
nor (n1774,n1775,n1396);
and (n1775,n71,n809);
nand (n1776,n1777,n1778,n1779);
nand (n1777,n1368,n1372);
nand (n1778,n1376,n1372);
nand (n1779,n1368,n1376);
nand (n1780,n1781,n1782,n1783);
nand (n1781,n1388,n1392);
nand (n1782,n1401,n1392);
nand (n1783,n1388,n1401);
nand (n1784,n1785,n1786,n1787);
nand (n1785,n1362,n1366);
nand (n1786,n1380,n1366);
nand (n1787,n1362,n1380);
nand (n1788,n1789,n1790,n1791);
nand (n1789,n1386,n1402);
nand (n1790,n1406,n1402);
nand (n1791,n1386,n1406);
xor (n1792,n1793,n1856);
xor (n1793,n1794,n1832);
xor (n1794,n1795,n1817);
xor (n1795,n1796,n1810);
xor (n1796,n1797,n1806);
xor (n1797,n1798,n1802);
xor (n1798,n1799,n103);
or (n1799,n1800,n1801);
and (n1800,n48,n183);
and (n1801,n52,n187);
xor (n1802,n1803,n74);
or (n1803,n1804,n1805);
and (n1804,n59,n101);
and (n1805,n63,n105);
xor (n1806,n1807,n15);
or (n1807,n1808,n1809);
and (n1808,n88,n72);
and (n1809,n175,n76);
xor (n1810,n1811,n1813);
xor (n1811,n66,n1812);
and (n1812,n1393,n1397);
xor (n1813,n1814,n42);
or (n1814,n1815,n1816);
and (n1815,n475,n36);
and (n1816,n609,n40);
xor (n1817,n1818,n1827);
xor (n1818,n1819,n1823);
xor (n1819,n1820,n20);
or (n1820,n1821,n1822);
and (n1821,n221,n13);
and (n1822,n293,n18);
xor (n1823,n1824,n31);
or (n1824,n1825,n1826);
and (n1825,n469,n25);
and (n1826,n473,n29);
xor (n1827,n66,n1828);
xor (n1828,n1829,n185);
or (n1829,n1830,n1831);
and (n1830,n35,n322);
and (n1831,n39,n326);
xor (n1832,n1833,n1842);
xor (n1833,n1834,n1838);
nand (n1834,n1835,n1836,n1837);
nand (n1835,n1408,n1412);
nand (n1836,n1416,n1412);
nand (n1837,n1408,n1416);
nand (n1838,n1839,n1840,n1841);
nand (n1839,n1424,n1428);
nand (n1840,n1442,n1428);
nand (n1841,n1424,n1442);
xor (n1842,n1843,n1852);
xor (n1843,n1844,n1848);
xor (n1844,n1845,n55);
or (n1845,n1846,n1847);
and (n1846,n794,n49);
and (n1847,n798,n53);
xor (n1848,n1849,n66);
or (n1849,n1850,n1851);
and (n1850,n800,n60);
and (n1851,n823,n64);
nand (n1852,n1853,n1854,n1855);
nand (n1853,n1430,n1434);
nand (n1854,n1438,n1434);
nand (n1855,n1430,n1438);
nand (n1856,n1857,n1858,n1859);
nand (n1857,n1422,n1446);
nand (n1858,n1450,n1446);
nand (n1859,n1422,n1450);
nand (n1860,n1861,n1862,n1863);
nand (n1861,n1360,n1384);
nand (n1862,n1420,n1384);
nand (n1863,n1360,n1420);
nor (n1864,n1865,n1869);
nand (n1865,n1866,n1867,n1868);
nand (n1866,n1759,n1792);
nand (n1867,n1860,n1792);
nand (n1868,n1759,n1860);
xor (n1869,n1870,n1879);
xor (n1870,n1871,n1875);
nand (n1871,n1872,n1873,n1874);
nand (n1872,n1761,n1784);
nand (n1873,n1788,n1784);
nand (n1874,n1761,n1788);
nand (n1875,n1876,n1877,n1878);
nand (n1876,n1794,n1832);
nand (n1877,n1856,n1832);
nand (n1878,n1794,n1856);
xor (n1879,n1880,n1937);
xor (n1880,n1881,n1912);
xor (n1881,n1882,n1898);
xor (n1882,n1883,n1887);
nand (n1883,n1884,n1885,n1886);
nand (n1884,n66,n1812);
nand (n1885,n1813,n1812);
nand (n1886,n66,n1813);
xor (n1887,n1888,n1894);
xor (n1888,n1889,n1893);
xor (n1889,n1890,n31);
or (n1890,n1891,n1892);
and (n1891,n293,n25);
and (n1892,n469,n29);
and (n1893,n66,n1828);
xor (n1894,n1895,n42);
or (n1895,n1896,n1897);
and (n1896,n473,n36);
and (n1897,n475,n40);
xor (n1898,n1899,n1908);
xor (n1899,n1900,n1904);
xor (n1900,n1901,n55);
or (n1901,n1902,n1903);
and (n1902,n609,n49);
and (n1903,n794,n53);
xor (n1904,n1905,n66);
or (n1905,n1906,n1907);
and (n1906,n798,n60);
and (n1907,n800,n64);
nand (n1908,n1909,n1910,n1911);
nand (n1909,n1765,n1769);
nand (n1910,n1773,n1769);
nand (n1911,n1765,n1773);
xor (n1912,n1913,n1922);
xor (n1913,n1914,n1918);
nand (n1914,n1915,n1916,n1917);
nand (n1915,n1844,n1848);
nand (n1916,n1852,n1848);
nand (n1917,n1844,n1852);
nand (n1918,n1919,n1920,n1921);
nand (n1919,n1763,n1776);
nand (n1920,n1780,n1776);
nand (n1921,n1763,n1780);
xor (n1922,n1923,n66);
xor (n1923,n1924,n1928);
nand (n1924,n1925,n1926,n1927);
nand (n1925,n1798,n1802);
nand (n1926,n1806,n1802);
nand (n1927,n1798,n1806);
xor (n1928,n1929,n1934);
not (n1929,n1930);
xor (n1930,n1931,n185);
or (n1931,n1932,n1933);
and (n1932,n28,n322);
and (n1933,n35,n326);
xor (n1934,n1935,n502);
or (n1935,n624,n1936);
and (n1936,n12,n629);
xor (n1937,n1938,n1974);
xor (n1938,n1939,n1943);
nand (n1939,n1940,n1941,n1942);
nand (n1940,n1796,n1810);
nand (n1941,n1817,n1810);
nand (n1942,n1796,n1817);
xor (n1943,n1944,n1963);
xor (n1944,n1945,n1949);
nand (n1945,n1946,n1947,n1948);
nand (n1946,n1819,n1823);
nand (n1947,n1827,n1823);
nand (n1948,n1819,n1827);
xor (n1949,n1950,n1959);
xor (n1950,n1951,n1955);
xor (n1951,n1952,n74);
or (n1952,n1953,n1954);
and (n1953,n52,n101);
and (n1954,n59,n105);
xor (n1955,n1956,n15);
or (n1956,n1957,n1958);
and (n1957,n63,n72);
and (n1958,n88,n76);
xor (n1959,n1960,n20);
or (n1960,n1961,n1962);
and (n1961,n175,n13);
and (n1962,n221,n18);
xor (n1963,n1964,n1970);
xor (n1964,n1965,n1969);
xor (n1965,n1966,n324);
or (n1966,n1967,n1968);
and (n1967,n17,n500);
and (n1968,n24,n504);
not (n1969,n1773);
xor (n1970,n1971,n103);
or (n1971,n1972,n1973);
and (n1972,n39,n183);
and (n1973,n48,n187);
nand (n1974,n1975,n1976,n1977);
nand (n1975,n1834,n1838);
nand (n1976,n1842,n1838);
nand (n1977,n1834,n1842);
nor (n1978,n1979,n2086);
nor (n1979,n1980,n1984);
nand (n1980,n1981,n1982,n1983);
nand (n1981,n1871,n1875);
nand (n1982,n1879,n1875);
nand (n1983,n1871,n1879);
xor (n1984,n1985,n2082);
xor (n1985,n1986,n2026);
xor (n1986,n1987,n2022);
xor (n1987,n1988,n2018);
xor (n1988,n1989,n2014);
xor (n1989,n1990,n2004);
xor (n1990,n1991,n2000);
xor (n1991,n1992,n1996);
xor (n1992,n1993,n74);
or (n1993,n1994,n1995);
and (n1994,n48,n101);
and (n1995,n52,n105);
xor (n1996,n1997,n15);
or (n1997,n1998,n1999);
and (n1998,n59,n72);
and (n1999,n63,n76);
xor (n2000,n2001,n31);
or (n2001,n2002,n2003);
and (n2002,n221,n25);
and (n2003,n293,n29);
xor (n2004,n2005,n2010);
xor (n2005,n2006,n622);
xor (n2006,n2007,n185);
or (n2007,n2008,n2009);
and (n2008,n24,n322);
and (n2009,n28,n326);
xor (n2010,n2011,n103);
or (n2011,n2012,n2013);
and (n2012,n35,n183);
and (n2013,n39,n187);
nand (n2014,n2015,n2016,n2017);
nand (n2015,n1889,n1893);
nand (n2016,n1894,n1893);
nand (n2017,n1889,n1894);
nand (n2018,n2019,n2020,n2021);
nand (n2019,n1883,n1887);
nand (n2020,n1898,n1887);
nand (n2021,n1883,n1898);
nand (n2022,n2023,n2024,n2025);
nand (n2023,n1914,n1918);
nand (n2024,n1922,n1918);
nand (n2025,n1914,n1922);
xor (n2026,n2027,n2078);
xor (n2027,n2028,n2049);
xor (n2028,n2029,n2045);
xor (n2029,n2030,n2041);
xor (n2030,n2031,n2037);
xor (n2031,n2032,n2033);
not (n2032,n663);
xor (n2033,n2034,n20);
or (n2034,n2035,n2036);
and (n2035,n88,n13);
and (n2036,n175,n18);
xor (n2037,n2038,n42);
or (n2038,n2039,n2040);
and (n2039,n469,n36);
and (n2040,n473,n40);
nand (n2041,n2042,n2043,n2044);
nand (n2042,n1900,n1904);
nand (n2043,n1908,n1904);
nand (n2044,n1900,n1908);
nand (n2045,n2046,n2047,n2048);
nand (n2046,n1924,n1928);
nand (n2047,n66,n1928);
nand (n2048,n1924,n66);
xor (n2049,n2050,n2074);
xor (n2050,n2051,n2064);
xor (n2051,n2052,n2061);
xor (n2052,n2053,n2057);
xor (n2053,n2054,n55);
or (n2054,n2055,n2056);
and (n2055,n475,n49);
and (n2056,n609,n53);
xor (n2057,n2058,n66);
or (n2058,n2059,n2060);
and (n2059,n794,n60);
and (n2060,n798,n64);
nand (n2061,n1929,n2062,n2063);
nand (n2062,n1934,n1930);
not (n2063,n1934);
xor (n2064,n2065,n2070);
xor (n2065,n66,n2066);
nand (n2066,n2067,n2068,n2069);
nand (n2067,n1965,n1969);
nand (n2068,n1970,n1969);
nand (n2069,n1965,n1970);
nand (n2070,n2071,n2072,n2073);
nand (n2071,n1951,n1955);
nand (n2072,n1959,n1955);
nand (n2073,n1951,n1959);
nand (n2074,n2075,n2076,n2077);
nand (n2075,n1945,n1949);
nand (n2076,n1963,n1949);
nand (n2077,n1945,n1963);
nand (n2078,n2079,n2080,n2081);
nand (n2079,n1939,n1943);
nand (n2080,n1974,n1943);
nand (n2081,n1939,n1974);
nand (n2082,n2083,n2084,n2085);
nand (n2083,n1881,n1912);
nand (n2084,n1937,n1912);
nand (n2085,n1881,n1937);
nor (n2086,n2087,n2091);
nand (n2087,n2088,n2089,n2090);
nand (n2088,n1986,n2026);
nand (n2089,n2082,n2026);
nand (n2090,n1986,n2082);
xor (n2091,n2092,n2101);
xor (n2092,n2093,n2097);
nand (n2093,n2094,n2095,n2096);
nand (n2094,n1988,n2018);
nand (n2095,n2022,n2018);
nand (n2096,n1988,n2022);
nand (n2097,n2098,n2099,n2100);
nand (n2098,n2028,n2049);
nand (n2099,n2078,n2049);
nand (n2100,n2028,n2078);
xor (n2101,n2102,n2133);
xor (n2102,n2103,n2107);
nand (n2103,n2104,n2105,n2106);
nand (n2104,n2051,n2064);
nand (n2105,n2074,n2064);
nand (n2106,n2051,n2074);
xor (n2107,n2108,n2121);
xor (n2108,n2109,n2113);
nand (n2109,n2110,n2111,n2112);
nand (n2110,n66,n2066);
nand (n2111,n2070,n2066);
nand (n2112,n66,n2070);
xor (n2113,n2114,n2117);
xor (n2114,n2115,n66);
xor (n2115,n2116,n621);
xor (n2116,n613,n616);
nand (n2117,n2118,n2119,n2120);
nand (n2118,n2006,n622);
nand (n2119,n2010,n622);
nand (n2120,n2006,n2010);
xor (n2121,n2122,n2129);
xor (n2122,n2123,n2125);
xor (n2123,n2124,n649);
xor (n2124,n640,n644);
nand (n2125,n2126,n2127,n2128);
nand (n2126,n1992,n1996);
nand (n2127,n2000,n1996);
nand (n2128,n1992,n2000);
nand (n2129,n2130,n2131,n2132);
nand (n2130,n2053,n2057);
nand (n2131,n2061,n2057);
nand (n2132,n2053,n2061);
xor (n2133,n2134,n2143);
xor (n2134,n2135,n2139);
nand (n2135,n2136,n2137,n2138);
nand (n2136,n1990,n2004);
nand (n2137,n2014,n2004);
nand (n2138,n1990,n2014);
nand (n2139,n2140,n2141,n2142);
nand (n2140,n2030,n2041);
nand (n2141,n2045,n2041);
nand (n2142,n2030,n2045);
xor (n2143,n2144,n2151);
xor (n2144,n2145,n2149);
nand (n2145,n2146,n2147,n2148);
nand (n2146,n2032,n2033);
nand (n2147,n2037,n2033);
nand (n2148,n2032,n2037);
xor (n2149,n2150,n668);
xor (n2150,n659,n663);
xor (n2151,n2152,n2161);
xor (n2152,n2153,n2157);
xor (n2153,n2154,n42);
or (n2154,n2155,n2156);
and (n2155,n293,n36);
and (n2156,n469,n40);
xor (n2157,n2158,n55);
or (n2158,n2159,n2160);
and (n2159,n473,n49);
and (n2160,n475,n53);
xor (n2161,n2162,n66);
or (n2162,n2163,n2164);
and (n2163,n609,n60);
and (n2164,n794,n64);
nand (n2165,n2166,n2250);
nor (n2166,n2167,n2217);
nor (n2167,n2168,n2172);
nand (n2168,n2169,n2170,n2171);
nand (n2169,n2093,n2097);
nand (n2170,n2101,n2097);
nand (n2171,n2093,n2101);
xor (n2172,n2173,n2213);
xor (n2173,n2174,n2194);
xor (n2174,n2175,n2182);
xor (n2175,n2176,n2178);
xor (n2176,n2177,n657);
xor (n2177,n638,n654);
nand (n2178,n2179,n2180,n2181);
nand (n2179,n2145,n2149);
nand (n2180,n2151,n2149);
nand (n2181,n2145,n2151);
xor (n2182,n2183,n2190);
xor (n2183,n2184,n2188);
nand (n2184,n2185,n2186,n2187);
nand (n2185,n2153,n2157);
nand (n2186,n2161,n2157);
nand (n2187,n2153,n2161);
xor (n2188,n2189,n567);
xor (n2189,n561,n565);
nand (n2190,n2191,n2192,n2193);
nand (n2191,n2115,n66);
nand (n2192,n2117,n66);
nand (n2193,n2115,n2117);
xor (n2194,n2195,n2209);
xor (n2195,n2196,n2200);
nand (n2196,n2197,n2198,n2199);
nand (n2197,n2109,n2113);
nand (n2198,n2121,n2113);
nand (n2199,n2109,n2121);
xor (n2200,n2201,n2205);
xor (n2201,n2202,n2204);
xor (n2202,n2203,n583);
xor (n2203,n574,n578);
xor (n2204,n606,n611);
nand (n2205,n2206,n2207,n2208);
nand (n2206,n2123,n2125);
nand (n2207,n2129,n2125);
nand (n2208,n2123,n2129);
nand (n2209,n2210,n2211,n2212);
nand (n2210,n2135,n2139);
nand (n2211,n2143,n2139);
nand (n2212,n2135,n2143);
nand (n2213,n2214,n2215,n2216);
nand (n2214,n2103,n2107);
nand (n2215,n2133,n2107);
nand (n2216,n2103,n2133);
nor (n2217,n2218,n2222);
nand (n2218,n2219,n2220,n2221);
nand (n2219,n2174,n2194);
nand (n2220,n2213,n2194);
nand (n2221,n2174,n2213);
xor (n2222,n2223,n2246);
xor (n2223,n2224,n2234);
xor (n2224,n2225,n2232);
xor (n2225,n2226,n2228);
xor (n2226,n2227,n554);
xor (n2227,n539,n551);
nand (n2228,n2229,n2230,n2231);
nand (n2229,n2184,n2188);
nand (n2230,n2190,n2188);
nand (n2231,n2184,n2190);
xor (n2232,n2233,n589);
xor (n2233,n559,n572);
xor (n2234,n2235,n2242);
xor (n2235,n2236,n2238);
xor (n2236,n2237,n636);
xor (n2237,n603,n633);
nand (n2238,n2239,n2240,n2241);
nand (n2239,n2202,n2204);
nand (n2240,n2205,n2204);
nand (n2241,n2202,n2205);
nand (n2242,n2243,n2244,n2245);
nand (n2243,n2176,n2178);
nand (n2244,n2182,n2178);
nand (n2245,n2176,n2182);
nand (n2246,n2247,n2248,n2249);
nand (n2247,n2196,n2200);
nand (n2248,n2209,n2200);
nand (n2249,n2196,n2209);
nor (n2250,n2251,n2268);
nor (n2251,n2252,n2256);
nand (n2252,n2253,n2254,n2255);
nand (n2253,n2224,n2234);
nand (n2254,n2246,n2234);
nand (n2255,n2224,n2246);
xor (n2256,n2257,n2264);
xor (n2257,n2258,n2262);
nand (n2258,n2259,n2260,n2261);
nand (n2259,n2226,n2228);
nand (n2260,n2232,n2228);
nand (n2261,n2226,n2232);
xor (n2262,n2263,n676);
xor (n2263,n599,n601);
nand (n2264,n2265,n2266,n2267);
nand (n2265,n2236,n2238);
nand (n2266,n2242,n2238);
nand (n2267,n2236,n2242);
nor (n2268,n2269,n2273);
nand (n2269,n2270,n2271,n2272);
nand (n2270,n2258,n2262);
nand (n2271,n2264,n2262);
nand (n2272,n2258,n2264);
xor (n2273,n2274,n597);
xor (n2274,n375,n459);
not (n2275,n2276);
nor (n2276,n2277,n2292);
nor (n2277,n2165,n2278);
nor (n2278,n2279,n2286);
nor (n2279,n2280,n2285);
nor (n2280,n2281,n2283);
nor (n2281,n2282,n1864);
nand (n2282,n1753,n1757);
not (n2283,n2284);
nand (n2284,n1865,n1869);
not (n2285,n1978);
not (n2286,n2287);
nor (n2287,n2288,n2290);
nor (n2288,n2289,n2086);
nand (n2289,n1980,n1984);
not (n2290,n2291);
nand (n2291,n2087,n2091);
not (n2292,n2293);
nor (n2293,n2294,n2301);
nor (n2294,n2295,n2300);
nor (n2295,n2296,n2298);
nor (n2296,n2297,n2217);
nand (n2297,n2168,n2172);
not (n2298,n2299);
nand (n2299,n2218,n2222);
not (n2300,n2250);
not (n2301,n2302);
nor (n2302,n2303,n2305);
nor (n2303,n2304,n2268);
nand (n2304,n2252,n2256);
not (n2305,n2306);
nand (n2306,n2269,n2273);
nand (n2307,n2308,n2727);
nand (n2308,n2309,n2620);
nor (n2309,n2310,n2605);
nor (n2310,n2311,n2476);
nand (n2311,n2312,n2453);
nor (n2312,n2313,n2430);
nor (n2313,n2314,n2403);
nand (n2314,n2315,n2360,n2402);
nand (n2315,n2316,n2328);
xor (n2316,n2317,n2323);
xor (n2317,n2318,n2319);
xor (n2318,n1621,n1625);
xor (n2319,n2320,n74);
or (n2320,n2321,n2322);
and (n2321,n823,n101);
and (n2322,n837,n105);
and (n2323,n74,n2324);
xor (n2324,n2325,n502);
or (n2325,n2326,n2327);
and (n2326,n469,n625);
and (n2327,n473,n629);
nand (n2328,n2329,n2346,n2359);
nand (n2329,n2330,n2331);
xor (n2330,n74,n2324);
nand (n2331,n2332,n2341,n2345);
nand (n2332,n2333,n2337);
xor (n2333,n2334,n185);
or (n2334,n2335,n2336);
and (n2335,n798,n322);
and (n2336,n800,n326);
xor (n2337,n2338,n324);
or (n2338,n2339,n2340);
and (n2339,n609,n500);
and (n2340,n794,n504);
nand (n2341,n2342,n2337);
and (n2342,n103,n2343);
xnor (n2343,n2344,n103);
nand (n2344,n837,n183);
nand (n2345,n2333,n2342);
nand (n2346,n2347,n2331);
xor (n2347,n2348,n2355);
xor (n2348,n2349,n2353);
xnor (n2349,n2350,n627);
nor (n2350,n2351,n2352);
and (n2351,n293,n809);
and (n2352,n221,n811);
xnor (n2353,n2354,n74);
nand (n2354,n837,n101);
xor (n2355,n2356,n185);
or (n2356,n2357,n2358);
and (n2357,n794,n322);
and (n2358,n798,n326);
nand (n2359,n2330,n2347);
nand (n2360,n2361,n2328);
xor (n2361,n2362,n2381);
xor (n2362,n2363,n2367);
nand (n2363,n2364,n2365,n2366);
nand (n2364,n2349,n2353);
nand (n2365,n2355,n2353);
nand (n2366,n2349,n2355);
xor (n2367,n2368,n2377);
xor (n2368,n2369,n2373);
xor (n2369,n2370,n185);
or (n2370,n2371,n2372);
and (n2371,n609,n322);
and (n2372,n794,n326);
xor (n2373,n2374,n324);
or (n2374,n2375,n2376);
and (n2375,n473,n500);
and (n2376,n475,n504);
xor (n2377,n2378,n103);
or (n2378,n2379,n2380);
and (n2379,n798,n183);
and (n2380,n800,n187);
nand (n2381,n2382,n2396,n2401);
nand (n2382,n2383,n2387);
xor (n2383,n2384,n324);
or (n2384,n2385,n2386);
and (n2385,n475,n500);
and (n2386,n609,n504);
and (n2387,n2388,n2392);
xnor (n2388,n2389,n627);
nor (n2389,n2390,n2391);
and (n2390,n469,n809);
and (n2391,n293,n811);
xor (n2392,n2393,n502);
or (n2393,n2394,n2395);
and (n2394,n473,n625);
and (n2395,n475,n629);
nand (n2396,n2397,n2387);
xor (n2397,n2398,n103);
or (n2398,n2399,n2400);
and (n2399,n800,n183);
and (n2400,n823,n187);
nand (n2401,n2383,n2397);
nand (n2402,n2316,n2361);
xor (n2403,n2404,n2418);
xor (n2404,n2405,n2414);
xor (n2405,n2406,n2412);
xor (n2406,n2407,n2411);
xor (n2407,n2408,n74);
or (n2408,n2409,n2410);
and (n2409,n800,n101);
and (n2410,n823,n105);
xor (n2411,n1565,n15);
xor (n2412,n2413,n1608);
xor (n2413,n1601,n1605);
nand (n2414,n2415,n2416,n2417);
nand (n2415,n2363,n2367);
nand (n2416,n2381,n2367);
nand (n2417,n2363,n2381);
xor (n2418,n2419,n2428);
xor (n2419,n2420,n2424);
nand (n2420,n2421,n2422,n2423);
nand (n2421,n2318,n2319);
nand (n2422,n2323,n2319);
nand (n2423,n2318,n2323);
nand (n2424,n2425,n2426,n2427);
nand (n2425,n2369,n2373);
nand (n2426,n2377,n2373);
nand (n2427,n2369,n2377);
xor (n2428,n2429,n1630);
xor (n2429,n1616,n1620);
nor (n2430,n2431,n2435);
nand (n2431,n2432,n2433,n2434);
nand (n2432,n2405,n2414);
nand (n2433,n2418,n2414);
nand (n2434,n2405,n2418);
xor (n2435,n2436,n2443);
xor (n2436,n2437,n2439);
xor (n2437,n2438,n1614);
xor (n2438,n1595,n1599);
nand (n2439,n2440,n2441,n2442);
nand (n2440,n2420,n2424);
nand (n2441,n2428,n2424);
nand (n2442,n2420,n2428);
xor (n2443,n2444,n2449);
xor (n2444,n2445,n2447);
xor (n2445,n2446,n1564);
xor (n2446,n1555,n1559);
xor (n2447,n2448,n1579);
xor (n2448,n1573,n1577);
nand (n2449,n2450,n2451,n2452);
nand (n2450,n2407,n2411);
nand (n2451,n2412,n2411);
nand (n2452,n2407,n2412);
nor (n2453,n2454,n2469);
nor (n2454,n2455,n2459);
nand (n2455,n2456,n2457,n2458);
nand (n2456,n2437,n2439);
nand (n2457,n2443,n2439);
nand (n2458,n2437,n2443);
xor (n2459,n2460,n2467);
xor (n2460,n2461,n2463);
xor (n2461,n2462,n1571);
xor (n2462,n1551,n1553);
nand (n2463,n2464,n2465,n2466);
nand (n2464,n2445,n2447);
nand (n2465,n2449,n2447);
nand (n2466,n2445,n2449);
xor (n2467,n2468,n1593);
xor (n2468,n1588,n1590);
nor (n2469,n2470,n2474);
nand (n2470,n2471,n2472,n2473);
nand (n2471,n2461,n2463);
nand (n2472,n2467,n2463);
nand (n2473,n2461,n2467);
xor (n2474,n2475,n1586);
xor (n2475,n1461,n1512);
nor (n2476,n2477,n2599);
nor (n2477,n2478,n2575);
nor (n2478,n2479,n2572);
nor (n2479,n2480,n2548);
nand (n2480,n2481,n2520);
or (n2481,n2482,n2506,n2519);
and (n2482,n2483,n2492);
xor (n2483,n2484,n2488);
xnor (n2484,n2485,n627);
nor (n2485,n2486,n2487);
and (n2486,n475,n809);
and (n2487,n473,n811);
xnor (n2488,n2489,n502);
nor (n2489,n2490,n2491);
and (n2490,n794,n629);
and (n2491,n609,n625);
or (n2492,n2493,n2500,n2505);
and (n2493,n2494,n2496);
not (n2494,n2495);
nand (n2495,n837,n322);
xnor (n2496,n2497,n627);
nor (n2497,n2498,n2499);
and (n2498,n609,n809);
and (n2499,n475,n811);
and (n2500,n2496,n2501);
xnor (n2501,n2502,n502);
nor (n2502,n2503,n2504);
and (n2503,n798,n629);
and (n2504,n794,n625);
and (n2505,n2494,n2501);
and (n2506,n2492,n2507);
xor (n2507,n2508,n2515);
xor (n2508,n2509,n2511);
and (n2509,n185,n2510);
xnor (n2510,n2495,n185);
xnor (n2511,n2512,n324);
nor (n2512,n2513,n2514);
and (n2513,n800,n504);
and (n2514,n798,n500);
xnor (n2515,n2516,n185);
nor (n2516,n2517,n2518);
and (n2517,n837,n326);
and (n2518,n823,n322);
and (n2519,n2483,n2507);
xor (n2520,n2521,n2537);
xor (n2521,n2522,n2526);
or (n2522,n2523,n2524,n2525);
and (n2523,n2509,n2511);
and (n2524,n2511,n2515);
and (n2525,n2509,n2515);
xor (n2526,n2527,n2533);
xor (n2527,n2528,n2529);
and (n2528,n2484,n2488);
xnor (n2529,n2530,n324);
nor (n2530,n2531,n2532);
and (n2531,n798,n504);
and (n2532,n794,n500);
xnor (n2533,n2534,n185);
nor (n2534,n2535,n2536);
and (n2535,n823,n326);
and (n2536,n800,n322);
xor (n2537,n2538,n2544);
xor (n2538,n2539,n2540);
not (n2539,n2344);
xnor (n2540,n2541,n627);
nor (n2541,n2542,n2543);
and (n2542,n473,n809);
and (n2543,n469,n811);
xnor (n2544,n2545,n502);
nor (n2545,n2546,n2547);
and (n2546,n609,n629);
and (n2547,n475,n625);
nor (n2548,n2549,n2553);
or (n2549,n2550,n2551,n2552);
and (n2550,n2522,n2526);
and (n2551,n2526,n2537);
and (n2552,n2522,n2537);
xor (n2553,n2554,n2561);
xor (n2554,n2555,n2559);
or (n2555,n2556,n2557,n2558);
and (n2556,n2528,n2529);
and (n2557,n2529,n2533);
and (n2558,n2528,n2533);
xor (n2559,n2560,n2342);
xor (n2560,n2333,n2337);
xor (n2561,n2562,n2568);
xor (n2562,n2563,n2567);
xor (n2563,n2564,n103);
or (n2564,n2565,n2566);
and (n2565,n823,n183);
and (n2566,n837,n187);
xor (n2567,n2388,n2392);
or (n2568,n2569,n2570,n2571);
and (n2569,n2539,n2540);
and (n2570,n2540,n2544);
and (n2571,n2539,n2544);
not (n2572,n2573);
not (n2573,n2574);
and (n2574,n2549,n2553);
not (n2575,n2576);
nor (n2576,n2577,n2592);
nor (n2577,n2578,n2582);
nand (n2578,n2579,n2580,n2581);
nand (n2579,n2555,n2559);
nand (n2580,n2561,n2559);
nand (n2581,n2555,n2561);
xor (n2582,n2583,n2590);
xor (n2583,n2584,n2586);
xor (n2584,n2585,n2397);
xor (n2585,n2383,n2387);
nand (n2586,n2587,n2588,n2589);
nand (n2587,n2563,n2567);
nand (n2588,n2568,n2567);
nand (n2589,n2563,n2568);
xor (n2590,n2591,n2347);
xor (n2591,n2330,n2331);
nor (n2592,n2593,n2597);
nand (n2593,n2594,n2595,n2596);
nand (n2594,n2584,n2586);
nand (n2595,n2590,n2586);
nand (n2596,n2584,n2590);
xor (n2597,n2598,n2361);
xor (n2598,n2316,n2328);
not (n2599,n2600);
nor (n2600,n2601,n2603);
nor (n2601,n2602,n2592);
nand (n2602,n2578,n2582);
not (n2603,n2604);
nand (n2604,n2593,n2597);
not (n2605,n2606);
nor (n2606,n2607,n2614);
nor (n2607,n2608,n2613);
nor (n2608,n2609,n2611);
nor (n2609,n2610,n2430);
nand (n2610,n2314,n2403);
not (n2611,n2612);
nand (n2612,n2431,n2435);
not (n2613,n2453);
not (n2614,n2615);
nor (n2615,n2616,n2618);
nor (n2616,n2617,n2469);
nand (n2617,n2455,n2459);
not (n2618,n2619);
nand (n2619,n2470,n2474);
nand (n2620,n2621,n2625);
nor (n2621,n2622,n2311);
nand (n2622,n2623,n2576);
nor (n2623,n2624,n2548);
nor (n2624,n2481,n2520);
or (n2625,n2626,n2648);
and (n2626,n2627,n2629);
xor (n2627,n2628,n2507);
xor (n2628,n2483,n2492);
or (n2629,n2630,n2644,n2647);
and (n2630,n2631,n2640);
and (n2631,n2632,n2636);
xnor (n2632,n2633,n627);
nor (n2633,n2634,n2635);
and (n2634,n794,n809);
and (n2635,n609,n811);
xnor (n2636,n2637,n502);
nor (n2637,n2638,n2639);
and (n2638,n800,n629);
and (n2639,n798,n625);
xnor (n2640,n2641,n324);
nor (n2641,n2642,n2643);
and (n2642,n823,n504);
and (n2643,n800,n500);
and (n2644,n2640,n2645);
xor (n2645,n2646,n2501);
xor (n2646,n2494,n2496);
and (n2647,n2631,n2645);
and (n2648,n2649,n2650);
xor (n2649,n2627,n2629);
or (n2650,n2651,n2666);
and (n2651,n2652,n2664);
or (n2652,n2653,n2658,n2663);
and (n2653,n2654,n2655);
xor (n2654,n2632,n2636);
and (n2655,n324,n2656);
xnor (n2656,n2657,n324);
nand (n2657,n837,n500);
and (n2658,n2655,n2659);
xnor (n2659,n2660,n324);
nor (n2660,n2661,n2662);
and (n2661,n837,n504);
and (n2662,n823,n500);
and (n2663,n2654,n2659);
xor (n2664,n2665,n2645);
xor (n2665,n2631,n2640);
and (n2666,n2667,n2668);
xor (n2667,n2652,n2664);
or (n2668,n2669,n2685);
and (n2669,n2670,n2672);
xor (n2670,n2671,n2659);
xor (n2671,n2654,n2655);
or (n2672,n2673,n2679,n2684);
and (n2673,n2674,n2675);
not (n2674,n2657);
xnor (n2675,n2676,n627);
nor (n2676,n2677,n2678);
and (n2677,n798,n809);
and (n2678,n794,n811);
and (n2679,n2675,n2680);
xnor (n2680,n2681,n502);
nor (n2681,n2682,n2683);
and (n2682,n823,n629);
and (n2683,n800,n625);
and (n2684,n2674,n2680);
and (n2685,n2686,n2687);
xor (n2686,n2670,n2672);
or (n2687,n2688,n2699);
and (n2688,n2689,n2691);
xor (n2689,n2690,n2680);
xor (n2690,n2674,n2675);
and (n2691,n2692,n2695);
and (n2692,n502,n2693);
xnor (n2693,n2694,n502);
nand (n2694,n837,n625);
xnor (n2695,n2696,n627);
nor (n2696,n2697,n2698);
and (n2697,n800,n809);
and (n2698,n798,n811);
and (n2699,n2700,n2701);
xor (n2700,n2689,n2691);
or (n2701,n2702,n2708);
and (n2702,n2703,n2707);
xnor (n2703,n2704,n502);
nor (n2704,n2705,n2706);
and (n2705,n837,n629);
and (n2706,n823,n625);
xor (n2707,n2692,n2695);
and (n2708,n2709,n2710);
xor (n2709,n2703,n2707);
or (n2710,n2711,n2717);
and (n2711,n2712,n2716);
xnor (n2712,n2713,n627);
nor (n2713,n2714,n2715);
and (n2714,n823,n809);
and (n2715,n800,n811);
not (n2716,n2694);
and (n2717,n2718,n2719);
xor (n2718,n2712,n2716);
and (n2719,n2720,n2724);
xnor (n2720,n2721,n627);
nor (n2721,n2722,n2723);
and (n2722,n837,n809);
and (n2723,n823,n811);
and (n2724,n2725,n627);
xnor (n2725,n2726,n627);
nand (n2726,n837,n811);
not (n2727,n2728);
nand (n2728,n2729,n1749);
nor (n2729,n2730,n781);
nand (n2730,n2731,n1704);
nor (n2731,n2732,n1676);
nor (n2732,n1459,n1638);
not (n2733,n2734);
nand (n2734,n2735,n746);
nor (n2735,n2736,n718);
nor (n2736,n373,n680);
not (n2737,n2738);
nor (n2738,n3,n243);
nand (n2739,n2740,n2796);
not (n2740,n2741);
nor (n2741,n2742,n2746);
nand (n2742,n2743,n2744,n2745);
nand (n2743,n5,n91);
nand (n2744,n200,n91);
nand (n2745,n5,n200);
xor (n2746,n2747,n2792);
xor (n2747,n2748,n2752);
nand (n2748,n2749,n2750,n2751);
nand (n2749,n7,n43);
nand (n2750,n78,n43);
nand (n2751,n7,n78);
xor (n2752,n2753,n2766);
xor (n2753,n2754,n2758);
nand (n2754,n2755,n2756,n2757);
nand (n2755,n66,n95);
nand (n2756,n116,n95);
nand (n2757,n66,n116);
xor (n2758,n2759,n2762);
or (n2759,n2760,n2761);
and (n2760,n52,n60);
and (n2761,n59,n64);
nand (n2762,n2763,n2764,n2765);
nand (n2763,n9,n21);
nand (n2764,n32,n21);
nand (n2765,n9,n32);
xor (n2766,n2767,n2782);
xor (n2767,n2768,n2772);
nand (n2768,n2769,n2770,n2771);
nand (n2769,n45,n56);
nand (n2770,n67,n56);
nand (n2771,n45,n67);
xor (n2772,n2773,n2778);
xor (n2773,n67,n2774);
xor (n2774,n2775,n20);
or (n2775,n2776,n2777);
and (n2776,n71,n13);
and (n2777,n12,n18);
xor (n2778,n2779,n31);
or (n2779,n2780,n2781);
and (n2780,n17,n25);
and (n2781,n24,n29);
xor (n2782,n2783,n2788);
xor (n2783,n2784,n68);
xor (n2784,n2785,n42);
or (n2785,n2786,n2787);
and (n2786,n28,n36);
and (n2787,n35,n40);
xor (n2788,n2789,n55);
or (n2789,n2790,n2791);
and (n2790,n39,n49);
and (n2791,n48,n53);
nand (n2792,n2793,n2794,n2795);
nand (n2793,n93,n128);
nand (n2794,n162,n128);
nand (n2795,n93,n162);
nand (n2796,n2742,n2746);
xor (n2797,n2798,n2954);
xor (n2798,n2799,n2883);
xor (n2799,n2800,n2860);
or (n2800,n2801,n2844,n2859);
and (n2801,n2802,n2810);
xor (n2802,n2803,n2809);
xor (n2803,n2804,n2805);
not (n2804,n79);
or (n2805,n2806,n2807,n2808);
not (n2806,n96);
and (n2807,n107,n118);
and (n2808,n97,n118);
not (n2809,n6);
or (n2810,n2811,n2832,n2843);
and (n2811,n2812,n2819);
xor (n2812,n2813,n2818);
xor (n2813,n132,n2814);
or (n2814,n2815,n2816,n2817);
and (n2815,n98,n151);
not (n2816,n155);
and (n2817,n98,n156);
xor (n2818,n131,n118);
or (n2819,n2820,n2826,n2831);
and (n2820,n280,n2821);
and (n2821,n2822,n296);
or (n2822,n2823,n2824,n2825);
and (n2823,n180,n285);
not (n2824,n284);
and (n2825,n180,n289);
and (n2826,n2821,n2827);
or (n2827,n2828,n2829,n2830);
not (n2828,n230);
and (n2829,n231,n256);
and (n2830,n226,n256);
and (n2831,n280,n2827);
and (n2832,n2819,n2833);
xor (n2833,n2834,n2841);
xor (n2834,n2835,n2836);
not (n2835,n203);
or (n2836,n2837,n2839,n2840);
and (n2837,n171,n2838);
not (n2838,n247);
and (n2839,n2838,n177);
not (n2840,n198);
xor (n2841,n2842,n165);
xor (n2842,n111,n123);
and (n2843,n2812,n2833);
and (n2844,n2810,n2845);
xor (n2845,n2846,n2855);
xor (n2846,n2847,n2851);
or (n2847,n2848,n2849,n2850);
and (n2848,n111,n123);
and (n2849,n123,n165);
and (n2850,n111,n165);
or (n2851,n2852,n2853,n2854);
and (n2852,n132,n2814);
and (n2853,n2814,n2818);
and (n2854,n132,n2818);
or (n2855,n2856,n2857,n2858);
and (n2856,n2835,n2836);
and (n2857,n2836,n2841);
and (n2858,n2835,n2841);
and (n2859,n2802,n2845);
xor (n2860,n2861,n2879);
xor (n2861,n2862,n2866);
or (n2862,n2863,n2864,n2865);
and (n2863,n2804,n2805);
and (n2864,n2805,n2809);
and (n2865,n2804,n2809);
xor (n2866,n2867,n2873);
xor (n2867,n2868,n2871);
xor (n2868,n2869,n2870);
xor (n2869,n2784,n2788);
xor (n2870,n2759,n66);
and (n2871,n7,n2872);
not (n2872,n43);
xor (n2873,n2874,n2772);
xor (n2874,n2762,n2875);
or (n2875,n2876,n2877,n2878);
and (n2876,n68,n45);
not (n2877,n2769);
and (n2878,n68,n56);
or (n2879,n2880,n2881,n2882);
and (n2880,n2847,n2851);
and (n2881,n2851,n2855);
and (n2882,n2847,n2855);
or (n2883,n2884,n2886);
xor (n2884,n2885,n2845);
xor (n2885,n2802,n2810);
or (n2886,n2887,n2918,n2953);
and (n2887,n2888,n2916);
or (n2888,n2889,n2898,n2915);
and (n2889,n2890,n2892);
xor (n2890,n2891,n177);
xor (n2891,n171,n2838);
or (n2892,n2893,n2895,n2897);
and (n2893,n2894,n253);
not (n2894,n306);
and (n2895,n253,n2896);
xor (n2896,n2822,n296);
and (n2897,n2894,n2896);
and (n2898,n2892,n2899);
or (n2899,n2900,n2911,n2914);
and (n2900,n2901,n2906);
or (n2901,n2902,n2904,n2905);
and (n2902,n340,n2903);
not (n2903,n700);
and (n2904,n2903,n699);
and (n2905,n340,n699);
or (n2906,n2907,n2909,n2910);
and (n2907,n343,n2908);
not (n2908,n695);
and (n2909,n2908,n316);
and (n2910,n343,n316);
and (n2911,n2906,n2912);
xor (n2912,n2913,n256);
xor (n2913,n226,n231);
and (n2914,n2901,n2912);
and (n2915,n2890,n2899);
xor (n2916,n2917,n2833);
xor (n2917,n2812,n2819);
and (n2918,n2916,n2919);
or (n2919,n2920,n2949,n2952);
and (n2920,n2921,n2923);
xor (n2921,n2922,n2827);
xor (n2922,n280,n2821);
or (n2923,n2924,n2945,n2948);
and (n2924,n2925,n2943);
or (n2925,n2926,n2939,n2942);
and (n2926,n2927,n2931);
or (n2927,n2928,n2929,n2930);
and (n2928,n379,n453);
and (n2929,n453,n522);
and (n2930,n379,n522);
or (n2931,n2932,n2933,n2938);
and (n2932,n383,n455);
and (n2933,n455,n2934);
or (n2934,n2935,n2936,n2937);
and (n2935,n319,n484);
not (n2936,n520);
and (n2937,n319,n480);
and (n2938,n383,n2934);
and (n2939,n2931,n2940);
xor (n2940,n2941,n699);
xor (n2941,n340,n2903);
and (n2942,n2927,n2940);
xor (n2943,n2944,n2896);
xor (n2944,n2894,n253);
and (n2945,n2943,n2946);
xor (n2946,n2947,n2912);
xor (n2947,n2901,n2906);
and (n2948,n2925,n2946);
and (n2949,n2923,n2950);
xor (n2950,n2951,n2899);
xor (n2951,n2890,n2892);
and (n2952,n2921,n2950);
and (n2953,n2888,n2919);
and (n2954,n2955,n2956);
xnor (n2955,n2884,n2886);
or (n2956,n2957,n3037);
and (n2957,n2958,n2960);
xor (n2958,n2959,n2919);
xor (n2959,n2888,n2916);
or (n2960,n2961,n2963);
xor (n2961,n2962,n2950);
xor (n2962,n2921,n2923);
or (n2963,n2964,n2987,n3036);
and (n2964,n2965,n2985);
or (n2965,n2966,n2981,n2984);
and (n2966,n2967,n2969);
xor (n2967,n2968,n316);
xor (n2968,n343,n2908);
or (n2969,n2970,n2977,n2980);
and (n2970,n451,n2971);
or (n2971,n2972,n2974,n2976);
and (n2972,n512,n2973);
not (n2973,n478);
and (n2974,n2973,n2975);
not (n2975,n464);
and (n2976,n512,n2975);
and (n2977,n2971,n2978);
xor (n2978,n2979,n522);
xor (n2979,n379,n453);
and (n2980,n451,n2978);
and (n2981,n2969,n2982);
xor (n2982,n2983,n2940);
xor (n2983,n2927,n2931);
and (n2984,n2967,n2982);
xor (n2985,n2986,n2946);
xor (n2986,n2925,n2943);
and (n2987,n2985,n2988);
or (n2988,n2989,n3000,n3035);
and (n2989,n2990,n2998);
or (n2990,n2991,n2994,n2997);
and (n2991,n2992,n399);
xor (n2992,n2993,n2934);
xor (n2993,n383,n455);
and (n2994,n399,n2995);
xor (n2995,n2996,n2978);
xor (n2996,n451,n2971);
and (n2997,n2992,n2995);
xor (n2998,n2999,n2982);
xor (n2999,n2967,n2969);
and (n3000,n2998,n3001);
or (n3001,n3002,n3031,n3034);
and (n3002,n3003,n3016);
or (n3003,n3004,n3014,n3015);
and (n3004,n3005,n557);
or (n3005,n3006,n3011,n3013);
and (n3006,n3007,n551);
or (n3007,n3008,n3009,n3010);
and (n3008,n496,n541);
not (n3009,n545);
and (n3010,n496,n546);
and (n3011,n551,n3012);
not (n3012,n554);
and (n3013,n3007,n3012);
not (n3014,n592);
and (n3015,n3005,n593);
or (n3016,n3017,n3024,n3030);
and (n3017,n3018,n3022);
or (n3018,n3019,n3020,n3021);
and (n3019,n497,n493);
not (n3020,n511);
and (n3021,n497,n507);
xor (n3022,n3023,n2975);
xor (n3023,n512,n2973);
and (n3024,n3022,n3025);
or (n3025,n3026,n3027,n3029);
and (n3026,n496,n634);
and (n3027,n634,n3028);
not (n3028,n2229);
and (n3029,n496,n3028);
and (n3030,n3018,n3025);
and (n3031,n3016,n3032);
xor (n3032,n3033,n2995);
xor (n3033,n2992,n399);
and (n3034,n3003,n3032);
and (n3035,n2990,n3001);
and (n3036,n2965,n2988);
and (n3037,n3038,n3039);
xor (n3038,n2958,n2960);
and (n3039,n3040,n3041);
xnor (n3040,n2961,n2963);
or (n3041,n3042,n3127);
and (n3042,n3043,n3045);
xor (n3043,n3044,n2988);
xor (n3044,n2965,n2985);
or (n3045,n3046,n3048);
xor (n3046,n3047,n3001);
xor (n3047,n2990,n2998);
or (n3048,n3049,n3071,n3126);
and (n3049,n3050,n3069);
or (n3050,n3051,n3065,n3068);
and (n3051,n3052,n3054);
xor (n3052,n3053,n593);
xor (n3053,n3005,n557);
or (n3054,n3055,n3058,n3064);
and (n3055,n3056,n2232);
xor (n3056,n3057,n3012);
xor (n3057,n3007,n551);
and (n3058,n2232,n3059);
or (n3059,n3060,n3061,n3063);
not (n3060,n673);
and (n3061,n657,n3062);
not (n3062,n654);
and (n3063,n638,n3062);
and (n3064,n3056,n3059);
and (n3065,n3054,n3066);
xor (n3066,n3067,n3025);
xor (n3067,n3018,n3022);
and (n3068,n3052,n3066);
xor (n3069,n3070,n3032);
xor (n3070,n3003,n3016);
and (n3071,n3069,n3072);
or (n3072,n3073,n3088,n3125);
and (n3073,n3074,n3086);
or (n3074,n3075,n3082,n3085);
and (n3075,n3076,n3080);
or (n3076,n3077,n3078,n3079);
and (n3077,n605,n2202);
and (n3078,n2202,n2183);
and (n3079,n605,n2183);
xor (n3080,n3081,n3028);
xor (n3081,n496,n634);
and (n3082,n3080,n3083);
and (n3083,n2178,n3084);
not (n3084,n2176);
and (n3085,n3076,n3083);
xor (n3086,n3087,n3066);
xor (n3087,n3052,n3054);
and (n3088,n3086,n3089);
or (n3089,n3090,n3110,n3124);
and (n3090,n3091,n3108);
or (n3091,n3092,n3097,n3107);
and (n3092,n3093,n2205);
or (n3093,n3094,n3095,n3096);
and (n3094,n622,n613);
not (n3095,n612);
and (n3096,n622,n616);
and (n3097,n2205,n3098);
or (n3098,n3099,n3104,n3106);
and (n3099,n621,n3100);
or (n3100,n3101,n3102,n3103);
and (n3101,n621,n2006);
not (n3102,n2120);
and (n3103,n621,n2010);
and (n3104,n3100,n3105);
not (n3105,n2115);
and (n3106,n621,n3105);
and (n3107,n3093,n3098);
xor (n3108,n3109,n3059);
xor (n3109,n3056,n2232);
and (n3110,n3108,n3111);
or (n3111,n3112,n3116,n3123);
and (n3112,n3113,n3115);
xor (n3113,n3114,n2183);
xor (n3114,n605,n2202);
not (n3115,n2175);
and (n3116,n3115,n3117);
or (n3117,n3118,n3121,n3122);
and (n3118,n3119,n2121);
and (n3119,n1990,n3120);
not (n3120,n2004);
and (n3121,n2121,n2143);
and (n3122,n3119,n2143);
and (n3123,n3113,n3117);
and (n3124,n3091,n3111);
and (n3125,n3074,n3089);
and (n3126,n3050,n3072);
and (n3127,n3128,n3129);
xor (n3128,n3043,n3045);
and (n3129,n3130,n3131);
xnor (n3130,n3046,n3048);
or (n3131,n3132,n3336);
and (n3132,n3133,n3135);
xor (n3133,n3134,n3072);
xor (n3134,n3050,n3069);
or (n3135,n3136,n3211,n3335);
and (n3136,n3137,n3209);
or (n3137,n3138,n3205,n3208);
and (n3138,n3139,n3141);
xor (n3139,n3140,n3083);
xor (n3140,n3076,n3080);
or (n3141,n3142,n3176,n3204);
and (n3142,n3143,n3174);
or (n3143,n3144,n3162,n3173);
and (n3144,n3145,n3154);
and (n3145,n3146,n2030);
or (n3146,n3147,n3152,n3153);
and (n3147,n3148,n1900);
or (n3148,n3149,n3150,n3151);
and (n3149,n1969,n1765);
not (n3150,n1909);
and (n3151,n1969,n1769);
not (n3152,n2042);
and (n3153,n3148,n1904);
or (n3154,n3155,n3160,n3161);
and (n3155,n2070,n3156);
or (n3156,n3157,n3158,n3159);
and (n3157,n1969,n1889);
not (n3158,n2017);
and (n3159,n1969,n1894);
and (n3160,n3156,n2051);
and (n3161,n2070,n2051);
and (n3162,n3154,n3163);
or (n3163,n3164,n3170,n3172);
and (n3164,n3165,n3166);
not (n3165,n1989);
or (n3166,n3167,n3168,n3169);
and (n3167,n1773,n1965);
not (n3168,n2069);
and (n3169,n1773,n1970);
and (n3170,n3166,n3171);
not (n3171,n2046);
and (n3172,n3165,n3171);
and (n3173,n3145,n3163);
xor (n3174,n3175,n3098);
xor (n3175,n3093,n2205);
and (n3176,n3174,n3177);
or (n3177,n3178,n3200,n3203);
and (n3178,n3179,n3181);
xor (n3179,n3180,n3105);
xor (n3180,n621,n3100);
or (n3181,n3182,n3191,n3199);
and (n3182,n3183,n3190);
or (n3183,n3184,n3186,n3189);
and (n3184,n1949,n3185);
not (n3185,n1946);
and (n3186,n3185,n3187);
xor (n3187,n3188,n1894);
xor (n3188,n1969,n1889);
and (n3189,n1949,n3187);
xor (n3190,n3146,n2030);
and (n3191,n3190,n3192);
or (n3192,n3193,n3197,n3198);
and (n3193,n3194,n3195);
not (n3194,n1963);
xor (n3195,n3196,n1904);
xor (n3196,n3148,n1900);
and (n3197,n3195,n1923);
and (n3198,n3194,n1923);
and (n3199,n3183,n3192);
and (n3200,n3181,n3201);
xor (n3201,n3202,n2143);
xor (n3202,n3119,n2121);
and (n3203,n3179,n3201);
and (n3204,n3143,n3177);
and (n3205,n3141,n3206);
xor (n3206,n3207,n3111);
xor (n3207,n3091,n3108);
and (n3208,n3139,n3206);
xor (n3209,n3210,n3089);
xor (n3210,n3074,n3086);
and (n3211,n3209,n3212);
or (n3212,n3213,n3246,n3334);
and (n3213,n3214,n3244);
or (n3214,n3215,n3240,n3243);
and (n3215,n3216,n3218);
xor (n3216,n3217,n3117);
xor (n3217,n3113,n3115);
or (n3218,n3219,n3236,n3239);
and (n3219,n3220,n3222);
xor (n3220,n3221,n3163);
xor (n3221,n3145,n3154);
or (n3222,n3223,n3228,n3235);
and (n3223,n3224,n3226);
xor (n3224,n3225,n2051);
xor (n3225,n2070,n3156);
xor (n3226,n3227,n3171);
xor (n3227,n3165,n3166);
and (n3228,n3226,n3229);
and (n3229,n1914,n3230);
or (n3230,n3231,n3232,n3234);
not (n3231,n1920);
and (n3232,n1780,n3233);
not (n3233,n1763);
and (n3234,n1776,n3233);
and (n3235,n3224,n3229);
and (n3236,n3222,n3237);
xor (n3237,n3238,n3201);
xor (n3238,n3179,n3181);
and (n3239,n3220,n3237);
and (n3240,n3218,n3241);
xor (n3241,n3242,n3177);
xor (n3242,n3143,n3174);
and (n3243,n3216,n3241);
xor (n3244,n3245,n3206);
xor (n3245,n3139,n3141);
and (n3246,n3244,n3247);
or (n3247,n3248,n3305,n3333);
and (n3248,n3249,n3251);
xor (n3249,n3250,n3241);
xor (n3250,n3216,n3218);
or (n3251,n3252,n3284,n3304);
and (n3252,n3253,n3282);
or (n3253,n3254,n3267,n3281);
and (n3254,n3255,n3265);
or (n3255,n3256,n3263,n3264);
and (n3256,n3257,n3261);
or (n3257,n3258,n3259,n3260);
and (n3258,n1828,n1813);
and (n3259,n1813,n1796);
and (n3260,n1828,n1796);
xor (n3261,n3262,n3187);
xor (n3262,n1949,n3185);
and (n3263,n3261,n1974);
and (n3264,n3257,n1974);
xor (n3265,n3266,n3192);
xor (n3266,n3183,n3190);
and (n3267,n3265,n3268);
or (n3268,n3269,n3278,n3280);
and (n3269,n3270,n3276);
or (n3270,n3271,n3272,n3275);
and (n3271,n1818,n1812);
and (n3272,n1812,n3273);
xor (n3273,n3274,n1796);
xor (n3274,n1828,n1813);
and (n3275,n1818,n3273);
xor (n3276,n3277,n1923);
xor (n3277,n3194,n3195);
and (n3278,n3276,n3279);
xor (n3279,n1914,n3230);
and (n3280,n3270,n3279);
and (n3281,n3255,n3268);
xor (n3282,n3283,n3237);
xor (n3283,n3220,n3222);
and (n3284,n3282,n3285);
or (n3285,n3286,n3300,n3303);
and (n3286,n3287,n3289);
xor (n3287,n3288,n3229);
xor (n3288,n3224,n3226);
or (n3289,n3290,n3298,n3299);
and (n3290,n3291,n3293);
xor (n3291,n3292,n1974);
xor (n3292,n3257,n3261);
or (n3293,n3294,n3295,n3297);
not (n3294,n1873);
and (n3295,n1788,n3296);
not (n3296,n1761);
and (n3297,n1784,n3296);
and (n3298,n3293,n1875);
and (n3299,n3291,n1875);
and (n3300,n3289,n3301);
xor (n3301,n3302,n3268);
xor (n3302,n3255,n3265);
and (n3303,n3287,n3301);
and (n3304,n3253,n3285);
and (n3305,n3251,n3306);
or (n3306,n3307,n3309);
xor (n3307,n3308,n3285);
xor (n3308,n3253,n3282);
or (n3309,n3310,n3326,n3332);
and (n3310,n3311,n3324);
or (n3311,n3312,n3320,n3323);
and (n3312,n3313,n3315);
xor (n3313,n3314,n3279);
xor (n3314,n3270,n3276);
or (n3315,n3316,n3318,n3319);
and (n3316,n3317,n1860);
not (n3317,n1759);
not (n3318,n1867);
and (n3319,n3317,n1792);
and (n3320,n3315,n3321);
xor (n3321,n3322,n1875);
xor (n3322,n3291,n3293);
and (n3323,n3313,n3321);
xor (n3324,n3325,n3301);
xor (n3325,n3287,n3289);
and (n3326,n3324,n3327);
or (n3327,n3328,n3330);
or (n3328,n1753,n3329);
not (n3329,n1757);
xor (n3330,n3331,n3321);
xor (n3331,n3313,n3315);
and (n3332,n3311,n3327);
and (n3333,n3249,n3306);
and (n3334,n3214,n3247);
and (n3335,n3137,n3212);
and (n3336,n3337,n3338);
xor (n3337,n3133,n3135);
and (n3338,n3339,n3341);
xor (n3339,n3340,n3212);
xor (n3340,n3137,n3209);
or (n3341,n3342,n3344);
xor (n3342,n3343,n3247);
xor (n3343,n3214,n3244);
and (n3344,n3345,n3346);
not (n3345,n3342);
and (n3346,n3347,n3349);
xor (n3347,n3348,n3306);
xor (n3348,n3249,n3251);
and (n3349,n3350,n3351);
xnor (n3350,n3307,n3309);
and (n3351,n3352,n3354);
xor (n3352,n3353,n3327);
xor (n3353,n3311,n3324);
and (n3354,n3355,n3356);
xnor (n3355,n3328,n3330);
and (n3356,n3357,n3360);
not (n3357,n3358);
nand (n3358,n3359,n2282);
not (n3359,n1752);
nand (n3360,n779,n3361);
nand (n3361,n2729,n2308);
endmodule
