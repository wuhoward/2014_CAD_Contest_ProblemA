module top (out,n3,n6,n7,n25,n29,n33,n36,n43,n45
        ,n52,n53,n62,n69,n71,n77,n83,n89,n98,n100
        ,n107,n114,n124,n130,n139,n150,n151,n155,n160,n182
        ,n188,n229,n238,n243,n256,n301,n363,n436);
output out;
input n3;
input n6;
input n7;
input n25;
input n29;
input n33;
input n36;
input n43;
input n45;
input n52;
input n53;
input n62;
input n69;
input n71;
input n77;
input n83;
input n89;
input n98;
input n100;
input n107;
input n114;
input n124;
input n130;
input n139;
input n150;
input n151;
input n155;
input n160;
input n182;
input n188;
input n229;
input n238;
input n243;
input n256;
input n301;
input n363;
input n436;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n239;
wire n240;
wire n241;
wire n242;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
xor (out,n0,n1465);
nand (n0,n1,n8);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nor (n5,n6,n7);
nand (n8,n9,n1462);
nand (n9,n10,n1461);
or (n10,n11,n520);
not (n11,n12);
nor (n12,n13,n519);
not (n13,n14);
nand (n14,n15,n448);
or (n15,n16,n447);
and (n16,n17,n373);
xor (n17,n18,n191);
xor (n18,n19,n164);
xor (n19,n20,n92);
xor (n20,n21,n64);
xor (n21,n22,n37);
nand (n22,n23,n35);
or (n23,n24,n26);
not (n24,n25);
not (n26,n27);
nor (n27,n28,n30);
not (n28,n29);
nand (n30,n31,n34);
or (n31,n32,n29);
not (n32,n33);
nand (n34,n29,n32);
nand (n35,n30,n36);
nand (n37,n38,n58);
or (n38,n39,n47);
not (n39,n40);
nor (n40,n41,n46);
and (n41,n42,n44);
not (n42,n43);
not (n44,n45);
and (n46,n43,n45);
nand (n47,n48,n55);
not (n48,n49);
nand (n49,n50,n54);
or (n50,n51,n53);
not (n51,n52);
nand (n54,n53,n51);
nand (n55,n56,n57);
nand (n56,n51,n45);
nand (n57,n52,n44);
nand (n58,n49,n59);
nor (n59,n60,n63);
and (n60,n61,n44);
not (n61,n62);
and (n63,n62,n45);
nand (n64,n65,n85);
or (n65,n66,n79);
nand (n66,n67,n73);
nand (n67,n68,n72);
or (n68,n69,n70);
not (n70,n71);
nand (n72,n70,n69);
not (n73,n74);
nand (n74,n75,n78);
or (n75,n76,n69);
not (n76,n77);
nand (n78,n69,n76);
not (n79,n80);
nor (n80,n81,n84);
and (n81,n82,n70);
not (n82,n83);
and (n84,n83,n71);
or (n85,n73,n86);
not (n86,n87);
nor (n87,n88,n90);
and (n88,n89,n71);
and (n90,n91,n70);
not (n91,n89);
xor (n92,n93,n141);
xor (n93,n94,n118);
nand (n94,n95,n110);
or (n95,n96,n103);
nor (n96,n97,n101);
and (n97,n98,n99);
not (n99,n100);
and (n101,n102,n100);
not (n102,n98);
nand (n103,n104,n109);
nor (n104,n105,n108);
and (n105,n106,n45);
not (n106,n107);
and (n108,n107,n44);
xor (n109,n106,n102);
nand (n110,n111,n117);
not (n111,n112);
nor (n112,n113,n115);
and (n113,n102,n114);
and (n115,n116,n98);
not (n116,n114);
not (n117,n104);
nand (n118,n119,n135);
or (n119,n120,n126);
not (n120,n121);
nor (n121,n122,n125);
and (n122,n123,n32);
not (n123,n124);
and (n125,n124,n33);
nand (n126,n127,n132);
not (n127,n128);
nand (n128,n129,n131);
or (n129,n102,n130);
nand (n131,n102,n130);
nand (n132,n133,n134);
or (n133,n130,n32);
nand (n134,n32,n130);
nand (n135,n128,n136);
nand (n136,n137,n140);
or (n137,n33,n138);
not (n138,n139);
or (n140,n32,n139);
not (n141,n142);
nor (n142,n143,n163);
and (n143,n144,n157);
not (n144,n145);
nand (n145,n146,n153);
not (n146,n147);
nand (n147,n148,n152);
or (n148,n149,n151);
not (n149,n150);
nand (n152,n149,n151);
nand (n153,n154,n156);
or (n154,n155,n149);
nand (n156,n149,n155);
nor (n157,n158,n162);
and (n158,n159,n161);
not (n159,n160);
not (n161,n155);
and (n162,n160,n155);
nor (n163,n146,n161);
or (n164,n165,n190);
and (n165,n166,n175);
xor (n166,n167,n142);
nand (n167,n168,n174);
or (n168,n169,n126);
not (n169,n170);
nor (n170,n171,n173);
and (n171,n172,n32);
not (n172,n36);
and (n173,n36,n33);
nand (n174,n128,n121);
nand (n175,n176,n151);
nor (n176,n177,n184);
and (n177,n178,n179);
not (n178,n66);
nor (n179,n180,n183);
and (n180,n181,n70);
not (n181,n182);
and (n183,n182,n71);
and (n184,n74,n185);
nor (n185,n186,n189);
and (n186,n187,n70);
not (n187,n188);
and (n189,n188,n71);
and (n190,n167,n142);
xor (n191,n192,n338);
xor (n192,n193,n285);
xor (n193,n194,n267);
xor (n194,n195,n216);
or (n195,n196,n215);
and (n196,n197,n209);
xor (n197,n198,n205);
nand (n198,n199,n204);
or (n199,n200,n47);
not (n200,n201);
nand (n201,n202,n203);
or (n202,n114,n44);
nand (n203,n44,n114);
nand (n204,n40,n49);
nand (n205,n206,n208);
or (n206,n207,n66);
not (n207,n185);
nand (n208,n74,n80);
nand (n209,n210,n214);
or (n210,n103,n211);
nor (n211,n212,n213);
and (n212,n139,n102);
and (n213,n98,n138);
or (n214,n96,n104);
and (n215,n198,n205);
or (n216,n217,n266);
and (n217,n218,n245);
xor (n218,n219,n240);
nand (n219,n220,n235);
or (n220,n221,n225);
not (n221,n222);
nor (n222,n223,n224);
and (n223,n91,n76);
and (n224,n89,n77);
not (n225,n226);
nor (n226,n227,n231);
nand (n227,n228,n230);
or (n228,n161,n229);
nand (n230,n229,n161);
nor (n231,n232,n234);
and (n232,n233,n77);
not (n233,n229);
and (n234,n229,n76);
nand (n235,n236,n227);
nand (n236,n237,n239);
or (n237,n238,n76);
nand (n239,n76,n238);
nand (n240,n241,n244);
or (n241,n242,n26);
not (n242,n243);
nand (n244,n30,n25);
nand (n245,n246,n262);
or (n246,n247,n252);
not (n247,n248);
nor (n248,n249,n251);
and (n249,n61,n250);
not (n250,n53);
and (n251,n62,n53);
not (n252,n253);
nor (n253,n254,n259);
nor (n254,n255,n257);
and (n255,n256,n250);
and (n257,n53,n258);
not (n258,n256);
nand (n259,n260,n261);
or (n260,n70,n256);
nand (n261,n256,n70);
nand (n262,n259,n263);
nand (n263,n264,n265);
or (n264,n53,n181);
or (n265,n250,n182);
and (n266,n219,n240);
xor (n267,n268,n278);
xor (n268,n269,n271);
nand (n269,n270,n155);
or (n270,n147,n144);
nand (n271,n272,n274);
or (n272,n273,n225);
not (n273,n236);
nand (n274,n275,n227);
nor (n275,n276,n277);
and (n276,n160,n77);
and (n277,n159,n76);
nand (n278,n279,n281);
or (n279,n280,n252);
not (n280,n263);
nand (n281,n259,n282);
nor (n282,n283,n284);
and (n283,n187,n250);
and (n284,n188,n53);
or (n285,n286,n337);
and (n286,n287,n336);
xor (n287,n288,n313);
or (n288,n289,n312);
and (n289,n290,n303);
xor (n290,n291,n298);
nand (n291,n292,n297);
or (n292,n293,n126);
not (n293,n294);
nor (n294,n295,n296);
and (n295,n24,n32);
and (n296,n25,n33);
nand (n297,n170,n128);
nand (n298,n299,n302);
or (n299,n300,n26);
not (n300,n301);
nand (n302,n30,n243);
nand (n303,n304,n306);
or (n304,n305,n146);
not (n305,n157);
or (n306,n145,n307);
not (n307,n308);
or (n308,n309,n311);
and (n309,n310,n155);
not (n310,n238);
and (n311,n238,n161);
and (n312,n291,n298);
or (n313,n314,n335);
and (n314,n315,n329);
xor (n315,n316,n323);
nand (n316,n317,n322);
or (n317,n318,n252);
not (n318,n319);
nor (n319,n320,n321);
and (n320,n42,n250);
and (n321,n43,n53);
nand (n322,n259,n248);
nand (n323,n324,n328);
or (n324,n325,n225);
nor (n325,n326,n327);
and (n326,n82,n77);
and (n327,n83,n76);
nand (n328,n222,n227);
nand (n329,n330,n334);
or (n330,n47,n331);
nor (n331,n332,n333);
and (n332,n44,n100);
and (n333,n45,n99);
or (n334,n48,n200);
and (n335,n316,n323);
xor (n336,n197,n209);
and (n337,n288,n313);
or (n338,n339,n372);
and (n339,n340,n343);
xor (n340,n341,n342);
xor (n341,n218,n245);
xor (n342,n166,n175);
and (n343,n344,n366);
or (n344,n345,n365);
and (n345,n346,n360);
xor (n346,n347,n353);
nand (n347,n348,n352);
or (n348,n349,n66);
nor (n349,n350,n351);
and (n350,n61,n71);
and (n351,n62,n70);
nand (n352,n179,n74);
nand (n353,n354,n359);
or (n354,n355,n126);
not (n355,n356);
nand (n356,n357,n358);
or (n357,n33,n242);
or (n358,n32,n243);
nand (n359,n128,n294);
nand (n360,n361,n364);
or (n361,n362,n26);
not (n362,n363);
nand (n364,n30,n301);
and (n365,n347,n353);
nand (n366,n367,n371);
or (n367,n103,n368);
nor (n368,n369,n370);
and (n369,n102,n124);
and (n370,n98,n123);
or (n371,n104,n211);
and (n372,n341,n342);
or (n373,n374,n446);
and (n374,n375,n410);
xor (n375,n376,n377);
xor (n376,n287,n336);
or (n377,n378,n409);
and (n378,n379,n407);
xor (n379,n380,n406);
or (n380,n381,n405);
and (n381,n382,n397);
xor (n382,n383,n390);
nand (n383,n384,n389);
or (n384,n385,n145);
not (n385,n386);
nor (n386,n387,n388);
and (n387,n91,n161);
and (n388,n89,n155);
nand (n389,n147,n308);
nand (n390,n391,n396);
or (n391,n392,n252);
not (n392,n393);
nand (n393,n394,n395);
or (n394,n53,n116);
or (n395,n250,n114);
nand (n396,n259,n319);
nand (n397,n398,n403);
or (n398,n225,n399);
not (n399,n400);
nor (n400,n401,n402);
and (n401,n76,n187);
and (n402,n188,n77);
or (n403,n325,n404);
not (n404,n227);
and (n405,n383,n390);
xor (n406,n315,n329);
nand (n407,n408,n175);
or (n408,n151,n176);
and (n409,n380,n406);
or (n410,n411,n445);
and (n411,n412,n444);
xor (n412,n413,n414);
xor (n413,n290,n303);
or (n414,n415,n443);
and (n415,n416,n432);
xor (n416,n417,n425);
nand (n417,n418,n423);
or (n418,n419,n47);
not (n419,n420);
nor (n420,n421,n422);
and (n421,n138,n44);
and (n422,n139,n45);
nand (n423,n424,n49);
not (n424,n331);
nand (n425,n426,n431);
or (n426,n427,n103);
not (n427,n428);
nand (n428,n429,n430);
or (n429,n98,n172);
or (n430,n102,n36);
or (n431,n104,n368);
nand (n432,n433,n442);
or (n433,n434,n437);
nand (n434,n435,n151);
not (n435,n436);
not (n437,n438);
nor (n438,n439,n441);
and (n439,n159,n440);
not (n440,n151);
and (n441,n160,n151);
or (n442,n440,n435);
and (n443,n417,n425);
xor (n444,n344,n366);
and (n445,n413,n414);
and (n446,n376,n377);
and (n447,n18,n191);
xor (n448,n449,n516);
xor (n449,n450,n453);
or (n450,n451,n452);
and (n451,n19,n164);
and (n452,n20,n92);
xor (n453,n454,n471);
xor (n454,n455,n468);
xor (n455,n456,n465);
xor (n456,n457,n462);
not (n457,n458);
nand (n458,n459,n461);
or (n459,n460,n225);
not (n460,n275);
nand (n461,n227,n77);
or (n462,n463,n464);
and (n463,n268,n278);
and (n464,n269,n271);
or (n465,n466,n467);
and (n466,n21,n64);
and (n467,n22,n37);
or (n468,n469,n470);
and (n469,n194,n267);
and (n470,n195,n216);
xor (n471,n472,n513);
xor (n472,n473,n490);
xor (n473,n474,n487);
xor (n474,n475,n482);
nand (n475,n476,n478);
or (n476,n477,n252);
not (n477,n282);
nand (n478,n259,n479);
nor (n479,n480,n481);
and (n480,n82,n250);
and (n481,n83,n53);
nand (n482,n483,n485);
or (n483,n484,n126);
not (n484,n136);
nand (n485,n128,n486);
xnor (n486,n99,n33);
nand (n487,n488,n489);
or (n488,n172,n26);
nand (n489,n30,n124);
xor (n490,n491,n505);
xor (n491,n492,n498);
nand (n492,n493,n494);
or (n493,n86,n66);
nand (n494,n74,n495);
nor (n495,n496,n497);
and (n496,n310,n70);
and (n497,n238,n71);
nand (n498,n499,n501);
or (n499,n500,n47);
not (n500,n59);
or (n501,n48,n502);
nor (n502,n503,n504);
and (n503,n181,n45);
and (n504,n182,n44);
nand (n505,n506,n511);
or (n506,n507,n104);
not (n507,n508);
nand (n508,n509,n510);
or (n509,n42,n98);
or (n510,n43,n102);
nand (n511,n111,n512);
not (n512,n103);
or (n513,n514,n515);
and (n514,n93,n141);
and (n515,n94,n118);
or (n516,n517,n518);
and (n517,n192,n338);
and (n518,n193,n285);
nor (n519,n448,n15);
nand (n520,n521,n1460);
or (n521,n522,n611);
nor (n522,n523,n524);
xor (n523,n17,n373);
or (n524,n525,n610);
and (n525,n526,n609);
xor (n526,n527,n528);
xor (n527,n340,n343);
or (n528,n529,n608);
and (n529,n530,n607);
xor (n530,n531,n600);
or (n531,n532,n599);
and (n532,n533,n575);
xor (n533,n534,n552);
or (n534,n535,n551);
and (n535,n536,n544);
xor (n536,n537,n538);
and (n537,n30,n363);
nand (n538,n539,n540);
or (n539,n435,n437);
or (n540,n541,n434);
nor (n541,n542,n543);
and (n542,n440,n238);
and (n543,n151,n310);
nand (n544,n545,n550);
or (n545,n145,n546);
not (n546,n547);
nor (n547,n548,n549);
and (n548,n82,n161);
and (n549,n83,n155);
nand (n550,n147,n386);
and (n551,n537,n538);
or (n552,n553,n574);
and (n553,n554,n568);
xor (n554,n555,n562);
nand (n555,n556,n561);
or (n556,n557,n225);
not (n557,n558);
nand (n558,n559,n560);
or (n559,n77,n181);
or (n560,n76,n182);
nand (n561,n400,n227);
nand (n562,n563,n567);
or (n563,n564,n47);
nor (n564,n565,n566);
and (n565,n123,n45);
and (n566,n124,n44);
nand (n567,n420,n49);
nand (n568,n569,n570);
or (n569,n427,n104);
or (n570,n103,n571);
nor (n571,n572,n573);
and (n572,n25,n102);
and (n573,n98,n24);
and (n574,n555,n562);
or (n575,n576,n598);
and (n576,n577,n591);
xor (n577,n578,n585);
nand (n578,n579,n584);
or (n579,n580,n126);
not (n580,n581);
nand (n581,n582,n583);
or (n582,n33,n300);
or (n583,n32,n301);
nand (n584,n356,n128);
nand (n585,n586,n590);
or (n586,n66,n587);
nor (n587,n588,n589);
and (n588,n42,n71);
and (n589,n43,n70);
or (n590,n73,n349);
nand (n591,n592,n596);
or (n592,n252,n593);
nor (n593,n594,n595);
and (n594,n99,n53);
and (n595,n100,n250);
or (n596,n597,n392);
not (n597,n259);
and (n598,n578,n585);
and (n599,n534,n552);
or (n600,n601,n606);
and (n601,n602,n605);
xor (n602,n603,n604);
xor (n603,n346,n360);
xor (n604,n382,n397);
xor (n605,n416,n432);
and (n606,n603,n604);
xor (n607,n379,n407);
and (n608,n531,n600);
xor (n609,n375,n410);
and (n610,n527,n528);
not (n611,n612);
nand (n612,n613,n1445);
or (n613,n614,n1375);
not (n614,n615);
nand (n615,n616,n1362);
or (n616,n617,n1068);
not (n617,n618);
nand (n618,n619,n1057,n1067);
nand (n619,n620,n813,n917);
nand (n620,n621,n777);
not (n621,n622);
xor (n622,n623,n736);
xor (n623,n624,n665);
xor (n624,n625,n644);
xor (n625,n626,n635);
nand (n626,n627,n631);
or (n627,n47,n628);
nor (n628,n629,n630);
and (n629,n362,n45);
and (n630,n44,n363);
or (n631,n48,n632);
nor (n632,n633,n634);
and (n633,n44,n301);
and (n634,n45,n300);
nand (n635,n636,n640);
or (n636,n225,n637);
nor (n637,n638,n639);
and (n638,n76,n139);
and (n639,n77,n138);
or (n640,n641,n404);
nor (n641,n642,n643);
and (n642,n76,n100);
and (n643,n77,n99);
nand (n644,n645,n664);
or (n645,n646,n653);
not (n646,n647);
nand (n647,n648,n45);
nand (n648,n649,n650);
or (n649,n363,n52);
nand (n650,n651,n250);
not (n651,n652);
and (n652,n363,n52);
not (n653,n654);
nand (n654,n655,n660);
or (n655,n656,n145);
not (n656,n657);
nand (n657,n658,n659);
or (n658,n155,n116);
or (n659,n161,n114);
nand (n660,n147,n661);
nand (n661,n662,n663);
or (n662,n155,n42);
or (n663,n161,n43);
or (n664,n654,n647);
xor (n665,n666,n716);
xor (n666,n667,n688);
or (n667,n668,n687);
and (n668,n669,n677);
xor (n669,n670,n671);
and (n670,n49,n363);
nand (n671,n672,n676);
or (n672,n673,n145);
nor (n673,n674,n675);
and (n674,n99,n155);
and (n675,n100,n161);
nand (n676,n147,n657);
nand (n677,n678,n683);
or (n678,n66,n679);
not (n679,n680);
nor (n680,n681,n682);
and (n681,n24,n70);
and (n682,n25,n71);
or (n683,n73,n684);
nor (n684,n685,n686);
and (n685,n36,n70);
and (n686,n172,n71);
and (n687,n670,n671);
or (n688,n689,n715);
and (n689,n690,n709);
xor (n690,n691,n700);
nand (n691,n692,n696);
or (n692,n252,n693);
nor (n693,n694,n695);
and (n694,n300,n53);
and (n695,n301,n250);
or (n696,n597,n697);
nor (n697,n698,n699);
and (n698,n243,n250);
and (n699,n242,n53);
nand (n700,n701,n705);
or (n701,n702,n434);
nor (n702,n703,n704);
and (n703,n440,n43);
and (n704,n151,n42);
or (n705,n706,n435);
nor (n706,n707,n708);
and (n707,n440,n62);
and (n708,n151,n61);
nand (n709,n710,n714);
or (n710,n225,n711);
nor (n711,n712,n713);
and (n712,n76,n124);
and (n713,n77,n123);
or (n714,n637,n404);
and (n715,n691,n700);
xor (n716,n717,n730);
xor (n717,n718,n724);
nand (n718,n719,n720);
or (n719,n66,n684);
or (n720,n721,n73);
nor (n721,n722,n723);
and (n722,n123,n71);
and (n723,n124,n70);
nand (n724,n725,n726);
or (n725,n252,n697);
or (n726,n597,n727);
nor (n727,n728,n729);
and (n728,n24,n53);
and (n729,n25,n250);
nand (n730,n731,n732);
or (n731,n706,n434);
or (n732,n733,n435);
nor (n733,n734,n735);
and (n734,n440,n182);
and (n735,n151,n181);
or (n736,n737,n776);
and (n737,n738,n775);
xor (n738,n739,n752);
and (n739,n740,n746);
and (n740,n741,n53);
nand (n741,n742,n743);
or (n742,n363,n256);
nand (n743,n744,n70);
not (n744,n745);
and (n745,n363,n256);
nand (n746,n747,n751);
or (n747,n145,n748);
nor (n748,n749,n750);
and (n749,n161,n139);
and (n750,n155,n138);
or (n751,n146,n673);
or (n752,n753,n774);
and (n753,n754,n768);
xor (n754,n755,n762);
nand (n755,n756,n761);
or (n756,n757,n66);
not (n757,n758);
nor (n758,n759,n760);
and (n759,n243,n71);
and (n760,n242,n70);
nand (n761,n74,n680);
nand (n762,n763,n767);
or (n763,n252,n764);
nor (n764,n765,n766);
and (n765,n53,n362);
and (n766,n250,n363);
or (n767,n597,n693);
nand (n768,n769,n773);
or (n769,n434,n770);
nor (n770,n771,n772);
and (n771,n440,n114);
and (n772,n151,n116);
or (n773,n702,n435);
and (n774,n755,n762);
xor (n775,n669,n677);
and (n776,n739,n752);
not (n777,n778);
or (n778,n779,n812);
and (n779,n780,n811);
xor (n780,n781,n782);
xor (n781,n690,n709);
or (n782,n783,n810);
and (n783,n784,n792);
xor (n784,n785,n791);
nand (n785,n786,n790);
or (n786,n225,n787);
nor (n787,n788,n789);
and (n788,n76,n36);
and (n789,n77,n172);
or (n790,n711,n404);
xor (n791,n740,n746);
or (n792,n793,n809);
and (n793,n794,n802);
xor (n794,n795,n796);
and (n795,n259,n363);
nand (n796,n797,n801);
or (n797,n798,n434);
nor (n798,n799,n800);
and (n799,n440,n100);
and (n800,n151,n99);
or (n801,n770,n435);
nand (n802,n803,n808);
or (n803,n66,n804);
not (n804,n805);
nand (n805,n806,n807);
or (n806,n71,n300);
or (n807,n70,n301);
or (n808,n73,n757);
and (n809,n795,n796);
and (n810,n785,n791);
xor (n811,n738,n775);
and (n812,n781,n782);
nor (n813,n814,n854);
not (n814,n815);
or (n815,n816,n817);
xor (n816,n780,n811);
or (n817,n818,n853);
and (n818,n819,n852);
xor (n819,n820,n821);
xor (n820,n754,n768);
or (n821,n822,n851);
and (n822,n823,n836);
xor (n823,n824,n830);
nand (n824,n825,n829);
or (n825,n145,n826);
nor (n826,n827,n828);
and (n827,n161,n124);
and (n828,n155,n123);
or (n829,n146,n748);
nand (n830,n831,n835);
or (n831,n225,n832);
nor (n832,n833,n834);
and (n833,n76,n25);
and (n834,n77,n24);
or (n835,n787,n404);
and (n836,n837,n844);
nor (n837,n838,n70);
nor (n838,n839,n842);
and (n839,n840,n76);
not (n840,n841);
and (n841,n363,n69);
and (n842,n362,n843);
not (n843,n69);
nand (n844,n845,n850);
or (n845,n434,n846);
not (n846,n847);
nor (n847,n848,n849);
and (n848,n139,n151);
and (n849,n138,n440);
or (n850,n798,n435);
and (n851,n824,n830);
xor (n852,n784,n792);
and (n853,n820,n821);
nand (n854,n855,n911);
not (n855,n856);
nor (n856,n857,n886);
xor (n857,n858,n885);
xor (n858,n859,n884);
or (n859,n860,n883);
and (n860,n861,n877);
xor (n861,n862,n869);
nand (n862,n863,n868);
or (n863,n864,n66);
not (n864,n865);
nand (n865,n866,n867);
or (n866,n70,n363);
or (n867,n71,n362);
nand (n868,n74,n805);
nand (n869,n870,n875);
or (n870,n871,n145);
not (n871,n872);
nand (n872,n873,n874);
or (n873,n155,n172);
or (n874,n161,n36);
nand (n875,n876,n147);
not (n876,n826);
nand (n877,n878,n882);
or (n878,n225,n879);
nor (n879,n880,n881);
and (n880,n76,n243);
and (n881,n77,n242);
or (n882,n832,n404);
and (n883,n862,n869);
xor (n884,n794,n802);
xor (n885,n823,n836);
or (n886,n887,n910);
and (n887,n888,n909);
xor (n888,n889,n890);
xor (n889,n837,n844);
or (n890,n891,n908);
and (n891,n892,n901);
xor (n892,n893,n894);
and (n893,n74,n363);
nand (n894,n895,n896);
or (n895,n435,n846);
or (n896,n897,n434);
not (n897,n898);
nand (n898,n899,n900);
or (n899,n124,n440);
nand (n900,n440,n124);
nand (n901,n902,n907);
or (n902,n903,n145);
not (n903,n904);
nand (n904,n905,n906);
or (n905,n155,n24);
or (n906,n161,n25);
nand (n907,n147,n872);
and (n908,n893,n894);
xor (n909,n861,n877);
and (n910,n889,n890);
not (n911,n912);
nor (n912,n913,n914);
xor (n913,n819,n852);
or (n914,n915,n916);
and (n915,n858,n885);
and (n916,n859,n884);
or (n917,n918,n1056);
and (n918,n919,n946);
xor (n919,n920,n945);
or (n920,n921,n944);
and (n921,n922,n943);
xor (n922,n923,n929);
nand (n923,n924,n928);
or (n924,n225,n925);
nor (n925,n926,n927);
and (n926,n76,n301);
and (n927,n77,n300);
or (n928,n879,n404);
nor (n929,n930,n938);
not (n930,n931);
nand (n931,n932,n937);
or (n932,n434,n933);
not (n933,n934);
nor (n934,n935,n936);
and (n935,n36,n151);
and (n936,n172,n440);
nand (n937,n898,n436);
nand (n938,n939,n77);
nand (n939,n940,n942);
or (n940,n941,n155);
and (n941,n363,n229);
or (n942,n363,n229);
xor (n943,n892,n901);
and (n944,n923,n929);
xor (n945,n888,n909);
or (n946,n947,n1055);
and (n947,n948,n972);
xor (n948,n949,n971);
or (n949,n950,n970);
and (n950,n951,n966);
xor (n951,n952,n959);
nand (n952,n953,n958);
or (n953,n954,n145);
not (n954,n955);
nor (n955,n956,n957);
and (n956,n242,n161);
and (n957,n243,n155);
nand (n958,n147,n904);
nand (n959,n960,n965);
or (n960,n961,n225);
not (n961,n962);
nand (n962,n963,n964);
or (n963,n76,n363);
or (n964,n362,n77);
or (n965,n925,n404);
nand (n966,n967,n969);
or (n967,n968,n930);
not (n968,n938);
or (n969,n931,n938);
and (n970,n952,n959);
xor (n971,n922,n943);
or (n972,n973,n1054);
and (n973,n974,n995);
xor (n974,n975,n994);
or (n975,n976,n993);
and (n976,n977,n986);
xor (n977,n978,n979);
and (n978,n227,n363);
nand (n979,n980,n985);
or (n980,n981,n145);
not (n981,n982);
nor (n982,n983,n984);
and (n983,n300,n161);
and (n984,n301,n155);
nand (n985,n147,n955);
nand (n986,n987,n988);
or (n987,n435,n933);
or (n988,n434,n989);
not (n989,n990);
nor (n990,n991,n992);
and (n991,n24,n440);
and (n992,n25,n151);
and (n993,n978,n979);
xor (n994,n951,n966);
nand (n995,n996,n1053);
or (n996,n997,n1013);
nor (n997,n998,n999);
xor (n998,n977,n986);
and (n999,n1000,n1007);
nand (n1000,n1001,n1002);
nand (n1001,n990,n436);
nand (n1002,n1003,n1006);
nor (n1003,n1004,n1005);
and (n1004,n242,n440);
and (n1005,n243,n151);
not (n1006,n434);
not (n1007,n1008);
nand (n1008,n1009,n155);
nand (n1009,n1010,n1012);
or (n1010,n1011,n151);
and (n1011,n363,n150);
or (n1012,n363,n150);
nor (n1013,n1014,n1052);
and (n1014,n1015,n1026);
nand (n1015,n1016,n1020);
nor (n1016,n1017,n1019);
and (n1017,n1018,n1007);
not (n1018,n1000);
and (n1019,n1000,n1008);
nor (n1020,n1021,n1022);
and (n1021,n147,n982);
and (n1022,n144,n1023);
nand (n1023,n1024,n1025);
or (n1024,n161,n363);
or (n1025,n362,n155);
nand (n1026,n1027,n1050);
or (n1027,n1028,n1042);
not (n1028,n1029);
and (n1029,n1030,n1040);
nand (n1030,n1031,n1036);
or (n1031,n435,n1032);
not (n1032,n1033);
nor (n1033,n1034,n1035);
and (n1034,n300,n440);
and (n1035,n301,n151);
nand (n1036,n1037,n1006);
nand (n1037,n1038,n1039);
or (n1038,n440,n363);
or (n1039,n151,n362);
nor (n1040,n1041,n440);
and (n1041,n363,n436);
not (n1042,n1043);
nand (n1043,n1044,n1049);
not (n1044,n1045);
nand (n1045,n1046,n1048);
or (n1046,n435,n1047);
not (n1047,n1003);
nand (n1048,n1033,n1006);
nand (n1049,n147,n363);
nand (n1050,n1051,n1045);
not (n1051,n1049);
nor (n1052,n1016,n1020);
nand (n1053,n998,n999);
and (n1054,n975,n994);
and (n1055,n949,n971);
and (n1056,n920,n945);
nand (n1057,n1058,n620);
or (n1058,n1059,n1061);
not (n1059,n1060);
nand (n1060,n816,n817);
not (n1061,n1062);
nand (n1062,n815,n1063);
nand (n1063,n1064,n1066);
or (n1064,n912,n1065);
nand (n1065,n857,n886);
nand (n1066,n913,n914);
nand (n1067,n622,n778);
not (n1068,n1069);
nor (n1069,n1070,n1325);
nor (n1070,n1071,n1302);
xor (n1071,n1072,n1224);
xor (n1072,n1073,n1142);
xor (n1073,n1074,n1122);
xor (n1074,n1075,n1107);
or (n1075,n1076,n1106);
and (n1076,n1077,n1097);
xor (n1077,n1078,n1088);
nand (n1078,n1079,n1084);
or (n1079,n1080,n66);
not (n1080,n1081);
nand (n1081,n1082,n1083);
or (n1082,n71,n99);
or (n1083,n70,n100);
nand (n1084,n74,n1085);
nor (n1085,n1086,n1087);
and (n1086,n116,n70);
and (n1087,n114,n71);
nand (n1088,n1089,n1093);
or (n1089,n252,n1090);
nor (n1090,n1091,n1092);
and (n1091,n250,n124);
and (n1092,n53,n123);
nand (n1093,n259,n1094);
nor (n1094,n1095,n1096);
and (n1095,n138,n250);
and (n1096,n139,n53);
nand (n1097,n1098,n1102);
or (n1098,n225,n1099);
nor (n1099,n1100,n1101);
and (n1100,n76,n43);
and (n1101,n77,n42);
or (n1102,n1103,n404);
nor (n1103,n1104,n1105);
and (n1104,n76,n62);
and (n1105,n77,n61);
and (n1106,n1078,n1088);
xor (n1107,n1108,n1116);
xor (n1108,n1109,n1113);
nand (n1109,n1110,n1112);
or (n1110,n1111,n252);
not (n1111,n1094);
or (n1112,n593,n597);
nand (n1113,n1114,n1115);
or (n1114,n1103,n225);
nand (n1115,n227,n558);
nand (n1116,n1117,n1121);
or (n1117,n47,n1118);
nor (n1118,n1119,n1120);
and (n1119,n44,n36);
and (n1120,n45,n172);
or (n1121,n48,n564);
xor (n1122,n1123,n1138);
xor (n1123,n1124,n1131);
nand (n1124,n1125,n1130);
or (n1125,n1126,n145);
not (n1126,n1127);
nand (n1127,n1128,n1129);
or (n1128,n155,n187);
or (n1129,n161,n188);
nand (n1130,n147,n547);
nand (n1131,n1132,n1137);
or (n1132,n1133,n126);
not (n1133,n1134);
nand (n1134,n1135,n1136);
or (n1135,n32,n363);
or (n1136,n33,n362);
nand (n1137,n581,n128);
nand (n1138,n1139,n1141);
or (n1139,n66,n1140);
not (n1140,n1085);
or (n1141,n73,n587);
or (n1142,n1143,n1223);
and (n1143,n1144,n1180);
xor (n1144,n1145,n1146);
xor (n1145,n1077,n1097);
xor (n1146,n1147,n1164);
xor (n1147,n1148,n1155);
nand (n1148,n1149,n1153);
or (n1149,n1150,n47);
nor (n1150,n1151,n1152);
and (n1151,n24,n45);
and (n1152,n25,n44);
nand (n1153,n1154,n49);
not (n1154,n1118);
nand (n1155,n1156,n1160);
or (n1156,n1157,n103);
nor (n1157,n1158,n1159);
and (n1158,n102,n301);
and (n1159,n98,n300);
or (n1160,n104,n1161);
nor (n1161,n1162,n1163);
and (n1162,n102,n243);
and (n1163,n98,n242);
and (n1164,n1165,n1170);
nor (n1165,n1166,n102);
nor (n1166,n1167,n1169);
and (n1167,n1168,n44);
nand (n1168,n363,n107);
and (n1169,n362,n106);
nand (n1170,n1171,n1176);
or (n1171,n435,n1172);
not (n1172,n1173);
nor (n1173,n1174,n1175);
and (n1174,n82,n440);
and (n1175,n83,n151);
or (n1176,n1177,n434);
nor (n1177,n1178,n1179);
and (n1178,n187,n151);
and (n1179,n188,n440);
or (n1180,n1181,n1222);
and (n1181,n1182,n1203);
xor (n1182,n1183,n1184);
xor (n1183,n1165,n1170);
or (n1184,n1185,n1202);
and (n1185,n1186,n1195);
xor (n1186,n1187,n1188);
and (n1187,n117,n363);
nand (n1188,n1189,n1191);
or (n1189,n1190,n145);
not (n1190,n661);
nand (n1191,n147,n1192);
nor (n1192,n1193,n1194);
and (n1193,n61,n161);
and (n1194,n62,n155);
nand (n1195,n1196,n1201);
or (n1196,n1197,n73);
not (n1197,n1198);
nand (n1198,n1199,n1200);
or (n1199,n71,n138);
or (n1200,n70,n139);
or (n1201,n66,n721);
and (n1202,n1187,n1188);
or (n1203,n1204,n1221);
and (n1204,n1205,n1215);
xor (n1205,n1206,n1212);
nand (n1206,n1207,n1208);
or (n1207,n727,n252);
nand (n1208,n1209,n259);
nand (n1209,n1210,n1211);
or (n1210,n53,n172);
or (n1211,n250,n36);
nand (n1212,n1213,n1214);
or (n1213,n733,n434);
or (n1214,n1177,n435);
nand (n1215,n1216,n1217);
or (n1216,n632,n47);
or (n1217,n1218,n48);
nor (n1218,n1219,n1220);
and (n1219,n44,n243);
and (n1220,n45,n242);
and (n1221,n1206,n1212);
and (n1222,n1183,n1184);
and (n1223,n1145,n1146);
xor (n1224,n1225,n1263);
xor (n1225,n1226,n1229);
or (n1226,n1227,n1228);
and (n1227,n1147,n1164);
and (n1228,n1148,n1155);
xor (n1229,n1230,n1247);
xor (n1230,n1231,n1234);
nand (n1231,n1232,n1233);
or (n1232,n103,n1161);
or (n1233,n104,n571);
xor (n1234,n1235,n1241);
nor (n1235,n1236,n32);
nor (n1236,n1237,n1239);
and (n1237,n1238,n102);
nand (n1238,n363,n130);
and (n1239,n362,n1240);
not (n1240,n130);
nand (n1241,n1242,n1246);
or (n1242,n1243,n434);
nor (n1243,n1244,n1245);
and (n1244,n91,n151);
and (n1245,n89,n440);
or (n1246,n541,n435);
or (n1247,n1248,n1262);
and (n1248,n1249,n1255);
xor (n1249,n1250,n1251);
nor (n1250,n127,n362);
nand (n1251,n1252,n1253);
or (n1252,n434,n1172);
nand (n1253,n1254,n436);
not (n1254,n1243);
nand (n1255,n1256,n1261);
or (n1256,n145,n1257);
not (n1257,n1258);
nand (n1258,n1259,n1260);
or (n1259,n155,n181);
or (n1260,n161,n182);
or (n1261,n146,n1126);
and (n1262,n1250,n1251);
or (n1263,n1264,n1301);
and (n1264,n1265,n1300);
xor (n1265,n1266,n1281);
or (n1266,n1267,n1280);
and (n1267,n1268,n1276);
xor (n1268,n1269,n1273);
nand (n1269,n1270,n1272);
or (n1270,n1271,n145);
not (n1271,n1192);
nand (n1272,n1258,n147);
nand (n1273,n1274,n1275);
or (n1274,n1197,n66);
nand (n1275,n74,n1081);
nand (n1276,n1277,n1279);
or (n1277,n252,n1278);
not (n1278,n1209);
or (n1279,n597,n1090);
and (n1280,n1269,n1273);
or (n1281,n1282,n1299);
and (n1282,n1283,n1293);
xor (n1283,n1284,n1290);
nand (n1284,n1285,n1289);
or (n1285,n225,n1286);
nor (n1286,n1287,n1288);
and (n1287,n76,n114);
and (n1288,n77,n116);
or (n1289,n1099,n404);
nand (n1290,n1291,n1292);
or (n1291,n47,n1218);
or (n1292,n1150,n48);
nand (n1293,n1294,n1298);
or (n1294,n103,n1295);
nor (n1295,n1296,n1297);
and (n1296,n362,n98);
and (n1297,n363,n102);
or (n1298,n1157,n104);
and (n1299,n1284,n1290);
xor (n1300,n1249,n1255);
and (n1301,n1266,n1281);
or (n1302,n1303,n1324);
and (n1303,n1304,n1307);
xor (n1304,n1305,n1306);
xor (n1305,n1265,n1300);
xor (n1306,n1144,n1180);
or (n1307,n1308,n1323);
and (n1308,n1309,n1312);
xor (n1309,n1310,n1311);
xor (n1310,n1283,n1293);
xor (n1311,n1268,n1276);
or (n1312,n1313,n1322);
and (n1313,n1314,n1319);
xor (n1314,n1315,n1318);
nand (n1315,n1316,n1317);
or (n1316,n225,n641);
or (n1317,n1286,n404);
and (n1318,n654,n646);
or (n1319,n1320,n1321);
and (n1320,n717,n730);
and (n1321,n718,n724);
and (n1322,n1315,n1318);
and (n1323,n1310,n1311);
and (n1324,n1305,n1306);
nand (n1325,n1326,n1355);
nor (n1326,n1327,n1350);
nor (n1327,n1328,n1341);
xor (n1328,n1329,n1340);
xor (n1329,n1330,n1331);
xor (n1330,n1182,n1203);
or (n1331,n1332,n1339);
and (n1332,n1333,n1336);
xor (n1333,n1334,n1335);
xor (n1334,n1205,n1215);
xor (n1335,n1186,n1195);
or (n1336,n1337,n1338);
and (n1337,n625,n644);
and (n1338,n626,n635);
and (n1339,n1334,n1335);
xor (n1340,n1309,n1312);
or (n1341,n1342,n1349);
and (n1342,n1343,n1348);
xor (n1343,n1344,n1345);
xor (n1344,n1314,n1319);
or (n1345,n1346,n1347);
and (n1346,n666,n716);
and (n1347,n667,n688);
xor (n1348,n1333,n1336);
and (n1349,n1344,n1345);
nor (n1350,n1351,n1354);
or (n1351,n1352,n1353);
and (n1352,n623,n736);
and (n1353,n624,n665);
xor (n1354,n1343,n1348);
nand (n1355,n1356,n1358);
not (n1356,n1357);
xor (n1357,n1304,n1307);
not (n1358,n1359);
or (n1359,n1360,n1361);
and (n1360,n1329,n1340);
and (n1361,n1330,n1331);
nor (n1362,n1363,n1374);
and (n1363,n1364,n1365);
not (n1364,n1070);
nand (n1365,n1366,n1373);
or (n1366,n1367,n1368);
not (n1367,n1355);
not (n1368,n1369);
nand (n1369,n1370,n1372);
or (n1370,n1327,n1371);
nand (n1371,n1351,n1354);
nand (n1372,n1328,n1341);
nand (n1373,n1357,n1359);
and (n1374,n1071,n1302);
not (n1375,n1376);
and (n1376,n1377,n1428);
nor (n1377,n1378,n1409);
nor (n1378,n1379,n1380);
xor (n1379,n526,n609);
or (n1380,n1381,n1408);
and (n1381,n1382,n1407);
xor (n1382,n1383,n1384);
xor (n1383,n412,n444);
or (n1384,n1385,n1406);
and (n1385,n1386,n1399);
xor (n1386,n1387,n1398);
or (n1387,n1388,n1397);
and (n1388,n1389,n1394);
xor (n1389,n1390,n1391);
and (n1390,n1235,n1241);
or (n1391,n1392,n1393);
and (n1392,n1123,n1138);
and (n1393,n1124,n1131);
or (n1394,n1395,n1396);
and (n1395,n1108,n1116);
and (n1396,n1109,n1113);
and (n1397,n1390,n1391);
xor (n1398,n533,n575);
or (n1399,n1400,n1405);
and (n1400,n1401,n1404);
xor (n1401,n1402,n1403);
xor (n1402,n554,n568);
xor (n1403,n536,n544);
xor (n1404,n577,n591);
and (n1405,n1402,n1403);
and (n1406,n1387,n1398);
xor (n1407,n530,n607);
and (n1408,n1383,n1384);
nor (n1409,n1410,n1411);
xor (n1410,n1382,n1407);
or (n1411,n1412,n1427);
and (n1412,n1413,n1426);
xor (n1413,n1414,n1415);
xor (n1414,n602,n605);
or (n1415,n1416,n1425);
and (n1416,n1417,n1422);
xor (n1417,n1418,n1421);
or (n1418,n1419,n1420);
and (n1419,n1230,n1247);
and (n1420,n1231,n1234);
xor (n1421,n1389,n1394);
or (n1422,n1423,n1424);
and (n1423,n1074,n1122);
and (n1424,n1075,n1107);
and (n1425,n1418,n1421);
xor (n1426,n1386,n1399);
and (n1427,n1414,n1415);
nor (n1428,n1429,n1440);
nor (n1429,n1430,n1431);
xor (n1430,n1413,n1426);
or (n1431,n1432,n1439);
and (n1432,n1433,n1438);
xor (n1433,n1434,n1435);
xor (n1434,n1401,n1404);
or (n1435,n1436,n1437);
and (n1436,n1225,n1263);
and (n1437,n1226,n1229);
xor (n1438,n1417,n1422);
and (n1439,n1434,n1435);
nor (n1440,n1441,n1442);
xor (n1441,n1433,n1438);
or (n1442,n1443,n1444);
and (n1443,n1072,n1224);
and (n1444,n1073,n1142);
not (n1445,n1446);
nand (n1446,n1447,n1454);
or (n1447,n1448,n1453);
not (n1448,n1449);
nor (n1449,n1450,n1429);
and (n1450,n1451,n1452);
nand (n1451,n1430,n1431);
nand (n1452,n1441,n1442);
not (n1453,n1377);
nor (n1454,n1455,n1459);
and (n1455,n1456,n1457);
not (n1456,n1378);
not (n1457,n1458);
nand (n1458,n1410,n1411);
and (n1459,n1379,n1380);
nand (n1460,n523,n524);
nand (n1461,n11,n520);
not (n1462,n1463);
nand (n1463,n1464,n6);
not (n1464,n7);
wire s0n1465,s1n1465,notn1465;
or (n1465,s0n1465,s1n1465);
not(notn1465,n7);
and (s0n1465,notn1465,n1466);
and (s1n1465,n7,1'b0);
wire s0n1466,s1n1466,notn1466;
or (n1466,s0n1466,s1n1466);
not(notn1466,n6);
and (s0n1466,notn1466,n3);
and (s1n1466,n6,n1467);
xor (n1467,n1468,n2547);
xor (n1468,n1469,n2546);
xor (n1469,n1470,n2516);
xor (n1470,n1471,n2515);
xor (n1471,n1472,n2476);
xor (n1472,n1473,n2475);
xor (n1473,n1474,n2430);
xor (n1474,n1475,n2429);
xor (n1475,n1476,n2378);
xor (n1476,n1477,n2377);
xor (n1477,n1478,n2322);
xor (n1478,n1479,n63);
xor (n1479,n1480,n2260);
xor (n1480,n1481,n2259);
xor (n1481,n1482,n2193);
xor (n1482,n1483,n284);
xor (n1483,n1484,n2119);
xor (n1484,n1485,n2118);
xor (n1485,n1486,n2043);
xor (n1486,n1487,n88);
xor (n1487,n1488,n1957);
xor (n1488,n1489,n1956);
xor (n1489,n1490,n1865);
xor (n1490,n1491,n276);
or (n1491,n1492,n1771);
and (n1492,n1493,n1770);
or (n1493,n1494,n1680);
and (n1494,n1495,n162);
or (n1495,n1496,n1586);
and (n1496,n1497,n1585);
and (n1497,n441,n1498);
or (n1498,n1499,n1502);
and (n1499,n1500,n1501);
and (n1500,n160,n436);
and (n1501,n238,n151);
and (n1502,n1503,n1504);
xor (n1503,n1500,n1501);
or (n1504,n1505,n1508);
and (n1505,n1506,n1507);
and (n1506,n238,n436);
and (n1507,n89,n151);
and (n1508,n1509,n1510);
xor (n1509,n1506,n1507);
or (n1510,n1511,n1513);
and (n1511,n1512,n1175);
and (n1512,n89,n436);
and (n1513,n1514,n1515);
xor (n1514,n1512,n1175);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
and (n1517,n83,n436);
and (n1518,n188,n151);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
and (n1523,n188,n436);
and (n1524,n182,n151);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
and (n1529,n182,n436);
and (n1530,n62,n151);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
and (n1535,n62,n436);
and (n1536,n43,n151);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
and (n1541,n43,n436);
and (n1542,n114,n151);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
and (n1547,n114,n436);
and (n1548,n100,n151);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1554);
and (n1552,n1553,n848);
and (n1553,n100,n436);
and (n1554,n1555,n1556);
xor (n1555,n1553,n848);
or (n1556,n1557,n1560);
and (n1557,n1558,n1559);
and (n1558,n139,n436);
and (n1559,n124,n151);
and (n1560,n1561,n1562);
xor (n1561,n1558,n1559);
or (n1562,n1563,n1565);
and (n1563,n1564,n935);
and (n1564,n124,n436);
and (n1565,n1566,n1567);
xor (n1566,n1564,n935);
or (n1567,n1568,n1570);
and (n1568,n1569,n992);
and (n1569,n36,n436);
and (n1570,n1571,n1572);
xor (n1571,n1569,n992);
or (n1572,n1573,n1575);
and (n1573,n1574,n1005);
and (n1574,n25,n436);
and (n1575,n1576,n1577);
xor (n1576,n1574,n1005);
or (n1577,n1578,n1580);
and (n1578,n1579,n1035);
and (n1579,n243,n436);
and (n1580,n1581,n1582);
xor (n1581,n1579,n1035);
and (n1582,n1583,n1584);
and (n1583,n301,n436);
and (n1584,n363,n151);
and (n1585,n160,n150);
and (n1586,n1587,n1588);
xor (n1587,n1497,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n441,n1498);
and (n1591,n238,n150);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1503,n1504);
and (n1597,n89,n150);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1509,n1510);
and (n1603,n83,n150);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1514,n1515);
and (n1609,n188,n150);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1520,n1521);
and (n1615,n182,n150);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1526,n1527);
and (n1621,n62,n150);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1532,n1533);
and (n1627,n43,n150);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1538,n1539);
and (n1633,n114,n150);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1544,n1545);
and (n1639,n100,n150);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1550,n1551);
and (n1645,n139,n150);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1555,n1556);
and (n1651,n124,n150);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1561,n1562);
and (n1657,n36,n150);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1566,n1567);
and (n1663,n25,n150);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1571,n1572);
and (n1669,n243,n150);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1576,n1577);
and (n1675,n301,n150);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
and (n1678,n1679,n1011);
xor (n1679,n1581,n1582);
and (n1680,n1681,n1682);
xor (n1681,n1495,n162);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1587,n1588);
and (n1685,n238,n155);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1691);
and (n1689,n1690,n388);
xor (n1690,n1593,n1594);
and (n1691,n1692,n1693);
xor (n1692,n1690,n388);
or (n1693,n1694,n1696);
and (n1694,n1695,n549);
xor (n1695,n1599,n1600);
and (n1696,n1697,n1698);
xor (n1697,n1695,n549);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
xor (n1700,n1605,n1606);
and (n1701,n188,n155);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1611,n1612);
and (n1707,n182,n155);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
or (n1710,n1711,n1713);
and (n1711,n1712,n1194);
xor (n1712,n1617,n1618);
and (n1713,n1714,n1715);
xor (n1714,n1712,n1194);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1623,n1624);
and (n1718,n43,n155);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1629,n1630);
and (n1724,n114,n155);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1635,n1636);
and (n1730,n100,n155);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1641,n1642);
and (n1736,n139,n155);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1647,n1648);
and (n1742,n124,n155);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
or (n1745,n1746,n1749);
and (n1746,n1747,n1748);
xor (n1747,n1653,n1654);
and (n1748,n36,n155);
and (n1749,n1750,n1751);
xor (n1750,n1747,n1748);
or (n1751,n1752,n1755);
and (n1752,n1753,n1754);
xor (n1753,n1659,n1660);
and (n1754,n25,n155);
and (n1755,n1756,n1757);
xor (n1756,n1753,n1754);
or (n1757,n1758,n1760);
and (n1758,n1759,n957);
xor (n1759,n1665,n1666);
and (n1760,n1761,n1762);
xor (n1761,n1759,n957);
or (n1762,n1763,n1765);
and (n1763,n1764,n984);
xor (n1764,n1671,n1672);
and (n1765,n1766,n1767);
xor (n1766,n1764,n984);
and (n1767,n1768,n1769);
xor (n1768,n1677,n1678);
and (n1769,n363,n155);
and (n1770,n160,n229);
and (n1771,n1772,n1773);
xor (n1772,n1493,n1770);
or (n1773,n1774,n1777);
and (n1774,n1775,n1776);
xor (n1775,n1681,n1682);
and (n1776,n238,n229);
and (n1777,n1778,n1779);
xor (n1778,n1775,n1776);
or (n1779,n1780,n1783);
and (n1780,n1781,n1782);
xor (n1781,n1687,n1688);
and (n1782,n89,n229);
and (n1783,n1784,n1785);
xor (n1784,n1781,n1782);
or (n1785,n1786,n1789);
and (n1786,n1787,n1788);
xor (n1787,n1692,n1693);
and (n1788,n83,n229);
and (n1789,n1790,n1791);
xor (n1790,n1787,n1788);
or (n1791,n1792,n1795);
and (n1792,n1793,n1794);
xor (n1793,n1697,n1698);
and (n1794,n188,n229);
and (n1795,n1796,n1797);
xor (n1796,n1793,n1794);
or (n1797,n1798,n1801);
and (n1798,n1799,n1800);
xor (n1799,n1703,n1704);
and (n1800,n182,n229);
and (n1801,n1802,n1803);
xor (n1802,n1799,n1800);
or (n1803,n1804,n1807);
and (n1804,n1805,n1806);
xor (n1805,n1709,n1710);
and (n1806,n62,n229);
and (n1807,n1808,n1809);
xor (n1808,n1805,n1806);
or (n1809,n1810,n1813);
and (n1810,n1811,n1812);
xor (n1811,n1714,n1715);
and (n1812,n43,n229);
and (n1813,n1814,n1815);
xor (n1814,n1811,n1812);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1720,n1721);
and (n1818,n114,n229);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1825);
and (n1822,n1823,n1824);
xor (n1823,n1726,n1727);
and (n1824,n100,n229);
and (n1825,n1826,n1827);
xor (n1826,n1823,n1824);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1732,n1733);
and (n1830,n139,n229);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
or (n1833,n1834,n1837);
and (n1834,n1835,n1836);
xor (n1835,n1738,n1739);
and (n1836,n124,n229);
and (n1837,n1838,n1839);
xor (n1838,n1835,n1836);
or (n1839,n1840,n1843);
and (n1840,n1841,n1842);
xor (n1841,n1744,n1745);
and (n1842,n36,n229);
and (n1843,n1844,n1845);
xor (n1844,n1841,n1842);
or (n1845,n1846,n1849);
and (n1846,n1847,n1848);
xor (n1847,n1750,n1751);
and (n1848,n25,n229);
and (n1849,n1850,n1851);
xor (n1850,n1847,n1848);
or (n1851,n1852,n1855);
and (n1852,n1853,n1854);
xor (n1853,n1756,n1757);
and (n1854,n243,n229);
and (n1855,n1856,n1857);
xor (n1856,n1853,n1854);
or (n1857,n1858,n1861);
and (n1858,n1859,n1860);
xor (n1859,n1761,n1762);
and (n1860,n301,n229);
and (n1861,n1862,n1863);
xor (n1862,n1859,n1860);
and (n1863,n1864,n941);
xor (n1864,n1766,n1767);
or (n1865,n1866,n1869);
and (n1866,n1867,n1868);
xor (n1867,n1772,n1773);
and (n1868,n238,n77);
and (n1869,n1870,n1871);
xor (n1870,n1867,n1868);
or (n1871,n1872,n1874);
and (n1872,n1873,n224);
xor (n1873,n1778,n1779);
and (n1874,n1875,n1876);
xor (n1875,n1873,n224);
or (n1876,n1877,n1880);
and (n1877,n1878,n1879);
xor (n1878,n1784,n1785);
and (n1879,n83,n77);
and (n1880,n1881,n1882);
xor (n1881,n1878,n1879);
or (n1882,n1883,n1885);
and (n1883,n1884,n402);
xor (n1884,n1790,n1791);
and (n1885,n1886,n1887);
xor (n1886,n1884,n402);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
xor (n1889,n1796,n1797);
and (n1890,n182,n77);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
or (n1893,n1894,n1897);
and (n1894,n1895,n1896);
xor (n1895,n1802,n1803);
and (n1896,n62,n77);
and (n1897,n1898,n1899);
xor (n1898,n1895,n1896);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1808,n1809);
and (n1902,n43,n77);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1814,n1815);
and (n1908,n114,n77);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
or (n1911,n1912,n1915);
and (n1912,n1913,n1914);
xor (n1913,n1820,n1821);
and (n1914,n100,n77);
and (n1915,n1916,n1917);
xor (n1916,n1913,n1914);
or (n1917,n1918,n1921);
and (n1918,n1919,n1920);
xor (n1919,n1826,n1827);
and (n1920,n139,n77);
and (n1921,n1922,n1923);
xor (n1922,n1919,n1920);
or (n1923,n1924,n1927);
and (n1924,n1925,n1926);
xor (n1925,n1832,n1833);
and (n1926,n124,n77);
and (n1927,n1928,n1929);
xor (n1928,n1925,n1926);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1838,n1839);
and (n1932,n36,n77);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1844,n1845);
and (n1938,n25,n77);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1850,n1851);
and (n1944,n243,n77);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1856,n1857);
and (n1950,n301,n77);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
and (n1953,n1954,n1955);
xor (n1954,n1862,n1863);
and (n1955,n363,n77);
and (n1956,n238,n69);
or (n1957,n1958,n1961);
and (n1958,n1959,n1960);
xor (n1959,n1870,n1871);
and (n1960,n89,n69);
and (n1961,n1962,n1963);
xor (n1962,n1959,n1960);
or (n1963,n1964,n1967);
and (n1964,n1965,n1966);
xor (n1965,n1875,n1876);
and (n1966,n83,n69);
and (n1967,n1968,n1969);
xor (n1968,n1965,n1966);
or (n1969,n1970,n1973);
and (n1970,n1971,n1972);
xor (n1971,n1881,n1882);
and (n1972,n188,n69);
and (n1973,n1974,n1975);
xor (n1974,n1971,n1972);
or (n1975,n1976,n1979);
and (n1976,n1977,n1978);
xor (n1977,n1886,n1887);
and (n1978,n182,n69);
and (n1979,n1980,n1981);
xor (n1980,n1977,n1978);
or (n1981,n1982,n1985);
and (n1982,n1983,n1984);
xor (n1983,n1892,n1893);
and (n1984,n62,n69);
and (n1985,n1986,n1987);
xor (n1986,n1983,n1984);
or (n1987,n1988,n1991);
and (n1988,n1989,n1990);
xor (n1989,n1898,n1899);
and (n1990,n43,n69);
and (n1991,n1992,n1993);
xor (n1992,n1989,n1990);
or (n1993,n1994,n1997);
and (n1994,n1995,n1996);
xor (n1995,n1904,n1905);
and (n1996,n114,n69);
and (n1997,n1998,n1999);
xor (n1998,n1995,n1996);
or (n1999,n2000,n2003);
and (n2000,n2001,n2002);
xor (n2001,n1910,n1911);
and (n2002,n100,n69);
and (n2003,n2004,n2005);
xor (n2004,n2001,n2002);
or (n2005,n2006,n2009);
and (n2006,n2007,n2008);
xor (n2007,n1916,n1917);
and (n2008,n139,n69);
and (n2009,n2010,n2011);
xor (n2010,n2007,n2008);
or (n2011,n2012,n2015);
and (n2012,n2013,n2014);
xor (n2013,n1922,n1923);
and (n2014,n124,n69);
and (n2015,n2016,n2017);
xor (n2016,n2013,n2014);
or (n2017,n2018,n2021);
and (n2018,n2019,n2020);
xor (n2019,n1928,n1929);
and (n2020,n36,n69);
and (n2021,n2022,n2023);
xor (n2022,n2019,n2020);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
xor (n2025,n1934,n1935);
and (n2026,n25,n69);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1940,n1941);
and (n2032,n243,n69);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1946,n1947);
and (n2038,n301,n69);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
and (n2041,n2042,n841);
xor (n2042,n1952,n1953);
or (n2043,n2044,n2046);
and (n2044,n2045,n84);
xor (n2045,n1962,n1963);
and (n2046,n2047,n2048);
xor (n2047,n2045,n84);
or (n2048,n2049,n2051);
and (n2049,n2050,n189);
xor (n2050,n1968,n1969);
and (n2051,n2052,n2053);
xor (n2052,n2050,n189);
or (n2053,n2054,n2056);
and (n2054,n2055,n183);
xor (n2055,n1974,n1975);
and (n2056,n2057,n2058);
xor (n2057,n2055,n183);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n1980,n1981);
and (n2061,n62,n71);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n1986,n1987);
and (n2067,n43,n71);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2073);
and (n2071,n2072,n1087);
xor (n2072,n1992,n1993);
and (n2073,n2074,n2075);
xor (n2074,n2072,n1087);
or (n2075,n2076,n2079);
and (n2076,n2077,n2078);
xor (n2077,n1998,n1999);
and (n2078,n100,n71);
and (n2079,n2080,n2081);
xor (n2080,n2077,n2078);
or (n2081,n2082,n2085);
and (n2082,n2083,n2084);
xor (n2083,n2004,n2005);
and (n2084,n139,n71);
and (n2085,n2086,n2087);
xor (n2086,n2083,n2084);
or (n2087,n2088,n2091);
and (n2088,n2089,n2090);
xor (n2089,n2010,n2011);
and (n2090,n124,n71);
and (n2091,n2092,n2093);
xor (n2092,n2089,n2090);
or (n2093,n2094,n2097);
and (n2094,n2095,n2096);
xor (n2095,n2016,n2017);
and (n2096,n36,n71);
and (n2097,n2098,n2099);
xor (n2098,n2095,n2096);
or (n2099,n2100,n2102);
and (n2100,n2101,n682);
xor (n2101,n2022,n2023);
and (n2102,n2103,n2104);
xor (n2103,n2101,n682);
or (n2104,n2105,n2107);
and (n2105,n2106,n759);
xor (n2106,n2028,n2029);
and (n2107,n2108,n2109);
xor (n2108,n2106,n759);
or (n2109,n2110,n2113);
and (n2110,n2111,n2112);
xor (n2111,n2034,n2035);
and (n2112,n301,n71);
and (n2113,n2114,n2115);
xor (n2114,n2111,n2112);
and (n2115,n2116,n2117);
xor (n2116,n2040,n2041);
and (n2117,n363,n71);
and (n2118,n83,n256);
or (n2119,n2120,n2123);
and (n2120,n2121,n2122);
xor (n2121,n2047,n2048);
and (n2122,n188,n256);
and (n2123,n2124,n2125);
xor (n2124,n2121,n2122);
or (n2125,n2126,n2129);
and (n2126,n2127,n2128);
xor (n2127,n2052,n2053);
and (n2128,n182,n256);
and (n2129,n2130,n2131);
xor (n2130,n2127,n2128);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2057,n2058);
and (n2134,n62,n256);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2063,n2064);
and (n2140,n43,n256);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2069,n2070);
and (n2146,n114,n256);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2074,n2075);
and (n2152,n100,n256);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2080,n2081);
and (n2158,n139,n256);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2086,n2087);
and (n2164,n124,n256);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
or (n2167,n2168,n2171);
and (n2168,n2169,n2170);
xor (n2169,n2092,n2093);
and (n2170,n36,n256);
and (n2171,n2172,n2173);
xor (n2172,n2169,n2170);
or (n2173,n2174,n2177);
and (n2174,n2175,n2176);
xor (n2175,n2098,n2099);
and (n2176,n25,n256);
and (n2177,n2178,n2179);
xor (n2178,n2175,n2176);
or (n2179,n2180,n2183);
and (n2180,n2181,n2182);
xor (n2181,n2103,n2104);
and (n2182,n243,n256);
and (n2183,n2184,n2185);
xor (n2184,n2181,n2182);
or (n2185,n2186,n2189);
and (n2186,n2187,n2188);
xor (n2187,n2108,n2109);
and (n2188,n301,n256);
and (n2189,n2190,n2191);
xor (n2190,n2187,n2188);
and (n2191,n2192,n745);
xor (n2192,n2114,n2115);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
xor (n2195,n2124,n2125);
and (n2196,n182,n53);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2202);
and (n2200,n2201,n251);
xor (n2201,n2130,n2131);
and (n2202,n2203,n2204);
xor (n2203,n2201,n251);
or (n2204,n2205,n2207);
and (n2205,n2206,n321);
xor (n2206,n2136,n2137);
and (n2207,n2208,n2209);
xor (n2208,n2206,n321);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2142,n2143);
and (n2212,n114,n53);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
or (n2215,n2216,n2219);
and (n2216,n2217,n2218);
xor (n2217,n2148,n2149);
and (n2218,n100,n53);
and (n2219,n2220,n2221);
xor (n2220,n2217,n2218);
or (n2221,n2222,n2224);
and (n2222,n2223,n1096);
xor (n2223,n2154,n2155);
and (n2224,n2225,n2226);
xor (n2225,n2223,n1096);
or (n2226,n2227,n2230);
and (n2227,n2228,n2229);
xor (n2228,n2160,n2161);
and (n2229,n124,n53);
and (n2230,n2231,n2232);
xor (n2231,n2228,n2229);
or (n2232,n2233,n2236);
and (n2233,n2234,n2235);
xor (n2234,n2166,n2167);
and (n2235,n36,n53);
and (n2236,n2237,n2238);
xor (n2237,n2234,n2235);
or (n2238,n2239,n2242);
and (n2239,n2240,n2241);
xor (n2240,n2172,n2173);
and (n2241,n25,n53);
and (n2242,n2243,n2244);
xor (n2243,n2240,n2241);
or (n2244,n2245,n2248);
and (n2245,n2246,n2247);
xor (n2246,n2178,n2179);
and (n2247,n243,n53);
and (n2248,n2249,n2250);
xor (n2249,n2246,n2247);
or (n2250,n2251,n2254);
and (n2251,n2252,n2253);
xor (n2252,n2184,n2185);
and (n2253,n301,n53);
and (n2254,n2255,n2256);
xor (n2255,n2252,n2253);
and (n2256,n2257,n2258);
xor (n2257,n2190,n2191);
and (n2258,n363,n53);
and (n2259,n182,n52);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2198,n2199);
and (n2263,n62,n52);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2203,n2204);
and (n2269,n43,n52);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2208,n2209);
and (n2275,n114,n52);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2282);
and (n2279,n2280,n2281);
xor (n2280,n2214,n2215);
and (n2281,n100,n52);
and (n2282,n2283,n2284);
xor (n2283,n2280,n2281);
or (n2284,n2285,n2288);
and (n2285,n2286,n2287);
xor (n2286,n2220,n2221);
and (n2287,n139,n52);
and (n2288,n2289,n2290);
xor (n2289,n2286,n2287);
or (n2290,n2291,n2294);
and (n2291,n2292,n2293);
xor (n2292,n2225,n2226);
and (n2293,n124,n52);
and (n2294,n2295,n2296);
xor (n2295,n2292,n2293);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2231,n2232);
and (n2299,n36,n52);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
or (n2302,n2303,n2306);
and (n2303,n2304,n2305);
xor (n2304,n2237,n2238);
and (n2305,n25,n52);
and (n2306,n2307,n2308);
xor (n2307,n2304,n2305);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2243,n2244);
and (n2311,n243,n52);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2249,n2250);
and (n2317,n301,n52);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
and (n2320,n2321,n652);
xor (n2321,n2255,n2256);
or (n2322,n2323,n2325);
and (n2323,n2324,n46);
xor (n2324,n2265,n2266);
and (n2325,n2326,n2327);
xor (n2326,n2324,n46);
or (n2327,n2328,n2331);
and (n2328,n2329,n2330);
xor (n2329,n2271,n2272);
and (n2330,n114,n45);
and (n2331,n2332,n2333);
xor (n2332,n2329,n2330);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2277,n2278);
and (n2336,n100,n45);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
or (n2339,n2340,n2342);
and (n2340,n2341,n422);
xor (n2341,n2283,n2284);
and (n2342,n2343,n2344);
xor (n2343,n2341,n422);
or (n2344,n2345,n2348);
and (n2345,n2346,n2347);
xor (n2346,n2289,n2290);
and (n2347,n124,n45);
and (n2348,n2349,n2350);
xor (n2349,n2346,n2347);
or (n2350,n2351,n2354);
and (n2351,n2352,n2353);
xor (n2352,n2295,n2296);
and (n2353,n36,n45);
and (n2354,n2355,n2356);
xor (n2355,n2352,n2353);
or (n2356,n2357,n2360);
and (n2357,n2358,n2359);
xor (n2358,n2301,n2302);
and (n2359,n25,n45);
and (n2360,n2361,n2362);
xor (n2361,n2358,n2359);
or (n2362,n2363,n2366);
and (n2363,n2364,n2365);
xor (n2364,n2307,n2308);
and (n2365,n243,n45);
and (n2366,n2367,n2368);
xor (n2367,n2364,n2365);
or (n2368,n2369,n2372);
and (n2369,n2370,n2371);
xor (n2370,n2313,n2314);
and (n2371,n301,n45);
and (n2372,n2373,n2374);
xor (n2373,n2370,n2371);
and (n2374,n2375,n2376);
xor (n2375,n2319,n2320);
and (n2376,n363,n45);
and (n2377,n43,n107);
or (n2378,n2379,n2382);
and (n2379,n2380,n2381);
xor (n2380,n2326,n2327);
and (n2381,n114,n107);
and (n2382,n2383,n2384);
xor (n2383,n2380,n2381);
or (n2384,n2385,n2388);
and (n2385,n2386,n2387);
xor (n2386,n2332,n2333);
and (n2387,n100,n107);
and (n2388,n2389,n2390);
xor (n2389,n2386,n2387);
or (n2390,n2391,n2394);
and (n2391,n2392,n2393);
xor (n2392,n2338,n2339);
and (n2393,n139,n107);
and (n2394,n2395,n2396);
xor (n2395,n2392,n2393);
or (n2396,n2397,n2400);
and (n2397,n2398,n2399);
xor (n2398,n2343,n2344);
and (n2399,n124,n107);
and (n2400,n2401,n2402);
xor (n2401,n2398,n2399);
or (n2402,n2403,n2406);
and (n2403,n2404,n2405);
xor (n2404,n2349,n2350);
and (n2405,n36,n107);
and (n2406,n2407,n2408);
xor (n2407,n2404,n2405);
or (n2408,n2409,n2412);
and (n2409,n2410,n2411);
xor (n2410,n2355,n2356);
and (n2411,n25,n107);
and (n2412,n2413,n2414);
xor (n2413,n2410,n2411);
or (n2414,n2415,n2418);
and (n2415,n2416,n2417);
xor (n2416,n2361,n2362);
and (n2417,n243,n107);
and (n2418,n2419,n2420);
xor (n2419,n2416,n2417);
or (n2420,n2421,n2424);
and (n2421,n2422,n2423);
xor (n2422,n2367,n2368);
and (n2423,n301,n107);
and (n2424,n2425,n2426);
xor (n2425,n2422,n2423);
and (n2426,n2427,n2428);
xor (n2427,n2373,n2374);
not (n2428,n1168);
and (n2429,n114,n98);
or (n2430,n2431,n2434);
and (n2431,n2432,n2433);
xor (n2432,n2383,n2384);
and (n2433,n100,n98);
and (n2434,n2435,n2436);
xor (n2435,n2432,n2433);
or (n2436,n2437,n2440);
and (n2437,n2438,n2439);
xor (n2438,n2389,n2390);
and (n2439,n139,n98);
and (n2440,n2441,n2442);
xor (n2441,n2438,n2439);
or (n2442,n2443,n2446);
and (n2443,n2444,n2445);
xor (n2444,n2395,n2396);
and (n2445,n124,n98);
and (n2446,n2447,n2448);
xor (n2447,n2444,n2445);
or (n2448,n2449,n2452);
and (n2449,n2450,n2451);
xor (n2450,n2401,n2402);
and (n2451,n36,n98);
and (n2452,n2453,n2454);
xor (n2453,n2450,n2451);
or (n2454,n2455,n2458);
and (n2455,n2456,n2457);
xor (n2456,n2407,n2408);
and (n2457,n25,n98);
and (n2458,n2459,n2460);
xor (n2459,n2456,n2457);
or (n2460,n2461,n2464);
and (n2461,n2462,n2463);
xor (n2462,n2413,n2414);
and (n2463,n243,n98);
and (n2464,n2465,n2466);
xor (n2465,n2462,n2463);
or (n2466,n2467,n2470);
and (n2467,n2468,n2469);
xor (n2468,n2419,n2420);
and (n2469,n301,n98);
and (n2470,n2471,n2472);
xor (n2471,n2468,n2469);
and (n2472,n2473,n2474);
xor (n2473,n2425,n2426);
and (n2474,n363,n98);
and (n2475,n100,n130);
or (n2476,n2477,n2480);
and (n2477,n2478,n2479);
xor (n2478,n2435,n2436);
and (n2479,n139,n130);
and (n2480,n2481,n2482);
xor (n2481,n2478,n2479);
or (n2482,n2483,n2486);
and (n2483,n2484,n2485);
xor (n2484,n2441,n2442);
and (n2485,n124,n130);
and (n2486,n2487,n2488);
xor (n2487,n2484,n2485);
or (n2488,n2489,n2492);
and (n2489,n2490,n2491);
xor (n2490,n2447,n2448);
and (n2491,n36,n130);
and (n2492,n2493,n2494);
xor (n2493,n2490,n2491);
or (n2494,n2495,n2498);
and (n2495,n2496,n2497);
xor (n2496,n2453,n2454);
and (n2497,n25,n130);
and (n2498,n2499,n2500);
xor (n2499,n2496,n2497);
or (n2500,n2501,n2504);
and (n2501,n2502,n2503);
xor (n2502,n2459,n2460);
and (n2503,n243,n130);
and (n2504,n2505,n2506);
xor (n2505,n2502,n2503);
or (n2506,n2507,n2510);
and (n2507,n2508,n2509);
xor (n2508,n2465,n2466);
and (n2509,n301,n130);
and (n2510,n2511,n2512);
xor (n2511,n2508,n2509);
and (n2512,n2513,n2514);
xor (n2513,n2471,n2472);
not (n2514,n1238);
and (n2515,n139,n33);
or (n2516,n2517,n2519);
and (n2517,n2518,n125);
xor (n2518,n2481,n2482);
and (n2519,n2520,n2521);
xor (n2520,n2518,n125);
or (n2521,n2522,n2524);
and (n2522,n2523,n173);
xor (n2523,n2487,n2488);
and (n2524,n2525,n2526);
xor (n2525,n2523,n173);
or (n2526,n2527,n2529);
and (n2527,n2528,n296);
xor (n2528,n2493,n2494);
and (n2529,n2530,n2531);
xor (n2530,n2528,n296);
or (n2531,n2532,n2535);
and (n2532,n2533,n2534);
xor (n2533,n2499,n2500);
and (n2534,n243,n33);
and (n2535,n2536,n2537);
xor (n2536,n2533,n2534);
or (n2537,n2538,n2541);
and (n2538,n2539,n2540);
xor (n2539,n2505,n2506);
and (n2540,n301,n33);
and (n2541,n2542,n2543);
xor (n2542,n2539,n2540);
and (n2543,n2544,n2545);
xor (n2544,n2511,n2512);
and (n2545,n363,n33);
and (n2546,n124,n29);
or (n2547,n2548,n2551);
and (n2548,n2549,n2550);
xor (n2549,n2520,n2521);
and (n2550,n36,n29);
and (n2551,n2552,n2553);
xor (n2552,n2549,n2550);
or (n2553,n2554,n2557);
and (n2554,n2555,n2556);
xor (n2555,n2525,n2526);
and (n2556,n25,n29);
and (n2557,n2558,n2559);
xor (n2558,n2555,n2556);
or (n2559,n2560,n2563);
and (n2560,n2561,n2562);
xor (n2561,n2530,n2531);
and (n2562,n243,n29);
and (n2563,n2564,n2565);
xor (n2564,n2561,n2562);
or (n2565,n2566,n2569);
and (n2566,n2567,n2568);
xor (n2567,n2536,n2537);
and (n2568,n301,n29);
and (n2569,n2570,n2571);
xor (n2570,n2567,n2568);
and (n2571,n2572,n2573);
xor (n2572,n2542,n2543);
and (n2573,n363,n29);
endmodule
