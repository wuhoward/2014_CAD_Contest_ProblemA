module top (out,n15,n18,n20,n21,n23,n27,n36,n38,n39
        ,n41,n46,n49,n51,n56,n60,n68,n72,n73,n74
        ,n86,n90,n91,n92,n107,n108,n109,n110,n111,n115
        ,n116,n117,n122,n124,n126,n163,n165,n166,n167,n178
        ,n179,n180,n181,n193,n194,n195,n196,n210,n216,n218
        ,n219,n223,n224,n227,n229,n230,n231,n304,n359,n362
        ,n364,n452,n454,n455,n569,n572,n574,n576,n580,n583
        ,n585,n587,n591,n594,n596,n598,n600,n660,n663,n665
        ,n667,n671,n674,n676,n678,n682,n685,n687,n689,n693
        ,n696,n698,n700,n733,n736,n738,n740,n744,n747,n749
        ,n751,n755,n758,n760,n762,n766,n769,n771,n773,n801
        ,n802,n803,n807,n809,n810,n811,n829,n831,n833,n835
        ,n837,n839,n841,n843,n845,n847,n849,n851,n853,n855
        ,n857,n859,n864,n916,n928,n935,n937,n939,n941,n943
        ,n945,n947,n949,n951,n953,n955,n957,n959,n961,n963
        ,n965,n969,n971,n973,n975,n977,n979,n981,n983,n985
        ,n987,n989,n991,n993,n995,n997,n999,n1003,n1005,n1007
        ,n1009,n1011,n1013,n1015,n1017,n1019,n1021,n1023,n1025,n1027
        ,n1029,n1031,n1033,n1036,n1037,n1044,n1045,n1067,n1101,n1114
        ,n1117,n1119,n1121,n1125,n1128,n1130,n1132,n1136,n1139,n1141
        ,n1143,n1147,n1150,n1152,n1154,n1196,n1200,n1202,n1207,n1209
        ,n1251,n1262,n1267,n1272,n1277,n1285,n1288,n1297,n1301,n1307
        ,n1309,n1311,n1313,n1315,n1323,n1326,n1328,n1330,n1332,n1339
        ,n1340,n1350,n1353,n1357,n1362,n1365,n1368,n1371,n1376,n1378
        ,n1380,n1382,n1384,n1389,n1391,n1398,n1401,n1403,n1413,n1415
        ,n1417,n1419,n1421,n1426,n1428,n1431,n1433,n1435,n1439,n1441
        ,n1444,n1447,n1451,n1453,n1456,n1458,n1459,n1467,n1472,n1476
        ,n1480,n1484,n1489,n1491,n1494,n1496,n1498,n1502,n1504,n1507
        ,n1510,n1514,n1518,n1523,n1527,n1528,n1538,n1540,n1542,n1544
        ,n1546,n1552,n1554,n1556,n1558,n1563,n1564,n1567,n1570,n1573
        ,n1578,n1581,n1584,n1587,n1588,n1595,n1596,n1599,n1602,n1605
        ,n1610,n1613,n1616,n1619,n1624,n1626,n1629,n1633,n1635,n1640
        ,n1642,n1648,n1651,n1652,n1662,n1664,n1666,n1668,n1670,n1673
        ,n1675,n1681,n1683,n1685,n1687,n1689,n1694,n1697,n1699,n1701
        ,n1704,n1706,n1707,n1714,n1715,n1718,n1721,n1724,n1729,n1732
        ,n1735,n1738,n1743,n1745,n1747,n1749,n1751,n1756,n1758,n1764
        ,n1766,n1767,n1777,n1779,n1781,n1783,n1785,n1791,n1793,n1795
        ,n1797,n1802,n1803,n1806,n1809,n1812,n1817,n1820,n1823,n1826
        ,n1827,n1834,n1835,n1838,n1841,n1844,n1849,n1852,n1855,n1858
        ,n1863,n1865,n1868,n1872,n1874,n1879,n1881,n1887,n1890,n1891
        ,n1901,n1903,n1905,n1907,n1909,n1915,n1917,n1919,n1921,n1926
        ,n1927,n1930,n1933,n1936,n1941,n1944,n1947,n1950,n1951,n1958
        ,n1959,n1962,n1965,n1968,n1973,n1976,n1979,n1982,n1987,n1989
        ,n1992,n1996,n1998,n2003,n2005,n2008,n2013,n2014,n2023,n2025
        ,n2028,n2030,n2032,n2036,n2038,n2042,n2044,n2049,n2050,n2053
        ,n2056,n2059,n2064,n2067,n2070,n2073,n2074,n2081,n2082,n2085
        ,n2088,n2091,n2096,n2099,n2102,n2105,n2111,n2113,n2115,n2117
        ,n2119,n2128,n2130,n2132,n2134,n2135,n2144,n2146,n2148,n2150
        ,n2152,n2157,n2160,n2162,n2164,n2169,n2170,n2173,n2176,n2179
        ,n2184,n2187,n2190,n2193,n2194,n2201,n2202,n2205,n2208,n2211
        ,n2216,n2219,n2222,n2225,n2230,n2232,n2235,n2239,n2241,n2246
        ,n2248,n2251,n2256,n2257,n2273,n2275,n2285,n2287,n2289,n2291
        ,n2293,n2298,n2301,n2303,n2305,n2308,n2311,n2313,n2315,n2317
        ,n2320,n2322,n2325,n2327,n2328,n2335,n2337,n2339,n2341,n2343
        ,n2349,n2351,n2353,n2355,n2357,n2362,n2365,n2367,n2369,n2372
        ,n2374,n2377,n2379,n2380,n2391,n2393,n2395,n2397,n2399,n2404
        ,n2407,n2409,n2411,n2414,n2418,n2420,n2422,n2424,n2427,n2429
        ,n2432,n2434,n2435,n2442,n2444,n2449,n2451,n2454,n2459,n2461
        ,n2467,n2470,n2475,n2476,n2479,n2482,n2485,n2490,n2493,n2496
        ,n2499,n2500,n2508,n2512,n2515,n2517,n2519,n2524,n2526,n2529
        ,n2531,n2533,n2537,n2539,n2542,n2545,n2548,n2550,n2553,n2555
        ,n2556,n2561,n2564,n2567,n2569,n2571,n2577,n2579,n2581,n2583
        ,n2585,n2587,n2594,n2596,n2598,n2600,n2602,n2605,n2607,n2608
        ,n2618,n2620,n2625,n2627,n2630,n2635,n2637,n2643,n2646,n2651
        ,n2652,n2655,n2658,n2661,n2666,n2669,n2672,n2675,n2676,n2683
        ,n2685,n2687,n2689,n2691,n2696,n2698,n2704,n2706,n2711,n2712
        ,n2715,n2718,n2721,n2726,n2729,n2732,n2735,n2736,n2746,n2748
        ,n2753,n2755,n2758,n2763,n2765,n2771,n2774,n2779,n2780,n2783
        ,n2786,n2789,n2794,n2797,n2800,n2803,n2804,n2810,n2812,n2815
        ,n2817,n2819,n2823,n2825,n2829,n2831,n2836,n2837,n2840,n2843
        ,n2846,n2851,n2854,n2857,n2860,n2861,n2871,n2873,n2875,n2877
        ,n2879,n2885,n2887,n2889,n2891,n2896,n2897,n2900,n2903,n2906
        ,n2911,n2914,n2917,n2920,n2921,n2928,n2930,n2932,n2934,n2936
        ,n2941,n2944,n2946,n2948,n2953,n2954,n2957,n2960,n2963,n2968
        ,n2971,n2974,n2977,n2978,n2988,n2989,n2992,n2995,n2998,n3003
        ,n3005,n3009,n3011,n3016,n3017,n3020,n3023,n3026,n3031,n3034
        ,n3037,n3040,n3041,n3051,n3053,n3055,n3057,n3059,n3066,n3068
        ,n3070,n3072,n3077,n3078,n3081,n3084,n3087,n3092,n3095,n3098
        ,n3101,n3102,n3112,n3114,n3117,n3119,n3121,n3126,n3128,n3132
        ,n3134,n3139,n3140,n3143,n3146,n3149,n3154,n3157,n3160,n3163
        ,n3164,n3171,n3173,n3176,n3180,n3182,n3187,n3189,n3192,n3197
        ,n3202,n3203,n3206,n3209,n3212,n3217,n3220,n3223,n3226,n3227
        ,n3241,n3243,n3263,n3264,n3267,n3270,n3273,n3278,n3281,n3284
        ,n3287,n3288,n3291,n3296,n3298,n3301,n3303,n3305,n3311,n3313
        ,n3317,n3319,n3331,n3332,n3335,n3338,n3341,n3346,n3349,n3352
        ,n3355,n3356,n3366,n3368,n3370,n3372,n3374,n3380,n3382,n3384
        ,n3386,n3387,n3397,n3399,n3402,n3404,n3421,n3422,n3425,n3428
        ,n3431,n3436,n3439,n3442,n3445,n3446,n3450,n3457,n3459,n3461
        ,n3463,n3465,n3471,n3474,n3476,n3478,n3488,n3489,n3492,n3495
        ,n3498,n3503,n3506,n3509,n3512,n3513,n3520,n3522,n3525,n3527
        ,n3529,n3535,n3537,n3541,n3543,n3545,n3557,n3558,n3561,n3564
        ,n3567,n3572,n3575,n3578,n3581,n3582,n3589,n3591,n3596,n3598
        ,n3601,n3608,n3611,n3613,n3615,n3616,n3630,n3631,n3634,n3637
        ,n3640,n3645,n3648,n3651,n3654,n3655,n3658,n3664,n3666,n3668
        ,n3670,n3672,n3680,n3682,n3684,n3686,n3703,n3704,n3707,n3710
        ,n3713,n3718,n3721,n3724,n3727,n3728,n3736,n3738,n3740,n3742
        ,n3744,n3752,n3754,n3756,n3758,n3759,n3770,n3771,n3774,n3777
        ,n3780,n3785,n3788,n3791,n3794,n3795,n3800,n3809,n3811,n3813
        ,n3815,n3817,n3824,n3826,n3828,n3830,n4126,n4128,n4132,n4134
        ,n4139,n4141,n4159,n4161,n4167,n4169,n4184,n4186,n4252,n4254
        ,n4266,n4268,n4286,n4288,n4307,n4313,n4329,n4336,n4355,n4362
        ,n4368,n4370,n4795,n4797,n5728,n5729,n5732,n5733,n5740,n5741
        ,n5744,n5745,n5779,n5780,n5785,n5786,n5823,n5824,n5827,n5828
        ,n5856,n5857,n5861,n5862,n5893,n5894,n5897,n5898,n5935,n5936
        ,n5940,n5941,n5983,n5984,n5987,n5988,n6019,n6020,n6023,n6024
        ,n6062,n6063,n6066,n6067,n6098,n6099,n6102,n6103,n6140,n6141
        ,n6144,n6145,n6165,n6166,n6171,n6172,n6201,n6202,n6205,n6206
        ,n6237,n6238,n6243,n6244,n6273,n6274,n6277,n6278,n6437,n6440
        ,n6456,n6460,n6470,n6481,n6485,n6489,n6501,n6511,n6514,n6516
        ,n6520,n6522,n6536,n6538,n6550,n6560,n6563,n6565,n6569,n6571
        ,n6585,n6587,n6601,n6609,n6612,n6614,n6630,n6632,n6635,n6637
        ,n6652,n6663,n6666,n6668,n6674,n6689,n6691,n6693,n6705,n6715
        ,n6718,n6720,n6736,n6738,n6741,n6743,n6758,n6768,n6771,n6773
        ,n6779,n6794,n6796,n6798,n6815,n6817,n6819,n6829,n6850,n6852
        ,n6855,n6857,n7035,n7038,n7151,n7154,n7245,n7248,n7373,n7376
        ,n7630,n7633,n7649,n7652,n7783,n7786,n7892,n7895,n8006,n8016
        ,n8019,n8021,n8023,n8027,n8030,n8032,n8034,n8038,n8041,n8043
        ,n8045,n8049,n8052,n8054,n8056,n8064,n8067,n8069,n8071,n8075
        ,n8078,n8080,n8082,n8086,n8089,n8091,n8093,n8097,n8100,n8102
        ,n8104,n8147,n8174,n8189,n8204,n8219,n8234,n8253,n8331,n8342
        ,n8362,n8377,n8392,n8412,n8427,n8436,n8531,n8544,n8550,n8568
        ,n8588,n8598,n8612,n8664,n8671,n8690,n8721,n8782,n8796,n8806
        ,n8826,n8840,n9996,n9999,n10008,n10011,n10030,n10039,n10054,n10059
        ,n10081,n10083,n10086,n10088,n10099,n10101,n10104,n10106,n10116,n10118
        ,n10121,n10123,n10134,n10141,n10142,n10143,n10144,n10152,n10153,n10154
        ,n10155,n10171,n10176,n10187,n10192,n10199,n10202,n10204,n10247,n10248
        ,n10249,n10250,n10253,n10280,n10282,n10291,n10293,n10295,n10305,n10308
        ,n10315,n10318,n10323,n10330,n10343,n10344,n10363,n10404,n10405,n10430
        ,n10434,n10437,n10448,n10451,n10453,n10456,n10461,n10467,n10473,n10476
        ,n10483,n10487,n10492,n10498,n10502,n10540,n10543,n10546,n10548,n10558
        ,n10560,n10563,n10565,n10574,n10576,n10579,n10581,n10590,n10592,n10595
        ,n10597,n10606,n10608,n10611,n10613,n10623,n10626,n10628,n10635,n10637
        ,n10643,n10649,n10652,n10661,n10680,n10682,n10687,n10689,n10691,n10700
        ,n10703,n10705,n10707,n10709,n10711,n10715,n10716,n10729,n10747,n10748
        ,n10771,n10775,n10778,n10789,n10792,n10794,n10799,n10802,n10809,n10817
        ,n10821,n10828,n10831,n10836,n10842,n10846,n10883,n10886,n10889,n10891
        ,n10901,n10903,n10906,n10908,n10917,n10919,n10922,n10924,n10933,n10935
        ,n10938,n10940,n10949,n10951,n10954,n10956,n10966,n10969,n10971,n10975
        ,n10980,n10986,n10992,n10995,n11004,n11023,n11025,n11030,n11032,n11034
        ,n11043,n11046,n11048,n11050,n11052,n11054,n11058,n11059,n11072,n11090
        ,n11091,n11114,n11117,n11119,n11130,n11133,n11135,n11139,n11142,n11146
        ,n11152,n11156,n11167,n11171,n11175,n11181,n11185,n11223,n11226,n11229
        ,n11231,n11241,n11243,n11246,n11248,n11257,n11259,n11262,n11264,n11273
        ,n11275,n11278,n11280,n11289,n11291,n11294,n11296,n11306,n11309,n11311
        ,n11314,n11319,n11325,n11334,n11337,n11346,n11365,n11367,n11372,n11374
        ,n11376,n11385,n11388,n11390,n11392,n11394,n11396,n11400,n11401,n11414
        ,n11432,n11433,n11456,n11459,n11461,n11472,n11475,n11477,n11481,n11484
        ,n11488,n11494,n11498,n11511,n11515,n11519,n11525,n11529,n11567,n11570
        ,n11573,n11575,n11585,n11587,n11590,n11592,n11601,n11603,n11606,n11608
        ,n11617,n11619,n11622,n11624,n11633,n11635,n11638,n11640,n11650,n11653
        ,n11655,n11659,n11662,n11666,n11672,n11676,n11689,n11708,n11710,n11715
        ,n11717,n11719,n11728,n11731,n11733,n11735,n11737,n11739,n11743,n11744
        ,n11757,n11775,n11776,n11798,n11800,n11802,n11813,n11816,n11818,n11822
        ,n11829,n11832,n11835,n11840,n11849,n11851,n11853,n11862,n11866,n11901
        ,n11904,n11907,n11909,n11919,n11921,n11924,n11926,n11935,n11937,n11940
        ,n11942,n11951,n11953,n11956,n11958,n11967,n11969,n11972,n11974,n11984
        ,n11988,n11991,n11996,n12000,n12003,n12005,n12011,n12028,n12047,n12049
        ,n12054,n12056,n12058,n12067,n12070,n12072,n12074,n12076,n12078,n12082
        ,n12083,n12096,n12114,n12115,n12137,n12139,n12141,n12152,n12155,n12157
        ,n12162,n12165,n12170,n12172,n12174,n12189,n12191,n12193,n12203,n12207
        ,n12248,n12251,n12254,n12256,n12266,n12268,n12271,n12273,n12282,n12284
        ,n12287,n12289,n12298,n12300,n12303,n12305,n12314,n12316,n12319,n12321
        ,n12331,n12334,n12336,n12341,n12345,n12349,n12354,n12356,n12370,n12389
        ,n12391,n12396,n12398,n12400,n12409,n12412,n12414,n12416,n12418,n12420
        ,n12424,n12425,n12438,n12456,n12457,n12479,n12481,n12483,n12493,n12495
        ,n12497,n12502,n12506,n12509,n12515,n12517,n12529,n12531,n12533,n12539
        ,n12543,n12582,n12585,n12588,n12590,n12600,n12602,n12605,n12607,n12616
        ,n12618,n12621,n12623,n12632,n12634,n12637,n12639,n12648,n12650,n12653
        ,n12655,n12664,n12666,n12668,n12673,n12677,n12681,n12687,n12691,n12704
        ,n12723,n12725,n12730,n12732,n12734,n12743,n12746,n12748,n12750,n12752
        ,n12754,n12758,n12759,n12772,n12790,n12791,n12813,n12815,n12817,n12827
        ,n12829,n12831,n12835,n12837,n12842,n12846,n12854,n12865,n12867,n12869
        ,n12875,n12879,n12951,n12985,n12988,n12990,n13004,n13017,n13042,n13045
        ,n13047,n13050,n13063,n13086,n13089,n13091,n13094,n13107,n13130,n13133
        ,n13135,n13140,n13153,n13176,n13179,n13181,n13185,n13198,n13220,n13222
        ,n13224,n13230,n13261,n13274,n13276,n13278,n13282,n13298,n13308,n13311
        ,n13313,n13317,n13464,n13480,n13483,n13486,n13488,n13503,n13513,n13525
        ,n13530,n13550,n13553,n13556,n13559,n13561,n13566,n13568,n13579,n13584
        ,n13602,n13605,n13608,n13611,n13613,n13618,n13620,n13631,n13636,n13659
        ,n13662,n13665,n13668,n13670,n13679,n13681,n13692,n13697,n13715,n13718
        ,n13721,n13724,n13726,n13741,n13746,n13765,n13768,n13771,n13774,n13776
        ,n13791,n13796,n13814,n13817,n13820,n13823,n13825,n13840,n13845,n13877
        ,n13880,n13883,n13886,n13888,n13904,n13909);
output out;
input n15;
input n18;
input n20;
input n21;
input n23;
input n27;
input n36;
input n38;
input n39;
input n41;
input n46;
input n49;
input n51;
input n56;
input n60;
input n68;
input n72;
input n73;
input n74;
input n86;
input n90;
input n91;
input n92;
input n107;
input n108;
input n109;
input n110;
input n111;
input n115;
input n116;
input n117;
input n122;
input n124;
input n126;
input n163;
input n165;
input n166;
input n167;
input n178;
input n179;
input n180;
input n181;
input n193;
input n194;
input n195;
input n196;
input n210;
input n216;
input n218;
input n219;
input n223;
input n224;
input n227;
input n229;
input n230;
input n231;
input n304;
input n359;
input n362;
input n364;
input n452;
input n454;
input n455;
input n569;
input n572;
input n574;
input n576;
input n580;
input n583;
input n585;
input n587;
input n591;
input n594;
input n596;
input n598;
input n600;
input n660;
input n663;
input n665;
input n667;
input n671;
input n674;
input n676;
input n678;
input n682;
input n685;
input n687;
input n689;
input n693;
input n696;
input n698;
input n700;
input n733;
input n736;
input n738;
input n740;
input n744;
input n747;
input n749;
input n751;
input n755;
input n758;
input n760;
input n762;
input n766;
input n769;
input n771;
input n773;
input n801;
input n802;
input n803;
input n807;
input n809;
input n810;
input n811;
input n829;
input n831;
input n833;
input n835;
input n837;
input n839;
input n841;
input n843;
input n845;
input n847;
input n849;
input n851;
input n853;
input n855;
input n857;
input n859;
input n864;
input n916;
input n928;
input n935;
input n937;
input n939;
input n941;
input n943;
input n945;
input n947;
input n949;
input n951;
input n953;
input n955;
input n957;
input n959;
input n961;
input n963;
input n965;
input n969;
input n971;
input n973;
input n975;
input n977;
input n979;
input n981;
input n983;
input n985;
input n987;
input n989;
input n991;
input n993;
input n995;
input n997;
input n999;
input n1003;
input n1005;
input n1007;
input n1009;
input n1011;
input n1013;
input n1015;
input n1017;
input n1019;
input n1021;
input n1023;
input n1025;
input n1027;
input n1029;
input n1031;
input n1033;
input n1036;
input n1037;
input n1044;
input n1045;
input n1067;
input n1101;
input n1114;
input n1117;
input n1119;
input n1121;
input n1125;
input n1128;
input n1130;
input n1132;
input n1136;
input n1139;
input n1141;
input n1143;
input n1147;
input n1150;
input n1152;
input n1154;
input n1196;
input n1200;
input n1202;
input n1207;
input n1209;
input n1251;
input n1262;
input n1267;
input n1272;
input n1277;
input n1285;
input n1288;
input n1297;
input n1301;
input n1307;
input n1309;
input n1311;
input n1313;
input n1315;
input n1323;
input n1326;
input n1328;
input n1330;
input n1332;
input n1339;
input n1340;
input n1350;
input n1353;
input n1357;
input n1362;
input n1365;
input n1368;
input n1371;
input n1376;
input n1378;
input n1380;
input n1382;
input n1384;
input n1389;
input n1391;
input n1398;
input n1401;
input n1403;
input n1413;
input n1415;
input n1417;
input n1419;
input n1421;
input n1426;
input n1428;
input n1431;
input n1433;
input n1435;
input n1439;
input n1441;
input n1444;
input n1447;
input n1451;
input n1453;
input n1456;
input n1458;
input n1459;
input n1467;
input n1472;
input n1476;
input n1480;
input n1484;
input n1489;
input n1491;
input n1494;
input n1496;
input n1498;
input n1502;
input n1504;
input n1507;
input n1510;
input n1514;
input n1518;
input n1523;
input n1527;
input n1528;
input n1538;
input n1540;
input n1542;
input n1544;
input n1546;
input n1552;
input n1554;
input n1556;
input n1558;
input n1563;
input n1564;
input n1567;
input n1570;
input n1573;
input n1578;
input n1581;
input n1584;
input n1587;
input n1588;
input n1595;
input n1596;
input n1599;
input n1602;
input n1605;
input n1610;
input n1613;
input n1616;
input n1619;
input n1624;
input n1626;
input n1629;
input n1633;
input n1635;
input n1640;
input n1642;
input n1648;
input n1651;
input n1652;
input n1662;
input n1664;
input n1666;
input n1668;
input n1670;
input n1673;
input n1675;
input n1681;
input n1683;
input n1685;
input n1687;
input n1689;
input n1694;
input n1697;
input n1699;
input n1701;
input n1704;
input n1706;
input n1707;
input n1714;
input n1715;
input n1718;
input n1721;
input n1724;
input n1729;
input n1732;
input n1735;
input n1738;
input n1743;
input n1745;
input n1747;
input n1749;
input n1751;
input n1756;
input n1758;
input n1764;
input n1766;
input n1767;
input n1777;
input n1779;
input n1781;
input n1783;
input n1785;
input n1791;
input n1793;
input n1795;
input n1797;
input n1802;
input n1803;
input n1806;
input n1809;
input n1812;
input n1817;
input n1820;
input n1823;
input n1826;
input n1827;
input n1834;
input n1835;
input n1838;
input n1841;
input n1844;
input n1849;
input n1852;
input n1855;
input n1858;
input n1863;
input n1865;
input n1868;
input n1872;
input n1874;
input n1879;
input n1881;
input n1887;
input n1890;
input n1891;
input n1901;
input n1903;
input n1905;
input n1907;
input n1909;
input n1915;
input n1917;
input n1919;
input n1921;
input n1926;
input n1927;
input n1930;
input n1933;
input n1936;
input n1941;
input n1944;
input n1947;
input n1950;
input n1951;
input n1958;
input n1959;
input n1962;
input n1965;
input n1968;
input n1973;
input n1976;
input n1979;
input n1982;
input n1987;
input n1989;
input n1992;
input n1996;
input n1998;
input n2003;
input n2005;
input n2008;
input n2013;
input n2014;
input n2023;
input n2025;
input n2028;
input n2030;
input n2032;
input n2036;
input n2038;
input n2042;
input n2044;
input n2049;
input n2050;
input n2053;
input n2056;
input n2059;
input n2064;
input n2067;
input n2070;
input n2073;
input n2074;
input n2081;
input n2082;
input n2085;
input n2088;
input n2091;
input n2096;
input n2099;
input n2102;
input n2105;
input n2111;
input n2113;
input n2115;
input n2117;
input n2119;
input n2128;
input n2130;
input n2132;
input n2134;
input n2135;
input n2144;
input n2146;
input n2148;
input n2150;
input n2152;
input n2157;
input n2160;
input n2162;
input n2164;
input n2169;
input n2170;
input n2173;
input n2176;
input n2179;
input n2184;
input n2187;
input n2190;
input n2193;
input n2194;
input n2201;
input n2202;
input n2205;
input n2208;
input n2211;
input n2216;
input n2219;
input n2222;
input n2225;
input n2230;
input n2232;
input n2235;
input n2239;
input n2241;
input n2246;
input n2248;
input n2251;
input n2256;
input n2257;
input n2273;
input n2275;
input n2285;
input n2287;
input n2289;
input n2291;
input n2293;
input n2298;
input n2301;
input n2303;
input n2305;
input n2308;
input n2311;
input n2313;
input n2315;
input n2317;
input n2320;
input n2322;
input n2325;
input n2327;
input n2328;
input n2335;
input n2337;
input n2339;
input n2341;
input n2343;
input n2349;
input n2351;
input n2353;
input n2355;
input n2357;
input n2362;
input n2365;
input n2367;
input n2369;
input n2372;
input n2374;
input n2377;
input n2379;
input n2380;
input n2391;
input n2393;
input n2395;
input n2397;
input n2399;
input n2404;
input n2407;
input n2409;
input n2411;
input n2414;
input n2418;
input n2420;
input n2422;
input n2424;
input n2427;
input n2429;
input n2432;
input n2434;
input n2435;
input n2442;
input n2444;
input n2449;
input n2451;
input n2454;
input n2459;
input n2461;
input n2467;
input n2470;
input n2475;
input n2476;
input n2479;
input n2482;
input n2485;
input n2490;
input n2493;
input n2496;
input n2499;
input n2500;
input n2508;
input n2512;
input n2515;
input n2517;
input n2519;
input n2524;
input n2526;
input n2529;
input n2531;
input n2533;
input n2537;
input n2539;
input n2542;
input n2545;
input n2548;
input n2550;
input n2553;
input n2555;
input n2556;
input n2561;
input n2564;
input n2567;
input n2569;
input n2571;
input n2577;
input n2579;
input n2581;
input n2583;
input n2585;
input n2587;
input n2594;
input n2596;
input n2598;
input n2600;
input n2602;
input n2605;
input n2607;
input n2608;
input n2618;
input n2620;
input n2625;
input n2627;
input n2630;
input n2635;
input n2637;
input n2643;
input n2646;
input n2651;
input n2652;
input n2655;
input n2658;
input n2661;
input n2666;
input n2669;
input n2672;
input n2675;
input n2676;
input n2683;
input n2685;
input n2687;
input n2689;
input n2691;
input n2696;
input n2698;
input n2704;
input n2706;
input n2711;
input n2712;
input n2715;
input n2718;
input n2721;
input n2726;
input n2729;
input n2732;
input n2735;
input n2736;
input n2746;
input n2748;
input n2753;
input n2755;
input n2758;
input n2763;
input n2765;
input n2771;
input n2774;
input n2779;
input n2780;
input n2783;
input n2786;
input n2789;
input n2794;
input n2797;
input n2800;
input n2803;
input n2804;
input n2810;
input n2812;
input n2815;
input n2817;
input n2819;
input n2823;
input n2825;
input n2829;
input n2831;
input n2836;
input n2837;
input n2840;
input n2843;
input n2846;
input n2851;
input n2854;
input n2857;
input n2860;
input n2861;
input n2871;
input n2873;
input n2875;
input n2877;
input n2879;
input n2885;
input n2887;
input n2889;
input n2891;
input n2896;
input n2897;
input n2900;
input n2903;
input n2906;
input n2911;
input n2914;
input n2917;
input n2920;
input n2921;
input n2928;
input n2930;
input n2932;
input n2934;
input n2936;
input n2941;
input n2944;
input n2946;
input n2948;
input n2953;
input n2954;
input n2957;
input n2960;
input n2963;
input n2968;
input n2971;
input n2974;
input n2977;
input n2978;
input n2988;
input n2989;
input n2992;
input n2995;
input n2998;
input n3003;
input n3005;
input n3009;
input n3011;
input n3016;
input n3017;
input n3020;
input n3023;
input n3026;
input n3031;
input n3034;
input n3037;
input n3040;
input n3041;
input n3051;
input n3053;
input n3055;
input n3057;
input n3059;
input n3066;
input n3068;
input n3070;
input n3072;
input n3077;
input n3078;
input n3081;
input n3084;
input n3087;
input n3092;
input n3095;
input n3098;
input n3101;
input n3102;
input n3112;
input n3114;
input n3117;
input n3119;
input n3121;
input n3126;
input n3128;
input n3132;
input n3134;
input n3139;
input n3140;
input n3143;
input n3146;
input n3149;
input n3154;
input n3157;
input n3160;
input n3163;
input n3164;
input n3171;
input n3173;
input n3176;
input n3180;
input n3182;
input n3187;
input n3189;
input n3192;
input n3197;
input n3202;
input n3203;
input n3206;
input n3209;
input n3212;
input n3217;
input n3220;
input n3223;
input n3226;
input n3227;
input n3241;
input n3243;
input n3263;
input n3264;
input n3267;
input n3270;
input n3273;
input n3278;
input n3281;
input n3284;
input n3287;
input n3288;
input n3291;
input n3296;
input n3298;
input n3301;
input n3303;
input n3305;
input n3311;
input n3313;
input n3317;
input n3319;
input n3331;
input n3332;
input n3335;
input n3338;
input n3341;
input n3346;
input n3349;
input n3352;
input n3355;
input n3356;
input n3366;
input n3368;
input n3370;
input n3372;
input n3374;
input n3380;
input n3382;
input n3384;
input n3386;
input n3387;
input n3397;
input n3399;
input n3402;
input n3404;
input n3421;
input n3422;
input n3425;
input n3428;
input n3431;
input n3436;
input n3439;
input n3442;
input n3445;
input n3446;
input n3450;
input n3457;
input n3459;
input n3461;
input n3463;
input n3465;
input n3471;
input n3474;
input n3476;
input n3478;
input n3488;
input n3489;
input n3492;
input n3495;
input n3498;
input n3503;
input n3506;
input n3509;
input n3512;
input n3513;
input n3520;
input n3522;
input n3525;
input n3527;
input n3529;
input n3535;
input n3537;
input n3541;
input n3543;
input n3545;
input n3557;
input n3558;
input n3561;
input n3564;
input n3567;
input n3572;
input n3575;
input n3578;
input n3581;
input n3582;
input n3589;
input n3591;
input n3596;
input n3598;
input n3601;
input n3608;
input n3611;
input n3613;
input n3615;
input n3616;
input n3630;
input n3631;
input n3634;
input n3637;
input n3640;
input n3645;
input n3648;
input n3651;
input n3654;
input n3655;
input n3658;
input n3664;
input n3666;
input n3668;
input n3670;
input n3672;
input n3680;
input n3682;
input n3684;
input n3686;
input n3703;
input n3704;
input n3707;
input n3710;
input n3713;
input n3718;
input n3721;
input n3724;
input n3727;
input n3728;
input n3736;
input n3738;
input n3740;
input n3742;
input n3744;
input n3752;
input n3754;
input n3756;
input n3758;
input n3759;
input n3770;
input n3771;
input n3774;
input n3777;
input n3780;
input n3785;
input n3788;
input n3791;
input n3794;
input n3795;
input n3800;
input n3809;
input n3811;
input n3813;
input n3815;
input n3817;
input n3824;
input n3826;
input n3828;
input n3830;
input n4126;
input n4128;
input n4132;
input n4134;
input n4139;
input n4141;
input n4159;
input n4161;
input n4167;
input n4169;
input n4184;
input n4186;
input n4252;
input n4254;
input n4266;
input n4268;
input n4286;
input n4288;
input n4307;
input n4313;
input n4329;
input n4336;
input n4355;
input n4362;
input n4368;
input n4370;
input n4795;
input n4797;
input n5728;
input n5729;
input n5732;
input n5733;
input n5740;
input n5741;
input n5744;
input n5745;
input n5779;
input n5780;
input n5785;
input n5786;
input n5823;
input n5824;
input n5827;
input n5828;
input n5856;
input n5857;
input n5861;
input n5862;
input n5893;
input n5894;
input n5897;
input n5898;
input n5935;
input n5936;
input n5940;
input n5941;
input n5983;
input n5984;
input n5987;
input n5988;
input n6019;
input n6020;
input n6023;
input n6024;
input n6062;
input n6063;
input n6066;
input n6067;
input n6098;
input n6099;
input n6102;
input n6103;
input n6140;
input n6141;
input n6144;
input n6145;
input n6165;
input n6166;
input n6171;
input n6172;
input n6201;
input n6202;
input n6205;
input n6206;
input n6237;
input n6238;
input n6243;
input n6244;
input n6273;
input n6274;
input n6277;
input n6278;
input n6437;
input n6440;
input n6456;
input n6460;
input n6470;
input n6481;
input n6485;
input n6489;
input n6501;
input n6511;
input n6514;
input n6516;
input n6520;
input n6522;
input n6536;
input n6538;
input n6550;
input n6560;
input n6563;
input n6565;
input n6569;
input n6571;
input n6585;
input n6587;
input n6601;
input n6609;
input n6612;
input n6614;
input n6630;
input n6632;
input n6635;
input n6637;
input n6652;
input n6663;
input n6666;
input n6668;
input n6674;
input n6689;
input n6691;
input n6693;
input n6705;
input n6715;
input n6718;
input n6720;
input n6736;
input n6738;
input n6741;
input n6743;
input n6758;
input n6768;
input n6771;
input n6773;
input n6779;
input n6794;
input n6796;
input n6798;
input n6815;
input n6817;
input n6819;
input n6829;
input n6850;
input n6852;
input n6855;
input n6857;
input n7035;
input n7038;
input n7151;
input n7154;
input n7245;
input n7248;
input n7373;
input n7376;
input n7630;
input n7633;
input n7649;
input n7652;
input n7783;
input n7786;
input n7892;
input n7895;
input n8006;
input n8016;
input n8019;
input n8021;
input n8023;
input n8027;
input n8030;
input n8032;
input n8034;
input n8038;
input n8041;
input n8043;
input n8045;
input n8049;
input n8052;
input n8054;
input n8056;
input n8064;
input n8067;
input n8069;
input n8071;
input n8075;
input n8078;
input n8080;
input n8082;
input n8086;
input n8089;
input n8091;
input n8093;
input n8097;
input n8100;
input n8102;
input n8104;
input n8147;
input n8174;
input n8189;
input n8204;
input n8219;
input n8234;
input n8253;
input n8331;
input n8342;
input n8362;
input n8377;
input n8392;
input n8412;
input n8427;
input n8436;
input n8531;
input n8544;
input n8550;
input n8568;
input n8588;
input n8598;
input n8612;
input n8664;
input n8671;
input n8690;
input n8721;
input n8782;
input n8796;
input n8806;
input n8826;
input n8840;
input n9996;
input n9999;
input n10008;
input n10011;
input n10030;
input n10039;
input n10054;
input n10059;
input n10081;
input n10083;
input n10086;
input n10088;
input n10099;
input n10101;
input n10104;
input n10106;
input n10116;
input n10118;
input n10121;
input n10123;
input n10134;
input n10141;
input n10142;
input n10143;
input n10144;
input n10152;
input n10153;
input n10154;
input n10155;
input n10171;
input n10176;
input n10187;
input n10192;
input n10199;
input n10202;
input n10204;
input n10247;
input n10248;
input n10249;
input n10250;
input n10253;
input n10280;
input n10282;
input n10291;
input n10293;
input n10295;
input n10305;
input n10308;
input n10315;
input n10318;
input n10323;
input n10330;
input n10343;
input n10344;
input n10363;
input n10404;
input n10405;
input n10430;
input n10434;
input n10437;
input n10448;
input n10451;
input n10453;
input n10456;
input n10461;
input n10467;
input n10473;
input n10476;
input n10483;
input n10487;
input n10492;
input n10498;
input n10502;
input n10540;
input n10543;
input n10546;
input n10548;
input n10558;
input n10560;
input n10563;
input n10565;
input n10574;
input n10576;
input n10579;
input n10581;
input n10590;
input n10592;
input n10595;
input n10597;
input n10606;
input n10608;
input n10611;
input n10613;
input n10623;
input n10626;
input n10628;
input n10635;
input n10637;
input n10643;
input n10649;
input n10652;
input n10661;
input n10680;
input n10682;
input n10687;
input n10689;
input n10691;
input n10700;
input n10703;
input n10705;
input n10707;
input n10709;
input n10711;
input n10715;
input n10716;
input n10729;
input n10747;
input n10748;
input n10771;
input n10775;
input n10778;
input n10789;
input n10792;
input n10794;
input n10799;
input n10802;
input n10809;
input n10817;
input n10821;
input n10828;
input n10831;
input n10836;
input n10842;
input n10846;
input n10883;
input n10886;
input n10889;
input n10891;
input n10901;
input n10903;
input n10906;
input n10908;
input n10917;
input n10919;
input n10922;
input n10924;
input n10933;
input n10935;
input n10938;
input n10940;
input n10949;
input n10951;
input n10954;
input n10956;
input n10966;
input n10969;
input n10971;
input n10975;
input n10980;
input n10986;
input n10992;
input n10995;
input n11004;
input n11023;
input n11025;
input n11030;
input n11032;
input n11034;
input n11043;
input n11046;
input n11048;
input n11050;
input n11052;
input n11054;
input n11058;
input n11059;
input n11072;
input n11090;
input n11091;
input n11114;
input n11117;
input n11119;
input n11130;
input n11133;
input n11135;
input n11139;
input n11142;
input n11146;
input n11152;
input n11156;
input n11167;
input n11171;
input n11175;
input n11181;
input n11185;
input n11223;
input n11226;
input n11229;
input n11231;
input n11241;
input n11243;
input n11246;
input n11248;
input n11257;
input n11259;
input n11262;
input n11264;
input n11273;
input n11275;
input n11278;
input n11280;
input n11289;
input n11291;
input n11294;
input n11296;
input n11306;
input n11309;
input n11311;
input n11314;
input n11319;
input n11325;
input n11334;
input n11337;
input n11346;
input n11365;
input n11367;
input n11372;
input n11374;
input n11376;
input n11385;
input n11388;
input n11390;
input n11392;
input n11394;
input n11396;
input n11400;
input n11401;
input n11414;
input n11432;
input n11433;
input n11456;
input n11459;
input n11461;
input n11472;
input n11475;
input n11477;
input n11481;
input n11484;
input n11488;
input n11494;
input n11498;
input n11511;
input n11515;
input n11519;
input n11525;
input n11529;
input n11567;
input n11570;
input n11573;
input n11575;
input n11585;
input n11587;
input n11590;
input n11592;
input n11601;
input n11603;
input n11606;
input n11608;
input n11617;
input n11619;
input n11622;
input n11624;
input n11633;
input n11635;
input n11638;
input n11640;
input n11650;
input n11653;
input n11655;
input n11659;
input n11662;
input n11666;
input n11672;
input n11676;
input n11689;
input n11708;
input n11710;
input n11715;
input n11717;
input n11719;
input n11728;
input n11731;
input n11733;
input n11735;
input n11737;
input n11739;
input n11743;
input n11744;
input n11757;
input n11775;
input n11776;
input n11798;
input n11800;
input n11802;
input n11813;
input n11816;
input n11818;
input n11822;
input n11829;
input n11832;
input n11835;
input n11840;
input n11849;
input n11851;
input n11853;
input n11862;
input n11866;
input n11901;
input n11904;
input n11907;
input n11909;
input n11919;
input n11921;
input n11924;
input n11926;
input n11935;
input n11937;
input n11940;
input n11942;
input n11951;
input n11953;
input n11956;
input n11958;
input n11967;
input n11969;
input n11972;
input n11974;
input n11984;
input n11988;
input n11991;
input n11996;
input n12000;
input n12003;
input n12005;
input n12011;
input n12028;
input n12047;
input n12049;
input n12054;
input n12056;
input n12058;
input n12067;
input n12070;
input n12072;
input n12074;
input n12076;
input n12078;
input n12082;
input n12083;
input n12096;
input n12114;
input n12115;
input n12137;
input n12139;
input n12141;
input n12152;
input n12155;
input n12157;
input n12162;
input n12165;
input n12170;
input n12172;
input n12174;
input n12189;
input n12191;
input n12193;
input n12203;
input n12207;
input n12248;
input n12251;
input n12254;
input n12256;
input n12266;
input n12268;
input n12271;
input n12273;
input n12282;
input n12284;
input n12287;
input n12289;
input n12298;
input n12300;
input n12303;
input n12305;
input n12314;
input n12316;
input n12319;
input n12321;
input n12331;
input n12334;
input n12336;
input n12341;
input n12345;
input n12349;
input n12354;
input n12356;
input n12370;
input n12389;
input n12391;
input n12396;
input n12398;
input n12400;
input n12409;
input n12412;
input n12414;
input n12416;
input n12418;
input n12420;
input n12424;
input n12425;
input n12438;
input n12456;
input n12457;
input n12479;
input n12481;
input n12483;
input n12493;
input n12495;
input n12497;
input n12502;
input n12506;
input n12509;
input n12515;
input n12517;
input n12529;
input n12531;
input n12533;
input n12539;
input n12543;
input n12582;
input n12585;
input n12588;
input n12590;
input n12600;
input n12602;
input n12605;
input n12607;
input n12616;
input n12618;
input n12621;
input n12623;
input n12632;
input n12634;
input n12637;
input n12639;
input n12648;
input n12650;
input n12653;
input n12655;
input n12664;
input n12666;
input n12668;
input n12673;
input n12677;
input n12681;
input n12687;
input n12691;
input n12704;
input n12723;
input n12725;
input n12730;
input n12732;
input n12734;
input n12743;
input n12746;
input n12748;
input n12750;
input n12752;
input n12754;
input n12758;
input n12759;
input n12772;
input n12790;
input n12791;
input n12813;
input n12815;
input n12817;
input n12827;
input n12829;
input n12831;
input n12835;
input n12837;
input n12842;
input n12846;
input n12854;
input n12865;
input n12867;
input n12869;
input n12875;
input n12879;
input n12951;
input n12985;
input n12988;
input n12990;
input n13004;
input n13017;
input n13042;
input n13045;
input n13047;
input n13050;
input n13063;
input n13086;
input n13089;
input n13091;
input n13094;
input n13107;
input n13130;
input n13133;
input n13135;
input n13140;
input n13153;
input n13176;
input n13179;
input n13181;
input n13185;
input n13198;
input n13220;
input n13222;
input n13224;
input n13230;
input n13261;
input n13274;
input n13276;
input n13278;
input n13282;
input n13298;
input n13308;
input n13311;
input n13313;
input n13317;
input n13464;
input n13480;
input n13483;
input n13486;
input n13488;
input n13503;
input n13513;
input n13525;
input n13530;
input n13550;
input n13553;
input n13556;
input n13559;
input n13561;
input n13566;
input n13568;
input n13579;
input n13584;
input n13602;
input n13605;
input n13608;
input n13611;
input n13613;
input n13618;
input n13620;
input n13631;
input n13636;
input n13659;
input n13662;
input n13665;
input n13668;
input n13670;
input n13679;
input n13681;
input n13692;
input n13697;
input n13715;
input n13718;
input n13721;
input n13724;
input n13726;
input n13741;
input n13746;
input n13765;
input n13768;
input n13771;
input n13774;
input n13776;
input n13791;
input n13796;
input n13814;
input n13817;
input n13820;
input n13823;
input n13825;
input n13840;
input n13845;
input n13877;
input n13880;
input n13883;
input n13886;
input n13888;
input n13904;
input n13909;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n19;
wire n22;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n112;
wire n113;
wire n114;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n217;
wire n220;
wire n221;
wire n222;
wire n225;
wire n226;
wire n228;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n360;
wire n361;
wire n363;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n453;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n570;
wire n571;
wire n573;
wire n575;
wire n577;
wire n578;
wire n579;
wire n581;
wire n582;
wire n584;
wire n586;
wire n588;
wire n589;
wire n590;
wire n592;
wire n593;
wire n595;
wire n597;
wire n599;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n661;
wire n662;
wire n664;
wire n666;
wire n668;
wire n669;
wire n670;
wire n672;
wire n673;
wire n675;
wire n677;
wire n679;
wire n680;
wire n681;
wire n683;
wire n684;
wire n686;
wire n688;
wire n690;
wire n691;
wire n692;
wire n694;
wire n695;
wire n697;
wire n699;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n734;
wire n735;
wire n737;
wire n739;
wire n741;
wire n742;
wire n743;
wire n745;
wire n746;
wire n748;
wire n750;
wire n752;
wire n753;
wire n754;
wire n756;
wire n757;
wire n759;
wire n761;
wire n763;
wire n764;
wire n765;
wire n767;
wire n768;
wire n770;
wire n772;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n804;
wire n805;
wire n806;
wire n808;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n830;
wire n832;
wire n834;
wire n836;
wire n838;
wire n840;
wire n842;
wire n844;
wire n846;
wire n848;
wire n850;
wire n852;
wire n854;
wire n856;
wire n858;
wire n860;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n938;
wire n940;
wire n942;
wire n944;
wire n946;
wire n948;
wire n950;
wire n952;
wire n954;
wire n956;
wire n958;
wire n960;
wire n962;
wire n964;
wire n966;
wire n967;
wire n968;
wire n970;
wire n972;
wire n974;
wire n976;
wire n978;
wire n980;
wire n982;
wire n984;
wire n986;
wire n988;
wire n990;
wire n992;
wire n994;
wire n996;
wire n998;
wire n1000;
wire n1001;
wire n1002;
wire n1004;
wire n1006;
wire n1008;
wire n1010;
wire n1012;
wire n1014;
wire n1016;
wire n1018;
wire n1020;
wire n1022;
wire n1024;
wire n1026;
wire n1028;
wire n1030;
wire n1032;
wire n1034;
wire n1035;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1115;
wire n1116;
wire n1118;
wire n1120;
wire n1122;
wire n1123;
wire n1124;
wire n1126;
wire n1127;
wire n1129;
wire n1131;
wire n1133;
wire n1134;
wire n1135;
wire n1137;
wire n1138;
wire n1140;
wire n1142;
wire n1144;
wire n1145;
wire n1146;
wire n1148;
wire n1149;
wire n1151;
wire n1153;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1197;
wire n1198;
wire n1199;
wire n1201;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1208;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1286;
wire n1287;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1298;
wire n1299;
wire n1300;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1308;
wire n1310;
wire n1312;
wire n1314;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1324;
wire n1325;
wire n1327;
wire n1329;
wire n1331;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1351;
wire n1352;
wire n1354;
wire n1355;
wire n1356;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1363;
wire n1364;
wire n1366;
wire n1367;
wire n1369;
wire n1370;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1377;
wire n1379;
wire n1381;
wire n1383;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1390;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1399;
wire n1400;
wire n1402;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1414;
wire n1416;
wire n1418;
wire n1420;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1427;
wire n1429;
wire n1430;
wire n1432;
wire n1434;
wire n1436;
wire n1437;
wire n1438;
wire n1440;
wire n1442;
wire n1443;
wire n1445;
wire n1446;
wire n1448;
wire n1449;
wire n1450;
wire n1452;
wire n1454;
wire n1455;
wire n1457;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1473;
wire n1474;
wire n1475;
wire n1477;
wire n1478;
wire n1479;
wire n1481;
wire n1482;
wire n1483;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1490;
wire n1492;
wire n1493;
wire n1495;
wire n1497;
wire n1499;
wire n1500;
wire n1501;
wire n1503;
wire n1505;
wire n1506;
wire n1508;
wire n1509;
wire n1511;
wire n1512;
wire n1513;
wire n1515;
wire n1516;
wire n1517;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1524;
wire n1525;
wire n1526;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1539;
wire n1541;
wire n1543;
wire n1545;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1553;
wire n1555;
wire n1557;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1565;
wire n1566;
wire n1568;
wire n1569;
wire n1571;
wire n1572;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1579;
wire n1580;
wire n1582;
wire n1583;
wire n1585;
wire n1586;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1597;
wire n1598;
wire n1600;
wire n1601;
wire n1603;
wire n1604;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1611;
wire n1612;
wire n1614;
wire n1615;
wire n1617;
wire n1618;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1625;
wire n1627;
wire n1628;
wire n1630;
wire n1631;
wire n1632;
wire n1634;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1641;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1649;
wire n1650;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1663;
wire n1665;
wire n1667;
wire n1669;
wire n1671;
wire n1672;
wire n1674;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1682;
wire n1684;
wire n1686;
wire n1688;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1695;
wire n1696;
wire n1698;
wire n1700;
wire n1702;
wire n1703;
wire n1705;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1716;
wire n1717;
wire n1719;
wire n1720;
wire n1722;
wire n1723;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1730;
wire n1731;
wire n1733;
wire n1734;
wire n1736;
wire n1737;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1744;
wire n1746;
wire n1748;
wire n1750;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1757;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1765;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1778;
wire n1780;
wire n1782;
wire n1784;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1792;
wire n1794;
wire n1796;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1804;
wire n1805;
wire n1807;
wire n1808;
wire n1810;
wire n1811;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1818;
wire n1819;
wire n1821;
wire n1822;
wire n1824;
wire n1825;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1836;
wire n1837;
wire n1839;
wire n1840;
wire n1842;
wire n1843;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1850;
wire n1851;
wire n1853;
wire n1854;
wire n1856;
wire n1857;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1864;
wire n1866;
wire n1867;
wire n1869;
wire n1870;
wire n1871;
wire n1873;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1880;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1888;
wire n1889;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1902;
wire n1904;
wire n1906;
wire n1908;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1916;
wire n1918;
wire n1920;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1928;
wire n1929;
wire n1931;
wire n1932;
wire n1934;
wire n1935;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1942;
wire n1943;
wire n1945;
wire n1946;
wire n1948;
wire n1949;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1960;
wire n1961;
wire n1963;
wire n1964;
wire n1966;
wire n1967;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1974;
wire n1975;
wire n1977;
wire n1978;
wire n1980;
wire n1981;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1988;
wire n1990;
wire n1991;
wire n1993;
wire n1994;
wire n1995;
wire n1997;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2004;
wire n2006;
wire n2007;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2024;
wire n2026;
wire n2027;
wire n2029;
wire n2031;
wire n2033;
wire n2034;
wire n2035;
wire n2037;
wire n2039;
wire n2040;
wire n2041;
wire n2043;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2051;
wire n2052;
wire n2054;
wire n2055;
wire n2057;
wire n2058;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2065;
wire n2066;
wire n2068;
wire n2069;
wire n2071;
wire n2072;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2083;
wire n2084;
wire n2086;
wire n2087;
wire n2089;
wire n2090;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2097;
wire n2098;
wire n2100;
wire n2101;
wire n2103;
wire n2104;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2112;
wire n2114;
wire n2116;
wire n2118;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2129;
wire n2131;
wire n2133;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2145;
wire n2147;
wire n2149;
wire n2151;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2158;
wire n2159;
wire n2161;
wire n2163;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2171;
wire n2172;
wire n2174;
wire n2175;
wire n2177;
wire n2178;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2185;
wire n2186;
wire n2188;
wire n2189;
wire n2191;
wire n2192;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2203;
wire n2204;
wire n2206;
wire n2207;
wire n2209;
wire n2210;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2217;
wire n2218;
wire n2220;
wire n2221;
wire n2223;
wire n2224;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2231;
wire n2233;
wire n2234;
wire n2236;
wire n2237;
wire n2238;
wire n2240;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2247;
wire n2249;
wire n2250;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2274;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2286;
wire n2288;
wire n2290;
wire n2292;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2299;
wire n2300;
wire n2302;
wire n2304;
wire n2306;
wire n2307;
wire n2309;
wire n2310;
wire n2312;
wire n2314;
wire n2316;
wire n2318;
wire n2319;
wire n2321;
wire n2323;
wire n2324;
wire n2326;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2336;
wire n2338;
wire n2340;
wire n2342;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2350;
wire n2352;
wire n2354;
wire n2356;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2363;
wire n2364;
wire n2366;
wire n2368;
wire n2370;
wire n2371;
wire n2373;
wire n2375;
wire n2376;
wire n2378;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2392;
wire n2394;
wire n2396;
wire n2398;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2405;
wire n2406;
wire n2408;
wire n2410;
wire n2412;
wire n2413;
wire n2415;
wire n2416;
wire n2417;
wire n2419;
wire n2421;
wire n2423;
wire n2425;
wire n2426;
wire n2428;
wire n2430;
wire n2431;
wire n2433;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2443;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2450;
wire n2452;
wire n2453;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2460;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2468;
wire n2469;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2477;
wire n2478;
wire n2480;
wire n2481;
wire n2483;
wire n2484;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2491;
wire n2492;
wire n2494;
wire n2495;
wire n2497;
wire n2498;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2509;
wire n2510;
wire n2511;
wire n2513;
wire n2514;
wire n2516;
wire n2518;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2525;
wire n2527;
wire n2528;
wire n2530;
wire n2532;
wire n2534;
wire n2535;
wire n2536;
wire n2538;
wire n2540;
wire n2541;
wire n2543;
wire n2544;
wire n2546;
wire n2547;
wire n2549;
wire n2551;
wire n2552;
wire n2554;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2562;
wire n2563;
wire n2565;
wire n2566;
wire n2568;
wire n2570;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2578;
wire n2580;
wire n2582;
wire n2584;
wire n2586;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2595;
wire n2597;
wire n2599;
wire n2601;
wire n2603;
wire n2604;
wire n2606;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2619;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2626;
wire n2628;
wire n2629;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2636;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2644;
wire n2645;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2653;
wire n2654;
wire n2656;
wire n2657;
wire n2659;
wire n2660;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2667;
wire n2668;
wire n2670;
wire n2671;
wire n2673;
wire n2674;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2684;
wire n2686;
wire n2688;
wire n2690;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2697;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2705;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2713;
wire n2714;
wire n2716;
wire n2717;
wire n2719;
wire n2720;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2727;
wire n2728;
wire n2730;
wire n2731;
wire n2733;
wire n2734;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2747;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2754;
wire n2756;
wire n2757;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2764;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2772;
wire n2773;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2781;
wire n2782;
wire n2784;
wire n2785;
wire n2787;
wire n2788;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2795;
wire n2796;
wire n2798;
wire n2799;
wire n2801;
wire n2802;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2811;
wire n2813;
wire n2814;
wire n2816;
wire n2818;
wire n2820;
wire n2821;
wire n2822;
wire n2824;
wire n2826;
wire n2827;
wire n2828;
wire n2830;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2838;
wire n2839;
wire n2841;
wire n2842;
wire n2844;
wire n2845;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2852;
wire n2853;
wire n2855;
wire n2856;
wire n2858;
wire n2859;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2872;
wire n2874;
wire n2876;
wire n2878;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2886;
wire n2888;
wire n2890;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2898;
wire n2899;
wire n2901;
wire n2902;
wire n2904;
wire n2905;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2912;
wire n2913;
wire n2915;
wire n2916;
wire n2918;
wire n2919;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2929;
wire n2931;
wire n2933;
wire n2935;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2942;
wire n2943;
wire n2945;
wire n2947;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2955;
wire n2956;
wire n2958;
wire n2959;
wire n2961;
wire n2962;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2969;
wire n2970;
wire n2972;
wire n2973;
wire n2975;
wire n2976;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2990;
wire n2991;
wire n2993;
wire n2994;
wire n2996;
wire n2997;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3004;
wire n3006;
wire n3007;
wire n3008;
wire n3010;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3018;
wire n3019;
wire n3021;
wire n3022;
wire n3024;
wire n3025;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3032;
wire n3033;
wire n3035;
wire n3036;
wire n3038;
wire n3039;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3052;
wire n3054;
wire n3056;
wire n3058;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3067;
wire n3069;
wire n3071;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3079;
wire n3080;
wire n3082;
wire n3083;
wire n3085;
wire n3086;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3093;
wire n3094;
wire n3096;
wire n3097;
wire n3099;
wire n3100;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3113;
wire n3115;
wire n3116;
wire n3118;
wire n3120;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3127;
wire n3129;
wire n3130;
wire n3131;
wire n3133;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3141;
wire n3142;
wire n3144;
wire n3145;
wire n3147;
wire n3148;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3155;
wire n3156;
wire n3158;
wire n3159;
wire n3161;
wire n3162;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3172;
wire n3174;
wire n3175;
wire n3177;
wire n3178;
wire n3179;
wire n3181;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3188;
wire n3190;
wire n3191;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3204;
wire n3205;
wire n3207;
wire n3208;
wire n3210;
wire n3211;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3218;
wire n3219;
wire n3221;
wire n3222;
wire n3224;
wire n3225;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3242;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3265;
wire n3266;
wire n3268;
wire n3269;
wire n3271;
wire n3272;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3279;
wire n3280;
wire n3282;
wire n3283;
wire n3285;
wire n3286;
wire n3289;
wire n3290;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3297;
wire n3299;
wire n3300;
wire n3302;
wire n3304;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3312;
wire n3314;
wire n3315;
wire n3316;
wire n3318;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3333;
wire n3334;
wire n3336;
wire n3337;
wire n3339;
wire n3340;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3347;
wire n3348;
wire n3350;
wire n3351;
wire n3353;
wire n3354;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3367;
wire n3369;
wire n3371;
wire n3373;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3381;
wire n3383;
wire n3385;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3398;
wire n3400;
wire n3401;
wire n3403;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3423;
wire n3424;
wire n3426;
wire n3427;
wire n3429;
wire n3430;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3437;
wire n3438;
wire n3440;
wire n3441;
wire n3443;
wire n3444;
wire n3447;
wire n3448;
wire n3449;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3458;
wire n3460;
wire n3462;
wire n3464;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3472;
wire n3473;
wire n3475;
wire n3477;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3490;
wire n3491;
wire n3493;
wire n3494;
wire n3496;
wire n3497;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3504;
wire n3505;
wire n3507;
wire n3508;
wire n3510;
wire n3511;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3521;
wire n3523;
wire n3524;
wire n3526;
wire n3528;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3536;
wire n3538;
wire n3539;
wire n3540;
wire n3542;
wire n3544;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3559;
wire n3560;
wire n3562;
wire n3563;
wire n3565;
wire n3566;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3573;
wire n3574;
wire n3576;
wire n3577;
wire n3579;
wire n3580;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3590;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3597;
wire n3599;
wire n3600;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3609;
wire n3610;
wire n3612;
wire n3614;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3632;
wire n3633;
wire n3635;
wire n3636;
wire n3638;
wire n3639;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3646;
wire n3647;
wire n3649;
wire n3650;
wire n3652;
wire n3653;
wire n3656;
wire n3657;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3665;
wire n3667;
wire n3669;
wire n3671;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3681;
wire n3683;
wire n3685;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3705;
wire n3706;
wire n3708;
wire n3709;
wire n3711;
wire n3712;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3719;
wire n3720;
wire n3722;
wire n3723;
wire n3725;
wire n3726;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3737;
wire n3739;
wire n3741;
wire n3743;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3753;
wire n3755;
wire n3757;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3772;
wire n3773;
wire n3775;
wire n3776;
wire n3778;
wire n3779;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3786;
wire n3787;
wire n3789;
wire n3790;
wire n3792;
wire n3793;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3810;
wire n3812;
wire n3814;
wire n3816;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3825;
wire n3827;
wire n3829;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4127;
wire n4129;
wire n4130;
wire n4131;
wire n4133;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4140;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4160;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4168;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4185;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4253;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4267;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4287;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4369;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4796;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5730;
wire n5731;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5742;
wire n5743;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5825;
wire n5826;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5858;
wire n5859;
wire n5860;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5895;
wire n5896;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5937;
wire n5938;
wire n5939;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5985;
wire n5986;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6021;
wire n6022;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6064;
wire n6065;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6100;
wire n6101;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6142;
wire n6143;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6203;
wire n6204;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6275;
wire n6276;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6438;
wire n6439;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6457;
wire n6458;
wire n6459;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6482;
wire n6483;
wire n6484;
wire n6486;
wire n6487;
wire n6488;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6512;
wire n6513;
wire n6515;
wire n6517;
wire n6518;
wire n6519;
wire n6521;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6537;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6561;
wire n6562;
wire n6564;
wire n6566;
wire n6567;
wire n6568;
wire n6570;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6586;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6610;
wire n6611;
wire n6613;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6631;
wire n6633;
wire n6634;
wire n6636;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6664;
wire n6665;
wire n6667;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6690;
wire n6692;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6716;
wire n6717;
wire n6719;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6737;
wire n6739;
wire n6740;
wire n6742;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6769;
wire n6770;
wire n6772;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6795;
wire n6797;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6816;
wire n6818;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6851;
wire n6853;
wire n6854;
wire n6856;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7036;
wire n7037;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7152;
wire n7153;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7246;
wire n7247;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7374;
wire n7375;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7631;
wire n7632;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7650;
wire n7651;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7784;
wire n7785;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7893;
wire n7894;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8017;
wire n8018;
wire n8020;
wire n8022;
wire n8024;
wire n8025;
wire n8026;
wire n8028;
wire n8029;
wire n8031;
wire n8033;
wire n8035;
wire n8036;
wire n8037;
wire n8039;
wire n8040;
wire n8042;
wire n8044;
wire n8046;
wire n8047;
wire n8048;
wire n8050;
wire n8051;
wire n8053;
wire n8055;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8065;
wire n8066;
wire n8068;
wire n8070;
wire n8072;
wire n8073;
wire n8074;
wire n8076;
wire n8077;
wire n8079;
wire n8081;
wire n8083;
wire n8084;
wire n8085;
wire n8087;
wire n8088;
wire n8090;
wire n8092;
wire n8094;
wire n8095;
wire n8096;
wire n8098;
wire n8099;
wire n8101;
wire n8103;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9997;
wire n9998;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10009;
wire n10010;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10082;
wire n10084;
wire n10085;
wire n10087;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10100;
wire n10102;
wire n10103;
wire n10105;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10117;
wire n10119;
wire n10120;
wire n10122;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10200;
wire n10201;
wire n10203;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10251;
wire n10252;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10281;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10292;
wire n10294;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10306;
wire n10307;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10316;
wire n10317;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10429;
wire n10431;
wire n10432;
wire n10433;
wire n10435;
wire n10436;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10449;
wire n10450;
wire n10452;
wire n10454;
wire n10455;
wire n10457;
wire n10458;
wire n10459;
wire n10460;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10468;
wire n10469;
wire n10470;
wire n10471;
wire n10472;
wire n10474;
wire n10475;
wire n10477;
wire n10478;
wire n10479;
wire n10480;
wire n10481;
wire n10482;
wire n10484;
wire n10485;
wire n10486;
wire n10488;
wire n10489;
wire n10490;
wire n10491;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10499;
wire n10500;
wire n10501;
wire n10503;
wire n10504;
wire n10505;
wire n10506;
wire n10507;
wire n10508;
wire n10509;
wire n10510;
wire n10511;
wire n10512;
wire n10513;
wire n10514;
wire n10515;
wire n10516;
wire n10517;
wire n10518;
wire n10519;
wire n10520;
wire n10521;
wire n10522;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10538;
wire n10539;
wire n10541;
wire n10542;
wire n10544;
wire n10545;
wire n10547;
wire n10549;
wire n10550;
wire n10551;
wire n10552;
wire n10553;
wire n10554;
wire n10555;
wire n10556;
wire n10557;
wire n10559;
wire n10561;
wire n10562;
wire n10564;
wire n10566;
wire n10567;
wire n10568;
wire n10569;
wire n10570;
wire n10571;
wire n10572;
wire n10573;
wire n10575;
wire n10577;
wire n10578;
wire n10580;
wire n10582;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10589;
wire n10591;
wire n10593;
wire n10594;
wire n10596;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10602;
wire n10603;
wire n10604;
wire n10605;
wire n10607;
wire n10609;
wire n10610;
wire n10612;
wire n10614;
wire n10615;
wire n10616;
wire n10617;
wire n10618;
wire n10619;
wire n10620;
wire n10621;
wire n10622;
wire n10624;
wire n10625;
wire n10627;
wire n10629;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10636;
wire n10638;
wire n10639;
wire n10640;
wire n10641;
wire n10642;
wire n10644;
wire n10645;
wire n10646;
wire n10647;
wire n10648;
wire n10650;
wire n10651;
wire n10653;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n10670;
wire n10671;
wire n10672;
wire n10673;
wire n10674;
wire n10675;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10681;
wire n10683;
wire n10684;
wire n10685;
wire n10686;
wire n10688;
wire n10690;
wire n10692;
wire n10693;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n10701;
wire n10702;
wire n10704;
wire n10706;
wire n10708;
wire n10710;
wire n10712;
wire n10713;
wire n10714;
wire n10717;
wire n10718;
wire n10719;
wire n10720;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10730;
wire n10731;
wire n10732;
wire n10733;
wire n10734;
wire n10735;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10766;
wire n10767;
wire n10768;
wire n10769;
wire n10770;
wire n10772;
wire n10773;
wire n10774;
wire n10776;
wire n10777;
wire n10779;
wire n10780;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10790;
wire n10791;
wire n10793;
wire n10795;
wire n10796;
wire n10797;
wire n10798;
wire n10800;
wire n10801;
wire n10803;
wire n10804;
wire n10805;
wire n10806;
wire n10807;
wire n10808;
wire n10810;
wire n10811;
wire n10812;
wire n10813;
wire n10814;
wire n10815;
wire n10816;
wire n10818;
wire n10819;
wire n10820;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10829;
wire n10830;
wire n10832;
wire n10833;
wire n10834;
wire n10835;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10843;
wire n10844;
wire n10845;
wire n10847;
wire n10848;
wire n10849;
wire n10850;
wire n10851;
wire n10852;
wire n10853;
wire n10854;
wire n10855;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n10869;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10877;
wire n10878;
wire n10879;
wire n10880;
wire n10881;
wire n10882;
wire n10884;
wire n10885;
wire n10887;
wire n10888;
wire n10890;
wire n10892;
wire n10893;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10899;
wire n10900;
wire n10902;
wire n10904;
wire n10905;
wire n10907;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10918;
wire n10920;
wire n10921;
wire n10923;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10930;
wire n10931;
wire n10932;
wire n10934;
wire n10936;
wire n10937;
wire n10939;
wire n10941;
wire n10942;
wire n10943;
wire n10944;
wire n10945;
wire n10946;
wire n10947;
wire n10948;
wire n10950;
wire n10952;
wire n10953;
wire n10955;
wire n10957;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10963;
wire n10964;
wire n10965;
wire n10967;
wire n10968;
wire n10970;
wire n10972;
wire n10973;
wire n10974;
wire n10976;
wire n10977;
wire n10978;
wire n10979;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10993;
wire n10994;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11005;
wire n11006;
wire n11007;
wire n11008;
wire n11009;
wire n11010;
wire n11011;
wire n11012;
wire n11013;
wire n11014;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n11020;
wire n11021;
wire n11022;
wire n11024;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11031;
wire n11033;
wire n11035;
wire n11036;
wire n11037;
wire n11038;
wire n11039;
wire n11040;
wire n11041;
wire n11042;
wire n11044;
wire n11045;
wire n11047;
wire n11049;
wire n11051;
wire n11053;
wire n11055;
wire n11056;
wire n11057;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11071;
wire n11073;
wire n11074;
wire n11075;
wire n11076;
wire n11077;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11087;
wire n11088;
wire n11089;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11097;
wire n11098;
wire n11099;
wire n11100;
wire n11101;
wire n11102;
wire n11103;
wire n11104;
wire n11105;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11115;
wire n11116;
wire n11118;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11131;
wire n11132;
wire n11134;
wire n11136;
wire n11137;
wire n11138;
wire n11140;
wire n11141;
wire n11143;
wire n11144;
wire n11145;
wire n11147;
wire n11148;
wire n11149;
wire n11150;
wire n11151;
wire n11153;
wire n11154;
wire n11155;
wire n11157;
wire n11158;
wire n11159;
wire n11160;
wire n11161;
wire n11162;
wire n11163;
wire n11164;
wire n11165;
wire n11166;
wire n11168;
wire n11169;
wire n11170;
wire n11172;
wire n11173;
wire n11174;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11180;
wire n11182;
wire n11183;
wire n11184;
wire n11186;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11224;
wire n11225;
wire n11227;
wire n11228;
wire n11230;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11239;
wire n11240;
wire n11242;
wire n11244;
wire n11245;
wire n11247;
wire n11249;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11258;
wire n11260;
wire n11261;
wire n11263;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11274;
wire n11276;
wire n11277;
wire n11279;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11290;
wire n11292;
wire n11293;
wire n11295;
wire n11297;
wire n11298;
wire n11299;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11307;
wire n11308;
wire n11310;
wire n11312;
wire n11313;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11335;
wire n11336;
wire n11338;
wire n11339;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11347;
wire n11348;
wire n11349;
wire n11350;
wire n11351;
wire n11352;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11364;
wire n11366;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11373;
wire n11375;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11386;
wire n11387;
wire n11389;
wire n11391;
wire n11393;
wire n11395;
wire n11397;
wire n11398;
wire n11399;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n11450;
wire n11451;
wire n11452;
wire n11453;
wire n11454;
wire n11455;
wire n11457;
wire n11458;
wire n11460;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11469;
wire n11470;
wire n11471;
wire n11473;
wire n11474;
wire n11476;
wire n11478;
wire n11479;
wire n11480;
wire n11482;
wire n11483;
wire n11485;
wire n11486;
wire n11487;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11493;
wire n11495;
wire n11496;
wire n11497;
wire n11499;
wire n11500;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11506;
wire n11507;
wire n11508;
wire n11509;
wire n11510;
wire n11512;
wire n11513;
wire n11514;
wire n11516;
wire n11517;
wire n11518;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11526;
wire n11527;
wire n11528;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11563;
wire n11564;
wire n11565;
wire n11566;
wire n11568;
wire n11569;
wire n11571;
wire n11572;
wire n11574;
wire n11576;
wire n11577;
wire n11578;
wire n11579;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11586;
wire n11588;
wire n11589;
wire n11591;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11597;
wire n11598;
wire n11599;
wire n11600;
wire n11602;
wire n11604;
wire n11605;
wire n11607;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11618;
wire n11620;
wire n11621;
wire n11623;
wire n11625;
wire n11626;
wire n11627;
wire n11628;
wire n11629;
wire n11630;
wire n11631;
wire n11632;
wire n11634;
wire n11636;
wire n11637;
wire n11639;
wire n11641;
wire n11642;
wire n11643;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11649;
wire n11651;
wire n11652;
wire n11654;
wire n11656;
wire n11657;
wire n11658;
wire n11660;
wire n11661;
wire n11663;
wire n11664;
wire n11665;
wire n11667;
wire n11668;
wire n11669;
wire n11670;
wire n11671;
wire n11673;
wire n11674;
wire n11675;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11709;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11716;
wire n11718;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11729;
wire n11730;
wire n11732;
wire n11734;
wire n11736;
wire n11738;
wire n11740;
wire n11741;
wire n11742;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11758;
wire n11759;
wire n11760;
wire n11761;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11766;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11771;
wire n11772;
wire n11773;
wire n11774;
wire n11777;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11789;
wire n11790;
wire n11791;
wire n11792;
wire n11793;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11799;
wire n11801;
wire n11803;
wire n11804;
wire n11805;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11814;
wire n11815;
wire n11817;
wire n11819;
wire n11820;
wire n11821;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11830;
wire n11831;
wire n11833;
wire n11834;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11850;
wire n11852;
wire n11854;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11863;
wire n11864;
wire n11865;
wire n11867;
wire n11868;
wire n11869;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11874;
wire n11875;
wire n11876;
wire n11877;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11887;
wire n11888;
wire n11889;
wire n11890;
wire n11891;
wire n11892;
wire n11893;
wire n11894;
wire n11895;
wire n11896;
wire n11897;
wire n11898;
wire n11899;
wire n11900;
wire n11902;
wire n11903;
wire n11905;
wire n11906;
wire n11908;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11920;
wire n11922;
wire n11923;
wire n11925;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11936;
wire n11938;
wire n11939;
wire n11941;
wire n11943;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11949;
wire n11950;
wire n11952;
wire n11954;
wire n11955;
wire n11957;
wire n11959;
wire n11960;
wire n11961;
wire n11962;
wire n11963;
wire n11964;
wire n11965;
wire n11966;
wire n11968;
wire n11970;
wire n11971;
wire n11973;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11985;
wire n11986;
wire n11987;
wire n11989;
wire n11990;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11997;
wire n11998;
wire n11999;
wire n12001;
wire n12002;
wire n12004;
wire n12006;
wire n12007;
wire n12008;
wire n12009;
wire n12010;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12024;
wire n12025;
wire n12026;
wire n12027;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12043;
wire n12044;
wire n12045;
wire n12046;
wire n12048;
wire n12050;
wire n12051;
wire n12052;
wire n12053;
wire n12055;
wire n12057;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12068;
wire n12069;
wire n12071;
wire n12073;
wire n12075;
wire n12077;
wire n12079;
wire n12080;
wire n12081;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12095;
wire n12097;
wire n12098;
wire n12099;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12122;
wire n12123;
wire n12124;
wire n12125;
wire n12126;
wire n12127;
wire n12128;
wire n12129;
wire n12130;
wire n12131;
wire n12132;
wire n12133;
wire n12134;
wire n12135;
wire n12136;
wire n12138;
wire n12140;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12146;
wire n12147;
wire n12148;
wire n12149;
wire n12150;
wire n12151;
wire n12153;
wire n12154;
wire n12156;
wire n12158;
wire n12159;
wire n12160;
wire n12161;
wire n12163;
wire n12164;
wire n12166;
wire n12167;
wire n12168;
wire n12169;
wire n12171;
wire n12173;
wire n12175;
wire n12176;
wire n12177;
wire n12178;
wire n12179;
wire n12180;
wire n12181;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12190;
wire n12192;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n12200;
wire n12201;
wire n12202;
wire n12204;
wire n12205;
wire n12206;
wire n12208;
wire n12209;
wire n12210;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12228;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12233;
wire n12234;
wire n12235;
wire n12236;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12244;
wire n12245;
wire n12246;
wire n12247;
wire n12249;
wire n12250;
wire n12252;
wire n12253;
wire n12255;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12267;
wire n12269;
wire n12270;
wire n12272;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12281;
wire n12283;
wire n12285;
wire n12286;
wire n12288;
wire n12290;
wire n12291;
wire n12292;
wire n12293;
wire n12294;
wire n12295;
wire n12296;
wire n12297;
wire n12299;
wire n12301;
wire n12302;
wire n12304;
wire n12306;
wire n12307;
wire n12308;
wire n12309;
wire n12310;
wire n12311;
wire n12312;
wire n12313;
wire n12315;
wire n12317;
wire n12318;
wire n12320;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12326;
wire n12327;
wire n12328;
wire n12329;
wire n12330;
wire n12332;
wire n12333;
wire n12335;
wire n12337;
wire n12338;
wire n12339;
wire n12340;
wire n12342;
wire n12343;
wire n12344;
wire n12346;
wire n12347;
wire n12348;
wire n12350;
wire n12351;
wire n12352;
wire n12353;
wire n12355;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12390;
wire n12392;
wire n12393;
wire n12394;
wire n12395;
wire n12397;
wire n12399;
wire n12401;
wire n12402;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12410;
wire n12411;
wire n12413;
wire n12415;
wire n12417;
wire n12419;
wire n12421;
wire n12422;
wire n12423;
wire n12426;
wire n12427;
wire n12428;
wire n12429;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12439;
wire n12440;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12455;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12480;
wire n12482;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12494;
wire n12496;
wire n12498;
wire n12499;
wire n12500;
wire n12501;
wire n12503;
wire n12504;
wire n12505;
wire n12507;
wire n12508;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12516;
wire n12518;
wire n12519;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12527;
wire n12528;
wire n12530;
wire n12532;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12540;
wire n12541;
wire n12542;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12558;
wire n12559;
wire n12560;
wire n12561;
wire n12562;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12583;
wire n12584;
wire n12586;
wire n12587;
wire n12589;
wire n12591;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n12601;
wire n12603;
wire n12604;
wire n12606;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12617;
wire n12619;
wire n12620;
wire n12622;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12633;
wire n12635;
wire n12636;
wire n12638;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12649;
wire n12651;
wire n12652;
wire n12654;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12665;
wire n12667;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12674;
wire n12675;
wire n12676;
wire n12678;
wire n12679;
wire n12680;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12688;
wire n12689;
wire n12690;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12724;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12731;
wire n12733;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12744;
wire n12745;
wire n12747;
wire n12749;
wire n12751;
wire n12753;
wire n12755;
wire n12756;
wire n12757;
wire n12760;
wire n12761;
wire n12762;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12777;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12814;
wire n12816;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12825;
wire n12826;
wire n12828;
wire n12830;
wire n12832;
wire n12833;
wire n12834;
wire n12836;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12843;
wire n12844;
wire n12845;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12866;
wire n12868;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12874;
wire n12876;
wire n12877;
wire n12878;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12946;
wire n12947;
wire n12948;
wire n12949;
wire n12950;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12986;
wire n12987;
wire n12989;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13043;
wire n13044;
wire n13046;
wire n13048;
wire n13049;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13087;
wire n13088;
wire n13090;
wire n13092;
wire n13093;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n13100;
wire n13101;
wire n13102;
wire n13103;
wire n13104;
wire n13105;
wire n13106;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13131;
wire n13132;
wire n13134;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n13150;
wire n13151;
wire n13152;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13177;
wire n13178;
wire n13180;
wire n13182;
wire n13183;
wire n13184;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13221;
wire n13223;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13275;
wire n13277;
wire n13279;
wire n13280;
wire n13281;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13303;
wire n13304;
wire n13305;
wire n13306;
wire n13307;
wire n13309;
wire n13310;
wire n13312;
wire n13314;
wire n13315;
wire n13316;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13365;
wire n13366;
wire n13367;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13394;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13404;
wire n13405;
wire n13406;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13425;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n13481;
wire n13482;
wire n13484;
wire n13485;
wire n13487;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n13531;
wire n13532;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13551;
wire n13552;
wire n13554;
wire n13555;
wire n13557;
wire n13558;
wire n13560;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13567;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13597;
wire n13598;
wire n13599;
wire n13600;
wire n13601;
wire n13603;
wire n13604;
wire n13606;
wire n13607;
wire n13609;
wire n13610;
wire n13612;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13619;
wire n13621;
wire n13622;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n13630;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13660;
wire n13661;
wire n13663;
wire n13664;
wire n13666;
wire n13667;
wire n13669;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13680;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13716;
wire n13717;
wire n13719;
wire n13720;
wire n13722;
wire n13723;
wire n13725;
wire n13727;
wire n13728;
wire n13729;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13766;
wire n13767;
wire n13769;
wire n13770;
wire n13772;
wire n13773;
wire n13775;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13815;
wire n13816;
wire n13818;
wire n13819;
wire n13821;
wire n13822;
wire n13824;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13831;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13851;
wire n13852;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13868;
wire n13869;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13878;
wire n13879;
wire n13881;
wire n13882;
wire n13884;
wire n13885;
wire n13887;
wire n13889;
wire n13890;
wire n13891;
wire n13892;
wire n13893;
wire n13894;
wire n13895;
wire n13896;
wire n13897;
wire n13898;
wire n13899;
wire n13900;
wire n13901;
wire n13902;
wire n13903;
wire n13905;
wire n13906;
wire n13907;
wire n13908;
wire n13910;
wire n13911;
wire n13912;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13919;
wire n13920;
wire n13921;
wire n13922;
wire n13923;
wire n13924;
wire n13925;
wire n13926;
wire n13927;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13934;
wire n13935;
wire n13936;
wire n13937;
wire n13938;
wire n13939;
wire n13940;
wire n13941;
wire n13942;
wire n13943;
wire n13944;
wire n13945;
wire n13946;
wire n13947;
wire n13948;
wire n13949;
wire n13950;
wire n13951;
wire n13952;
wire n13953;
wire n13954;
wire n13955;
wire n13956;
wire n13957;
wire n13958;
wire n13959;
wire n13960;
wire n13961;
wire n13962;
wire n13963;
wire n13964;
wire n13965;
wire n13966;
wire n13967;
wire n13968;
wire n13969;
wire n13970;
wire n13971;
wire n13972;
wire n13973;
wire n13974;
wire n13975;
wire n13976;
wire n13977;
wire n13978;
wire n13979;
wire n13980;
wire n13981;
wire n13982;
wire n13983;
wire n13984;
wire n13985;
wire n13986;
wire n13987;
wire n13988;
wire n13989;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13997;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14002;
wire n14003;
wire n14004;
wire n14005;
wire n14006;
wire n14007;
wire n14008;
wire n14009;
wire n14010;
wire n14011;
wire n14012;
wire n14013;
wire n14014;
wire n14015;
wire n14016;
wire n14017;
wire n14018;
wire n14019;
wire n14020;
wire n14021;
wire n14022;
wire n14023;
wire n14024;
wire n14025;
wire n14026;
wire n14027;
wire n14028;
wire n14029;
wire n14030;
wire n14031;
wire n14032;
wire n14033;
wire n14034;
wire n14035;
wire n14036;
wire n14037;
wire n14038;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14043;
wire n14044;
wire n14045;
wire n14046;
wire n14047;
wire n14048;
wire n14049;
wire n14050;
wire n14051;
wire n14052;
wire n14053;
wire n14054;
wire n14055;
wire n14056;
wire n14057;
wire n14058;
wire n14059;
wire n14060;
wire n14061;
wire n14062;
wire n14063;
wire n14064;
wire n14065;
wire n14066;
wire n14067;
wire n14068;
wire n14069;
wire n14070;
wire n14071;
wire n14072;
wire n14073;
wire n14074;
wire n14075;
wire n14076;
wire n14077;
wire n14078;
wire n14079;
wire n14080;
wire n14081;
wire n14082;
wire n14083;
wire n14084;
wire n14085;
wire n14086;
wire n14087;
wire n14088;
wire n14089;
wire n14090;
wire n14091;
wire n14092;
wire n14093;
wire n14094;
wire n14095;
wire n14096;
wire n14097;
wire n14098;
wire n14099;
wire n14100;
wire n14101;
wire n14102;
wire n14103;
wire n14104;
wire n14105;
wire n14106;
wire n14107;
wire n14108;
wire n14109;
wire n14110;
wire n14111;
wire n14112;
wire n14113;
wire n14114;
wire n14115;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14121;
wire n14122;
wire n14123;
wire n14124;
wire n14125;
wire n14126;
wire n14127;
wire n14128;
wire n14129;
wire n14130;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14135;
wire n14136;
wire n14137;
wire n14138;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14146;
wire n14147;
wire n14148;
wire n14149;
wire n14150;
wire n14151;
wire n14152;
wire n14153;
wire n14154;
wire n14155;
wire n14156;
wire n14157;
wire n14158;
wire n14159;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14164;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14170;
wire n14171;
wire n14172;
wire n14173;
wire n14174;
wire n14175;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14192;
wire n14193;
wire n14194;
wire n14195;
wire n14196;
wire n14197;
wire n14198;
wire n14199;
wire n14200;
wire n14201;
wire n14202;
wire n14203;
wire n14204;
wire n14205;
wire n14206;
wire n14207;
wire n14208;
wire n14209;
wire n14210;
wire n14211;
wire n14212;
wire n14213;
wire n14214;
wire n14215;
wire n14216;
wire n14217;
wire n14218;
wire n14219;
wire n14220;
wire n14221;
wire n14222;
wire n14223;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14233;
wire n14234;
wire n14235;
wire n14236;
wire n14237;
wire n14238;
wire n14239;
wire n14240;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n14250;
wire n14251;
wire n14252;
wire n14253;
wire n14254;
wire n14255;
wire n14256;
wire n14257;
wire n14258;
wire n14259;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14265;
wire n14266;
wire n14267;
wire n14268;
wire n14269;
wire n14270;
wire n14271;
wire n14272;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14278;
wire n14279;
wire n14280;
wire n14281;
wire n14282;
wire n14283;
wire n14284;
wire n14285;
wire n14286;
wire n14287;
wire n14288;
wire n14289;
wire n14290;
wire n14291;
wire n14292;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n14300;
wire n14301;
wire n14302;
wire n14303;
wire n14304;
wire n14305;
wire n14306;
wire n14307;
wire n14308;
wire n14309;
wire n14310;
wire n14311;
wire n14312;
wire n14313;
wire n14314;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14320;
wire n14321;
wire n14322;
wire n14323;
wire n14324;
wire n14325;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14332;
wire n14333;
wire n14334;
wire n14335;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14341;
wire n14342;
wire n14343;
wire n14344;
wire n14345;
wire n14346;
wire n14347;
wire n14348;
wire n14349;
wire n14350;
wire n14351;
wire n14352;
wire n14353;
wire n14354;
wire n14355;
wire n14356;
wire n14357;
wire n14358;
wire n14359;
wire n14360;
wire n14361;
wire n14362;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14369;
wire n14370;
wire n14371;
wire n14372;
wire n14373;
wire n14374;
wire n14375;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14390;
wire n14391;
wire n14392;
wire n14393;
wire n14394;
wire n14395;
wire n14396;
wire n14397;
wire n14398;
wire n14399;
wire n14400;
wire n14401;
wire n14402;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14407;
wire n14408;
wire n14409;
wire n14410;
wire n14411;
wire n14412;
wire n14413;
wire n14414;
wire n14415;
wire n14416;
wire n14417;
wire n14418;
wire n14419;
wire n14420;
wire n14421;
wire n14422;
wire n14423;
wire n14424;
wire n14425;
wire n14426;
wire n14427;
wire n14428;
wire n14429;
wire n14430;
wire n14431;
wire n14432;
wire n14433;
wire n14434;
wire n14435;
wire n14436;
wire n14437;
wire n14438;
wire n14439;
wire n14440;
wire n14441;
wire n14442;
wire n14443;
wire n14444;
wire n14445;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14453;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n14460;
wire n14461;
wire n14462;
wire n14463;
wire n14464;
wire n14465;
wire n14466;
wire n14467;
wire n14468;
wire n14469;
wire n14470;
wire n14471;
wire n14472;
wire n14473;
wire n14474;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14480;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14486;
wire n14487;
wire n14488;
wire n14489;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14501;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14507;
wire n14508;
wire n14509;
wire n14510;
wire n14511;
wire n14512;
wire n14513;
wire n14514;
wire n14515;
wire n14516;
wire n14517;
wire n14518;
wire n14519;
wire n14520;
wire n14521;
wire n14522;
wire n14523;
wire n14524;
wire n14525;
wire n14526;
wire n14527;
wire n14528;
wire n14529;
wire n14530;
wire n14531;
wire n14532;
wire n14533;
wire n14534;
wire n14535;
wire n14536;
wire n14537;
wire n14538;
wire n14539;
wire n14540;
wire n14541;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14546;
wire n14547;
wire n14548;
wire n14549;
wire n14550;
wire n14551;
wire n14552;
wire n14553;
wire n14554;
wire n14555;
wire n14556;
wire n14557;
wire n14558;
wire n14559;
wire n14560;
wire n14561;
wire n14562;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14568;
wire n14569;
wire n14570;
wire n14571;
wire n14572;
wire n14573;
wire n14574;
wire n14575;
wire n14576;
wire n14577;
wire n14578;
wire n14579;
wire n14580;
wire n14581;
wire n14582;
wire n14583;
wire n14584;
wire n14585;
wire n14586;
wire n14587;
wire n14588;
wire n14589;
wire n14590;
wire n14591;
wire n14592;
wire n14593;
wire n14594;
wire n14595;
wire n14596;
wire n14597;
wire n14598;
wire n14599;
wire n14600;
wire n14601;
wire n14602;
wire n14603;
wire n14604;
wire n14605;
wire n14606;
wire n14607;
wire n14608;
wire n14609;
wire n14610;
wire n14611;
wire n14612;
wire n14613;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14618;
wire n14619;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14624;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n14640;
wire n14641;
wire n14642;
wire n14643;
wire n14644;
wire n14645;
wire n14646;
wire n14647;
wire n14648;
wire n14649;
wire n14650;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14657;
wire n14658;
wire n14659;
wire n14660;
wire n14661;
wire n14662;
wire n14663;
wire n14664;
wire n14665;
wire n14666;
wire n14667;
wire n14668;
wire n14669;
wire n14670;
wire n14671;
wire n14672;
wire n14673;
wire n14674;
wire n14675;
wire n14676;
wire n14677;
wire n14678;
wire n14679;
wire n14680;
wire n14681;
wire n14682;
wire n14683;
wire n14684;
wire n14685;
wire n14686;
wire n14687;
wire n14688;
wire n14689;
wire n14690;
wire n14691;
wire n14692;
wire n14693;
wire n14694;
wire n14695;
wire n14696;
wire n14697;
wire n14698;
wire n14699;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14707;
xor (out,n0,n13935);
or (n0,n1,n1068);
and (n1,n2,n1067);
and (n2,n3,n1058);
nor (n3,n4,n812);
and (n4,n5,n804,n807);
and (n5,n6,n799,n803);
and (n6,n7,n652,n726);
wire s0n7,s1n7,notn7;
or (n7,s0n7,s1n7);
not(notn7,n651);
and (s0n7,notn7,1'b0);
and (s1n7,n651,n9);
wire s0n9,s1n9,notn9;
or (n9,s0n9,s1n9);
not(notn9,n651);
and (s0n9,notn9,n10);
and (s1n9,n651,n603);
wire s0n10,s1n10,notn10;
or (n10,s0n10,s1n10);
not(notn10,n601);
and (s0n10,notn10,1'b0);
and (s1n10,n601,n11);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n600);
and (s0n11,notn11,n12);
and (s1n11,n600,n591);
or (n12,n13,n567,n578,n589);
and (n13,n14,n37);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n31);
and (s0n14,notn14,n15);
and (s1n14,n31,n16);
or (n16,n17,n22,n26,n29);
and (n17,n18,n19);
nor (n19,n20,n21);
and (n22,n23,n24);
and (n24,n20,n25);
not (n25,n21);
and (n26,n27,n28);
nor (n28,n20,n25);
and (n29,n15,n30);
and (n30,n20,n21);
nor (n31,n32,n65);
nor (n32,n33,n52);
and (n33,n34,n51);
or (n34,n35,n40,n45,n48);
and (n35,n36,n37);
and (n37,n38,n39);
and (n40,n41,n42);
not (n42,n43);
nand (n43,n44,n39);
not (n44,n38);
and (n45,n46,n47);
nor (n47,n44,n39);
and (n48,n49,n50);
nor (n50,n38,n39);
nor (n52,n53,n61,n51);
and (n53,n54,n59);
nand (n54,n55,n57);
or (n55,n56,n49);
or (n57,n58,n41);
not (n58,n56);
not (n59,n60);
and (n61,n62,n60);
nand (n62,n63,n64);
or (n63,n56,n46);
or (n64,n58,n36);
nand (n65,n66,n75);
or (n66,n67,n69);
not (n67,n68);
not (n69,n70);
nand (n70,n71,n74);
nor (n71,n72,n73);
nand (n75,n76,n531);
nand (n76,n77,n523);
or (n77,n78,n447);
not (n78,n79);
or (n79,1'b0,n80,n367,n445);
and (n80,n81,n366);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n357);
and (s0n81,notn81,n82);
and (s1n81,n357,1'b0);
wire s0n82,s1n82,notn82;
or (n82,s0n82,s1n82);
not(notn82,n293);
and (s0n82,notn82,1'b0);
and (s1n82,n293,n83);
or (n83,n84,n267,n273,n279,n284,1'b0,1'b0,1'b0);
and (n84,n85,n93);
xnor (n85,n86,n87);
not (n87,n88);
nor (n88,n89,n92);
or (n89,n90,n91);
and (n93,n94,n236,n255,n263);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n127);
and (s0n94,notn94,n95);
and (s1n94,n127,1'b0);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n125);
and (s0n95,notn95,n96);
and (s1n95,n125,n123);
wire s0n96,s1n96,notn96;
or (n96,s0n96,s1n96);
not(notn96,n118);
and (s0n96,notn96,n97);
and (s1n96,n118,n112);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n111);
and (s0n97,notn97,n98);
and (s1n97,n111,1'b0);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n110);
and (s0n98,notn98,n99);
and (s1n98,n110,1'b1);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n109);
and (s0n99,notn99,n100);
and (s1n99,n109,1'b0);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n108);
and (s0n100,notn100,n101);
and (s1n100,n108,1'b1);
wire s0n101,s1n101,notn101;
or (n101,s0n101,s1n101);
not(notn101,n107);
and (s0n101,notn101,n102);
and (s1n101,n107,1'b0);
wire s0n102,s1n102,notn102;
or (n102,s0n102,s1n102);
not(notn102,n86);
and (s0n102,notn102,n103);
and (s1n102,n86,1'b1);
wire s0n103,s1n103,notn103;
or (n103,s0n103,s1n103);
not(notn103,n92);
and (s0n103,notn103,n104);
and (s1n103,n92,1'b0);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n90);
and (s0n104,notn104,n105);
and (s1n104,n90,1'b1);
not (n105,n91);
wire s0n112,s1n112,notn112;
or (n112,s0n112,s1n112);
not(notn112,n117);
and (s0n112,notn112,n113);
and (s1n112,n117,1'b0);
wire s0n113,s1n113,notn113;
or (n113,s0n113,s1n113);
not(notn113,n116);
and (s0n113,notn113,n114);
and (s1n113,n116,1'b1);
not (n114,n115);
or (n118,n119,n122);
or (n119,n117,n120);
not (n120,n121);
nor (n121,n116,n115);
not (n123,n124);
or (n125,n124,n126);
not (n127,n128);
or (n128,n129,n234);
or (n129,n130,n232);
or (n130,n131,n226);
or (n131,n132,n225);
or (n132,n133,n221);
or (n133,n134,n220);
or (n134,n135,n215);
or (n135,n136,n214);
or (n136,n137,n213);
or (n137,n138,n211);
or (n138,n139,n208);
or (n139,n140,n207);
or (n140,n141,n206);
or (n141,n142,n205);
or (n142,n143,n204);
or (n143,n144,n202);
or (n144,n145,n200);
or (n145,n146,n199);
or (n146,n147,n197);
or (n147,n148,n191);
or (n148,n149,n190);
or (n149,n150,n189);
or (n150,n151,n188);
or (n151,n152,n187);
or (n152,n153,n186);
or (n153,n154,n184);
or (n154,n155,n182);
or (n155,n156,n176);
or (n156,n157,n175);
or (n157,n158,n174);
or (n158,n159,n173);
or (n159,n160,n172);
or (n160,n161,n170);
or (n161,n162,n168);
nor (n162,n163,n164,n166,n167);
not (n164,n165);
nor (n168,n163,n164,n169,n167);
not (n169,n166);
and (n170,n163,n165,n166,n171);
not (n171,n167);
and (n172,n163,n164,n166,n171);
nor (n173,n163,n165,n169,n167);
and (n174,n163,n164,n166,n167);
and (n175,n163,n165,n166,n167);
nor (n176,n177,n179,n180,n181);
not (n177,n178);
nor (n182,n177,n183,n180,n181);
not (n183,n179);
and (n184,n177,n179,n180,n185);
not (n185,n181);
and (n186,n178,n179,n180,n185);
and (n187,n178,n183,n180,n185);
and (n188,n177,n183,n180,n181);
and (n189,n178,n183,n180,n181);
and (n190,n178,n179,n180,n181);
nor (n191,n192,n194,n195,n196);
not (n192,n193);
nor (n197,n192,n198,n195,n196);
not (n198,n194);
nor (n199,n193,n198,n195,n196);
nor (n200,n192,n198,n201,n196);
not (n201,n195);
nor (n202,n193,n194,n201,n203);
not (n203,n196);
and (n204,n192,n194,n195,n196);
and (n205,n192,n194,n201,n196);
and (n206,n193,n194,n201,n196);
and (n207,n193,n198,n201,n196);
nor (n208,n209,n74,n72,n73);
not (n209,n210);
nor (n211,n210,n212,n72,n73);
not (n212,n74);
and (n213,n209,n212,n72,n73);
and (n214,n210,n212,n72,n73);
nor (n215,n216,n217,n219);
not (n217,n218);
and (n220,n216,n218,n219);
nor (n221,n222,n224);
not (n222,n223);
and (n225,n222,n224);
nor (n226,n227,n228,n230,n231);
not (n228,n229);
and (n232,n227,n229,n230,n233);
not (n233,n231);
and (n234,n235,n228,n230,n233);
not (n235,n227);
not (n236,n237);
or (n237,n127,n238);
nand (n238,n239,n254);
or (n239,n240,n253);
nor (n240,n241,n251);
nor (n241,n242,n248);
and (n242,n243,n247);
nand (n243,n244,n245);
or (n244,n90,n92);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n107);
and (s0n245,notn245,n246);
and (s1n245,n107,1'b0);
not (n246,n86);
nor (n247,n108,n109);
not (n248,n249);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n111);
and (s0n249,notn249,n250);
and (s1n249,n111,1'b0);
not (n250,n110);
nand (n251,n252,n114);
not (n252,n122);
or (n253,n117,n116);
not (n254,n125);
wire s0n255,s1n255,notn255;
or (n255,s0n255,s1n255);
not(notn255,n127);
and (s0n255,notn255,n256);
and (s1n255,n127,1'b0);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n125);
and (s0n256,notn256,n257);
and (s1n256,n125,1'b0);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n118);
and (s0n257,notn257,n258);
and (s1n257,n118,n262);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n111);
and (s0n258,notn258,n259);
and (s1n258,n111,1'b1);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n110);
and (s0n259,notn259,n260);
and (s1n259,n110,1'b1);
wire s0n260,s1n260,notn260;
or (n260,s0n260,s1n260);
not(notn260,n109);
and (s0n260,notn260,n261);
and (s1n260,n109,1'b0);
wire s0n261,s1n261,notn261;
or (n261,s0n261,s1n261);
not(notn261,n108);
and (s0n261,notn261,n245);
and (s1n261,n108,1'b0);
not (n262,n253);
not (n263,n264);
wire s0n264,s1n264,notn264;
or (n264,s0n264,s1n264);
not(notn264,n127);
and (s0n264,notn264,n265);
and (s1n264,n127,1'b0);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n125);
and (s0n265,notn265,n266);
and (s1n265,n125,1'b0);
wire s0n266,s1n266,notn266;
or (n266,s0n266,s1n266);
not(notn266,n118);
and (s0n266,notn266,n249);
and (s1n266,n118,1'b0);
and (n267,n268,n271);
xnor (n268,n108,n269);
or (n269,n107,n270);
or (n270,n86,n92);
and (n271,n272,n236,n255,n263);
not (n272,n94);
and (n273,n274,n278);
xnor (n274,n110,n275);
not (n275,n276);
nor (n276,n277,n109);
or (n277,n108,n107);
and (n278,n94,n237,n255,n263);
and (n279,n280,n283);
xnor (n280,n122,n281);
or (n281,n111,n282);
or (n282,n110,n109);
and (n283,n272,n237,n255,n263);
and (n284,n285,n288);
not (n285,n286);
nand (n286,n287,n263,n94,n236);
not (n287,n255);
not (n288,n289);
nand (n289,n290,n116);
or (n290,n115,n291);
not (n291,n292);
nor (n292,n111,n122);
or (n293,n294,n340);
or (n294,n295,n316,n324,n330);
nand (n295,n296,n307);
or (n296,n297,n216);
nand (n297,n298,n305,n218);
nor (n298,n299,n73);
not (n299,n300);
and (n300,n301,n302,n203);
nor (n301,n195,n194);
nor (n302,n303,n193);
not (n303,n304);
nor (n305,n306,n210);
nand (n306,n212,n72);
nor (n307,n308,n310);
and (n308,n298,n309,n223);
nor (n309,n209,n306);
nand (n310,n311,n315);
or (n311,n312,n314);
nor (n312,n313,n301);
and (n313,n194,n203);
nand (n314,n193,n304);
nand (n315,n201,n302,n194);
nor (n316,n317,n322,n181);
nand (n317,n298,n318);
and (n318,n319,n321,n212);
not (n319,n320);
or (n320,n163,n165,n166,n167);
nor (n321,n72,n210);
nor (n322,n323,n178);
and (n323,n180,n179);
nor (n324,n325,n326,n327,n319);
not (n325,n321);
not (n326,n298);
nor (n327,n328,n329);
and (n328,n166,n163);
nor (n329,n163,n167);
nor (n330,n331,n338);
nor (n331,n332,n305);
and (n332,n333,n337);
not (n333,n334);
nor (n334,n335,n336);
and (n335,n321,n74);
and (n336,n210,n212);
not (n337,n73);
nand (n338,n339,n300);
or (n339,n306,n73);
wire s0n340,s1n340,notn340;
or (n340,s0n340,s1n340);
not(notn340,n303);
and (s0n340,notn340,n341);
and (s1n340,n303,1'b0);
wire s0n341,s1n341,notn341;
or (n341,s0n341,s1n341);
not(notn341,n356);
and (s0n341,notn341,n342);
and (s1n341,n356,n355);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n354);
and (s0n342,notn342,n343);
and (s1n342,n354,n346);
wire s0n343,s1n343,notn343;
or (n343,s0n343,s1n343);
not(notn343,n320);
and (s0n343,notn343,n344);
and (s1n343,n320,1'b0);
or (n344,n345,n190);
or (n345,n188,n189);
or (n346,1'b0,n214,n347,n352,1'b0);
and (n347,n348,n351);
or (n348,1'b0,n220,n349,1'b0);
and (n349,n350,n218,n219);
not (n350,n216);
and (n351,n209,n212,n72,n337);
and (n352,n224,n353);
and (n353,n210,n212,n72,n337);
or (n354,n210,n74,n72,n73);
or (n355,n204,n206);
or (n356,n193,n194,n195,n196);
nor (n357,n358,n360,n363);
not (n358,n359);
not (n360,n361);
xor (n361,n362,n359);
xor (n363,n364,n365);
and (n365,n362,n359);
and (n366,n294,n340);
and (n367,n368,n443);
wire s0n368,s1n368,notn368;
or (n368,s0n368,s1n368);
not(notn368,n428);
and (s0n368,notn368,n369);
and (s1n368,n428,n424);
xor (n369,n370,n386);
not (n370,n371);
wire s0n371,s1n371,notn371;
or (n371,s0n371,s1n371);
not(notn371,n293);
and (s0n371,notn371,1'b0);
and (s1n371,n293,n372);
or (n372,n373,n376,n379,n383,1'b0,1'b0,1'b0,1'b0);
and (n373,n374,n93);
xnor (n374,n107,n375);
or (n375,n89,n270);
and (n376,n377,n271);
xnor (n377,n109,n378);
or (n378,n108,n269);
and (n379,n380,n278);
xnor (n380,n111,n381);
not (n381,n382);
and (n382,n276,n250);
and (n383,n384,n283);
xnor (n384,n115,n385);
or (n385,n122,n281);
and (n386,n387,n388);
not (n387,n82);
and (n388,n389,n406);
not (n389,n390);
wire s0n390,s1n390,notn390;
or (n390,s0n390,s1n390);
not(notn390,n293);
and (s0n390,notn390,1'b0);
and (s1n390,n293,n391);
or (n391,n392,n394,n396,n398,n400,n403,1'b0,1'b0);
and (n392,n393,n93);
xnor (n393,n92,n89);
and (n394,n395,n271);
xnor (n395,n107,n270);
and (n396,n397,n278);
xnor (n397,n109,n277);
and (n398,n399,n283);
xnor (n399,n111,n282);
nor (n400,n401,n286);
not (n401,n402);
xnor (n402,n115,n291);
and (n403,n404,n405);
xnor (n404,n117,n120);
nor (n405,n94,n237,n255,n264);
not (n406,n407);
wire s0n407,s1n407,notn407;
or (n407,s0n407,s1n407);
not(notn407,n293);
and (s0n407,notn407,1'b0);
and (s1n407,n293,n408);
or (n408,n409,n411,n413,n415,n417,n419,n421,1'b0);
and (n409,n410,n93);
xnor (n410,n90,n91);
and (n411,n412,n271);
xnor (n412,n86,n92);
and (n413,n414,n278);
xnor (n414,n108,n107);
and (n415,n416,n283);
xnor (n416,n110,n109);
and (n417,n418,n285);
xnor (n418,n122,n111);
and (n419,n420,n405);
xnor (n420,n116,n115);
and (n421,n422,n423);
xnor (n422,n126,n117);
nor (n423,n272,n236,n255,n264);
xor (n424,n371,n425);
and (n425,n82,n426);
and (n426,n390,n427);
and (n427,n407,n428);
wire s0n428,s1n428,notn428;
or (n428,s0n428,s1n428);
not(notn428,n293);
and (s0n428,notn428,1'b0);
and (s1n428,n293,n429);
or (n429,n430,n431,n433,n435,n437,n440,n441,1'b0);
and (n430,n105,n93);
and (n431,n432,n271);
not (n432,n92);
and (n433,n434,n278);
not (n434,n107);
and (n435,n436,n283);
not (n436,n109);
not (n437,n438);
nand (n438,n285,n439);
not (n439,n111);
and (n440,n114,n405);
and (n441,n442,n423);
not (n442,n117);
nor (n443,n444,n294);
not (n444,n340);
and (n445,n82,n446);
and (n446,n294,n444);
not (n447,n448);
nand (n448,n449,n473);
or (n449,n450,n457);
or (n450,n451,n456);
nor (n451,n452,n453,n455);
not (n453,n454);
and (n456,n452,n454,n455);
not (n457,n458);
nand (n458,n459,n467);
or (n459,1'b0,n460,n462,n466);
and (n460,n461,n366);
wire s0n461,s1n461,notn461;
or (n461,s0n461,s1n461);
not(notn461,n357);
and (s0n461,notn461,n390);
and (s1n461,n357,1'b0);
and (n462,n463,n443);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n428);
and (s0n463,notn463,n464);
and (s1n463,n428,n465);
xor (n464,n387,n388);
xor (n465,n82,n426);
and (n466,n390,n446);
or (n467,1'b0,n468,n470,n472);
and (n468,n469,n366);
wire s0n469,s1n469,notn469;
or (n469,s0n469,s1n469);
not(notn469,n357);
and (s0n469,notn469,n407);
and (s1n469,n357,1'b0);
and (n470,n471,n443);
xor (n471,n389,n406);
and (n472,n407,n446);
nor (n473,n474,n497);
not (n474,n475);
or (n475,1'b0,n476,n478,n496);
and (n476,n477,n366);
wire s0n477,s1n477,notn477;
or (n477,s0n477,s1n477);
not(notn477,n357);
and (s0n477,notn477,n371);
and (s1n477,n357,1'b0);
and (n478,n479,n443);
wire s0n479,s1n479,notn479;
or (n479,s0n479,s1n479);
not(notn479,n428);
and (s0n479,notn479,n480);
and (s1n479,n428,n494);
xor (n480,n481,n493);
not (n481,n482);
wire s0n482,s1n482,notn482;
or (n482,s0n482,s1n482);
not(notn482,n293);
and (s0n482,notn482,1'b0);
and (s1n482,n293,n483);
or (n483,n484,n487,n490,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n484,n485,n93);
xnor (n485,n108,n486);
or (n486,n375,n107);
and (n487,n488,n271);
xnor (n488,n110,n489);
or (n489,n109,n378);
and (n490,n491,n278);
xnor (n491,n122,n492);
or (n492,n111,n381);
and (n493,n370,n386);
xor (n494,n482,n495);
and (n495,n371,n425);
and (n496,n371,n446);
nor (n497,n498,n501);
nand (n498,n499,n500);
not (n499,n459);
not (n500,n467);
or (n501,1'b0,n502,n520,n522);
and (n502,n503,n366);
wire s0n503,s1n503,notn503;
or (n503,s0n503,s1n503);
not(notn503,n357);
and (s0n503,notn503,n428);
and (s1n503,n357,n504);
not (n504,n505);
nor (n505,n428,n407,n390,n82,n371,n482,n506,n517);
wire s0n506,s1n506,notn506;
or (n506,s0n506,s1n506);
not(notn506,n293);
and (s0n506,notn506,1'b0);
and (s1n506,n293,n507);
or (n507,n508,n514,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n508,n509,n93);
nand (n509,n510,n512);
or (n510,n511,n436);
nor (n511,n375,n277);
nand (n512,n513,n276);
not (n513,n375);
and (n514,n515,n271);
xnor (n515,n111,n516);
or (n516,n110,n489);
wire s0n517,s1n517,notn517;
or (n517,s0n517,s1n517);
not(notn517,n293);
and (s0n517,notn517,1'b0);
and (s1n517,n293,n518);
and (n518,n519,n93);
xnor (n519,n110,n512);
and (n520,n521,n443);
xor (n521,n407,n428);
and (n522,n428,n446);
nand (n523,n524,n78);
or (n524,n525,n527);
not (n525,n526);
nor (n526,n475,n450);
not (n527,n528);
nand (n528,n529,n459);
nand (n529,n530,n500);
not (n530,n501);
nor (n531,n532,n566);
nand (n532,n533,n548,n557);
not (n533,n534);
or (n534,1'b0,n535,n537,n547);
and (n535,n536,n366);
wire s0n536,s1n536,notn536;
or (n536,s0n536,s1n536);
not(notn536,n357);
and (s0n536,notn536,n506);
and (s1n536,n357,1'b0);
and (n537,n538,n443);
wire s0n538,s1n538,notn538;
or (n538,s0n538,s1n538);
not(notn538,n428);
and (s0n538,notn538,n539);
and (s1n538,n428,n544);
xor (n539,n540,n541);
not (n540,n517);
and (n541,n542,n543);
not (n542,n506);
and (n543,n481,n493);
xor (n544,n517,n545);
and (n545,n506,n546);
and (n546,n482,n495);
and (n547,n506,n446);
not (n548,n549);
or (n549,1'b0,n550,n552,n556);
and (n550,n551,n366);
wire s0n551,s1n551,notn551;
or (n551,s0n551,s1n551);
not(notn551,n357);
and (s0n551,notn551,n482);
and (s1n551,n357,1'b0);
and (n552,n553,n443);
wire s0n553,s1n553,notn553;
or (n553,s0n553,s1n553);
not(notn553,n428);
and (s0n553,notn553,n554);
and (s1n553,n428,n555);
xor (n554,n542,n543);
xor (n555,n506,n546);
and (n556,n482,n446);
not (n557,n558);
or (n558,1'b0,n559,n561,n565);
and (n559,n560,n366);
wire s0n560,s1n560,notn560;
or (n560,s0n560,s1n560);
not(notn560,n357);
and (s0n560,notn560,n517);
and (s1n560,n357,1'b0);
and (n561,n562,n443);
wire s0n562,s1n562,notn562;
or (n562,s0n562,s1n562);
not(notn562,n428);
and (s0n562,notn562,n563);
and (s1n562,n428,1'b0);
not (n563,n564);
and (n564,n540,n541);
and (n565,n517,n446);
not (n566,n211);
and (n567,n568,n42);
wire s0n568,s1n568,notn568;
or (n568,s0n568,s1n568);
not(notn568,n31);
and (s0n568,notn568,n569);
and (s1n568,n31,n570);
or (n570,n571,n573,n575,n577);
and (n571,n572,n19);
and (n573,n574,n24);
and (n575,n576,n28);
and (n577,n569,n30);
and (n578,n579,n47);
wire s0n579,s1n579,notn579;
or (n579,s0n579,s1n579);
not(notn579,n31);
and (s0n579,notn579,n580);
and (s1n579,n31,n581);
or (n581,n582,n584,n586,n588);
and (n582,n583,n19);
and (n584,n585,n24);
and (n586,n587,n28);
and (n588,n580,n30);
and (n589,n590,n50);
wire s0n590,s1n590,notn590;
or (n590,s0n590,s1n590);
not(notn590,n31);
and (s0n590,notn590,n591);
and (s1n590,n31,n592);
or (n592,n593,n595,n597,n599);
and (n593,n594,n19);
and (n595,n596,n24);
and (n597,n598,n28);
and (n599,n591,n30);
and (n601,n602,n51);
not (n602,n65);
wire s0n603,s1n603,notn603;
or (n603,s0n603,s1n603);
not(notn603,n600);
and (s0n603,notn603,n604);
and (s1n603,n600,n591);
wire s0n604,s1n604,notn604;
or (n604,s0n604,s1n604);
not(notn604,n31);
and (s0n604,notn604,n605);
and (s1n604,n31,n616);
or (n605,n606,n608,n610,n613);
and (n606,n15,n607);
and (n607,n60,n56);
and (n608,n569,n609);
and (n609,n59,n56);
and (n610,n580,n611);
not (n611,n612);
or (n612,n56,n59);
and (n613,n591,n614);
not (n614,n615);
or (n615,n60,n56);
or (n616,1'b0,n617,n620,n622,n625,n627,n629,n631,n633,n635,n637,n639,n641,n643,n645,n647,n649);
and (n617,n18,n618);
and (n618,n38,n39,n60,n56,n619);
not (n619,n51);
and (n620,n23,n621);
and (n621,n44,n39,n60,n56,n619);
and (n622,n27,n623);
and (n623,n38,n624,n60,n56,n619);
not (n624,n39);
and (n625,n15,n626);
and (n626,n44,n624,n60,n56,n619);
and (n627,n572,n628);
and (n628,n38,n39,n59,n56,n619);
and (n629,n574,n630);
and (n630,n44,n39,n59,n56,n619);
and (n631,n576,n632);
and (n632,n38,n624,n59,n56,n619);
and (n633,n569,n634);
and (n634,n44,n624,n59,n56,n619);
and (n635,n583,n636);
nor (n636,n44,n624,n59,n56,n51);
and (n637,n585,n638);
nor (n638,n38,n624,n59,n56,n51);
and (n639,n587,n640);
nor (n640,n44,n39,n59,n56,n51);
and (n641,n580,n642);
nor (n642,n38,n39,n59,n56,n51);
and (n643,n594,n644);
nor (n644,n44,n624,n60,n56,n51);
and (n645,n596,n646);
nor (n646,n38,n624,n60,n56,n51);
and (n647,n598,n648);
nor (n648,n44,n39,n60,n56,n51);
and (n649,n591,n650);
nor (n650,n38,n39,n60,n56,n51);
and (n651,n602,n619);
not (n652,n653);
wire s0n653,s1n653,notn653;
or (n653,s0n653,s1n653);
not(notn653,n651);
and (s0n653,notn653,1'b0);
and (s1n653,n651,n654);
wire s0n654,s1n654,notn654;
or (n654,s0n654,s1n654);
not(notn654,n651);
and (s0n654,notn654,n655);
and (s1n654,n651,n702);
wire s0n655,s1n655,notn655;
or (n655,s0n655,s1n655);
not(notn655,n601);
and (s0n655,notn655,1'b0);
and (s1n655,n601,n656);
wire s0n656,s1n656,notn656;
or (n656,s0n656,s1n656);
not(notn656,n600);
and (s0n656,notn656,n657);
and (s1n656,n600,n693);
or (n657,n658,n669,n680,n691);
and (n658,n659,n37);
wire s0n659,s1n659,notn659;
or (n659,s0n659,s1n659);
not(notn659,n31);
and (s0n659,notn659,n660);
and (s1n659,n31,n661);
or (n661,n662,n664,n666,n668);
and (n662,n663,n19);
and (n664,n665,n24);
and (n666,n667,n28);
and (n668,n660,n30);
and (n669,n670,n42);
wire s0n670,s1n670,notn670;
or (n670,s0n670,s1n670);
not(notn670,n31);
and (s0n670,notn670,n671);
and (s1n670,n31,n672);
or (n672,n673,n675,n677,n679);
and (n673,n674,n19);
and (n675,n676,n24);
and (n677,n678,n28);
and (n679,n671,n30);
and (n680,n681,n47);
wire s0n681,s1n681,notn681;
or (n681,s0n681,s1n681);
not(notn681,n31);
and (s0n681,notn681,n682);
and (s1n681,n31,n683);
or (n683,n684,n686,n688,n690);
and (n684,n685,n19);
and (n686,n687,n24);
and (n688,n689,n28);
and (n690,n682,n30);
and (n691,n692,n50);
wire s0n692,s1n692,notn692;
or (n692,s0n692,s1n692);
not(notn692,n31);
and (s0n692,notn692,n693);
and (s1n692,n31,n694);
or (n694,n695,n697,n699,n701);
and (n695,n696,n19);
and (n697,n698,n24);
and (n699,n700,n28);
and (n701,n693,n30);
wire s0n702,s1n702,notn702;
or (n702,s0n702,s1n702);
not(notn702,n600);
and (s0n702,notn702,n703);
and (s1n702,n600,n693);
wire s0n703,s1n703,notn703;
or (n703,s0n703,s1n703);
not(notn703,n31);
and (s0n703,notn703,n704);
and (s1n703,n31,n709);
or (n704,n705,n706,n707,n708);
and (n705,n660,n607);
and (n706,n671,n609);
and (n707,n682,n611);
and (n708,n693,n614);
or (n709,1'b0,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725);
and (n710,n663,n618);
and (n711,n665,n621);
and (n712,n667,n623);
and (n713,n660,n626);
and (n714,n674,n628);
and (n715,n676,n630);
and (n716,n678,n632);
and (n717,n671,n634);
and (n718,n685,n636);
and (n719,n687,n638);
and (n720,n689,n640);
and (n721,n682,n642);
and (n722,n696,n644);
and (n723,n698,n646);
and (n724,n700,n648);
and (n725,n693,n650);
wire s0n726,s1n726,notn726;
or (n726,s0n726,s1n726);
not(notn726,n651);
and (s0n726,notn726,1'b0);
and (s1n726,n651,n727);
wire s0n727,s1n727,notn727;
or (n727,s0n727,s1n727);
not(notn727,n651);
and (s0n727,notn727,n728);
and (s1n727,n651,n775);
wire s0n728,s1n728,notn728;
or (n728,s0n728,s1n728);
not(notn728,n601);
and (s0n728,notn728,1'b0);
and (s1n728,n601,n729);
wire s0n729,s1n729,notn729;
or (n729,s0n729,s1n729);
not(notn729,n600);
and (s0n729,notn729,n730);
and (s1n729,n600,n766);
or (n730,n731,n742,n753,n764);
and (n731,n732,n37);
wire s0n732,s1n732,notn732;
or (n732,s0n732,s1n732);
not(notn732,n31);
and (s0n732,notn732,n733);
and (s1n732,n31,n734);
or (n734,n735,n737,n739,n741);
and (n735,n736,n19);
and (n737,n738,n24);
and (n739,n740,n28);
and (n741,n733,n30);
and (n742,n743,n42);
wire s0n743,s1n743,notn743;
or (n743,s0n743,s1n743);
not(notn743,n31);
and (s0n743,notn743,n744);
and (s1n743,n31,n745);
or (n745,n746,n748,n750,n752);
and (n746,n747,n19);
and (n748,n749,n24);
and (n750,n751,n28);
and (n752,n744,n30);
and (n753,n754,n47);
wire s0n754,s1n754,notn754;
or (n754,s0n754,s1n754);
not(notn754,n31);
and (s0n754,notn754,n755);
and (s1n754,n31,n756);
or (n756,n757,n759,n761,n763);
and (n757,n758,n19);
and (n759,n760,n24);
and (n761,n762,n28);
and (n763,n755,n30);
and (n764,n765,n50);
wire s0n765,s1n765,notn765;
or (n765,s0n765,s1n765);
not(notn765,n31);
and (s0n765,notn765,n766);
and (s1n765,n31,n767);
or (n767,n768,n770,n772,n774);
and (n768,n769,n19);
and (n770,n771,n24);
and (n772,n773,n28);
and (n774,n766,n30);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n600);
and (s0n775,notn775,n776);
and (s1n775,n600,n766);
wire s0n776,s1n776,notn776;
or (n776,s0n776,s1n776);
not(notn776,n31);
and (s0n776,notn776,n777);
and (s1n776,n31,n782);
or (n777,n778,n779,n780,n781);
and (n778,n733,n607);
and (n779,n744,n609);
and (n780,n755,n611);
and (n781,n766,n614);
or (n782,1'b0,n783,n784,n785,n786,n787,n788,n789,n790,n791,n792,n793,n794,n795,n796,n797,n798);
and (n783,n736,n618);
and (n784,n738,n621);
and (n785,n740,n623);
and (n786,n733,n626);
and (n787,n747,n628);
and (n788,n749,n630);
and (n789,n751,n632);
and (n790,n744,n634);
and (n791,n758,n636);
and (n792,n760,n638);
and (n793,n762,n640);
and (n794,n755,n642);
and (n795,n769,n644);
and (n796,n771,n646);
and (n797,n773,n648);
and (n798,n766,n650);
nor (n799,n800,n802);
not (n800,n801);
and (n804,n805,n808);
and (n805,n651,n806);
or (n806,n803,n807,n801,n802);
nor (n808,n809,n810,n811);
nand (n812,n813,n818,n1046);
or (n813,n814,n816);
nand (n814,n815,n804);
not (n815,n6);
not (n816,n817);
nor (n817,n803,n807,n800,n802);
or (n818,n819,n820);
or (n819,n809,n810);
not (n820,n821);
nor (n821,n822,n808);
not (n822,n823);
nor (n823,n824,n1038);
or (n824,n825,n1034);
nor (n825,n826,n931,n966,n1000);
wire s0n826,s1n826,notn826;
or (n826,s0n826,s1n826);
not(notn826,n860);
and (s0n826,notn826,1'b1);
and (s1n826,n860,n827);
or (n827,n51,n828,n830,n832,n834,n836,n838,n840,n842,n844,n846,n848,n850,n852,n854,n856,n858);
and (n828,n829,n618);
and (n830,n831,n621);
and (n832,n833,n623);
and (n834,n835,n626);
and (n836,n837,n628);
and (n838,n839,n630);
and (n840,n841,n632);
and (n842,n843,n634);
and (n844,n845,n636);
and (n846,n847,n638);
and (n848,n849,n640);
and (n850,n851,n642);
and (n852,n853,n644);
and (n854,n855,n646);
and (n856,n857,n648);
and (n858,n859,n650);
and (n860,n861,n913,n926,n65);
not (n861,n862);
wire s0n862,s1n862,notn862;
or (n862,s0n862,s1n862);
not(notn862,n912);
and (s0n862,notn862,n863);
and (s1n862,n912,1'b1);
wire s0n863,s1n863,notn863;
or (n863,s0n863,s1n863);
not(notn863,n211);
and (s0n863,notn863,n864);
and (s1n863,n211,n865);
wire s0n865,s1n865,notn865;
or (n865,s0n865,s1n865);
not(notn865,n450);
and (s0n865,notn865,n866);
and (s1n865,n450,n905);
or (n866,n867,1'b0,1'b0,1'b0,n882,1'b0,n883,1'b0);
or (n867,n868,n881);
or (n868,n869,n880);
or (n869,n870,n879);
or (n870,n871,n878);
or (n871,n872,n877);
or (n872,n873,n876);
or (n873,n874,n875);
nor (n874,n501,n500,n459,n78,n475,n549,n534,n558);
nor (n875,n530,n500,n459,n78,n475,n549,n534,n558);
nor (n876,n501,n467,n499,n78,n475,n549,n534,n558);
nor (n877,n530,n467,n499,n78,n475,n549,n534,n558);
nor (n878,n501,n500,n499,n79,n474,n549,n534,n558);
nor (n879,n530,n500,n499,n79,n474,n549,n534,n558);
nor (n880,n501,n467,n459,n78,n474,n549,n534,n558);
nor (n881,n530,n467,n459,n78,n474,n549,n534,n558);
nor (n882,n530,n500,n459,n79,n475,n549,n534,n558);
or (n883,n884,n885);
nor (n884,n530,n467,n459,n79,n475,n549,n534,n558);
nor (n885,n505,n884,n886,n882,n887,n888,n889,n890,n891,n892,n893,n894,n895,n896,n874,n875,n876,n877,n878,n879,n880,n881,n897,n898,n899,n900,n901,n902,n903,n904);
nor (n886,n501,n500,n459,n79,n475,n549,n534,n558);
nor (n887,n501,n467,n499,n79,n475,n549,n534,n558);
nor (n888,n530,n467,n499,n79,n475,n549,n534,n558);
nor (n889,n501,n500,n499,n79,n475,n549,n534,n558);
nor (n890,n530,n500,n499,n79,n475,n549,n534,n558);
nor (n891,n501,n467,n459,n78,n475,n549,n534,n558);
nor (n892,n530,n467,n459,n78,n475,n549,n534,n558);
nor (n893,n501,n500,n459,n79,n474,n549,n534,n558);
nor (n894,n530,n500,n459,n79,n474,n549,n534,n558);
nor (n895,n501,n467,n499,n79,n474,n549,n534,n558);
nor (n896,n530,n467,n499,n79,n474,n549,n534,n558);
nor (n897,n501,n500,n499,n78,n475,n549,n534,n558);
nor (n898,n530,n500,n499,n78,n475,n549,n534,n558);
nor (n899,n501,n467,n459,n79,n474,n549,n534,n558);
nor (n900,n530,n467,n459,n79,n474,n549,n534,n558);
nor (n901,n501,n500,n459,n78,n474,n549,n534,n558);
nor (n902,n530,n500,n459,n78,n474,n549,n534,n558);
nor (n903,n501,n467,n499,n78,n474,n549,n534,n558);
nor (n904,n530,n467,n499,n78,n474,n549,n534,n558);
or (n905,n906,n895);
or (n906,n907,n894);
or (n907,n908,n893);
or (n908,n909,n900);
or (n909,n910,n891);
or (n910,n911,n890);
or (n911,n888,n889);
nor (n912,n209,n212,n72,n73);
not (n913,n914);
wire s0n914,s1n914,notn914;
or (n914,s0n914,s1n914);
not(notn914,n912);
and (s0n914,notn914,n915);
and (s1n914,n912,1'b0);
wire s0n915,s1n915,notn915;
or (n915,s0n915,s1n915);
not(notn915,n211);
and (s0n915,notn915,n916);
and (s1n915,n211,n917);
wire s0n917,s1n917,notn917;
or (n917,s0n917,s1n917);
not(notn917,n450);
and (s0n917,notn917,n918);
and (s1n917,n450,n919);
or (n918,1'b0,1'b0,1'b0,1'b0,n882,n886,1'b0,1'b0);
or (n919,n920,n880);
or (n920,n921,n879);
or (n921,n922,n878);
or (n922,n923,n896);
or (n923,n924,n876);
or (n924,n925,n875);
or (n925,n892,n874);
wire s0n926,s1n926,notn926;
or (n926,s0n926,s1n926);
not(notn926,n912);
and (s0n926,notn926,n927);
and (s1n926,n912,1'b1);
wire s0n927,s1n927,notn927;
or (n927,s0n927,s1n927);
not(notn927,n211);
and (s0n927,notn927,n928);
and (s1n927,n211,n929);
wire s0n929,s1n929,notn929;
or (n929,s0n929,s1n929);
not(notn929,n450);
and (s0n929,notn929,n930);
and (s1n929,n450,n505);
or (n930,1'b0,1'b0,n888,n887,1'b0,1'b0,1'b0,1'b0);
not (n931,n932);
wire s0n932,s1n932,notn932;
or (n932,s0n932,s1n932);
not(notn932,n860);
and (s0n932,notn932,1'b1);
and (s1n932,n860,n933);
or (n933,n51,n934,n936,n938,n940,n942,n944,n946,n948,n950,n952,n954,n956,n958,n960,n962,n964);
and (n934,n935,n618);
and (n936,n937,n621);
and (n938,n939,n623);
and (n940,n941,n626);
and (n942,n943,n628);
and (n944,n945,n630);
and (n946,n947,n632);
and (n948,n949,n634);
and (n950,n951,n636);
and (n952,n953,n638);
and (n954,n955,n640);
and (n956,n957,n642);
and (n958,n959,n644);
and (n960,n961,n646);
and (n962,n963,n648);
and (n964,n965,n650);
wire s0n966,s1n966,notn966;
or (n966,s0n966,s1n966);
not(notn966,n860);
and (s0n966,notn966,1'b1);
and (s1n966,n860,n967);
or (n967,n51,n968,n970,n972,n974,n976,n978,n980,n982,n984,n986,n988,n990,n992,n994,n996,n998);
and (n968,n969,n618);
and (n970,n971,n621);
and (n972,n973,n623);
and (n974,n975,n626);
and (n976,n977,n628);
and (n978,n979,n630);
and (n980,n981,n632);
and (n982,n983,n634);
and (n984,n985,n636);
and (n986,n987,n638);
and (n988,n989,n640);
and (n990,n991,n642);
and (n992,n993,n644);
and (n994,n995,n646);
and (n996,n997,n648);
and (n998,n999,n650);
wire s0n1000,s1n1000,notn1000;
or (n1000,s0n1000,s1n1000);
not(notn1000,n860);
and (s0n1000,notn1000,1'b1);
and (s1n1000,n860,n1001);
or (n1001,n51,n1002,n1004,n1006,n1008,n1010,n1012,n1014,n1016,n1018,n1020,n1022,n1024,n1026,n1028,n1030,n1032);
and (n1002,n1003,n618);
and (n1004,n1005,n621);
and (n1006,n1007,n623);
and (n1008,n1009,n626);
and (n1010,n1011,n628);
and (n1012,n1013,n630);
and (n1014,n1015,n632);
and (n1016,n1017,n634);
and (n1018,n1019,n636);
and (n1020,n1021,n638);
and (n1022,n1023,n640);
and (n1024,n1025,n642);
and (n1026,n1027,n644);
and (n1028,n1029,n646);
and (n1030,n1031,n648);
and (n1032,n1033,n650);
nor (n1034,n1035,n1036,n1037);
nand (n1035,n65,n51);
and (n1038,n1039,n1042);
and (n1039,n1040,n619);
and (n1040,n1041,n65);
not (n1041,n926);
and (n1042,n1043,n1045);
not (n1043,n1044);
nand (n1046,n1047,n1057);
nand (n1047,n1048,n1052);
or (n1048,n1049,n1050);
not (n1049,n824);
nand (n1050,n1051,n809,n810);
not (n1051,n811);
nand (n1052,n1053,n1038,n1055,n1056);
not (n1053,n1054);
or (n1054,n811,n810);
nor (n1055,n39,n60);
nor (n1056,n38,n56);
not (n1057,n808);
nand (n1058,n1059,n1064);
not (n1059,n1060);
nor (n1060,n1061,n1062);
and (n1061,n31,n21,n20);
and (n1062,n1063,n817);
not (n1063,n31);
nor (n1064,n1065,n805,n1057);
not (n1065,n1066);
and (n1066,n601,n806);
and (n1068,n1069,n1070);
not (n1069,n2);
nand (n1070,n1071,n9977);
or (n1071,n1072,n1074);
not (n1072,n1073);
or (n1073,n1064,n804);
not (n1074,n1075);
nand (n1075,n1076,n7997);
not (n1076,n1077);
nand (n1077,n1078,n7987);
or (n1078,n1079,n7984);
nor (n1079,n1080,n7978);
and (n1080,n1081,n7758);
nand (n1081,n1082,n7750);
or (n1082,n1083,n7237);
nand (n1083,n1084,n7125);
nand (n1084,n1085,n7031);
not (n1085,n1086);
or (n1086,1'b0,n1087,n4926,n4928,n4930);
and (n1087,n1088,n1189);
wire s0n1088,s1n1088,notn1088;
or (n1088,s0n1088,s1n1088);
not(notn1088,n4923);
and (s0n1088,notn1088,1'b0);
and (s1n1088,n4923,n1089);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n4903);
and (s0n1089,notn1089,n1090);
and (s1n1089,n4903,1'b0);
wire s0n1090,s1n1090,notn1090;
or (n1090,s0n1090,s1n1090);
not(notn1090,n4777);
and (s0n1090,notn1090,n1091);
and (s1n1090,n4777,1'b1);
wire s0n1091,s1n1091,notn1091;
or (n1091,s0n1091,s1n1091);
not(notn1091,n1102);
and (s0n1091,notn1091,n1092);
and (s1n1091,n1102,n4116);
wire s0n1092,s1n1092,notn1092;
or (n1092,s0n1092,s1n1092);
not(notn1092,n1102);
and (s0n1092,notn1092,n1093);
and (s1n1092,n1102,n4115);
xor (n1093,n1094,n4098);
xor (n1094,n1095,n4053);
xor (n1095,n1096,n3998);
xor (n1096,n1097,n3988);
xor (n1097,n1098,n2267);
xor (n1098,n1099,n1197);
xor (n1099,n1100,n1195);
wire s0n1100,s1n1100,notn1100;
or (n1100,s0n1100,s1n1100);
not(notn1100,n1102);
and (s0n1100,notn1100,1'b0);
and (s1n1100,n1102,n1101);
or (n1102,n1103,n1193);
or (n1103,n1104,n1188);
and (n1104,n1105,n1180);
and (n1105,n652,n726,n1106,n1107);
not (n1106,n7);
wire s0n1107,s1n1107,notn1107;
or (n1107,s0n1107,s1n1107);
not(notn1107,n651);
and (s0n1107,notn1107,1'b0);
and (s1n1107,n651,n1108);
wire s0n1108,s1n1108,notn1108;
or (n1108,s0n1108,s1n1108);
not(notn1108,n651);
and (s0n1108,notn1108,n1109);
and (s1n1108,n651,n1156);
wire s0n1109,s1n1109,notn1109;
or (n1109,s0n1109,s1n1109);
not(notn1109,n601);
and (s0n1109,notn1109,1'b0);
and (s1n1109,n601,n1110);
wire s0n1110,s1n1110,notn1110;
or (n1110,s0n1110,s1n1110);
not(notn1110,n600);
and (s0n1110,notn1110,n1111);
and (s1n1110,n600,n1147);
or (n1111,n1112,n1123,n1134,n1145);
and (n1112,n1113,n37);
wire s0n1113,s1n1113,notn1113;
or (n1113,s0n1113,s1n1113);
not(notn1113,n31);
and (s0n1113,notn1113,n1114);
and (s1n1113,n31,n1115);
or (n1115,n1116,n1118,n1120,n1122);
and (n1116,n1117,n19);
and (n1118,n1119,n24);
and (n1120,n1121,n28);
and (n1122,n1114,n30);
and (n1123,n1124,n42);
wire s0n1124,s1n1124,notn1124;
or (n1124,s0n1124,s1n1124);
not(notn1124,n31);
and (s0n1124,notn1124,n1125);
and (s1n1124,n31,n1126);
or (n1126,n1127,n1129,n1131,n1133);
and (n1127,n1128,n19);
and (n1129,n1130,n24);
and (n1131,n1132,n28);
and (n1133,n1125,n30);
and (n1134,n1135,n47);
wire s0n1135,s1n1135,notn1135;
or (n1135,s0n1135,s1n1135);
not(notn1135,n31);
and (s0n1135,notn1135,n1136);
and (s1n1135,n31,n1137);
or (n1137,n1138,n1140,n1142,n1144);
and (n1138,n1139,n19);
and (n1140,n1141,n24);
and (n1142,n1143,n28);
and (n1144,n1136,n30);
and (n1145,n1146,n50);
wire s0n1146,s1n1146,notn1146;
or (n1146,s0n1146,s1n1146);
not(notn1146,n31);
and (s0n1146,notn1146,n1147);
and (s1n1146,n31,n1148);
or (n1148,n1149,n1151,n1153,n1155);
and (n1149,n1150,n19);
and (n1151,n1152,n24);
and (n1153,n1154,n28);
and (n1155,n1147,n30);
wire s0n1156,s1n1156,notn1156;
or (n1156,s0n1156,s1n1156);
not(notn1156,n600);
and (s0n1156,notn1156,n1157);
and (s1n1156,n600,n1147);
wire s0n1157,s1n1157,notn1157;
or (n1157,s0n1157,s1n1157);
not(notn1157,n31);
and (s0n1157,notn1157,n1158);
and (s1n1157,n31,n1163);
or (n1158,n1159,n1160,n1161,n1162);
and (n1159,n1114,n607);
and (n1160,n1125,n609);
and (n1161,n1136,n611);
and (n1162,n1147,n614);
or (n1163,1'b0,n1164,n1165,n1166,n1167,n1168,n1169,n1170,n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179);
and (n1164,n1117,n618);
and (n1165,n1119,n621);
and (n1166,n1121,n623);
and (n1167,n1114,n626);
and (n1168,n1128,n628);
and (n1169,n1130,n630);
and (n1170,n1132,n632);
and (n1171,n1125,n634);
and (n1172,n1139,n636);
and (n1173,n1141,n638);
and (n1174,n1143,n640);
and (n1175,n1136,n642);
and (n1176,n1150,n644);
and (n1177,n1152,n646);
and (n1178,n1154,n648);
and (n1179,n1147,n650);
or (n1180,n1181,n1187);
or (n1181,n1182,n1186);
or (n1182,n817,n1183);
nor (n1183,n1184,n1185,n801,n802);
not (n1184,n803);
not (n1185,n807);
nor (n1186,n803,n1185,n801,n802);
nor (n1187,n1184,n807,n801,n802);
and (n1188,n1189,n1180);
or (n1189,n1190,n1192);
nor (n1190,n652,n726,n7,n1191);
not (n1191,n1107);
and (n1192,n653,n726,n1106,n1107);
and (n1193,n6,n651,n1194);
nor (n1194,n1184,n802);
wire s0n1195,s1n1195,notn1195;
or (n1195,s0n1195,s1n1195);
not(notn1195,n1102);
and (s0n1195,notn1195,1'b0);
and (s1n1195,n1102,n1196);
or (n1197,n1198,n1203,n2266);
and (n1198,n1199,n1201);
wire s0n1199,s1n1199,notn1199;
or (n1199,s0n1199,s1n1199);
not(notn1199,n1102);
and (s0n1199,notn1199,1'b0);
and (s1n1199,n1102,n1200);
wire s0n1201,s1n1201,notn1201;
or (n1201,s0n1201,s1n1201);
not(notn1201,n1102);
and (s0n1201,notn1201,1'b0);
and (s1n1201,n1102,n1202);
and (n1203,n1201,n1204);
or (n1204,n1205,n1210,n2265);
and (n1205,n1206,n1208);
wire s0n1206,s1n1206,notn1206;
or (n1206,s0n1206,s1n1206);
not(notn1206,n1102);
and (s0n1206,notn1206,1'b0);
and (s1n1206,n1102,n1207);
wire s0n1208,s1n1208,notn1208;
or (n1208,s0n1208,s1n1208);
not(notn1208,n1102);
and (s0n1208,notn1208,1'b0);
and (s1n1208,n1102,n1209);
and (n1210,n1208,n1211);
or (n1211,n1212,n1404,n2264);
and (n1212,n1213,n1333);
wire s0n1213,s1n1213,notn1213;
or (n1213,s0n1213,s1n1213);
not(notn1213,n1102);
and (s0n1213,notn1213,n1214);
and (s1n1213,n1102,n1332);
nand (n1214,n1215,n1278,n1290,n1302);
nor (n1215,n1216,n1273);
nand (n1216,n1217,n1263,n1268);
nor (n1217,n1218,n1252);
and (n1218,n1219,n1251);
and (n1219,n1220,n1246);
or (n1220,n1221,n1238);
not (n1221,n1222);
nand (n1222,n1223,n1233,n1191);
nand (n1223,n1224,n1231);
or (n1224,n1225,n1226);
not (n1225,n1187);
not (n1226,n1227);
nand (n1227,n1228,n1229);
nand (n1228,n1106,n1191,n726);
nand (n1229,n1230,n653);
or (n1230,n1191,n7);
not (n1231,n1232);
and (n1232,n7,n652,n726,n1186);
not (n1233,n1234);
nand (n1234,n1235,n1237);
or (n1235,n1236,n1226);
not (n1236,n1186);
nand (n1237,n7,n652,n726,n817);
not (n1238,n1239);
nand (n1239,n1240,n1234,n1242,n1107);
and (n1240,n1241,n1224);
nand (n1241,n1227,n1183);
and (n1242,n1231,n1243);
nand (n1243,n652,n7,n726,n1244);
and (n1244,n1184,n807,n801,n1245);
not (n1245,n802);
not (n1246,n1247);
nand (n1247,n1248,n1249,n651);
or (n1248,n31,n624);
not (n1249,n1250);
nor (n1250,n44,n31);
and (n1252,n1253,n1262);
not (n1253,n1254);
nand (n1254,n1255,n1246);
not (n1255,n1256);
nand (n1256,n1257,n1191);
nand (n1257,n1258,n1259);
or (n1258,n816,n1226);
not (n1259,n1260);
and (n1260,n6,n1261);
nor (n1261,n803,n807,n801,n1245);
nand (n1263,n1264,n1267);
and (n1264,n1220,n1265);
and (n1265,n1250,n1266);
and (n1266,n651,n624);
nand (n1268,n1269,n1272);
and (n1269,n1270,n1265);
and (n1270,n1271,n1223,n1233,n1107);
and (n1271,n1241,n1243);
and (n1273,n1274,n1277);
nand (n1274,n1275,n1276);
nand (n1275,n1270,n1246);
nand (n1276,n1255,n1265);
nor (n1278,n1279,n1286);
and (n1279,n1280,n1285);
not (n1280,n1281);
nand (n1281,n1282,n1265);
nand (n1282,n1283,n1284);
or (n1283,n1191,n1271);
nand (n1284,n1240,n1234,n1242,n1191);
nor (n1286,n1287,n1289);
not (n1287,n1288);
nand (n1289,n1282,n1246);
nor (n1290,n1291,n1298);
and (n1291,n1292,n1297);
not (n1292,n1293);
nand (n1293,n1294,n1265);
nand (n1294,n1295,n1296);
or (n1295,n1107,n1271);
nand (n1296,n1257,n1107);
and (n1298,n1299,n1301);
not (n1299,n1300);
nand (n1300,n1294,n1246);
nor (n1302,n1303,n1319);
and (n1303,n1304,n1316);
nand (n1304,n1305,n1310,n1312,n1314);
nor (n1305,n1306,n1308);
and (n1306,n1270,n1307);
and (n1308,n1255,n1309);
nand (n1310,n1220,n1311);
nand (n1312,n1282,n1313);
nand (n1314,n1294,n1315);
and (n1316,n1317,n1318);
and (n1317,n651,n39);
nor (n1318,n31,n38);
and (n1319,n1320,n1331);
nand (n1320,n1321,n1325,n1327,n1329);
nor (n1321,n1322,n1324);
and (n1322,n1270,n1323);
and (n1324,n1255,n1307);
nand (n1325,n1220,n1326);
nand (n1327,n1282,n1328);
nand (n1329,n1294,n1330);
and (n1331,n1317,n1250);
wire s0n1333,s1n1333,notn1333;
or (n1333,s0n1333,s1n1333);
not(notn1333,n1102);
and (s0n1333,notn1333,n1334);
and (s1n1333,n1102,n1403);
or (n1334,1'b0,n1335,n1358,n1372,n1385);
and (n1335,n1336,n1331);
or (n1336,1'b0,n1337,n1348,n1351,n1355);
and (n1337,n1338,n1223);
wire s0n1338,s1n1338,notn1338;
or (n1338,s0n1338,s1n1338);
not(notn1338,n1341);
and (s0n1338,notn1338,n1339);
and (s1n1338,n1341,n1340);
or (n1341,n1342,n1346);
or (n1342,n1343,n1345);
and (n1343,n653,n1344,n7,n1107);
not (n1344,n726);
and (n1345,n653,n726,n7,n1107);
not (n1346,n1347);
nand (n1347,n652,n726,n7,n1107);
and (n1348,n1349,n1234);
wire s0n1349,s1n1349,notn1349;
or (n1349,s0n1349,s1n1349);
not(notn1349,n1341);
and (s0n1349,notn1349,n1350);
and (s1n1349,n1341,n1339);
and (n1351,n1352,n1354);
wire s0n1352,s1n1352,notn1352;
or (n1352,s0n1352,s1n1352);
not(notn1352,n1341);
and (s0n1352,notn1352,n1353);
and (s1n1352,n1341,n1350);
not (n1354,n1271);
and (n1355,n1356,n1257);
wire s0n1356,s1n1356,notn1356;
or (n1356,s0n1356,s1n1356);
not(notn1356,n1341);
and (s0n1356,notn1356,n1357);
and (s1n1356,n1341,n1353);
and (n1358,n1359,n1316);
or (n1359,1'b0,n1360,n1363,n1366,n1369);
and (n1360,n1361,n1223);
wire s0n1361,s1n1361,notn1361;
or (n1361,s0n1361,s1n1361);
not(notn1361,n1341);
and (s0n1361,notn1361,n1362);
and (s1n1361,n1341,n1357);
and (n1363,n1364,n1234);
wire s0n1364,s1n1364,notn1364;
or (n1364,s0n1364,s1n1364);
not(notn1364,n1341);
and (s0n1364,notn1364,n1365);
and (s1n1364,n1341,n1362);
and (n1366,n1367,n1354);
wire s0n1367,s1n1367,notn1367;
or (n1367,s0n1367,s1n1367);
not(notn1367,n1341);
and (s0n1367,notn1367,n1368);
and (s1n1367,n1341,n1365);
and (n1369,n1370,n1257);
wire s0n1370,s1n1370,notn1370;
or (n1370,s0n1370,s1n1370);
not(notn1370,n1341);
and (s0n1370,notn1370,n1371);
and (s1n1370,n1341,n1368);
and (n1372,n1373,n1265);
nand (n1373,n1374,n1379,n1381,n1383);
nor (n1374,n1375,n1377);
and (n1375,n1270,n1376);
and (n1377,n1255,n1378);
nand (n1379,n1220,n1380);
nand (n1381,n1282,n1382);
nand (n1383,n1294,n1384);
and (n1385,n1386,n1246);
nand (n1386,n1387,n1392);
nor (n1387,n1388,n1390);
and (n1388,n1282,n1389);
and (n1390,n1294,n1391);
nor (n1392,n1393,n1399);
nand (n1393,n1394,n1397);
or (n1394,n1395,n1396);
not (n1395,n1378);
not (n1396,n1270);
nand (n1397,n1255,n1398);
nor (n1399,n1400,n1402);
not (n1400,n1401);
not (n1402,n1220);
and (n1404,n1333,n1405);
or (n1405,n1406,n1529,n2263);
and (n1406,n1407,n1460);
wire s0n1407,s1n1407,notn1407;
or (n1407,s0n1407,s1n1407);
not(notn1407,n1102);
and (s0n1407,notn1407,n1408);
and (s1n1407,n1102,n1459);
nand (n1408,n1409,n1422,n1448,n1454);
nor (n1409,n1410,n1420);
nand (n1410,n1411,n1416,n1418);
nor (n1411,n1412,n1414);
and (n1412,n1219,n1413);
and (n1414,n1253,n1415);
nand (n1416,n1264,n1417);
nand (n1418,n1269,n1419);
and (n1420,n1274,n1421);
nor (n1422,n1423,n1436);
and (n1423,n1424,n1316);
nand (n1424,n1425,n1427,n1429,n1434);
nand (n1425,n1282,n1426);
nand (n1427,n1294,n1428);
nor (n1429,n1430,n1432);
and (n1430,n1270,n1431);
and (n1432,n1255,n1433);
nand (n1434,n1220,n1435);
and (n1436,n1437,n1331);
nand (n1437,n1438,n1440,n1442,n1446);
nand (n1438,n1282,n1439);
nand (n1440,n1294,n1441);
nor (n1442,n1443,n1445);
and (n1443,n1270,n1444);
and (n1445,n1255,n1431);
nand (n1446,n1220,n1447);
nor (n1448,n1449,n1452);
and (n1449,n1450,n1451);
not (n1450,n1289);
and (n1452,n1280,n1453);
nor (n1454,n1455,n1457);
and (n1455,n1299,n1456);
and (n1457,n1292,n1458);
wire s0n1460,s1n1460,notn1460;
or (n1460,s0n1460,s1n1460);
not(notn1460,n1102);
and (s0n1460,notn1460,n1461);
and (s1n1460,n1102,n1528);
nand (n1461,n1462,n1485,n1511,n1519);
nor (n1462,n1463,n1468);
and (n1463,n1464,n1467);
nand (n1464,n1465,n1466);
nand (n1465,n1270,n1316);
nand (n1466,n1255,n1331);
nand (n1468,n1469,n1477,n1481);
nor (n1469,n1470,n1473);
and (n1470,n1471,n1472);
and (n1471,n1220,n1316);
and (n1473,n1474,n1476);
not (n1474,n1475);
nand (n1475,n1255,n1316);
nand (n1477,n1478,n1480);
not (n1478,n1479);
nand (n1479,n1220,n1331);
nand (n1481,n1482,n1484);
not (n1482,n1483);
nand (n1483,n1270,n1331);
nor (n1485,n1486,n1499);
and (n1486,n1487,n1246);
nand (n1487,n1488,n1490,n1492,n1497);
nand (n1488,n1282,n1489);
nand (n1490,n1294,n1491);
nor (n1492,n1493,n1495);
and (n1493,n1270,n1494);
and (n1495,n1255,n1496);
nand (n1497,n1220,n1498);
and (n1499,n1500,n1265);
nand (n1500,n1501,n1503,n1505,n1509);
nand (n1501,n1282,n1502);
nand (n1503,n1294,n1504);
nor (n1505,n1506,n1508);
and (n1506,n1270,n1507);
and (n1508,n1255,n1494);
nand (n1509,n1220,n1510);
nor (n1511,n1512,n1515);
and (n1512,n1513,n1514);
and (n1513,n1282,n1316);
and (n1515,n1516,n1518);
not (n1516,n1517);
nand (n1517,n1282,n1331);
nor (n1519,n1520,n1524);
and (n1520,n1521,n1523);
not (n1521,n1522);
nand (n1522,n1294,n1316);
and (n1524,n1525,n1527);
not (n1525,n1526);
nand (n1526,n1294,n1331);
and (n1529,n1460,n1530);
or (n1530,n1531,n1653,n2262);
and (n1531,n1532,n1589);
wire s0n1532,s1n1532,notn1532;
or (n1532,s0n1532,s1n1532);
not(notn1532,n1102);
and (s0n1532,notn1532,n1533);
and (s1n1532,n1102,n1588);
or (n1533,1'b0,n1534,n1547,n1559,n1574);
and (n1534,n1535,n1331);
nand (n1535,n1536,n1541,n1543,n1545);
nor (n1536,n1537,n1539);
and (n1537,n1270,n1538);
and (n1539,n1255,n1540);
nand (n1541,n1220,n1542);
nand (n1543,n1282,n1544);
nand (n1545,n1294,n1546);
and (n1547,n1548,n1316);
nand (n1548,n1549,n1553,n1555,n1557);
nor (n1549,n1550,n1551);
and (n1550,n1270,n1540);
and (n1551,n1255,n1552);
nand (n1553,n1220,n1554);
nand (n1555,n1282,n1556);
nand (n1557,n1294,n1558);
and (n1559,n1560,n1265);
or (n1560,1'b0,n1561,n1565,n1568,n1571);
and (n1561,n1562,n1223);
wire s0n1562,s1n1562,notn1562;
or (n1562,s0n1562,s1n1562);
not(notn1562,n1341);
and (s0n1562,notn1562,n1563);
and (s1n1562,n1341,n1564);
and (n1565,n1566,n1234);
wire s0n1566,s1n1566,notn1566;
or (n1566,s0n1566,s1n1566);
not(notn1566,n1341);
and (s0n1566,notn1566,n1567);
and (s1n1566,n1341,n1563);
and (n1568,n1569,n1354);
wire s0n1569,s1n1569,notn1569;
or (n1569,s0n1569,s1n1569);
not(notn1569,n1341);
and (s0n1569,notn1569,n1570);
and (s1n1569,n1341,n1567);
and (n1571,n1572,n1257);
wire s0n1572,s1n1572,notn1572;
or (n1572,s0n1572,s1n1572);
not(notn1572,n1341);
and (s0n1572,notn1572,n1573);
and (s1n1572,n1341,n1570);
and (n1574,n1575,n1246);
or (n1575,1'b0,n1576,n1579,n1582,n1585);
and (n1576,n1577,n1223);
wire s0n1577,s1n1577,notn1577;
or (n1577,s0n1577,s1n1577);
not(notn1577,n1341);
and (s0n1577,notn1577,n1578);
and (s1n1577,n1341,n1573);
and (n1579,n1580,n1234);
wire s0n1580,s1n1580,notn1580;
or (n1580,s0n1580,s1n1580);
not(notn1580,n1341);
and (s0n1580,notn1580,n1581);
and (s1n1580,n1341,n1578);
and (n1582,n1583,n1354);
wire s0n1583,s1n1583,notn1583;
or (n1583,s0n1583,s1n1583);
not(notn1583,n1341);
and (s0n1583,notn1583,n1584);
and (s1n1583,n1341,n1581);
and (n1585,n1586,n1257);
wire s0n1586,s1n1586,notn1586;
or (n1586,s0n1586,s1n1586);
not(notn1586,n1341);
and (s0n1586,notn1586,n1587);
and (s1n1586,n1341,n1584);
wire s0n1589,s1n1589,notn1589;
or (n1589,s0n1589,s1n1589);
not(notn1589,n1102);
and (s0n1589,notn1589,n1590);
and (s1n1589,n1102,n1652);
or (n1590,1'b0,n1591,n1606,n1620,n1636);
and (n1591,n1592,n1331);
or (n1592,1'b0,n1593,n1597,n1600,n1603);
and (n1593,n1594,n1223);
wire s0n1594,s1n1594,notn1594;
or (n1594,s0n1594,s1n1594);
not(notn1594,n1341);
and (s0n1594,notn1594,n1595);
and (s1n1594,n1341,n1596);
and (n1597,n1598,n1234);
wire s0n1598,s1n1598,notn1598;
or (n1598,s0n1598,s1n1598);
not(notn1598,n1341);
and (s0n1598,notn1598,n1599);
and (s1n1598,n1341,n1595);
and (n1600,n1601,n1354);
wire s0n1601,s1n1601,notn1601;
or (n1601,s0n1601,s1n1601);
not(notn1601,n1341);
and (s0n1601,notn1601,n1602);
and (s1n1601,n1341,n1599);
and (n1603,n1604,n1257);
wire s0n1604,s1n1604,notn1604;
or (n1604,s0n1604,s1n1604);
not(notn1604,n1341);
and (s0n1604,notn1604,n1605);
and (s1n1604,n1341,n1602);
and (n1606,n1607,n1316);
or (n1607,1'b0,n1608,n1611,n1614,n1617);
and (n1608,n1609,n1223);
wire s0n1609,s1n1609,notn1609;
or (n1609,s0n1609,s1n1609);
not(notn1609,n1341);
and (s0n1609,notn1609,n1610);
and (s1n1609,n1341,n1605);
and (n1611,n1612,n1234);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n1341);
and (s0n1612,notn1612,n1613);
and (s1n1612,n1341,n1610);
and (n1614,n1615,n1354);
wire s0n1615,s1n1615,notn1615;
or (n1615,s0n1615,s1n1615);
not(notn1615,n1341);
and (s0n1615,notn1615,n1616);
and (s1n1615,n1341,n1613);
and (n1617,n1618,n1257);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n1341);
and (s0n1618,notn1618,n1619);
and (s1n1618,n1341,n1616);
and (n1620,n1621,n1265);
nand (n1621,n1622,n1627);
nor (n1622,n1623,n1625);
and (n1623,n1282,n1624);
and (n1625,n1294,n1626);
nor (n1627,n1628,n1630);
and (n1628,n1220,n1629);
nand (n1630,n1631,n1634);
or (n1631,n1632,n1396);
not (n1632,n1633);
nand (n1634,n1255,n1635);
and (n1636,n1637,n1246);
nand (n1637,n1638,n1643);
nor (n1638,n1639,n1641);
and (n1639,n1282,n1640);
and (n1641,n1294,n1642);
nor (n1643,n1644,n1649);
nand (n1644,n1645,n1647);
or (n1645,n1646,n1396);
not (n1646,n1635);
nand (n1647,n1255,n1648);
nor (n1649,n1650,n1402);
not (n1650,n1651);
and (n1653,n1589,n1654);
or (n1654,n1655,n1768,n2261);
and (n1655,n1656,n1708);
wire s0n1656,s1n1656,notn1656;
or (n1656,s0n1656,s1n1656);
not(notn1656,n1102);
and (s0n1656,notn1656,n1657);
and (s1n1656,n1102,n1707);
nand (n1657,n1658,n1671,n1676,n1702);
nor (n1658,n1659,n1669);
nand (n1659,n1660,n1665,n1667);
nor (n1660,n1661,n1663);
and (n1661,n1219,n1662);
and (n1663,n1253,n1664);
nand (n1665,n1264,n1666);
nand (n1667,n1269,n1668);
and (n1669,n1274,n1670);
nor (n1671,n1672,n1674);
and (n1672,n1450,n1673);
and (n1674,n1280,n1675);
nor (n1676,n1677,n1690);
and (n1677,n1678,n1316);
nand (n1678,n1679,n1684,n1686,n1688);
nor (n1679,n1680,n1682);
and (n1680,n1270,n1681);
and (n1682,n1255,n1683);
nand (n1684,n1220,n1685);
nand (n1686,n1282,n1687);
nand (n1688,n1294,n1689);
and (n1690,n1691,n1331);
nand (n1691,n1692,n1696,n1698,n1700);
nor (n1692,n1693,n1695);
and (n1693,n1270,n1694);
and (n1695,n1255,n1681);
nand (n1696,n1220,n1697);
nand (n1698,n1282,n1699);
nand (n1700,n1294,n1701);
nor (n1702,n1703,n1705);
and (n1703,n1299,n1704);
and (n1705,n1292,n1706);
wire s0n1708,s1n1708,notn1708;
or (n1708,s0n1708,s1n1708);
not(notn1708,n1102);
and (s0n1708,notn1708,n1709);
and (s1n1708,n1102,n1767);
or (n1709,1'b0,n1710,n1725,n1739,n1752);
and (n1710,n1711,n1331);
or (n1711,1'b0,n1712,n1716,n1719,n1722);
and (n1712,n1713,n1223);
wire s0n1713,s1n1713,notn1713;
or (n1713,s0n1713,s1n1713);
not(notn1713,n1341);
and (s0n1713,notn1713,n1714);
and (s1n1713,n1341,n1715);
and (n1716,n1717,n1234);
wire s0n1717,s1n1717,notn1717;
or (n1717,s0n1717,s1n1717);
not(notn1717,n1341);
and (s0n1717,notn1717,n1718);
and (s1n1717,n1341,n1714);
and (n1719,n1720,n1354);
wire s0n1720,s1n1720,notn1720;
or (n1720,s0n1720,s1n1720);
not(notn1720,n1341);
and (s0n1720,notn1720,n1721);
and (s1n1720,n1341,n1718);
and (n1722,n1723,n1257);
wire s0n1723,s1n1723,notn1723;
or (n1723,s0n1723,s1n1723);
not(notn1723,n1341);
and (s0n1723,notn1723,n1724);
and (s1n1723,n1341,n1721);
and (n1725,n1726,n1316);
or (n1726,1'b0,n1727,n1730,n1733,n1736);
and (n1727,n1728,n1223);
wire s0n1728,s1n1728,notn1728;
or (n1728,s0n1728,s1n1728);
not(notn1728,n1341);
and (s0n1728,notn1728,n1729);
and (s1n1728,n1341,n1724);
and (n1730,n1731,n1234);
wire s0n1731,s1n1731,notn1731;
or (n1731,s0n1731,s1n1731);
not(notn1731,n1341);
and (s0n1731,notn1731,n1732);
and (s1n1731,n1341,n1729);
and (n1733,n1734,n1354);
wire s0n1734,s1n1734,notn1734;
or (n1734,s0n1734,s1n1734);
not(notn1734,n1341);
and (s0n1734,notn1734,n1735);
and (s1n1734,n1341,n1732);
and (n1736,n1737,n1257);
wire s0n1737,s1n1737,notn1737;
or (n1737,s0n1737,s1n1737);
not(notn1737,n1341);
and (s0n1737,notn1737,n1738);
and (s1n1737,n1341,n1735);
and (n1739,n1740,n1265);
nand (n1740,n1741,n1746,n1748,n1750);
nor (n1741,n1742,n1744);
and (n1742,n1255,n1743);
and (n1744,n1270,n1745);
nand (n1746,n1220,n1747);
nand (n1748,n1282,n1749);
nand (n1750,n1294,n1751);
and (n1752,n1753,n1246);
nand (n1753,n1754,n1759);
nor (n1754,n1755,n1757);
and (n1755,n1282,n1756);
and (n1757,n1294,n1758);
nor (n1759,n1760,n1765);
nand (n1760,n1761,n1763);
or (n1761,n1762,n1396);
not (n1762,n1743);
nand (n1763,n1255,n1764);
and (n1765,n1220,n1766);
and (n1768,n1708,n1769);
or (n1769,n1770,n1892,n2260);
and (n1770,n1771,n1828);
wire s0n1771,s1n1771,notn1771;
or (n1771,s0n1771,s1n1771);
not(notn1771,n1102);
and (s0n1771,notn1771,n1772);
and (s1n1771,n1102,n1827);
or (n1772,1'b0,n1773,n1786,n1798,n1813);
and (n1773,n1774,n1331);
nand (n1774,n1775,n1780,n1782,n1784);
nor (n1775,n1776,n1778);
and (n1776,n1270,n1777);
and (n1778,n1255,n1779);
nand (n1780,n1220,n1781);
nand (n1782,n1282,n1783);
nand (n1784,n1294,n1785);
and (n1786,n1787,n1316);
nand (n1787,n1788,n1792,n1794,n1796);
nor (n1788,n1789,n1790);
and (n1789,n1270,n1779);
and (n1790,n1255,n1791);
nand (n1792,n1220,n1793);
nand (n1794,n1282,n1795);
nand (n1796,n1294,n1797);
and (n1798,n1799,n1265);
or (n1799,1'b0,n1800,n1804,n1807,n1810);
and (n1800,n1801,n1223);
wire s0n1801,s1n1801,notn1801;
or (n1801,s0n1801,s1n1801);
not(notn1801,n1341);
and (s0n1801,notn1801,n1802);
and (s1n1801,n1341,n1803);
and (n1804,n1805,n1234);
wire s0n1805,s1n1805,notn1805;
or (n1805,s0n1805,s1n1805);
not(notn1805,n1341);
and (s0n1805,notn1805,n1806);
and (s1n1805,n1341,n1802);
and (n1807,n1808,n1354);
wire s0n1808,s1n1808,notn1808;
or (n1808,s0n1808,s1n1808);
not(notn1808,n1341);
and (s0n1808,notn1808,n1809);
and (s1n1808,n1341,n1806);
and (n1810,n1811,n1257);
wire s0n1811,s1n1811,notn1811;
or (n1811,s0n1811,s1n1811);
not(notn1811,n1341);
and (s0n1811,notn1811,n1812);
and (s1n1811,n1341,n1809);
and (n1813,n1814,n1246);
or (n1814,1'b0,n1815,n1818,n1821,n1824);
and (n1815,n1816,n1223);
wire s0n1816,s1n1816,notn1816;
or (n1816,s0n1816,s1n1816);
not(notn1816,n1341);
and (s0n1816,notn1816,n1817);
and (s1n1816,n1341,n1812);
and (n1818,n1819,n1234);
wire s0n1819,s1n1819,notn1819;
or (n1819,s0n1819,s1n1819);
not(notn1819,n1341);
and (s0n1819,notn1819,n1820);
and (s1n1819,n1341,n1817);
and (n1821,n1822,n1354);
wire s0n1822,s1n1822,notn1822;
or (n1822,s0n1822,s1n1822);
not(notn1822,n1341);
and (s0n1822,notn1822,n1823);
and (s1n1822,n1341,n1820);
and (n1824,n1825,n1257);
wire s0n1825,s1n1825,notn1825;
or (n1825,s0n1825,s1n1825);
not(notn1825,n1341);
and (s0n1825,notn1825,n1826);
and (s1n1825,n1341,n1823);
wire s0n1828,s1n1828,notn1828;
or (n1828,s0n1828,s1n1828);
not(notn1828,n1102);
and (s0n1828,notn1828,n1829);
and (s1n1828,n1102,n1891);
or (n1829,1'b0,n1830,n1845,n1859,n1875);
and (n1830,n1831,n1331);
or (n1831,1'b0,n1832,n1836,n1839,n1842);
and (n1832,n1833,n1223);
wire s0n1833,s1n1833,notn1833;
or (n1833,s0n1833,s1n1833);
not(notn1833,n1341);
and (s0n1833,notn1833,n1834);
and (s1n1833,n1341,n1835);
and (n1836,n1837,n1234);
wire s0n1837,s1n1837,notn1837;
or (n1837,s0n1837,s1n1837);
not(notn1837,n1341);
and (s0n1837,notn1837,n1838);
and (s1n1837,n1341,n1834);
and (n1839,n1840,n1354);
wire s0n1840,s1n1840,notn1840;
or (n1840,s0n1840,s1n1840);
not(notn1840,n1341);
and (s0n1840,notn1840,n1841);
and (s1n1840,n1341,n1838);
and (n1842,n1843,n1257);
wire s0n1843,s1n1843,notn1843;
or (n1843,s0n1843,s1n1843);
not(notn1843,n1341);
and (s0n1843,notn1843,n1844);
and (s1n1843,n1341,n1841);
and (n1845,n1846,n1316);
or (n1846,1'b0,n1847,n1850,n1853,n1856);
and (n1847,n1848,n1223);
wire s0n1848,s1n1848,notn1848;
or (n1848,s0n1848,s1n1848);
not(notn1848,n1341);
and (s0n1848,notn1848,n1849);
and (s1n1848,n1341,n1844);
and (n1850,n1851,n1234);
wire s0n1851,s1n1851,notn1851;
or (n1851,s0n1851,s1n1851);
not(notn1851,n1341);
and (s0n1851,notn1851,n1852);
and (s1n1851,n1341,n1849);
and (n1853,n1854,n1354);
wire s0n1854,s1n1854,notn1854;
or (n1854,s0n1854,s1n1854);
not(notn1854,n1341);
and (s0n1854,notn1854,n1855);
and (s1n1854,n1341,n1852);
and (n1856,n1857,n1257);
wire s0n1857,s1n1857,notn1857;
or (n1857,s0n1857,s1n1857);
not(notn1857,n1341);
and (s0n1857,notn1857,n1858);
and (s1n1857,n1341,n1855);
and (n1859,n1860,n1265);
nand (n1860,n1861,n1866);
nor (n1861,n1862,n1864);
and (n1862,n1282,n1863);
and (n1864,n1294,n1865);
nor (n1866,n1867,n1869);
and (n1867,n1220,n1868);
nand (n1869,n1870,n1873);
or (n1870,n1871,n1396);
not (n1871,n1872);
nand (n1873,n1255,n1874);
and (n1875,n1876,n1246);
nand (n1876,n1877,n1882);
nor (n1877,n1878,n1880);
and (n1878,n1282,n1879);
and (n1880,n1294,n1881);
nor (n1882,n1883,n1888);
nand (n1883,n1884,n1886);
or (n1884,n1885,n1396);
not (n1885,n1874);
nand (n1886,n1255,n1887);
nor (n1888,n1889,n1402);
not (n1889,n1890);
and (n1892,n1828,n1893);
or (n1893,n1894,n2015,n2259);
and (n1894,n1895,n1952);
wire s0n1895,s1n1895,notn1895;
or (n1895,s0n1895,s1n1895);
not(notn1895,n1102);
and (s0n1895,notn1895,n1896);
and (s1n1895,n1102,n1951);
or (n1896,1'b0,n1897,n1910,n1922,n1937);
and (n1897,n1898,n1331);
nand (n1898,n1899,n1904,n1906,n1908);
nor (n1899,n1900,n1902);
and (n1900,n1270,n1901);
and (n1902,n1255,n1903);
nand (n1904,n1220,n1905);
nand (n1906,n1282,n1907);
nand (n1908,n1294,n1909);
and (n1910,n1911,n1316);
nand (n1911,n1912,n1916,n1918,n1920);
nor (n1912,n1913,n1914);
and (n1913,n1270,n1903);
and (n1914,n1255,n1915);
nand (n1916,n1220,n1917);
nand (n1918,n1282,n1919);
nand (n1920,n1294,n1921);
and (n1922,n1923,n1265);
or (n1923,1'b0,n1924,n1928,n1931,n1934);
and (n1924,n1925,n1223);
wire s0n1925,s1n1925,notn1925;
or (n1925,s0n1925,s1n1925);
not(notn1925,n1341);
and (s0n1925,notn1925,n1926);
and (s1n1925,n1341,n1927);
and (n1928,n1929,n1234);
wire s0n1929,s1n1929,notn1929;
or (n1929,s0n1929,s1n1929);
not(notn1929,n1341);
and (s0n1929,notn1929,n1930);
and (s1n1929,n1341,n1926);
and (n1931,n1932,n1354);
wire s0n1932,s1n1932,notn1932;
or (n1932,s0n1932,s1n1932);
not(notn1932,n1341);
and (s0n1932,notn1932,n1933);
and (s1n1932,n1341,n1930);
and (n1934,n1935,n1257);
wire s0n1935,s1n1935,notn1935;
or (n1935,s0n1935,s1n1935);
not(notn1935,n1341);
and (s0n1935,notn1935,n1936);
and (s1n1935,n1341,n1933);
and (n1937,n1938,n1246);
or (n1938,1'b0,n1939,n1942,n1945,n1948);
and (n1939,n1940,n1223);
wire s0n1940,s1n1940,notn1940;
or (n1940,s0n1940,s1n1940);
not(notn1940,n1341);
and (s0n1940,notn1940,n1941);
and (s1n1940,n1341,n1936);
and (n1942,n1943,n1234);
wire s0n1943,s1n1943,notn1943;
or (n1943,s0n1943,s1n1943);
not(notn1943,n1341);
and (s0n1943,notn1943,n1944);
and (s1n1943,n1341,n1941);
and (n1945,n1946,n1354);
wire s0n1946,s1n1946,notn1946;
or (n1946,s0n1946,s1n1946);
not(notn1946,n1341);
and (s0n1946,notn1946,n1947);
and (s1n1946,n1341,n1944);
and (n1948,n1949,n1257);
wire s0n1949,s1n1949,notn1949;
or (n1949,s0n1949,s1n1949);
not(notn1949,n1341);
and (s0n1949,notn1949,n1950);
and (s1n1949,n1341,n1947);
wire s0n1952,s1n1952,notn1952;
or (n1952,s0n1952,s1n1952);
not(notn1952,n1102);
and (s0n1952,notn1952,n1953);
and (s1n1952,n1102,n2014);
or (n1953,1'b0,n1954,n1969,n1983,n1999);
and (n1954,n1955,n1331);
or (n1955,1'b0,n1956,n1960,n1963,n1966);
and (n1956,n1957,n1223);
wire s0n1957,s1n1957,notn1957;
or (n1957,s0n1957,s1n1957);
not(notn1957,n1341);
and (s0n1957,notn1957,n1958);
and (s1n1957,n1341,n1959);
and (n1960,n1961,n1234);
wire s0n1961,s1n1961,notn1961;
or (n1961,s0n1961,s1n1961);
not(notn1961,n1341);
and (s0n1961,notn1961,n1962);
and (s1n1961,n1341,n1958);
and (n1963,n1964,n1354);
wire s0n1964,s1n1964,notn1964;
or (n1964,s0n1964,s1n1964);
not(notn1964,n1341);
and (s0n1964,notn1964,n1965);
and (s1n1964,n1341,n1962);
and (n1966,n1967,n1257);
wire s0n1967,s1n1967,notn1967;
or (n1967,s0n1967,s1n1967);
not(notn1967,n1341);
and (s0n1967,notn1967,n1968);
and (s1n1967,n1341,n1965);
and (n1969,n1970,n1316);
or (n1970,1'b0,n1971,n1974,n1977,n1980);
and (n1971,n1972,n1223);
wire s0n1972,s1n1972,notn1972;
or (n1972,s0n1972,s1n1972);
not(notn1972,n1341);
and (s0n1972,notn1972,n1973);
and (s1n1972,n1341,n1968);
and (n1974,n1975,n1234);
wire s0n1975,s1n1975,notn1975;
or (n1975,s0n1975,s1n1975);
not(notn1975,n1341);
and (s0n1975,notn1975,n1976);
and (s1n1975,n1341,n1973);
and (n1977,n1978,n1354);
wire s0n1978,s1n1978,notn1978;
or (n1978,s0n1978,s1n1978);
not(notn1978,n1341);
and (s0n1978,notn1978,n1979);
and (s1n1978,n1341,n1976);
and (n1980,n1981,n1257);
wire s0n1981,s1n1981,notn1981;
or (n1981,s0n1981,s1n1981);
not(notn1981,n1341);
and (s0n1981,notn1981,n1982);
and (s1n1981,n1341,n1979);
and (n1983,n1984,n1265);
nand (n1984,n1985,n1990);
nor (n1985,n1986,n1988);
and (n1986,n1282,n1987);
and (n1988,n1294,n1989);
nor (n1990,n1991,n1993);
and (n1991,n1220,n1992);
nand (n1993,n1994,n1997);
or (n1994,n1995,n1396);
not (n1995,n1996);
nand (n1997,n1255,n1998);
and (n1999,n2000,n1246);
nand (n2000,n2001,n2006);
nor (n2001,n2002,n2004);
and (n2002,n1282,n2003);
and (n2004,n1294,n2005);
nor (n2006,n2007,n2009);
and (n2007,n1220,n2008);
nand (n2009,n2010,n2012);
or (n2010,n2011,n1396);
not (n2011,n1998);
nand (n2012,n1255,n2013);
and (n2015,n1952,n2016);
or (n2016,n2017,n2136,n2258);
and (n2017,n2018,n2075);
wire s0n2018,s1n2018,notn2018;
or (n2018,s0n2018,s1n2018);
not(notn2018,n1102);
and (s0n2018,notn2018,n2019);
and (s1n2018,n1102,n2074);
or (n2019,1'b0,n2020,n2033,n2045,n2060);
and (n2020,n2021,n1331);
nand (n2021,n2022,n2024,n2026,n2031);
nand (n2022,n1282,n2023);
nand (n2024,n1294,n2025);
nor (n2026,n2027,n2029);
and (n2027,n1270,n2028);
and (n2029,n1255,n2030);
nand (n2031,n1220,n2032);
and (n2033,n2034,n1316);
nand (n2034,n2035,n2037,n2039,n2043);
nand (n2035,n1282,n2036);
nand (n2037,n1294,n2038);
nor (n2039,n2040,n2041);
and (n2040,n1270,n2030);
and (n2041,n1255,n2042);
nand (n2043,n1220,n2044);
and (n2045,n2046,n1265);
or (n2046,1'b0,n2047,n2051,n2054,n2057);
and (n2047,n2048,n1223);
wire s0n2048,s1n2048,notn2048;
or (n2048,s0n2048,s1n2048);
not(notn2048,n1341);
and (s0n2048,notn2048,n2049);
and (s1n2048,n1341,n2050);
and (n2051,n2052,n1234);
wire s0n2052,s1n2052,notn2052;
or (n2052,s0n2052,s1n2052);
not(notn2052,n1341);
and (s0n2052,notn2052,n2053);
and (s1n2052,n1341,n2049);
and (n2054,n2055,n1354);
wire s0n2055,s1n2055,notn2055;
or (n2055,s0n2055,s1n2055);
not(notn2055,n1341);
and (s0n2055,notn2055,n2056);
and (s1n2055,n1341,n2053);
and (n2057,n2058,n1257);
wire s0n2058,s1n2058,notn2058;
or (n2058,s0n2058,s1n2058);
not(notn2058,n1341);
and (s0n2058,notn2058,n2059);
and (s1n2058,n1341,n2056);
and (n2060,n2061,n1246);
or (n2061,1'b0,n2062,n2065,n2068,n2071);
and (n2062,n2063,n1223);
wire s0n2063,s1n2063,notn2063;
or (n2063,s0n2063,s1n2063);
not(notn2063,n1341);
and (s0n2063,notn2063,n2064);
and (s1n2063,n1341,n2059);
and (n2065,n2066,n1234);
wire s0n2066,s1n2066,notn2066;
or (n2066,s0n2066,s1n2066);
not(notn2066,n1341);
and (s0n2066,notn2066,n2067);
and (s1n2066,n1341,n2064);
and (n2068,n2069,n1354);
wire s0n2069,s1n2069,notn2069;
or (n2069,s0n2069,s1n2069);
not(notn2069,n1341);
and (s0n2069,notn2069,n2070);
and (s1n2069,n1341,n2067);
and (n2071,n2072,n1257);
wire s0n2072,s1n2072,notn2072;
or (n2072,s0n2072,s1n2072);
not(notn2072,n1341);
and (s0n2072,notn2072,n2073);
and (s1n2072,n1341,n2070);
wire s0n2075,s1n2075,notn2075;
or (n2075,s0n2075,s1n2075);
not(notn2075,n1102);
and (s0n2075,notn2075,n2076);
and (s1n2075,n1102,n2135);
or (n2076,1'b0,n2077,n2092,n2106,n2120);
and (n2077,n2078,n1331);
or (n2078,1'b0,n2079,n2083,n2086,n2089);
and (n2079,n2080,n1223);
wire s0n2080,s1n2080,notn2080;
or (n2080,s0n2080,s1n2080);
not(notn2080,n1341);
and (s0n2080,notn2080,n2081);
and (s1n2080,n1341,n2082);
and (n2083,n2084,n1234);
wire s0n2084,s1n2084,notn2084;
or (n2084,s0n2084,s1n2084);
not(notn2084,n1341);
and (s0n2084,notn2084,n2085);
and (s1n2084,n1341,n2081);
and (n2086,n2087,n1354);
wire s0n2087,s1n2087,notn2087;
or (n2087,s0n2087,s1n2087);
not(notn2087,n1341);
and (s0n2087,notn2087,n2088);
and (s1n2087,n1341,n2085);
and (n2089,n2090,n1257);
wire s0n2090,s1n2090,notn2090;
or (n2090,s0n2090,s1n2090);
not(notn2090,n1341);
and (s0n2090,notn2090,n2091);
and (s1n2090,n1341,n2088);
and (n2092,n2093,n1316);
or (n2093,1'b0,n2094,n2097,n2100,n2103);
and (n2094,n2095,n1223);
wire s0n2095,s1n2095,notn2095;
or (n2095,s0n2095,s1n2095);
not(notn2095,n1341);
and (s0n2095,notn2095,n2096);
and (s1n2095,n1341,n2091);
and (n2097,n2098,n1234);
wire s0n2098,s1n2098,notn2098;
or (n2098,s0n2098,s1n2098);
not(notn2098,n1341);
and (s0n2098,notn2098,n2099);
and (s1n2098,n1341,n2096);
and (n2100,n2101,n1354);
wire s0n2101,s1n2101,notn2101;
or (n2101,s0n2101,s1n2101);
not(notn2101,n1341);
and (s0n2101,notn2101,n2102);
and (s1n2101,n1341,n2099);
and (n2103,n2104,n1257);
wire s0n2104,s1n2104,notn2104;
or (n2104,s0n2104,s1n2104);
not(notn2104,n1341);
and (s0n2104,notn2104,n2105);
and (s1n2104,n1341,n2102);
not (n2106,n2107);
nand (n2107,n2108,n1265);
nand (n2108,n2109,n2114,n2116,n2118);
nor (n2109,n2110,n2112);
and (n2110,n1270,n2111);
and (n2112,n1255,n2113);
nand (n2114,n1282,n2115);
nand (n2116,n1294,n2117);
nand (n2118,n1220,n2119);
not (n2120,n2121);
or (n2121,n1247,n2122);
not (n2122,n2123);
nand (n2123,n2124,n2129,n2131,n2133);
nor (n2124,n2125,n2126);
and (n2125,n1270,n2113);
nor (n2126,n2127,n1256);
not (n2127,n2128);
nand (n2129,n1282,n2130);
nand (n2131,n1294,n2132);
nand (n2133,n1220,n2134);
and (n2136,n2075,n2137);
and (n2137,n2138,n2195);
wire s0n2138,s1n2138,notn2138;
or (n2138,s0n2138,s1n2138);
not(notn2138,n1102);
and (s0n2138,notn2138,n2139);
and (s1n2138,n1102,n2194);
or (n2139,1'b0,n2140,n2153,n2165,n2180);
and (n2140,n2141,n1331);
nand (n2141,n2142,n2147,n2149,n2151);
nor (n2142,n2143,n2145);
and (n2143,n1255,n2144);
and (n2145,n1270,n2146);
nand (n2147,n1220,n2148);
nand (n2149,n1282,n2150);
nand (n2151,n1294,n2152);
and (n2153,n2154,n1316);
nand (n2154,n2155,n2159,n2161,n2163);
nor (n2155,n2156,n2158);
and (n2156,n1255,n2157);
and (n2158,n1270,n2144);
nand (n2159,n1220,n2160);
nand (n2161,n1282,n2162);
nand (n2163,n1294,n2164);
and (n2165,n2166,n1265);
or (n2166,1'b0,n2167,n2171,n2174,n2177);
and (n2167,n2168,n1223);
wire s0n2168,s1n2168,notn2168;
or (n2168,s0n2168,s1n2168);
not(notn2168,n1341);
and (s0n2168,notn2168,n2169);
and (s1n2168,n1341,n2170);
and (n2171,n2172,n1234);
wire s0n2172,s1n2172,notn2172;
or (n2172,s0n2172,s1n2172);
not(notn2172,n1341);
and (s0n2172,notn2172,n2173);
and (s1n2172,n1341,n2169);
and (n2174,n2175,n1354);
wire s0n2175,s1n2175,notn2175;
or (n2175,s0n2175,s1n2175);
not(notn2175,n1341);
and (s0n2175,notn2175,n2176);
and (s1n2175,n1341,n2173);
and (n2177,n2178,n1257);
wire s0n2178,s1n2178,notn2178;
or (n2178,s0n2178,s1n2178);
not(notn2178,n1341);
and (s0n2178,notn2178,n2179);
and (s1n2178,n1341,n2176);
and (n2180,n2181,n1246);
or (n2181,1'b0,n2182,n2185,n2188,n2191);
and (n2182,n2183,n1223);
wire s0n2183,s1n2183,notn2183;
or (n2183,s0n2183,s1n2183);
not(notn2183,n1341);
and (s0n2183,notn2183,n2184);
and (s1n2183,n1341,n2179);
and (n2185,n2186,n1234);
wire s0n2186,s1n2186,notn2186;
or (n2186,s0n2186,s1n2186);
not(notn2186,n1341);
and (s0n2186,notn2186,n2187);
and (s1n2186,n1341,n2184);
and (n2188,n2189,n1354);
wire s0n2189,s1n2189,notn2189;
or (n2189,s0n2189,s1n2189);
not(notn2189,n1341);
and (s0n2189,notn2189,n2190);
and (s1n2189,n1341,n2187);
and (n2191,n2192,n1257);
wire s0n2192,s1n2192,notn2192;
or (n2192,s0n2192,s1n2192);
not(notn2192,n1341);
and (s0n2192,notn2192,n2193);
and (s1n2192,n1341,n2190);
wire s0n2195,s1n2195,notn2195;
or (n2195,s0n2195,s1n2195);
not(notn2195,n1102);
and (s0n2195,notn2195,n2196);
and (s1n2195,n1102,n2257);
or (n2196,1'b0,n2197,n2212,n2226,n2242);
and (n2197,n2198,n1331);
or (n2198,1'b0,n2199,n2203,n2206,n2209);
and (n2199,n2200,n1223);
wire s0n2200,s1n2200,notn2200;
or (n2200,s0n2200,s1n2200);
not(notn2200,n1341);
and (s0n2200,notn2200,n2201);
and (s1n2200,n1341,n2202);
and (n2203,n2204,n1234);
wire s0n2204,s1n2204,notn2204;
or (n2204,s0n2204,s1n2204);
not(notn2204,n1341);
and (s0n2204,notn2204,n2205);
and (s1n2204,n1341,n2201);
and (n2206,n2207,n1354);
wire s0n2207,s1n2207,notn2207;
or (n2207,s0n2207,s1n2207);
not(notn2207,n1341);
and (s0n2207,notn2207,n2208);
and (s1n2207,n1341,n2205);
and (n2209,n2210,n1257);
wire s0n2210,s1n2210,notn2210;
or (n2210,s0n2210,s1n2210);
not(notn2210,n1341);
and (s0n2210,notn2210,n2211);
and (s1n2210,n1341,n2208);
and (n2212,n2213,n1316);
or (n2213,1'b0,n2214,n2217,n2220,n2223);
and (n2214,n2215,n1223);
wire s0n2215,s1n2215,notn2215;
or (n2215,s0n2215,s1n2215);
not(notn2215,n1341);
and (s0n2215,notn2215,n2216);
and (s1n2215,n1341,n2211);
and (n2217,n2218,n1234);
wire s0n2218,s1n2218,notn2218;
or (n2218,s0n2218,s1n2218);
not(notn2218,n1341);
and (s0n2218,notn2218,n2219);
and (s1n2218,n1341,n2216);
and (n2220,n2221,n1354);
wire s0n2221,s1n2221,notn2221;
or (n2221,s0n2221,s1n2221);
not(notn2221,n1341);
and (s0n2221,notn2221,n2222);
and (s1n2221,n1341,n2219);
and (n2223,n2224,n1257);
wire s0n2224,s1n2224,notn2224;
or (n2224,s0n2224,s1n2224);
not(notn2224,n1341);
and (s0n2224,notn2224,n2225);
and (s1n2224,n1341,n2222);
and (n2226,n2227,n1265);
nand (n2227,n2228,n2233);
nor (n2228,n2229,n2231);
and (n2229,n1294,n2230);
and (n2231,n1282,n2232);
nor (n2233,n2234,n2236);
and (n2234,n1220,n2235);
nand (n2236,n2237,n2240);
or (n2237,n2238,n1396);
not (n2238,n2239);
nand (n2240,n1255,n2241);
and (n2242,n2243,n1246);
nand (n2243,n2244,n2249);
nor (n2244,n2245,n2247);
and (n2245,n1294,n2246);
and (n2247,n1282,n2248);
nor (n2249,n2250,n2252);
and (n2250,n1220,n2251);
nand (n2252,n2253,n2255);
or (n2253,n2254,n1396);
not (n2254,n2241);
nand (n2255,n1255,n2256);
and (n2258,n2018,n2137);
and (n2259,n1895,n2016);
and (n2260,n1771,n1893);
and (n2261,n1656,n1769);
and (n2262,n1532,n1654);
and (n2263,n1407,n1530);
and (n2264,n1213,n1405);
and (n2265,n1206,n1211);
and (n2266,n1199,n1204);
xor (n2267,n2268,n3959);
xor (n2268,n2269,n3848);
xor (n2269,n2270,n3235);
xor (n2270,n2271,n2276);
xor (n2271,n2272,n2274);
wire s0n2272,s1n2272,notn2272;
or (n2272,s0n2272,s1n2272);
not(notn2272,n1102);
and (s0n2272,notn2272,1'b0);
and (s1n2272,n1102,n2273);
wire s0n2274,s1n2274,notn2274;
or (n2274,s0n2274,s1n2274);
not(notn2274,n1102);
and (s0n2274,notn2274,1'b0);
and (s1n2274,n1102,n2275);
or (n2276,n2277,n2381,n3234);
and (n2277,n2278,n2329);
wire s0n2278,s1n2278,notn2278;
or (n2278,s0n2278,s1n2278);
not(notn2278,n1102);
and (s0n2278,notn2278,n2279);
and (s1n2278,n1102,n2328);
nand (n2279,n2280,n2306,n2318,n2323);
nor (n2280,n2281,n2294);
and (n2281,n2282,n1316);
nand (n2282,n2283,n2288,n2290,n2292);
nor (n2283,n2284,n2286);
and (n2284,n1270,n2285);
and (n2286,n1255,n2287);
nand (n2288,n1220,n2289);
nand (n2290,n1282,n2291);
nand (n2292,n1294,n2293);
and (n2294,n2295,n1331);
nand (n2295,n2296,n2300,n2302,n2304);
nor (n2296,n2297,n2299);
and (n2297,n1270,n2298);
and (n2299,n1255,n2285);
nand (n2300,n1220,n2301);
nand (n2302,n1282,n2303);
nand (n2304,n1294,n2305);
nor (n2306,n2307,n2309);
and (n2307,n1274,n2308);
nand (n2309,n2310,n2312,n2314,n2316);
nand (n2310,n1264,n2311);
nand (n2312,n1219,n2313);
nand (n2314,n1269,n2315);
nand (n2316,n1253,n2317);
nor (n2318,n2319,n2321);
and (n2319,n1280,n2320);
and (n2321,n1292,n2322);
nor (n2323,n2324,n2326);
and (n2324,n1450,n2325);
and (n2326,n1299,n2327);
wire s0n2329,s1n2329,notn2329;
or (n2329,s0n2329,s1n2329);
not(notn2329,n1102);
and (s0n2329,notn2329,n2330);
and (s1n2329,n1102,n2380);
nand (n2330,n2331,n2344,n2370,n2375);
nor (n2331,n2332,n2342);
nand (n2332,n2333,n2338,n2340);
nor (n2333,n2334,n2336);
and (n2334,n1219,n2335);
and (n2336,n1253,n2337);
nand (n2338,n1264,n2339);
nand (n2340,n1269,n2341);
and (n2342,n1274,n2343);
nor (n2344,n2345,n2358);
and (n2345,n2346,n1316);
nand (n2346,n2347,n2352,n2354,n2356);
nor (n2347,n2348,n2350);
and (n2348,n1270,n2349);
and (n2350,n1255,n2351);
nand (n2352,n1220,n2353);
nand (n2354,n1282,n2355);
nand (n2356,n1294,n2357);
and (n2358,n2359,n1331);
nand (n2359,n2360,n2364,n2366,n2368);
nor (n2360,n2361,n2363);
and (n2361,n1270,n2362);
and (n2363,n1255,n2349);
nand (n2364,n1220,n2365);
nand (n2366,n1282,n2367);
nand (n2368,n1294,n2369);
nor (n2370,n2371,n2373);
and (n2371,n1450,n2372);
and (n2373,n1280,n2374);
nor (n2375,n2376,n2378);
and (n2376,n1299,n2377);
and (n2378,n1292,n2379);
and (n2381,n2329,n2382);
or (n2382,n2383,n2501,n3233);
and (n2383,n2384,n2436);
wire s0n2384,s1n2384,notn2384;
or (n2384,s0n2384,s1n2384);
not(notn2384,n1102);
and (s0n2384,notn2384,n2385);
and (s1n2384,n1102,n2435);
nand (n2385,n2386,n2412,n2425,n2430);
nor (n2386,n2387,n2400);
and (n2387,n2388,n1316);
nand (n2388,n2389,n2394,n2396,n2398);
nor (n2389,n2390,n2392);
and (n2390,n1270,n2391);
and (n2392,n1255,n2393);
nand (n2394,n1220,n2395);
nand (n2396,n1282,n2397);
nand (n2398,n1294,n2399);
and (n2400,n2401,n1331);
nand (n2401,n2402,n2406,n2408,n2410);
nor (n2402,n2403,n2405);
and (n2403,n1270,n2404);
and (n2405,n1255,n2391);
nand (n2406,n1220,n2407);
nand (n2408,n1282,n2409);
nand (n2410,n1294,n2411);
nor (n2412,n2413,n2415);
and (n2413,n1274,n2414);
nand (n2415,n2416,n2421,n2423);
nor (n2416,n2417,n2419);
and (n2417,n1253,n2418);
and (n2419,n1219,n2420);
nand (n2421,n1269,n2422);
nand (n2423,n1264,n2424);
nor (n2425,n2426,n2428);
and (n2426,n1450,n2427);
and (n2428,n1280,n2429);
nor (n2430,n2431,n2433);
and (n2431,n1299,n2432);
and (n2433,n1292,n2434);
wire s0n2436,s1n2436,notn2436;
or (n2436,s0n2436,s1n2436);
not(notn2436,n1102);
and (s0n2436,notn2436,n2437);
and (s1n2436,n1102,n2500);
or (n2437,1'b0,n2438,n2455,n2471,n2486);
and (n2438,n2439,n1331);
nand (n2439,n2440,n2445);
nor (n2440,n2441,n2443);
and (n2441,n1282,n2442);
and (n2443,n1294,n2444);
nor (n2445,n2446,n2452);
nand (n2446,n2447,n2450);
or (n2447,n2448,n1396);
not (n2448,n2449);
nand (n2450,n1255,n2451);
nor (n2452,n2453,n1402);
not (n2453,n2454);
and (n2455,n2456,n1316);
nand (n2456,n2457,n2462);
nor (n2457,n2458,n2460);
and (n2458,n1282,n2459);
and (n2460,n1294,n2461);
nor (n2462,n2463,n2468);
nand (n2463,n2464,n2466);
or (n2464,n2465,n1396);
not (n2465,n2451);
nand (n2466,n1255,n2467);
nor (n2468,n2469,n1402);
not (n2469,n2470);
and (n2471,n2472,n1265);
or (n2472,1'b0,n2473,n2477,n2480,n2483);
and (n2473,n2474,n1223);
wire s0n2474,s1n2474,notn2474;
or (n2474,s0n2474,s1n2474);
not(notn2474,n1341);
and (s0n2474,notn2474,n2475);
and (s1n2474,n1341,n2476);
and (n2477,n2478,n1234);
wire s0n2478,s1n2478,notn2478;
or (n2478,s0n2478,s1n2478);
not(notn2478,n1341);
and (s0n2478,notn2478,n2479);
and (s1n2478,n1341,n2475);
and (n2480,n2481,n1354);
wire s0n2481,s1n2481,notn2481;
or (n2481,s0n2481,s1n2481);
not(notn2481,n1341);
and (s0n2481,notn2481,n2482);
and (s1n2481,n1341,n2479);
and (n2483,n2484,n1257);
wire s0n2484,s1n2484,notn2484;
or (n2484,s0n2484,s1n2484);
not(notn2484,n1341);
and (s0n2484,notn2484,n2485);
and (s1n2484,n1341,n2482);
and (n2486,n2487,n1246);
or (n2487,1'b0,n2488,n2491,n2494,n2497);
and (n2488,n2489,n1223);
wire s0n2489,s1n2489,notn2489;
or (n2489,s0n2489,s1n2489);
not(notn2489,n1341);
and (s0n2489,notn2489,n2490);
and (s1n2489,n1341,n2485);
and (n2491,n2492,n1234);
wire s0n2492,s1n2492,notn2492;
or (n2492,s0n2492,s1n2492);
not(notn2492,n1341);
and (s0n2492,notn2492,n2493);
and (s1n2492,n1341,n2490);
and (n2494,n2495,n1354);
wire s0n2495,s1n2495,notn2495;
or (n2495,s0n2495,s1n2495);
not(notn2495,n1341);
and (s0n2495,notn2495,n2496);
and (s1n2495,n1341,n2493);
and (n2497,n2498,n1257);
wire s0n2498,s1n2498,notn2498;
or (n2498,s0n2498,s1n2498);
not(notn2498,n1341);
and (s0n2498,notn2498,n2499);
and (s1n2498,n1341,n2496);
and (n2501,n2436,n2502);
or (n2502,n2503,n2609,n3232);
and (n2503,n2504,n2557);
wire s0n2504,s1n2504,notn2504;
or (n2504,s0n2504,s1n2504);
not(notn2504,n1102);
and (s0n2504,notn2504,n2505);
and (s1n2504,n1102,n2556);
nand (n2505,n2506,n2520,n2546,n2551);
nor (n2506,n2507,n2509);
and (n2507,n1274,n2508);
nand (n2509,n2510,n2516,n2518);
nor (n2510,n2511,n2513);
and (n2511,n1219,n2512);
nor (n2513,n2514,n1254);
not (n2514,n2515);
nand (n2516,n1269,n2517);
nand (n2518,n1264,n2519);
nor (n2520,n2521,n2534);
and (n2521,n2522,n1316);
nand (n2522,n2523,n2525,n2527,n2532);
nand (n2523,n1282,n2524);
nand (n2525,n1294,n2526);
nor (n2527,n2528,n2530);
and (n2528,n1270,n2529);
and (n2530,n1255,n2531);
nand (n2532,n1220,n2533);
and (n2534,n2535,n1331);
nand (n2535,n2536,n2538,n2540,n2544);
nand (n2536,n1282,n2537);
nand (n2538,n1294,n2539);
nor (n2540,n2541,n2543);
and (n2541,n1270,n2542);
and (n2543,n1255,n2529);
nand (n2544,n1220,n2545);
nor (n2546,n2547,n2549);
and (n2547,n1450,n2548);
and (n2549,n1280,n2550);
nor (n2551,n2552,n2554);
and (n2552,n1299,n2553);
and (n2554,n1292,n2555);
wire s0n2557,s1n2557,notn2557;
or (n2557,s0n2557,s1n2557);
not(notn2557,n1102);
and (s0n2557,notn2557,n2558);
and (s1n2557,n1102,n2608);
nand (n2558,n2559,n2572,n2588,n2603);
nor (n2559,n2560,n2562);
and (n2560,n1274,n2561);
nand (n2562,n2563,n2565,n2570);
nand (n2563,n1219,n2564);
nor (n2565,n2566,n2568);
and (n2566,n1264,n2567);
and (n2568,n1253,n2569);
nand (n2570,n1269,n2571);
nor (n2572,n2573,n2586);
and (n2573,n2574,n1331);
nand (n2574,n2575,n2580,n2582,n2584);
nor (n2575,n2576,n2578);
and (n2576,n1270,n2577);
and (n2578,n1255,n2579);
nand (n2580,n1220,n2581);
nand (n2582,n1282,n2583);
nand (n2584,n1294,n2585);
and (n2586,n1450,n2587);
nor (n2588,n2589,n2601);
and (n2589,n2590,n1316);
nand (n2590,n2591,n2595,n2597,n2599);
nor (n2591,n2592,n2593);
and (n2592,n1270,n2579);
and (n2593,n1255,n2594);
nand (n2595,n1220,n2596);
nand (n2597,n1282,n2598);
nand (n2599,n1294,n2600);
and (n2601,n1292,n2602);
nor (n2603,n2604,n2606);
and (n2604,n1280,n2605);
and (n2606,n1299,n2607);
and (n2609,n2557,n2610);
or (n2610,n2611,n2737,n3231);
and (n2611,n2612,n2677);
wire s0n2612,s1n2612,notn2612;
or (n2612,s0n2612,s1n2612);
not(notn2612,n1102);
and (s0n2612,notn2612,n2613);
and (s1n2612,n1102,n2676);
or (n2613,1'b0,n2614,n2631,n2647,n2662);
and (n2614,n2615,n1331);
nand (n2615,n2616,n2621);
nor (n2616,n2617,n2619);
and (n2617,n1294,n2618);
and (n2619,n1282,n2620);
nor (n2621,n2622,n2628);
nand (n2622,n2623,n2626);
or (n2623,n2624,n1396);
not (n2624,n2625);
nand (n2626,n1255,n2627);
nor (n2628,n2629,n1402);
not (n2629,n2630);
and (n2631,n2632,n1316);
nand (n2632,n2633,n2638);
nor (n2633,n2634,n2636);
and (n2634,n1294,n2635);
and (n2636,n1282,n2637);
nor (n2638,n2639,n2644);
nand (n2639,n2640,n2642);
or (n2640,n2641,n1396);
not (n2641,n2627);
nand (n2642,n1255,n2643);
nor (n2644,n1402,n2645);
not (n2645,n2646);
and (n2647,n2648,n1265);
or (n2648,1'b0,n2649,n2653,n2656,n2659);
and (n2649,n2650,n1223);
wire s0n2650,s1n2650,notn2650;
or (n2650,s0n2650,s1n2650);
not(notn2650,n1341);
and (s0n2650,notn2650,n2651);
and (s1n2650,n1341,n2652);
and (n2653,n2654,n1234);
wire s0n2654,s1n2654,notn2654;
or (n2654,s0n2654,s1n2654);
not(notn2654,n1341);
and (s0n2654,notn2654,n2655);
and (s1n2654,n1341,n2651);
and (n2656,n2657,n1354);
wire s0n2657,s1n2657,notn2657;
or (n2657,s0n2657,s1n2657);
not(notn2657,n1341);
and (s0n2657,notn2657,n2658);
and (s1n2657,n1341,n2655);
and (n2659,n2660,n1257);
wire s0n2660,s1n2660,notn2660;
or (n2660,s0n2660,s1n2660);
not(notn2660,n1341);
and (s0n2660,notn2660,n2661);
and (s1n2660,n1341,n2658);
and (n2662,n2663,n1246);
or (n2663,1'b0,n2664,n2667,n2670,n2673);
and (n2664,n2665,n1223);
wire s0n2665,s1n2665,notn2665;
or (n2665,s0n2665,s1n2665);
not(notn2665,n1341);
and (s0n2665,notn2665,n2666);
and (s1n2665,n1341,n2661);
and (n2667,n2668,n1234);
wire s0n2668,s1n2668,notn2668;
or (n2668,s0n2668,s1n2668);
not(notn2668,n1341);
and (s0n2668,notn2668,n2669);
and (s1n2668,n1341,n2666);
and (n2670,n2671,n1354);
wire s0n2671,s1n2671,notn2671;
or (n2671,s0n2671,s1n2671);
not(notn2671,n1341);
and (s0n2671,notn2671,n2672);
and (s1n2671,n1341,n2669);
and (n2673,n2674,n1257);
wire s0n2674,s1n2674,notn2674;
or (n2674,s0n2674,s1n2674);
not(notn2674,n1341);
and (s0n2674,notn2674,n2675);
and (s1n2674,n1341,n2672);
wire s0n2677,s1n2677,notn2677;
or (n2677,s0n2677,s1n2677);
not(notn2677,n1102);
and (s0n2677,notn2677,n2678);
and (s1n2677,n1102,n2736);
or (n2678,1'b0,n2679,n2692,n2707,n2722);
and (n2679,n2680,n1331);
nand (n2680,n2681,n2686,n2688,n2690);
nor (n2681,n2682,n2684);
and (n2682,n1270,n2683);
and (n2684,n1255,n2685);
nand (n2686,n1220,n2687);
nand (n2688,n1282,n2689);
nand (n2690,n1294,n2691);
and (n2692,n2693,n1316);
nand (n2693,n2694,n2699);
nor (n2694,n2695,n2697);
and (n2695,n1282,n2696);
and (n2697,n1294,n2698);
nor (n2699,n2700,n2705);
nand (n2700,n2701,n2703);
or (n2701,n2702,n1396);
not (n2702,n2685);
nand (n2703,n1255,n2704);
and (n2705,n1220,n2706);
and (n2707,n2708,n1265);
or (n2708,1'b0,n2709,n2713,n2716,n2719);
and (n2709,n2710,n1223);
wire s0n2710,s1n2710,notn2710;
or (n2710,s0n2710,s1n2710);
not(notn2710,n1341);
and (s0n2710,notn2710,n2711);
and (s1n2710,n1341,n2712);
and (n2713,n2714,n1234);
wire s0n2714,s1n2714,notn2714;
or (n2714,s0n2714,s1n2714);
not(notn2714,n1341);
and (s0n2714,notn2714,n2715);
and (s1n2714,n1341,n2711);
and (n2716,n2717,n1354);
wire s0n2717,s1n2717,notn2717;
or (n2717,s0n2717,s1n2717);
not(notn2717,n1341);
and (s0n2717,notn2717,n2718);
and (s1n2717,n1341,n2715);
and (n2719,n2720,n1257);
wire s0n2720,s1n2720,notn2720;
or (n2720,s0n2720,s1n2720);
not(notn2720,n1341);
and (s0n2720,notn2720,n2721);
and (s1n2720,n1341,n2718);
and (n2722,n2723,n1246);
or (n2723,1'b0,n2724,n2727,n2730,n2733);
and (n2724,n2725,n1223);
wire s0n2725,s1n2725,notn2725;
or (n2725,s0n2725,s1n2725);
not(notn2725,n1341);
and (s0n2725,notn2725,n2726);
and (s1n2725,n1341,n2721);
and (n2727,n2728,n1234);
wire s0n2728,s1n2728,notn2728;
or (n2728,s0n2728,s1n2728);
not(notn2728,n1341);
and (s0n2728,notn2728,n2729);
and (s1n2728,n1341,n2726);
and (n2730,n2731,n1354);
wire s0n2731,s1n2731,notn2731;
or (n2731,s0n2731,s1n2731);
not(notn2731,n1341);
and (s0n2731,notn2731,n2732);
and (s1n2731,n1341,n2729);
and (n2733,n2734,n1257);
wire s0n2734,s1n2734,notn2734;
or (n2734,s0n2734,s1n2734);
not(notn2734,n1341);
and (s0n2734,notn2734,n2735);
and (s1n2734,n1341,n2732);
and (n2737,n2677,n2738);
or (n2738,n2739,n2862,n3230);
and (n2739,n2740,n2805);
wire s0n2740,s1n2740,notn2740;
or (n2740,s0n2740,s1n2740);
not(notn2740,n1102);
and (s0n2740,notn2740,n2741);
and (s1n2740,n1102,n2804);
or (n2741,1'b0,n2742,n2759,n2775,n2790);
and (n2742,n2743,n1331);
nand (n2743,n2744,n2749);
nor (n2744,n2745,n2747);
and (n2745,n1282,n2746);
and (n2747,n1294,n2748);
nor (n2749,n2750,n2756);
nand (n2750,n2751,n2754);
or (n2751,n2752,n1396);
not (n2752,n2753);
nand (n2754,n1255,n2755);
nor (n2756,n2757,n1402);
not (n2757,n2758);
and (n2759,n2760,n1316);
nand (n2760,n2761,n2766);
nor (n2761,n2762,n2764);
and (n2762,n1282,n2763);
and (n2764,n1294,n2765);
nor (n2766,n2767,n2772);
nand (n2767,n2768,n2770);
or (n2768,n2769,n1396);
not (n2769,n2755);
nand (n2770,n1255,n2771);
nor (n2772,n2773,n1402);
not (n2773,n2774);
and (n2775,n2776,n1265);
or (n2776,1'b0,n2777,n2781,n2784,n2787);
and (n2777,n2778,n1223);
wire s0n2778,s1n2778,notn2778;
or (n2778,s0n2778,s1n2778);
not(notn2778,n1341);
and (s0n2778,notn2778,n2779);
and (s1n2778,n1341,n2780);
and (n2781,n2782,n1234);
wire s0n2782,s1n2782,notn2782;
or (n2782,s0n2782,s1n2782);
not(notn2782,n1341);
and (s0n2782,notn2782,n2783);
and (s1n2782,n1341,n2779);
and (n2784,n2785,n1354);
wire s0n2785,s1n2785,notn2785;
or (n2785,s0n2785,s1n2785);
not(notn2785,n1341);
and (s0n2785,notn2785,n2786);
and (s1n2785,n1341,n2783);
and (n2787,n2788,n1257);
wire s0n2788,s1n2788,notn2788;
or (n2788,s0n2788,s1n2788);
not(notn2788,n1341);
and (s0n2788,notn2788,n2789);
and (s1n2788,n1341,n2786);
and (n2790,n2791,n1246);
or (n2791,1'b0,n2792,n2795,n2798,n2801);
and (n2792,n2793,n1223);
wire s0n2793,s1n2793,notn2793;
or (n2793,s0n2793,s1n2793);
not(notn2793,n1341);
and (s0n2793,notn2793,n2794);
and (s1n2793,n1341,n2789);
and (n2795,n2796,n1234);
wire s0n2796,s1n2796,notn2796;
or (n2796,s0n2796,s1n2796);
not(notn2796,n1341);
and (s0n2796,notn2796,n2797);
and (s1n2796,n1341,n2794);
and (n2798,n2799,n1354);
wire s0n2799,s1n2799,notn2799;
or (n2799,s0n2799,s1n2799);
not(notn2799,n1341);
and (s0n2799,notn2799,n2800);
and (s1n2799,n1341,n2797);
and (n2801,n2802,n1257);
wire s0n2802,s1n2802,notn2802;
or (n2802,s0n2802,s1n2802);
not(notn2802,n1341);
and (s0n2802,notn2802,n2803);
and (s1n2802,n1341,n2800);
wire s0n2805,s1n2805,notn2805;
or (n2805,s0n2805,s1n2805);
not(notn2805,n1102);
and (s0n2805,notn2805,n2806);
and (s1n2805,n1102,n2861);
or (n2806,1'b0,n2807,n2820,n2832,n2847);
and (n2807,n2808,n1331);
nand (n2808,n2809,n2811,n2813,n2818);
nand (n2809,n1282,n2810);
nand (n2811,n1294,n2812);
nor (n2813,n2814,n2816);
and (n2814,n1270,n2815);
and (n2816,n1255,n2817);
nand (n2818,n1220,n2819);
and (n2820,n2821,n1316);
nand (n2821,n2822,n2824,n2826,n2830);
nand (n2822,n1282,n2823);
nand (n2824,n1294,n2825);
nor (n2826,n2827,n2828);
and (n2827,n1270,n2817);
and (n2828,n1255,n2829);
nand (n2830,n1220,n2831);
and (n2832,n2833,n1265);
or (n2833,1'b0,n2834,n2838,n2841,n2844);
and (n2834,n2835,n1223);
wire s0n2835,s1n2835,notn2835;
or (n2835,s0n2835,s1n2835);
not(notn2835,n1341);
and (s0n2835,notn2835,n2836);
and (s1n2835,n1341,n2837);
and (n2838,n2839,n1234);
wire s0n2839,s1n2839,notn2839;
or (n2839,s0n2839,s1n2839);
not(notn2839,n1341);
and (s0n2839,notn2839,n2840);
and (s1n2839,n1341,n2836);
and (n2841,n2842,n1354);
wire s0n2842,s1n2842,notn2842;
or (n2842,s0n2842,s1n2842);
not(notn2842,n1341);
and (s0n2842,notn2842,n2843);
and (s1n2842,n1341,n2840);
and (n2844,n2845,n1257);
wire s0n2845,s1n2845,notn2845;
or (n2845,s0n2845,s1n2845);
not(notn2845,n1341);
and (s0n2845,notn2845,n2846);
and (s1n2845,n1341,n2843);
and (n2847,n2848,n1246);
or (n2848,1'b0,n2849,n2852,n2855,n2858);
and (n2849,n2850,n1223);
wire s0n2850,s1n2850,notn2850;
or (n2850,s0n2850,s1n2850);
not(notn2850,n1341);
and (s0n2850,notn2850,n2851);
and (s1n2850,n1341,n2846);
and (n2852,n2853,n1234);
wire s0n2853,s1n2853,notn2853;
or (n2853,s0n2853,s1n2853);
not(notn2853,n1341);
and (s0n2853,notn2853,n2854);
and (s1n2853,n1341,n2851);
and (n2855,n2856,n1354);
wire s0n2856,s1n2856,notn2856;
or (n2856,s0n2856,s1n2856);
not(notn2856,n1341);
and (s0n2856,notn2856,n2857);
and (s1n2856,n1341,n2854);
and (n2858,n2859,n1257);
wire s0n2859,s1n2859,notn2859;
or (n2859,s0n2859,s1n2859);
not(notn2859,n1341);
and (s0n2859,notn2859,n2860);
and (s1n2859,n1341,n2857);
and (n2862,n2805,n2863);
or (n2863,n2864,n2979,n3229);
and (n2864,n2865,n2922);
wire s0n2865,s1n2865,notn2865;
or (n2865,s0n2865,s1n2865);
not(notn2865,n1102);
and (s0n2865,notn2865,n2866);
and (s1n2865,n1102,n2921);
or (n2866,1'b0,n2867,n2880,n2892,n2907);
and (n2867,n2868,n1331);
nand (n2868,n2869,n2874,n2876,n2878);
nor (n2869,n2870,n2872);
and (n2870,n1270,n2871);
and (n2872,n1255,n2873);
nand (n2874,n1220,n2875);
nand (n2876,n1282,n2877);
nand (n2878,n1294,n2879);
and (n2880,n2881,n1316);
nand (n2881,n2882,n2886,n2888,n2890);
nor (n2882,n2883,n2884);
and (n2883,n1270,n2873);
and (n2884,n1255,n2885);
nand (n2886,n1220,n2887);
nand (n2888,n1282,n2889);
nand (n2890,n1294,n2891);
and (n2892,n2893,n1265);
or (n2893,1'b0,n2894,n2898,n2901,n2904);
and (n2894,n2895,n1223);
wire s0n2895,s1n2895,notn2895;
or (n2895,s0n2895,s1n2895);
not(notn2895,n1341);
and (s0n2895,notn2895,n2896);
and (s1n2895,n1341,n2897);
and (n2898,n2899,n1234);
wire s0n2899,s1n2899,notn2899;
or (n2899,s0n2899,s1n2899);
not(notn2899,n1341);
and (s0n2899,notn2899,n2900);
and (s1n2899,n1341,n2896);
and (n2901,n2902,n1354);
wire s0n2902,s1n2902,notn2902;
or (n2902,s0n2902,s1n2902);
not(notn2902,n1341);
and (s0n2902,notn2902,n2903);
and (s1n2902,n1341,n2900);
and (n2904,n2905,n1257);
wire s0n2905,s1n2905,notn2905;
or (n2905,s0n2905,s1n2905);
not(notn2905,n1341);
and (s0n2905,notn2905,n2906);
and (s1n2905,n1341,n2903);
and (n2907,n2908,n1246);
or (n2908,1'b0,n2909,n2912,n2915,n2918);
and (n2909,n2910,n1223);
wire s0n2910,s1n2910,notn2910;
or (n2910,s0n2910,s1n2910);
not(notn2910,n1341);
and (s0n2910,notn2910,n2911);
and (s1n2910,n1341,n2906);
and (n2912,n2913,n1234);
wire s0n2913,s1n2913,notn2913;
or (n2913,s0n2913,s1n2913);
not(notn2913,n1341);
and (s0n2913,notn2913,n2914);
and (s1n2913,n1341,n2911);
and (n2915,n2916,n1354);
wire s0n2916,s1n2916,notn2916;
or (n2916,s0n2916,s1n2916);
not(notn2916,n1341);
and (s0n2916,notn2916,n2917);
and (s1n2916,n1341,n2914);
and (n2918,n2919,n1257);
wire s0n2919,s1n2919,notn2919;
or (n2919,s0n2919,s1n2919);
not(notn2919,n1341);
and (s0n2919,notn2919,n2920);
and (s1n2919,n1341,n2917);
wire s0n2922,s1n2922,notn2922;
or (n2922,s0n2922,s1n2922);
not(notn2922,n1102);
and (s0n2922,notn2922,n2923);
and (s1n2922,n1102,n2978);
or (n2923,1'b0,n2924,n2937,n2949,n2964);
and (n2924,n2925,n1331);
nand (n2925,n2926,n2931,n2933,n2935);
nor (n2926,n2927,n2929);
and (n2927,n1270,n2928);
and (n2929,n1255,n2930);
nand (n2931,n1220,n2932);
nand (n2933,n1282,n2934);
nand (n2935,n1294,n2936);
and (n2937,n2938,n1316);
nand (n2938,n2939,n2943,n2945,n2947);
nor (n2939,n2940,n2942);
and (n2940,n1255,n2941);
and (n2942,n1270,n2930);
nand (n2943,n1220,n2944);
nand (n2945,n1282,n2946);
nand (n2947,n1294,n2948);
and (n2949,n2950,n1265);
or (n2950,1'b0,n2951,n2955,n2958,n2961);
and (n2951,n2952,n1223);
wire s0n2952,s1n2952,notn2952;
or (n2952,s0n2952,s1n2952);
not(notn2952,n1341);
and (s0n2952,notn2952,n2953);
and (s1n2952,n1341,n2954);
and (n2955,n2956,n1234);
wire s0n2956,s1n2956,notn2956;
or (n2956,s0n2956,s1n2956);
not(notn2956,n1341);
and (s0n2956,notn2956,n2957);
and (s1n2956,n1341,n2953);
and (n2958,n2959,n1354);
wire s0n2959,s1n2959,notn2959;
or (n2959,s0n2959,s1n2959);
not(notn2959,n1341);
and (s0n2959,notn2959,n2960);
and (s1n2959,n1341,n2957);
and (n2961,n2962,n1257);
wire s0n2962,s1n2962,notn2962;
or (n2962,s0n2962,s1n2962);
not(notn2962,n1341);
and (s0n2962,notn2962,n2963);
and (s1n2962,n1341,n2960);
and (n2964,n2965,n1246);
or (n2965,1'b0,n2966,n2969,n2972,n2975);
and (n2966,n2967,n1223);
wire s0n2967,s1n2967,notn2967;
or (n2967,s0n2967,s1n2967);
not(notn2967,n1341);
and (s0n2967,notn2967,n2968);
and (s1n2967,n1341,n2963);
and (n2969,n2970,n1234);
wire s0n2970,s1n2970,notn2970;
or (n2970,s0n2970,s1n2970);
not(notn2970,n1341);
and (s0n2970,notn2970,n2971);
and (s1n2970,n1341,n2968);
and (n2972,n2973,n1354);
wire s0n2973,s1n2973,notn2973;
or (n2973,s0n2973,s1n2973);
not(notn2973,n1341);
and (s0n2973,notn2973,n2974);
and (s1n2973,n1341,n2971);
and (n2975,n2976,n1257);
wire s0n2976,s1n2976,notn2976;
or (n2976,s0n2976,s1n2976);
not(notn2976,n1341);
and (s0n2976,notn2976,n2977);
and (s1n2976,n1341,n2974);
and (n2979,n2922,n2980);
or (n2980,n2981,n3103,n3228);
and (n2981,n2982,n3042);
wire s0n2982,s1n2982,notn2982;
or (n2982,s0n2982,s1n2982);
not(notn2982,n1102);
and (s0n2982,notn2982,n2983);
and (s1n2982,n1102,n3041);
or (n2983,1'b0,n2984,n2999,n3012,n3027);
and (n2984,n2985,n1331);
or (n2985,1'b0,n2986,n2990,n2993,n2996);
and (n2986,n2987,n1223);
wire s0n2987,s1n2987,notn2987;
or (n2987,s0n2987,s1n2987);
not(notn2987,n1341);
and (s0n2987,notn2987,n2988);
and (s1n2987,n1341,n2989);
and (n2990,n2991,n1234);
wire s0n2991,s1n2991,notn2991;
or (n2991,s0n2991,s1n2991);
not(notn2991,n1341);
and (s0n2991,notn2991,n2992);
and (s1n2991,n1341,n2988);
and (n2993,n2994,n1354);
wire s0n2994,s1n2994,notn2994;
or (n2994,s0n2994,s1n2994);
not(notn2994,n1341);
and (s0n2994,notn2994,n2995);
and (s1n2994,n1341,n2992);
and (n2996,n2997,n1257);
wire s0n2997,s1n2997,notn2997;
or (n2997,s0n2997,s1n2997);
not(notn2997,n1341);
and (s0n2997,notn2997,n2998);
and (s1n2997,n1341,n2995);
and (n2999,n3000,n1316);
nand (n3000,n3001,n3006);
nor (n3001,n3002,n3004);
and (n3002,n1294,n3003);
and (n3004,n1282,n3005);
and (n3006,n3007,n3008,n3010);
nand (n3007,n1270,n2998);
nand (n3008,n1220,n3009);
nand (n3010,n1255,n3011);
and (n3012,n3013,n1265);
or (n3013,1'b0,n3014,n3018,n3021,n3024);
and (n3014,n3015,n1223);
wire s0n3015,s1n3015,notn3015;
or (n3015,s0n3015,s1n3015);
not(notn3015,n1341);
and (s0n3015,notn3015,n3016);
and (s1n3015,n1341,n3017);
and (n3018,n3019,n1234);
wire s0n3019,s1n3019,notn3019;
or (n3019,s0n3019,s1n3019);
not(notn3019,n1341);
and (s0n3019,notn3019,n3020);
and (s1n3019,n1341,n3016);
and (n3021,n3022,n1354);
wire s0n3022,s1n3022,notn3022;
or (n3022,s0n3022,s1n3022);
not(notn3022,n1341);
and (s0n3022,notn3022,n3023);
and (s1n3022,n1341,n3020);
and (n3024,n3025,n1257);
wire s0n3025,s1n3025,notn3025;
or (n3025,s0n3025,s1n3025);
not(notn3025,n1341);
and (s0n3025,notn3025,n3026);
and (s1n3025,n1341,n3023);
and (n3027,n3028,n1246);
or (n3028,1'b0,n3029,n3032,n3035,n3038);
and (n3029,n3030,n1223);
wire s0n3030,s1n3030,notn3030;
or (n3030,s0n3030,s1n3030);
not(notn3030,n1341);
and (s0n3030,notn3030,n3031);
and (s1n3030,n1341,n3026);
and (n3032,n3033,n1234);
wire s0n3033,s1n3033,notn3033;
or (n3033,s0n3033,s1n3033);
not(notn3033,n1341);
and (s0n3033,notn3033,n3034);
and (s1n3033,n1341,n3031);
and (n3035,n3036,n1354);
wire s0n3036,s1n3036,notn3036;
or (n3036,s0n3036,s1n3036);
not(notn3036,n1341);
and (s0n3036,notn3036,n3037);
and (s1n3036,n1341,n3034);
and (n3038,n3039,n1257);
wire s0n3039,s1n3039,notn3039;
or (n3039,s0n3039,s1n3039);
not(notn3039,n1341);
and (s0n3039,notn3039,n3040);
and (s1n3039,n1341,n3037);
wire s0n3042,s1n3042,notn3042;
or (n3042,s0n3042,s1n3042);
not(notn3042,n1102);
and (s0n3042,notn3042,n3043);
and (s1n3042,n1102,n3102);
or (n3043,1'b0,n3044,n3060,n3073,n3088);
not (n3044,n3045);
or (n3045,n3046,n3047);
not (n3046,n1331);
not (n3047,n3048);
nand (n3048,n3049,n3054,n3056,n3058);
nor (n3049,n3050,n3052);
and (n3050,n1270,n3051);
and (n3052,n1255,n3053);
nand (n3054,n1220,n3055);
nand (n3056,n1282,n3057);
nand (n3058,n1294,n3059);
not (n3060,n3061);
nand (n3061,n3062,n1316);
nand (n3062,n3063,n3067,n3069,n3071);
nor (n3063,n3064,n3065);
and (n3064,n1270,n3053);
and (n3065,n1255,n3066);
nand (n3067,n1220,n3068);
nand (n3069,n1282,n3070);
nand (n3071,n1294,n3072);
and (n3073,n3074,n1265);
or (n3074,1'b0,n3075,n3079,n3082,n3085);
and (n3075,n3076,n1223);
wire s0n3076,s1n3076,notn3076;
or (n3076,s0n3076,s1n3076);
not(notn3076,n1341);
and (s0n3076,notn3076,n3077);
and (s1n3076,n1341,n3078);
and (n3079,n3080,n1234);
wire s0n3080,s1n3080,notn3080;
or (n3080,s0n3080,s1n3080);
not(notn3080,n1341);
and (s0n3080,notn3080,n3081);
and (s1n3080,n1341,n3077);
and (n3082,n3083,n1354);
wire s0n3083,s1n3083,notn3083;
or (n3083,s0n3083,s1n3083);
not(notn3083,n1341);
and (s0n3083,notn3083,n3084);
and (s1n3083,n1341,n3081);
and (n3085,n3086,n1257);
wire s0n3086,s1n3086,notn3086;
or (n3086,s0n3086,s1n3086);
not(notn3086,n1341);
and (s0n3086,notn3086,n3087);
and (s1n3086,n1341,n3084);
and (n3088,n3089,n1246);
or (n3089,1'b0,n3090,n3093,n3096,n3099);
and (n3090,n3091,n1223);
wire s0n3091,s1n3091,notn3091;
or (n3091,s0n3091,s1n3091);
not(notn3091,n1341);
and (s0n3091,notn3091,n3092);
and (s1n3091,n1341,n3087);
and (n3093,n3094,n1234);
wire s0n3094,s1n3094,notn3094;
or (n3094,s0n3094,s1n3094);
not(notn3094,n1341);
and (s0n3094,notn3094,n3095);
and (s1n3094,n1341,n3092);
and (n3096,n3097,n1354);
wire s0n3097,s1n3097,notn3097;
or (n3097,s0n3097,s1n3097);
not(notn3097,n1341);
and (s0n3097,notn3097,n3098);
and (s1n3097,n1341,n3095);
and (n3099,n3100,n1257);
wire s0n3100,s1n3100,notn3100;
or (n3100,s0n3100,s1n3100);
not(notn3100,n1341);
and (s0n3100,notn3100,n3101);
and (s1n3100,n1341,n3098);
and (n3103,n3042,n3104);
and (n3104,n3105,n3165);
wire s0n3105,s1n3105,notn3105;
or (n3105,s0n3105,s1n3105);
not(notn3105,n1102);
and (s0n3105,notn3105,n3106);
and (s1n3105,n1102,n3164);
or (n3106,1'b0,n3107,n3122,n3135,n3150);
not (n3107,n3108);
nand (n3108,n3109,n1331);
nand (n3109,n3110,n3115);
nor (n3110,n3111,n3113);
and (n3111,n1294,n3112);
and (n3113,n1282,n3114);
and (n3115,n3116,n3118,n3120);
nand (n3116,n1270,n3117);
nand (n3118,n1220,n3119);
nand (n3120,n1255,n3121);
and (n3122,n3123,n1316);
nand (n3123,n3124,n3129);
nor (n3124,n3125,n3127);
and (n3125,n1282,n3126);
and (n3127,n1294,n3128);
and (n3129,n3130,n3131,n3133);
nand (n3130,n1270,n3121);
nand (n3131,n1220,n3132);
nand (n3133,n1255,n3134);
and (n3135,n3136,n1265);
or (n3136,1'b0,n3137,n3141,n3144,n3147);
and (n3137,n3138,n1223);
wire s0n3138,s1n3138,notn3138;
or (n3138,s0n3138,s1n3138);
not(notn3138,n1341);
and (s0n3138,notn3138,n3139);
and (s1n3138,n1341,n3140);
and (n3141,n3142,n1234);
wire s0n3142,s1n3142,notn3142;
or (n3142,s0n3142,s1n3142);
not(notn3142,n1341);
and (s0n3142,notn3142,n3143);
and (s1n3142,n1341,n3139);
and (n3144,n3145,n1354);
wire s0n3145,s1n3145,notn3145;
or (n3145,s0n3145,s1n3145);
not(notn3145,n1341);
and (s0n3145,notn3145,n3146);
and (s1n3145,n1341,n3143);
and (n3147,n3148,n1257);
wire s0n3148,s1n3148,notn3148;
or (n3148,s0n3148,s1n3148);
not(notn3148,n1341);
and (s0n3148,notn3148,n3149);
and (s1n3148,n1341,n3146);
and (n3150,n3151,n1246);
or (n3151,1'b0,n3152,n3155,n3158,n3161);
and (n3152,n3153,n1223);
wire s0n3153,s1n3153,notn3153;
or (n3153,s0n3153,s1n3153);
not(notn3153,n1341);
and (s0n3153,notn3153,n3154);
and (s1n3153,n1341,n3149);
and (n3155,n3156,n1234);
wire s0n3156,s1n3156,notn3156;
or (n3156,s0n3156,s1n3156);
not(notn3156,n1341);
and (s0n3156,notn3156,n3157);
and (s1n3156,n1341,n3154);
and (n3158,n3159,n1354);
wire s0n3159,s1n3159,notn3159;
or (n3159,s0n3159,s1n3159);
not(notn3159,n1341);
and (s0n3159,notn3159,n3160);
and (s1n3159,n1341,n3157);
and (n3161,n3162,n1257);
wire s0n3162,s1n3162,notn3162;
or (n3162,s0n3162,s1n3162);
not(notn3162,n1341);
and (s0n3162,notn3162,n3163);
and (s1n3162,n1341,n3160);
wire s0n3165,s1n3165,notn3165;
or (n3165,s0n3165,s1n3165);
not(notn3165,n1102);
and (s0n3165,notn3165,n3166);
and (s1n3165,n1102,n3227);
or (n3166,1'b0,n3167,n3183,n3198,n3213);
and (n3167,n3168,n1331);
nand (n3168,n3169,n3174);
nor (n3169,n3170,n3172);
and (n3170,n1282,n3171);
and (n3172,n1294,n3173);
nor (n3174,n3175,n3177);
and (n3175,n1220,n3176);
nand (n3177,n3178,n3181);
or (n3178,n3179,n1396);
not (n3179,n3180);
nand (n3181,n1255,n3182);
and (n3183,n3184,n1316);
nand (n3184,n3185,n3190);
nor (n3185,n3186,n3188);
and (n3186,n1282,n3187);
and (n3188,n1294,n3189);
nor (n3190,n3191,n3193);
and (n3191,n1220,n3192);
nand (n3193,n3194,n3196);
or (n3194,n3195,n1396);
not (n3195,n3182);
nand (n3196,n1255,n3197);
and (n3198,n3199,n1265);
or (n3199,1'b0,n3200,n3204,n3207,n3210);
and (n3200,n3201,n1223);
wire s0n3201,s1n3201,notn3201;
or (n3201,s0n3201,s1n3201);
not(notn3201,n1341);
and (s0n3201,notn3201,n3202);
and (s1n3201,n1341,n3203);
and (n3204,n3205,n1234);
wire s0n3205,s1n3205,notn3205;
or (n3205,s0n3205,s1n3205);
not(notn3205,n1341);
and (s0n3205,notn3205,n3206);
and (s1n3205,n1341,n3202);
and (n3207,n3208,n1354);
wire s0n3208,s1n3208,notn3208;
or (n3208,s0n3208,s1n3208);
not(notn3208,n1341);
and (s0n3208,notn3208,n3209);
and (s1n3208,n1341,n3206);
and (n3210,n3211,n1257);
wire s0n3211,s1n3211,notn3211;
or (n3211,s0n3211,s1n3211);
not(notn3211,n1341);
and (s0n3211,notn3211,n3212);
and (s1n3211,n1341,n3209);
and (n3213,n3214,n1246);
or (n3214,1'b0,n3215,n3218,n3221,n3224);
and (n3215,n3216,n1223);
wire s0n3216,s1n3216,notn3216;
or (n3216,s0n3216,s1n3216);
not(notn3216,n1341);
and (s0n3216,notn3216,n3217);
and (s1n3216,n1341,n3212);
and (n3218,n3219,n1234);
wire s0n3219,s1n3219,notn3219;
or (n3219,s0n3219,s1n3219);
not(notn3219,n1341);
and (s0n3219,notn3219,n3220);
and (s1n3219,n1341,n3217);
and (n3221,n3222,n1354);
wire s0n3222,s1n3222,notn3222;
or (n3222,s0n3222,s1n3222);
not(notn3222,n1341);
and (s0n3222,notn3222,n3223);
and (s1n3222,n1341,n3220);
and (n3224,n3225,n1257);
wire s0n3225,s1n3225,notn3225;
or (n3225,s0n3225,s1n3225);
not(notn3225,n1341);
and (s0n3225,notn3225,n3226);
and (s1n3225,n1341,n3223);
and (n3228,n2982,n3104);
and (n3229,n2865,n2980);
and (n3230,n2740,n2863);
and (n3231,n2612,n2738);
and (n3232,n2504,n2610);
and (n3233,n2384,n2502);
and (n3234,n2278,n2382);
not (n3235,n3236);
nor (n3236,n3237,n3847);
and (n3237,n3238,n3244);
not (n3238,n3239);
xor (n3239,n3240,n3242);
wire s0n3240,s1n3240,notn3240;
or (n3240,s0n3240,s1n3240);
not(notn3240,n1102);
and (s0n3240,notn3240,1'b0);
and (s1n3240,n1102,n3241);
wire s0n3242,s1n3242,notn3242;
or (n3242,s0n3242,s1n3242);
not(notn3242,n1102);
and (s0n3242,notn3242,1'b0);
and (s1n3242,n1102,n3243);
not (n3244,n3245);
nand (n3245,n3246,n3839);
or (n3246,n3247,n3405);
not (n3247,n3248);
and (n3248,n3249,n3394);
nand (n3249,n3250,n3390);
not (n3250,n3251);
nand (n3251,n3252,n3388);
or (n3252,n3253,n3320);
not (n3253,n3254);
and (n3254,n3255,n3289);
wire s0n3255,s1n3255,notn3255;
or (n3255,s0n3255,s1n3255);
not(notn3255,n1102);
and (s0n3255,notn3255,n3256);
and (s1n3255,n1102,n3288);
or (n3256,1'b0,n3257,n3258,n3259,n3274);
and (n3257,n1500,n1331);
and (n3258,n1487,n1316);
and (n3259,n3260,n1265);
or (n3260,1'b0,n3261,n3265,n3268,n3271);
and (n3261,n3262,n1223);
wire s0n3262,s1n3262,notn3262;
or (n3262,s0n3262,s1n3262);
not(notn3262,n1341);
and (s0n3262,notn3262,n3263);
and (s1n3262,n1341,n3264);
and (n3265,n3266,n1234);
wire s0n3266,s1n3266,notn3266;
or (n3266,s0n3266,s1n3266);
not(notn3266,n1341);
and (s0n3266,notn3266,n3267);
and (s1n3266,n1341,n3263);
and (n3268,n3269,n1354);
wire s0n3269,s1n3269,notn3269;
or (n3269,s0n3269,s1n3269);
not(notn3269,n1341);
and (s0n3269,notn3269,n3270);
and (s1n3269,n1341,n3267);
and (n3271,n3272,n1257);
wire s0n3272,s1n3272,notn3272;
or (n3272,s0n3272,s1n3272);
not(notn3272,n1341);
and (s0n3272,notn3272,n3273);
and (s1n3272,n1341,n3270);
and (n3274,n3275,n1246);
or (n3275,1'b0,n3276,n3279,n3282,n3285);
and (n3276,n3277,n1223);
wire s0n3277,s1n3277,notn3277;
or (n3277,s0n3277,s1n3277);
not(notn3277,n1341);
and (s0n3277,notn3277,n3278);
and (s1n3277,n1341,n3273);
and (n3279,n3280,n1234);
wire s0n3280,s1n3280,notn3280;
or (n3280,s0n3280,s1n3280);
not(notn3280,n1341);
and (s0n3280,notn3280,n3281);
and (s1n3280,n1341,n3278);
and (n3282,n3283,n1354);
wire s0n3283,s1n3283,notn3283;
or (n3283,s0n3283,s1n3283);
not(notn3283,n1341);
and (s0n3283,notn3283,n3284);
and (s1n3283,n1341,n3281);
and (n3285,n3286,n1257);
wire s0n3286,s1n3286,notn3286;
or (n3286,s0n3286,s1n3286);
not(notn3286,n1341);
and (s0n3286,notn3286,n3287);
and (s1n3286,n1341,n3284);
or (n3289,n3290,n3292);
and (n3290,n1102,n3291);
nand (n3292,n3293,n3306,n3307,n3308);
nand (n3293,n3294,n1331);
nand (n3294,n3295,n3297,n3299,n3304);
nand (n3295,n1282,n3296);
nand (n3297,n1294,n3298);
nor (n3299,n3300,n3302);
and (n3300,n1270,n3301);
and (n3302,n1255,n3303);
nand (n3304,n1220,n3305);
nand (n3306,n1424,n1246);
nand (n3307,n1437,n1265);
nand (n3308,n3309,n1316);
nand (n3309,n3310,n3312,n3314,n3318);
nand (n3310,n1282,n3311);
nand (n3312,n1294,n3313);
nor (n3314,n3315,n3316);
and (n3315,n1270,n3303);
and (n3316,n1255,n3317);
nand (n3318,n1220,n3319);
not (n3320,n3321);
nand (n3321,n3322,n3357);
not (n3322,n3323);
wire s0n3323,s1n3323,notn3323;
or (n3323,s0n3323,s1n3323);
not(notn3323,n1102);
and (s0n3323,notn3323,n3324);
and (s1n3323,n1102,n3356);
or (n3324,1'b0,n3325,n3326,n3327,n3342);
and (n3325,n1373,n1331);
and (n3326,n1386,n1316);
and (n3327,n3328,n1265);
or (n3328,1'b0,n3329,n3333,n3336,n3339);
and (n3329,n3330,n1223);
wire s0n3330,s1n3330,notn3330;
or (n3330,s0n3330,s1n3330);
not(notn3330,n1341);
and (s0n3330,notn3330,n3331);
and (s1n3330,n1341,n3332);
and (n3333,n3334,n1234);
wire s0n3334,s1n3334,notn3334;
or (n3334,s0n3334,s1n3334);
not(notn3334,n1341);
and (s0n3334,notn3334,n3335);
and (s1n3334,n1341,n3331);
and (n3336,n3337,n1354);
wire s0n3337,s1n3337,notn3337;
or (n3337,s0n3337,s1n3337);
not(notn3337,n1341);
and (s0n3337,notn3337,n3338);
and (s1n3337,n1341,n3335);
and (n3339,n3340,n1257);
wire s0n3340,s1n3340,notn3340;
or (n3340,s0n3340,s1n3340);
not(notn3340,n1341);
and (s0n3340,notn3340,n3341);
and (s1n3340,n1341,n3338);
and (n3342,n3343,n1246);
or (n3343,1'b0,n3344,n3347,n3350,n3353);
and (n3344,n3345,n1223);
wire s0n3345,s1n3345,notn3345;
or (n3345,s0n3345,s1n3345);
not(notn3345,n1341);
and (s0n3345,notn3345,n3346);
and (s1n3345,n1341,n3341);
and (n3347,n3348,n1234);
wire s0n3348,s1n3348,notn3348;
or (n3348,s0n3348,s1n3348);
not(notn3348,n1341);
and (s0n3348,notn3348,n3349);
and (s1n3348,n1341,n3346);
and (n3350,n3351,n1354);
wire s0n3351,s1n3351,notn3351;
or (n3351,s0n3351,s1n3351);
not(notn3351,n1341);
and (s0n3351,notn3351,n3352);
and (s1n3351,n1341,n3349);
and (n3353,n3354,n1257);
wire s0n3354,s1n3354,notn3354;
or (n3354,s0n3354,s1n3354);
not(notn3354,n1341);
and (s0n3354,notn3354,n3355);
and (s1n3354,n1341,n3352);
not (n3357,n3358);
wire s0n3358,s1n3358,notn3358;
or (n3358,s0n3358,s1n3358);
not(notn3358,n1102);
and (s0n3358,notn3358,n3359);
and (s1n3358,n1102,n3387);
nand (n3359,n3360,n3361,n3362,n3375);
nand (n3360,n1304,n1246);
nand (n3361,n1320,n1265);
nand (n3362,n3363,n1331);
nand (n3363,n3364,n3369,n3371,n3373);
nor (n3364,n3365,n3367);
and (n3365,n1270,n3366);
and (n3367,n1255,n3368);
nand (n3369,n1220,n3370);
nand (n3371,n1282,n3372);
nand (n3373,n1294,n3374);
nand (n3375,n3376,n1316);
nand (n3376,n3377,n3381,n3383,n3385);
nor (n3377,n3378,n3379);
and (n3378,n1270,n3368);
and (n3379,n1255,n3380);
nand (n3381,n1220,n3382);
nand (n3383,n1282,n3384);
nand (n3385,n1294,n3386);
not (n3388,n3389);
and (n3389,n3323,n3358);
nand (n3390,n3391,n3321);
nand (n3391,n3392,n3393);
not (n3392,n3255);
not (n3393,n3289);
and (n3394,n3395,n3400);
or (n3395,n3396,n3398);
wire s0n3396,s1n3396,notn3396;
or (n3396,s0n3396,s1n3396);
not(notn3396,n1102);
and (s0n3396,notn3396,1'b0);
and (s1n3396,n1102,n3397);
wire s0n3398,s1n3398,notn3398;
or (n3398,s0n3398,s1n3398);
not(notn3398,n1102);
and (s0n3398,notn3398,1'b0);
and (s1n3398,n1102,n3399);
or (n3400,n3401,n3403);
wire s0n3401,s1n3401,notn3401;
or (n3401,s0n3401,s1n3401);
not(notn3401,n1102);
and (s0n3401,notn3401,1'b0);
and (s1n3401,n1102,n3402);
wire s0n3403,s1n3403,notn3403;
or (n3403,s0n3403,s1n3403);
not(notn3403,n1102);
and (s0n3403,notn3403,1'b0);
and (s1n3403,n1102,n3404);
not (n3405,n3406);
nand (n3406,n3407,n3831);
or (n3407,n3408,n3689);
not (n3408,n3409);
nand (n3409,n3410,n3619);
nand (n3410,n3411,n3479,n3546);
nand (n3411,n3412,n3447);
not (n3412,n3413);
wire s0n3413,s1n3413,notn3413;
or (n3413,s0n3413,s1n3413);
not(notn3413,n1102);
and (s0n3413,notn3413,n3414);
and (s1n3413,n1102,n3446);
or (n3414,1'b0,n3415,n3416,n3417,n3432);
and (n3415,n1984,n1331);
and (n3416,n2000,n1316);
and (n3417,n3418,n1265);
or (n3418,1'b0,n3419,n3423,n3426,n3429);
and (n3419,n3420,n1223);
wire s0n3420,s1n3420,notn3420;
or (n3420,s0n3420,s1n3420);
not(notn3420,n1341);
and (s0n3420,notn3420,n3421);
and (s1n3420,n1341,n3422);
and (n3423,n3424,n1234);
wire s0n3424,s1n3424,notn3424;
or (n3424,s0n3424,s1n3424);
not(notn3424,n1341);
and (s0n3424,notn3424,n3425);
and (s1n3424,n1341,n3421);
and (n3426,n3427,n1354);
wire s0n3427,s1n3427,notn3427;
or (n3427,s0n3427,s1n3427);
not(notn3427,n1341);
and (s0n3427,notn3427,n3428);
and (s1n3427,n1341,n3425);
and (n3429,n3430,n1257);
wire s0n3430,s1n3430,notn3430;
or (n3430,s0n3430,s1n3430);
not(notn3430,n1341);
and (s0n3430,notn3430,n3431);
and (s1n3430,n1341,n3428);
and (n3432,n3433,n1246);
or (n3433,1'b0,n3434,n3437,n3440,n3443);
and (n3434,n3435,n1223);
wire s0n3435,s1n3435,notn3435;
or (n3435,s0n3435,s1n3435);
not(notn3435,n1341);
and (s0n3435,notn3435,n3436);
and (s1n3435,n1341,n3431);
and (n3437,n3438,n1234);
wire s0n3438,s1n3438,notn3438;
or (n3438,s0n3438,s1n3438);
not(notn3438,n1341);
and (s0n3438,notn3438,n3439);
and (s1n3438,n1341,n3436);
and (n3440,n3441,n1354);
wire s0n3441,s1n3441,notn3441;
or (n3441,s0n3441,s1n3441);
not(notn3441,n1341);
and (s0n3441,notn3441,n3442);
and (s1n3441,n1341,n3439);
and (n3443,n3444,n1257);
wire s0n3444,s1n3444,notn3444;
or (n3444,s0n3444,s1n3444);
not(notn3444,n1341);
and (s0n3444,notn3444,n3445);
and (s1n3444,n1341,n3442);
not (n3447,n3448);
or (n3448,n3449,n3451);
and (n3449,n1102,n3450);
nand (n3451,n3452,n3453,n3466,n3467);
nand (n3452,n1898,n1265);
nand (n3453,n3454,n1316);
nand (n3454,n3455,n3460,n3462,n3464);
nor (n3455,n3456,n3458);
and (n3456,n1270,n3457);
and (n3458,n1255,n3459);
nand (n3460,n1220,n3461);
nand (n3462,n1282,n3463);
nand (n3464,n1294,n3465);
nand (n3466,n1911,n1246);
nand (n3467,n3468,n1331);
nand (n3468,n3469,n3473,n3475,n3477);
nor (n3469,n3470,n3472);
and (n3470,n1270,n3471);
and (n3472,n1255,n3457);
nand (n3473,n1220,n3474);
nand (n3475,n1282,n3476);
nand (n3477,n1294,n3478);
or (n3479,n3480,n3514);
wire s0n3480,s1n3480,notn3480;
or (n3480,s0n3480,s1n3480);
not(notn3480,n1102);
and (s0n3480,notn3480,n3481);
and (s1n3480,n1102,n3513);
or (n3481,1'b0,n3482,n3483,n3484,n3499);
and (n3482,n2108,n1331);
and (n3483,n2123,n1316);
and (n3484,n3485,n1265);
or (n3485,1'b0,n3486,n3490,n3493,n3496);
and (n3486,n3487,n1223);
wire s0n3487,s1n3487,notn3487;
or (n3487,s0n3487,s1n3487);
not(notn3487,n1341);
and (s0n3487,notn3487,n3488);
and (s1n3487,n1341,n3489);
and (n3490,n3491,n1234);
wire s0n3491,s1n3491,notn3491;
or (n3491,s0n3491,s1n3491);
not(notn3491,n1341);
and (s0n3491,notn3491,n3492);
and (s1n3491,n1341,n3488);
and (n3493,n3494,n1354);
wire s0n3494,s1n3494,notn3494;
or (n3494,s0n3494,s1n3494);
not(notn3494,n1341);
and (s0n3494,notn3494,n3495);
and (s1n3494,n1341,n3492);
and (n3496,n3497,n1257);
wire s0n3497,s1n3497,notn3497;
or (n3497,s0n3497,s1n3497);
not(notn3497,n1341);
and (s0n3497,notn3497,n3498);
and (s1n3497,n1341,n3495);
and (n3499,n3500,n1246);
or (n3500,1'b0,n3501,n3504,n3507,n3510);
and (n3501,n3502,n1223);
wire s0n3502,s1n3502,notn3502;
or (n3502,s0n3502,s1n3502);
not(notn3502,n1341);
and (s0n3502,notn3502,n3503);
and (s1n3502,n1341,n3498);
and (n3504,n3505,n1234);
wire s0n3505,s1n3505,notn3505;
or (n3505,s0n3505,s1n3505);
not(notn3505,n1341);
and (s0n3505,notn3505,n3506);
and (s1n3505,n1341,n3503);
and (n3507,n3508,n1354);
wire s0n3508,s1n3508,notn3508;
or (n3508,s0n3508,s1n3508);
not(notn3508,n1341);
and (s0n3508,notn3508,n3509);
and (s1n3508,n1341,n3506);
and (n3510,n3511,n1257);
wire s0n3511,s1n3511,notn3511;
or (n3511,s0n3511,s1n3511);
not(notn3511,n1341);
and (s0n3511,notn3511,n3512);
and (s1n3511,n1341,n3509);
not (n3514,n3515);
nor (n3515,n3516,n3544);
nand (n3516,n3517,n3530,n3531,n3532);
nand (n3517,n3518,n1331);
nand (n3518,n3519,n3521,n3523,n3528);
nand (n3519,n1282,n3520);
nand (n3521,n1294,n3522);
nor (n3523,n3524,n3526);
and (n3524,n1270,n3525);
and (n3526,n1255,n3527);
nand (n3528,n1220,n3529);
nand (n3530,n2034,n1246);
nand (n3531,n2021,n1265);
nand (n3532,n3533,n1316);
nand (n3533,n3534,n3536,n3538,n3542);
nand (n3534,n1282,n3535);
nand (n3536,n1294,n3537);
nor (n3538,n3539,n3540);
and (n3539,n1270,n3527);
and (n3540,n1255,n3541);
nand (n3542,n1220,n3543);
and (n3544,n1102,n3545);
nand (n3546,n3547,n3617);
not (n3547,n3548);
and (n3548,n3549,n3583);
wire s0n3549,s1n3549,notn3549;
or (n3549,s0n3549,s1n3549);
not(notn3549,n1102);
and (s0n3549,notn3549,n3550);
and (s1n3549,n1102,n3582);
or (n3550,1'b0,n3551,n3552,n3553,n3568);
and (n3551,n2227,n1331);
and (n3552,n2243,n1316);
and (n3553,n3554,n1265);
or (n3554,1'b0,n3555,n3559,n3562,n3565);
and (n3555,n3556,n1223);
wire s0n3556,s1n3556,notn3556;
or (n3556,s0n3556,s1n3556);
not(notn3556,n1341);
and (s0n3556,notn3556,n3557);
and (s1n3556,n1341,n3558);
and (n3559,n3560,n1234);
wire s0n3560,s1n3560,notn3560;
or (n3560,s0n3560,s1n3560);
not(notn3560,n1341);
and (s0n3560,notn3560,n3561);
and (s1n3560,n1341,n3557);
and (n3562,n3563,n1354);
wire s0n3563,s1n3563,notn3563;
or (n3563,s0n3563,s1n3563);
not(notn3563,n1341);
and (s0n3563,notn3563,n3564);
and (s1n3563,n1341,n3561);
and (n3565,n3566,n1257);
wire s0n3566,s1n3566,notn3566;
or (n3566,s0n3566,s1n3566);
not(notn3566,n1341);
and (s0n3566,notn3566,n3567);
and (s1n3566,n1341,n3564);
and (n3568,n3569,n1246);
or (n3569,1'b0,n3570,n3573,n3576,n3579);
and (n3570,n3571,n1223);
wire s0n3571,s1n3571,notn3571;
or (n3571,s0n3571,s1n3571);
not(notn3571,n1341);
and (s0n3571,notn3571,n3572);
and (s1n3571,n1341,n3567);
and (n3573,n3574,n1234);
wire s0n3574,s1n3574,notn3574;
or (n3574,s0n3574,s1n3574);
not(notn3574,n1341);
and (s0n3574,notn3574,n3575);
and (s1n3574,n1341,n3572);
and (n3576,n3577,n1354);
wire s0n3577,s1n3577,notn3577;
or (n3577,s0n3577,s1n3577);
not(notn3577,n1341);
and (s0n3577,notn3577,n3578);
and (s1n3577,n1341,n3575);
and (n3579,n3580,n1257);
wire s0n3580,s1n3580,notn3580;
or (n3580,s0n3580,s1n3580);
not(notn3580,n1341);
and (s0n3580,notn3580,n3581);
and (s1n3580,n1341,n3578);
wire s0n3583,s1n3583,notn3583;
or (n3583,s0n3583,s1n3583);
not(notn3583,n1102);
and (s0n3583,notn3583,n3584);
and (s1n3583,n1102,n3616);
nand (n3584,n3585,n3602,n3603,n3604);
nand (n3585,n3586,n1331);
nand (n3586,n3587,n3592);
nor (n3587,n3588,n3590);
and (n3588,n1282,n3589);
and (n3590,n1294,n3591);
nor (n3592,n3593,n3599);
nand (n3593,n3594,n3597);
or (n3594,n3595,n1396);
not (n3595,n3596);
nand (n3597,n1255,n3598);
nor (n3599,n3600,n1402);
not (n3600,n3601);
nand (n3602,n2141,n1265);
nand (n3603,n2154,n1246);
nand (n3604,n3605,n1316);
nand (n3605,n3606,n3610,n3612,n3614);
nor (n3606,n3607,n3609);
and (n3607,n1255,n3608);
and (n3609,n1270,n3598);
nand (n3610,n1220,n3611);
nand (n3612,n1282,n3613);
nand (n3614,n1294,n3615);
not (n3617,n3618);
and (n3618,n3480,n3514);
and (n3619,n3620,n3687);
not (n3620,n3621);
and (n3621,n3622,n3656);
wire s0n3622,s1n3622,notn3622;
or (n3622,s0n3622,s1n3622);
not(notn3622,n1102);
and (s0n3622,notn3622,n3623);
and (s1n3622,n1102,n3655);
or (n3623,1'b0,n3624,n3625,n3626,n3641);
and (n3624,n1860,n1331);
and (n3625,n1876,n1316);
and (n3626,n3627,n1265);
or (n3627,1'b0,n3628,n3632,n3635,n3638);
and (n3628,n3629,n1223);
wire s0n3629,s1n3629,notn3629;
or (n3629,s0n3629,s1n3629);
not(notn3629,n1341);
and (s0n3629,notn3629,n3630);
and (s1n3629,n1341,n3631);
and (n3632,n3633,n1234);
wire s0n3633,s1n3633,notn3633;
or (n3633,s0n3633,s1n3633);
not(notn3633,n1341);
and (s0n3633,notn3633,n3634);
and (s1n3633,n1341,n3630);
and (n3635,n3636,n1354);
wire s0n3636,s1n3636,notn3636;
or (n3636,s0n3636,s1n3636);
not(notn3636,n1341);
and (s0n3636,notn3636,n3637);
and (s1n3636,n1341,n3634);
and (n3638,n3639,n1257);
wire s0n3639,s1n3639,notn3639;
or (n3639,s0n3639,s1n3639);
not(notn3639,n1341);
and (s0n3639,notn3639,n3640);
and (s1n3639,n1341,n3637);
and (n3641,n3642,n1246);
or (n3642,1'b0,n3643,n3646,n3649,n3652);
and (n3643,n3644,n1223);
wire s0n3644,s1n3644,notn3644;
or (n3644,s0n3644,s1n3644);
not(notn3644,n1341);
and (s0n3644,notn3644,n3645);
and (s1n3644,n1341,n3640);
and (n3646,n3647,n1234);
wire s0n3647,s1n3647,notn3647;
or (n3647,s0n3647,s1n3647);
not(notn3647,n1341);
and (s0n3647,notn3647,n3648);
and (s1n3647,n1341,n3645);
and (n3649,n3650,n1354);
wire s0n3650,s1n3650,notn3650;
or (n3650,s0n3650,s1n3650);
not(notn3650,n1341);
and (s0n3650,notn3650,n3651);
and (s1n3650,n1341,n3648);
and (n3652,n3653,n1257);
wire s0n3653,s1n3653,notn3653;
or (n3653,s0n3653,s1n3653);
not(notn3653,n1341);
and (s0n3653,notn3653,n3654);
and (s1n3653,n1341,n3651);
or (n3656,n3657,n3659);
and (n3657,n1102,n3658);
nand (n3659,n3660,n3673,n3674,n3675);
nand (n3660,n3661,n1331);
nand (n3661,n3662,n3667,n3669,n3671);
nor (n3662,n3663,n3665);
and (n3663,n1270,n3664);
and (n3665,n1255,n3666);
nand (n3667,n1220,n3668);
nand (n3669,n1282,n3670);
nand (n3671,n1294,n3672);
nand (n3673,n1774,n1265);
nand (n3674,n1787,n1246);
nand (n3675,n3676,n1316);
nand (n3676,n3677,n3681,n3683,n3685);
nor (n3677,n3678,n3679);
and (n3678,n1270,n3666);
and (n3679,n1255,n3680);
nand (n3681,n1220,n3682);
nand (n3683,n1282,n3684);
nand (n3685,n1294,n3686);
not (n3687,n3688);
and (n3688,n3413,n3448);
not (n3689,n3690);
nor (n3690,n3691,n3692);
nor (n3691,n3622,n3656);
nand (n3692,n3693,n3760);
nand (n3693,n3694,n3729);
not (n3694,n3695);
wire s0n3695,s1n3695,notn3695;
or (n3695,s0n3695,s1n3695);
not(notn3695,n1102);
and (s0n3695,notn3695,n3696);
and (s1n3695,n1102,n3728);
or (n3696,1'b0,n3697,n3698,n3699,n3714);
and (n3697,n1621,n1331);
and (n3698,n1637,n1316);
and (n3699,n3700,n1265);
or (n3700,1'b0,n3701,n3705,n3708,n3711);
and (n3701,n3702,n1223);
wire s0n3702,s1n3702,notn3702;
or (n3702,s0n3702,s1n3702);
not(notn3702,n1341);
and (s0n3702,notn3702,n3703);
and (s1n3702,n1341,n3704);
and (n3705,n3706,n1234);
wire s0n3706,s1n3706,notn3706;
or (n3706,s0n3706,s1n3706);
not(notn3706,n1341);
and (s0n3706,notn3706,n3707);
and (s1n3706,n1341,n3703);
and (n3708,n3709,n1354);
wire s0n3709,s1n3709,notn3709;
or (n3709,s0n3709,s1n3709);
not(notn3709,n1341);
and (s0n3709,notn3709,n3710);
and (s1n3709,n1341,n3707);
and (n3711,n3712,n1257);
wire s0n3712,s1n3712,notn3712;
or (n3712,s0n3712,s1n3712);
not(notn3712,n1341);
and (s0n3712,notn3712,n3713);
and (s1n3712,n1341,n3710);
and (n3714,n3715,n1246);
or (n3715,1'b0,n3716,n3719,n3722,n3725);
and (n3716,n3717,n1223);
wire s0n3717,s1n3717,notn3717;
or (n3717,s0n3717,s1n3717);
not(notn3717,n1341);
and (s0n3717,notn3717,n3718);
and (s1n3717,n1341,n3713);
and (n3719,n3720,n1234);
wire s0n3720,s1n3720,notn3720;
or (n3720,s0n3720,s1n3720);
not(notn3720,n1341);
and (s0n3720,notn3720,n3721);
and (s1n3720,n1341,n3718);
and (n3722,n3723,n1354);
wire s0n3723,s1n3723,notn3723;
or (n3723,s0n3723,s1n3723);
not(notn3723,n1341);
and (s0n3723,notn3723,n3724);
and (s1n3723,n1341,n3721);
and (n3725,n3726,n1257);
wire s0n3726,s1n3726,notn3726;
or (n3726,s0n3726,s1n3726);
not(notn3726,n1341);
and (s0n3726,notn3726,n3727);
and (s1n3726,n1341,n3724);
not (n3729,n3730);
wire s0n3730,s1n3730,notn3730;
or (n3730,s0n3730,s1n3730);
not(notn3730,n1102);
and (s0n3730,notn3730,n3731);
and (s1n3730,n1102,n3759);
nand (n3731,n3732,n3745,n3746,n3747);
nand (n3732,n3733,n1331);
nand (n3733,n3734,n3739,n3741,n3743);
nor (n3734,n3735,n3737);
and (n3735,n1270,n3736);
and (n3737,n1255,n3738);
nand (n3739,n1220,n3740);
nand (n3741,n1282,n3742);
nand (n3743,n1294,n3744);
nand (n3745,n1535,n1265);
nand (n3746,n1548,n1246);
nand (n3747,n3748,n1316);
nand (n3748,n3749,n3753,n3755,n3757);
nor (n3749,n3750,n3751);
and (n3750,n1270,n3738);
and (n3751,n1255,n3752);
nand (n3753,n1220,n3754);
nand (n3755,n1282,n3756);
nand (n3757,n1294,n3758);
nand (n3760,n3761,n3796);
not (n3761,n3762);
wire s0n3762,s1n3762,notn3762;
or (n3762,s0n3762,s1n3762);
not(notn3762,n1102);
and (s0n3762,notn3762,n3763);
and (s1n3762,n1102,n3795);
or (n3763,1'b0,n3764,n3765,n3766,n3781);
and (n3764,n1740,n1331);
and (n3765,n1753,n1316);
and (n3766,n3767,n1265);
or (n3767,1'b0,n3768,n3772,n3775,n3778);
and (n3768,n3769,n1223);
wire s0n3769,s1n3769,notn3769;
or (n3769,s0n3769,s1n3769);
not(notn3769,n1341);
and (s0n3769,notn3769,n3770);
and (s1n3769,n1341,n3771);
and (n3772,n3773,n1234);
wire s0n3773,s1n3773,notn3773;
or (n3773,s0n3773,s1n3773);
not(notn3773,n1341);
and (s0n3773,notn3773,n3774);
and (s1n3773,n1341,n3770);
and (n3775,n3776,n1354);
wire s0n3776,s1n3776,notn3776;
or (n3776,s0n3776,s1n3776);
not(notn3776,n1341);
and (s0n3776,notn3776,n3777);
and (s1n3776,n1341,n3774);
and (n3778,n3779,n1257);
wire s0n3779,s1n3779,notn3779;
or (n3779,s0n3779,s1n3779);
not(notn3779,n1341);
and (s0n3779,notn3779,n3780);
and (s1n3779,n1341,n3777);
and (n3781,n3782,n1246);
or (n3782,1'b0,n3783,n3786,n3789,n3792);
and (n3783,n3784,n1223);
wire s0n3784,s1n3784,notn3784;
or (n3784,s0n3784,s1n3784);
not(notn3784,n1341);
and (s0n3784,notn3784,n3785);
and (s1n3784,n1341,n3780);
and (n3786,n3787,n1234);
wire s0n3787,s1n3787,notn3787;
or (n3787,s0n3787,s1n3787);
not(notn3787,n1341);
and (s0n3787,notn3787,n3788);
and (s1n3787,n1341,n3785);
and (n3789,n3790,n1354);
wire s0n3790,s1n3790,notn3790;
or (n3790,s0n3790,s1n3790);
not(notn3790,n1341);
and (s0n3790,notn3790,n3791);
and (s1n3790,n1341,n3788);
and (n3792,n3793,n1257);
wire s0n3793,s1n3793,notn3793;
or (n3793,s0n3793,s1n3793);
not(notn3793,n1341);
and (s0n3793,notn3793,n3794);
and (s1n3793,n1341,n3791);
not (n3796,n3797);
nand (n3797,n3798,n3802);
or (n3798,n3799,n3801);
not (n3799,n3800);
not (n3801,n1102);
not (n3802,n3803);
nand (n3803,n3804,n3805,n3818,n3819);
nand (n3804,n1678,n1246);
nand (n3805,n3806,n1331);
nand (n3806,n3807,n3812,n3814,n3816);
nor (n3807,n3808,n3810);
and (n3808,n1270,n3809);
and (n3810,n1255,n3811);
nand (n3812,n1220,n3813);
nand (n3814,n1282,n3815);
nand (n3816,n1294,n3817);
nand (n3818,n1691,n1265);
nand (n3819,n3820,n1316);
nand (n3820,n3821,n3825,n3827,n3829);
nor (n3821,n3822,n3823);
and (n3822,n1270,n3811);
and (n3823,n1255,n3824);
nand (n3825,n1220,n3826);
nand (n3827,n1282,n3828);
nand (n3829,n1294,n3830);
nor (n3831,n3251,n3832);
nand (n3832,n3833,n3837);
or (n3833,n3834,n3836);
not (n3834,n3835);
and (n3835,n3762,n3797);
not (n3836,n3693);
not (n3837,n3838);
and (n3838,n3695,n3730);
not (n3839,n3840);
nand (n3840,n3841,n3845);
or (n3841,n3842,n3843);
not (n3842,n3400);
not (n3843,n3844);
and (n3844,n3398,n3396);
not (n3845,n3846);
and (n3846,n3403,n3401);
and (n3847,n3239,n3245);
or (n3848,n3849,n3868,n3958);
and (n3849,n3850,n3852);
xor (n3850,n3851,n2382);
xor (n3851,n2278,n2329);
not (n3852,n3853);
nor (n3853,n3854,n3865);
and (n3854,n3855,n3856);
xor (n3855,n3403,n3401);
nand (n3856,n3857,n3862,n3864);
nand (n3857,n3409,n3858,n3860,n3861);
and (n3858,n3859,n3395);
not (n3859,n3691);
not (n3860,n3390);
not (n3861,n3692);
nor (n3862,n3863,n3844);
and (n3863,n3251,n3395);
nand (n3864,n3832,n3860,n3395);
and (n3865,n3866,n3867);
not (n3866,n3855);
not (n3867,n3856);
and (n3868,n3852,n3869);
or (n3869,n3870,n3883,n3957);
and (n3870,n3871,n3873);
xor (n3871,n3872,n2502);
xor (n3872,n2384,n2436);
not (n3873,n3874);
nand (n3874,n3875,n3882);
or (n3875,n3876,n3877);
xor (n3876,n3398,n3396);
not (n3877,n3878);
nand (n3878,n3879,n3881);
nor (n3879,n3880,n3251);
and (n3880,n3832,n3860);
nand (n3881,n3409,n3690,n3860);
nand (n3882,n3877,n3876);
and (n3883,n3873,n3884);
or (n3884,n3885,n3908,n3956);
and (n3885,n3886,n3888);
xor (n3886,n3887,n2610);
xor (n3887,n2504,n2557);
not (n3888,n3889);
xor (n3889,n3890,n3891);
xor (n3890,n3323,n3358);
nand (n3891,n3892,n3906);
or (n3892,n3893,n3896);
not (n3893,n3894);
nor (n3894,n3895,n3692);
not (n3895,n3391);
not (n3896,n3897);
or (n3897,n3621,n3898,n3905);
and (n3898,n3656,n3899);
or (n3899,n3688,n3900,n3904);
and (n3900,n3448,n3901);
or (n3901,n3618,n3902,n3903);
and (n3902,n3514,n3548);
and (n3903,n3480,n3548);
and (n3904,n3413,n3901);
and (n3905,n3622,n3899);
nor (n3906,n3907,n3254);
and (n3907,n3832,n3391);
and (n3908,n3888,n3909);
or (n3909,n3910,n3922,n3955);
and (n3910,n3911,n3913);
xor (n3911,n3912,n2738);
xor (n3912,n2612,n2677);
not (n3913,n3914);
xor (n3914,n3915,n3916);
xor (n3915,n3255,n3289);
or (n3916,n3838,n3917,n3921);
and (n3917,n3730,n3918);
or (n3918,n3835,n3919,n3920);
and (n3919,n3797,n3897);
and (n3920,n3762,n3897);
and (n3921,n3695,n3918);
and (n3922,n3913,n3923);
or (n3923,n3924,n3930,n3954);
and (n3924,n3925,n3927);
xor (n3925,n3926,n2863);
xor (n3926,n2740,n2805);
not (n3927,n3928);
xor (n3928,n3929,n3918);
xor (n3929,n3695,n3730);
and (n3930,n3927,n3931);
or (n3931,n3932,n3938,n3953);
and (n3932,n3933,n3935);
xor (n3933,n3934,n2980);
xor (n3934,n2865,n2922);
not (n3935,n3936);
xor (n3936,n3937,n3897);
xor (n3937,n3762,n3797);
and (n3938,n3935,n3939);
or (n3939,n3940,n3946,n3952);
and (n3940,n3941,n3943);
xor (n3941,n3942,n3104);
xor (n3942,n2982,n3042);
not (n3943,n3944);
xor (n3944,n3945,n3899);
xor (n3945,n3622,n3656);
and (n3946,n3943,n3947);
and (n3947,n3948,n3949);
xor (n3948,n3105,n3165);
not (n3949,n3950);
xor (n3950,n3951,n3901);
xor (n3951,n3413,n3448);
and (n3952,n3941,n3947);
and (n3953,n3933,n3939);
and (n3954,n3925,n3931);
and (n3955,n3911,n3923);
and (n3956,n3886,n3909);
and (n3957,n3871,n3884);
and (n3958,n3850,n3869);
and (n3959,n3960,n3962);
xor (n3960,n3961,n3869);
xor (n3961,n3850,n3852);
and (n3962,n3963,n3965);
xor (n3963,n3964,n3884);
xor (n3964,n3871,n3873);
and (n3965,n3966,n3968);
xor (n3966,n3967,n3909);
xor (n3967,n3886,n3888);
and (n3968,n3969,n3971);
xor (n3969,n3970,n3923);
xor (n3970,n3911,n3913);
and (n3971,n3972,n3974);
xor (n3972,n3973,n3931);
xor (n3973,n3925,n3927);
and (n3974,n3975,n3977);
xor (n3975,n3976,n3939);
xor (n3976,n3933,n3935);
and (n3977,n3978,n3980);
xor (n3978,n3979,n3947);
xor (n3979,n3941,n3943);
and (n3980,n3981,n3982);
xor (n3981,n3948,n3949);
and (n3982,n3983,n3986);
not (n3983,n3984);
xor (n3984,n3985,n3548);
xor (n3985,n3480,n3514);
not (n3986,n3987);
xor (n3987,n3549,n3583);
or (n3988,n3989,n3993,n4052);
and (n3989,n3990,n3992);
xor (n3990,n3991,n1204);
xor (n3991,n1199,n1201);
xor (n3992,n3960,n3962);
and (n3993,n3992,n3994);
or (n3994,n3995,n3999,n4051);
and (n3995,n3996,n3998);
xor (n3996,n3997,n1211);
xor (n3997,n1206,n1208);
xor (n3998,n3963,n3965);
and (n3999,n3998,n4000);
or (n4000,n4001,n4005,n4050);
and (n4001,n4002,n4004);
xor (n4002,n4003,n1405);
xor (n4003,n1213,n1333);
xor (n4004,n3966,n3968);
and (n4005,n4004,n4006);
or (n4006,n4007,n4011,n4049);
and (n4007,n4008,n4010);
xor (n4008,n4009,n1530);
xor (n4009,n1407,n1460);
xor (n4010,n3969,n3971);
and (n4011,n4010,n4012);
or (n4012,n4013,n4017,n4048);
and (n4013,n4014,n4016);
xor (n4014,n4015,n1654);
xor (n4015,n1532,n1589);
xor (n4016,n3972,n3974);
and (n4017,n4016,n4018);
or (n4018,n4019,n4023,n4047);
and (n4019,n4020,n4022);
xor (n4020,n4021,n1769);
xor (n4021,n1656,n1708);
xor (n4022,n3975,n3977);
and (n4023,n4022,n4024);
or (n4024,n4025,n4029,n4046);
and (n4025,n4026,n4028);
xor (n4026,n4027,n1893);
xor (n4027,n1771,n1828);
xor (n4028,n3978,n3980);
and (n4029,n4028,n4030);
or (n4030,n4031,n4035,n4045);
and (n4031,n4032,n4034);
xor (n4032,n4033,n2016);
xor (n4033,n1895,n1952);
xor (n4034,n3981,n3982);
and (n4035,n4034,n4036);
or (n4036,n4037,n4041,n4044);
and (n4037,n4038,n4040);
xor (n4038,n4039,n2137);
xor (n4039,n2018,n2075);
xor (n4040,n3983,n3986);
and (n4041,n4040,n4042);
and (n4042,n4043,n3987);
xor (n4043,n2138,n2195);
and (n4044,n4038,n4042);
and (n4045,n4032,n4036);
and (n4046,n4026,n4030);
and (n4047,n4020,n4024);
and (n4048,n4014,n4018);
and (n4049,n4008,n4012);
and (n4050,n4002,n4006);
and (n4051,n3996,n4000);
and (n4052,n3990,n3994);
or (n4053,n4054,n4057,n4097);
and (n4054,n4055,n4004);
xor (n4055,n4056,n3994);
xor (n4056,n3990,n3992);
and (n4057,n4004,n4058);
or (n4058,n4059,n4062,n4096);
and (n4059,n4060,n4010);
xor (n4060,n4061,n4000);
xor (n4061,n3996,n3998);
and (n4062,n4010,n4063);
or (n4063,n4064,n4067,n4095);
and (n4064,n4065,n4016);
xor (n4065,n4066,n4006);
xor (n4066,n4002,n4004);
and (n4067,n4016,n4068);
or (n4068,n4069,n4072,n4094);
and (n4069,n4070,n4022);
xor (n4070,n4071,n4012);
xor (n4071,n4008,n4010);
and (n4072,n4022,n4073);
or (n4073,n4074,n4077,n4093);
and (n4074,n4075,n4028);
xor (n4075,n4076,n4018);
xor (n4076,n4014,n4016);
and (n4077,n4028,n4078);
or (n4078,n4079,n4082,n4092);
and (n4079,n4080,n4034);
xor (n4080,n4081,n4024);
xor (n4081,n4020,n4022);
and (n4082,n4034,n4083);
or (n4083,n4084,n4087,n4091);
and (n4084,n4085,n4040);
xor (n4085,n4086,n4030);
xor (n4086,n4026,n4028);
and (n4087,n4040,n4088);
and (n4088,n4089,n3987);
xor (n4089,n4090,n4036);
xor (n4090,n4032,n4034);
and (n4091,n4085,n4088);
and (n4092,n4080,n4083);
and (n4093,n4075,n4078);
and (n4094,n4070,n4073);
and (n4095,n4065,n4068);
and (n4096,n4060,n4063);
and (n4097,n4055,n4058);
and (n4098,n4099,n4101);
xor (n4099,n4100,n4058);
xor (n4100,n4055,n4004);
and (n4101,n4102,n4104);
xor (n4102,n4103,n4063);
xor (n4103,n4060,n4010);
and (n4104,n4105,n4107);
xor (n4105,n4106,n4068);
xor (n4106,n4065,n4016);
and (n4107,n4108,n4110);
xor (n4108,n4109,n4073);
xor (n4109,n4070,n4022);
and (n4110,n4111,n4113);
xor (n4111,n4112,n4078);
xor (n4112,n4075,n4028);
xor (n4113,n4114,n4083);
xor (n4114,n4080,n4034);
xor (n4115,n1094,n4099);
wire s0n4116,s1n4116,notn4116;
or (n4116,s0n4116,s1n4116);
not(notn4116,n1102);
and (s0n4116,notn4116,n4117);
and (s1n4116,n1102,n4771);
xor (n4117,n4118,n4758);
xor (n4118,n4119,n4609);
xor (n4119,n4120,n4241);
xor (n4120,n4121,n4234);
xor (n4121,n4122,n4190);
xor (n4122,n4123,n4149);
xor (n4123,n4124,n4129);
xor (n4124,n4125,n4127);
wire s0n4125,s1n4125,notn4125;
or (n4125,s0n4125,s1n4125);
not(notn4125,n1102);
and (s0n4125,notn4125,1'b0);
and (s1n4125,n1102,n4126);
wire s0n4127,s1n4127,notn4127;
or (n4127,s0n4127,s1n4127);
not(notn4127,n1102);
and (s0n4127,notn4127,1'b0);
and (s1n4127,n1102,n4128);
or (n4129,n4130,n4135,n4148);
and (n4130,n4131,n4133);
wire s0n4131,s1n4131,notn4131;
or (n4131,s0n4131,s1n4131);
not(notn4131,n1102);
and (s0n4131,notn4131,1'b0);
and (s1n4131,n1102,n4132);
wire s0n4133,s1n4133,notn4133;
or (n4133,s0n4133,s1n4133);
not(notn4133,n1102);
and (s0n4133,notn4133,1'b0);
and (s1n4133,n1102,n4134);
and (n4135,n4133,n4136);
or (n4136,n4137,n4142,n4147);
and (n4137,n4138,n4140);
wire s0n4138,s1n4138,notn4138;
or (n4138,s0n4138,s1n4138);
not(notn4138,n1102);
and (s0n4138,notn4138,1'b0);
and (s1n4138,n1102,n4139);
wire s0n4140,s1n4140,notn4140;
or (n4140,s0n4140,s1n4140);
not(notn4140,n1102);
and (s0n4140,notn4140,1'b0);
and (s1n4140,n1102,n4141);
and (n4142,n4140,n4143);
or (n4143,n4144,n4145,n4146);
and (n4144,n2272,n2274);
and (n4145,n2274,n2276);
and (n4146,n2272,n2276);
and (n4147,n4138,n4143);
and (n4148,n4131,n4136);
not (n4149,n4150);
nor (n4150,n4151,n4187);
and (n4151,n4152,n4182);
nand (n4152,n4153,n4171);
or (n4153,n4154,n3877);
not (n4154,n4155);
nor (n4155,n4156,n4162);
not (n4156,n4157);
or (n4157,n4158,n4160);
wire s0n4158,s1n4158,notn4158;
or (n4158,s0n4158,s1n4158);
not(notn4158,n1102);
and (s0n4158,notn4158,1'b0);
and (s1n4158,n1102,n4159);
wire s0n4160,s1n4160,notn4160;
or (n4160,s0n4160,s1n4160);
not(notn4160,n1102);
and (s0n4160,notn4160,1'b0);
and (s1n4160,n1102,n4161);
not (n4162,n4163);
and (n4163,n3394,n4164);
nor (n4164,n4165,n4170);
nor (n4165,n4166,n4168);
wire s0n4166,s1n4166,notn4166;
or (n4166,s0n4166,s1n4166);
not(notn4166,n1102);
and (s0n4166,notn4166,1'b0);
and (s1n4166,n1102,n4167);
wire s0n4168,s1n4168,notn4168;
or (n4168,s0n4168,s1n4168);
not(notn4168,n1102);
and (s0n4168,notn4168,1'b0);
and (s1n4168,n1102,n4169);
nor (n4170,n3242,n3240);
nor (n4171,n4172,n4181);
and (n4172,n4173,n4157);
nand (n4173,n4174,n4176);
or (n4174,n4175,n3839);
not (n4175,n4164);
nor (n4176,n4177,n4180);
and (n4177,n4178,n4179);
not (n4178,n4165);
and (n4179,n3240,n3242);
and (n4180,n4168,n4166);
and (n4181,n4160,n4158);
xor (n4182,n4183,n4185);
wire s0n4183,s1n4183,notn4183;
or (n4183,s0n4183,s1n4183);
not(notn4183,n1102);
and (s0n4183,notn4183,1'b0);
and (s1n4183,n1102,n4184);
wire s0n4185,s1n4185,notn4185;
or (n4185,s0n4185,s1n4185);
not(notn4185,n1102);
and (s0n4185,notn4185,1'b0);
and (s1n4185,n1102,n4186);
and (n4187,n4188,n4189);
not (n4188,n4152);
not (n4189,n4182);
or (n4190,n4191,n4206,n4233);
and (n4191,n4192,n4194);
xor (n4192,n4193,n4136);
xor (n4193,n4131,n4133);
not (n4194,n4195);
nor (n4195,n4196,n4205);
and (n4196,n4197,n4199);
not (n4197,n4198);
xor (n4198,n4160,n4158);
not (n4199,n4200);
nand (n4200,n4201,n4204);
or (n4201,n4202,n3405);
not (n4202,n4203);
and (n4203,n3249,n4163);
not (n4204,n4173);
and (n4205,n4198,n4200);
and (n4206,n4194,n4207);
or (n4207,n4208,n4227,n4232);
and (n4208,n4209,n4211);
xor (n4209,n4210,n4143);
xor (n4210,n4138,n4140);
not (n4211,n4212);
nor (n4212,n4213,n4224);
and (n4213,n4214,n4215);
xor (n4214,n4168,n4166);
nand (n4215,n4216,n4221);
or (n4216,n4217,n3405);
not (n4217,n4218);
and (n4218,n3249,n4219);
nor (n4219,n4220,n4170);
not (n4220,n3394);
nor (n4221,n4222,n4179);
and (n4222,n3840,n4223);
not (n4223,n4170);
and (n4224,n4225,n4226);
not (n4225,n4214);
not (n4226,n4215);
and (n4227,n4211,n4228);
or (n4228,n4229,n4230,n4231);
and (n4229,n2270,n3235);
and (n4230,n3235,n3848);
and (n4231,n2270,n3848);
and (n4232,n4209,n4228);
and (n4233,n4192,n4207);
and (n4234,n4235,n4237);
xor (n4235,n4236,n4207);
xor (n4236,n4192,n4194);
and (n4237,n4238,n4240);
xor (n4238,n4239,n4228);
xor (n4239,n4209,n4211);
and (n4240,n2268,n3959);
nand (n4241,n4242,n4608);
or (n4242,n4243,n4342);
not (n4243,n4244);
nor (n4244,n4245,n4338);
not (n4245,n4246);
nand (n4246,n4247,n4315);
xor (n4247,n4248,n4302);
xor (n4248,n4249,n4281);
xor (n4249,n4250,n4255);
xor (n4250,n4251,n4253);
wire s0n4251,s1n4251,notn4251;
or (n4251,s0n4251,s1n4251);
not(notn4251,n1102);
and (s0n4251,notn4251,1'b0);
and (s1n4251,n1102,n4252);
wire s0n4253,s1n4253,notn4253;
or (n4253,s0n4253,s1n4253);
not(notn4253,n1102);
and (s0n4253,notn4253,1'b0);
and (s1n4253,n1102,n4254);
not (n4255,n4256);
nor (n4256,n4257,n4269);
and (n4257,n3878,n4258);
nor (n4258,n4162,n4259);
nand (n4259,n4260,n4263);
not (n4260,n4261);
nand (n4261,n4262,n4157);
or (n4262,n4185,n4183);
not (n4263,n4264);
and (n4264,n4265,n4267);
wire s0n4265,s1n4265,notn4265;
or (n4265,s0n4265,s1n4265);
not(notn4265,n1102);
and (s0n4265,notn4265,1'b0);
and (s1n4265,n1102,n4266);
wire s0n4267,s1n4267,notn4267;
or (n4267,s0n4267,s1n4267);
not(notn4267,n1102);
and (s0n4267,notn4267,1'b0);
and (s1n4267,n1102,n4268);
nand (n4269,n4270,n4271);
or (n4270,n4204,n4259);
nor (n4271,n4272,n4279);
and (n4272,n4273,n4263);
nand (n4273,n4274,n4277);
or (n4274,n4275,n4276);
not (n4275,n4181);
not (n4276,n4262);
not (n4277,n4278);
and (n4278,n4183,n4185);
not (n4279,n4280);
or (n4280,n4267,n4265);
not (n4281,n4282);
or (n4282,n4283,n4301);
and (n4283,n4284,n4289);
xor (n4284,n4285,n4287);
wire s0n4285,s1n4285,notn4285;
or (n4285,s0n4285,s1n4285);
not(notn4285,n1102);
and (s0n4285,notn4285,1'b0);
and (s1n4285,n1102,n4286);
wire s0n4287,s1n4287,notn4287;
or (n4287,s0n4287,s1n4287);
not(notn4287,n1102);
and (s0n4287,notn4287,1'b0);
and (s1n4287,n1102,n4288);
not (n4289,n4290);
nand (n4290,n4291,n4300);
or (n4291,n4292,n4294);
not (n4292,n4293);
xor (n4293,n4265,n4267);
nand (n4294,n4295,n4298);
or (n4295,n4296,n3877);
not (n4296,n4297);
nor (n4297,n4162,n4261);
nor (n4298,n4299,n4273);
and (n4299,n4173,n4260);
nand (n4300,n4294,n4292);
and (n4301,n4285,n4287);
nand (n4302,n4303,n4314);
nand (n4303,n4304,n4311);
or (n4304,n4305,n4308);
not (n4305,n4306);
wire s0n4306,s1n4306,notn4306;
or (n4306,s0n4306,s1n4306);
not(notn4306,n1102);
and (s0n4306,notn4306,1'b0);
and (s1n4306,n1102,n4307);
or (n4308,n4309,n4310);
and (n4309,n4124,n4149);
and (n4310,n4125,n4127);
not (n4311,n4312);
wire s0n4312,s1n4312,notn4312;
or (n4312,s0n4312,s1n4312);
not(notn4312,n1102);
and (s0n4312,notn4312,1'b0);
and (s1n4312,n1102,n4313);
nand (n4314,n4305,n4308);
or (n4315,n4316,n4337);
and (n4316,n4317,n4325);
xor (n4317,n4318,n4319);
xor (n4318,n4284,n4289);
nor (n4319,n4320,n4324);
and (n4320,n4321,n4323);
not (n4321,n4322);
xor (n4322,n4306,n4312);
not (n4323,n4308);
and (n4324,n4322,n4308);
nand (n4325,n4326,n4333);
or (n4326,n4327,n4330);
not (n4327,n4328);
wire s0n4328,s1n4328,notn4328;
or (n4328,s0n4328,s1n4328);
not(notn4328,n1102);
and (s0n4328,notn4328,1'b0);
and (s1n4328,n1102,n4329);
not (n4330,n4331);
or (n4331,n4332,n4130);
and (n4332,n4193,n4194);
nand (n4333,n4334,n4335);
or (n4334,n4328,n4331);
wire s0n4335,s1n4335,notn4335;
or (n4335,s0n4335,s1n4335);
not(notn4335,n1102);
and (s0n4335,notn4335,1'b0);
and (s1n4335,n1102,n4336);
and (n4337,n4318,n4319);
not (n4338,n4339);
nand (n4339,n4340,n4341);
not (n4340,n4247);
not (n4341,n4315);
nand (n4342,n4343,n4584,n4598);
nand (n4343,n4344,n4415,n4533);
and (n4344,n4345,n4408);
and (n4345,n4346,n4390);
nand (n4346,n4347,n4374);
not (n4347,n4348);
xor (n4348,n4349,n4363);
xor (n4349,n4350,n4351);
xor (n4350,n4193,n4194);
nand (n4351,n4352,n4359);
or (n4352,n4353,n4356);
not (n4353,n4354);
wire s0n4354,s1n4354,notn4354;
or (n4354,s0n4354,s1n4354);
not(notn4354,n1102);
and (s0n4354,notn4354,1'b0);
and (s1n4354,n1102,n4355);
not (n4356,n4357);
or (n4357,n4358,n4144);
and (n4358,n2271,n3235);
nand (n4359,n4360,n4361);
or (n4360,n4354,n4357);
wire s0n4361,s1n4361,notn4361;
or (n4361,s0n4361,s1n4361);
not(notn4361,n1102);
and (s0n4361,notn4361,1'b0);
and (s1n4361,n1102,n4362);
nand (n4363,n4364,n4373);
or (n4364,n4365,n4371);
not (n4365,n4366);
xor (n4366,n4367,n4369);
wire s0n4367,s1n4367,notn4367;
or (n4367,s0n4367,s1n4367);
not(notn4367,n1102);
and (s0n4367,notn4367,1'b0);
and (s1n4367,n1102,n4368);
wire s0n4369,s1n4369,notn4369;
or (n4369,s0n4369,s1n4369);
not(notn4369,n1102);
and (s0n4369,notn4369,1'b0);
and (s1n4369,n1102,n4370);
or (n4371,n4372,n4137);
and (n4372,n4210,n4211);
nand (n4373,n4365,n4371);
not (n4374,n4375);
or (n4375,n4376,n4389);
and (n4376,n4377,n4384);
xor (n4377,n4378,n4379);
xor (n4378,n4210,n4211);
or (n4379,n4380,n4383);
and (n4380,n1099,n4381);
or (n4381,n4382,n2277);
and (n4382,n3851,n3852);
and (n4383,n1100,n1195);
nand (n4384,n4385,n4388);
or (n4385,n4386,n4357);
not (n4386,n4387);
xor (n4387,n4354,n4361);
nand (n4388,n4386,n4357);
and (n4389,n4378,n4379);
nand (n4390,n4391,n4404);
not (n4391,n4392);
xor (n4392,n4393,n4400);
xor (n4393,n4394,n4395);
xor (n4394,n4124,n4149);
nand (n4395,n4396,n4399);
or (n4396,n4397,n4331);
not (n4397,n4398);
xor (n4398,n4328,n4335);
nand (n4399,n4397,n4331);
nand (n4400,n4401,n4403);
nand (n4401,n4402,n4369);
or (n4402,n4367,n4371);
nand (n4403,n4371,n4367);
not (n4404,n4405);
or (n4405,n4406,n4407);
and (n4406,n4349,n4363);
and (n4407,n4350,n4351);
nand (n4408,n4409,n4411);
not (n4409,n4410);
xor (n4410,n4317,n4325);
not (n4411,n4412);
or (n4412,n4413,n4414);
and (n4413,n4393,n4400);
and (n4414,n4394,n4395);
nand (n4415,n4416,n4526);
or (n4416,n4417,n4461);
not (n4417,n4418);
and (n4418,n4419,n4447);
nand (n4419,n4420,n4433);
not (n4420,n4421);
xor (n4421,n4422,n4430);
xor (n4422,n4423,n4424);
xor (n4423,n3912,n3913);
nand (n4424,n4425,n4429);
nand (n4425,n4426,n1589);
or (n4426,n1532,n4427);
or (n4427,n4428,n2864);
and (n4428,n3934,n3935);
nand (n4429,n4427,n1532);
xor (n4430,n4009,n4431);
or (n4431,n4432,n2739);
and (n4432,n3926,n3927);
not (n4433,n4434);
or (n4434,n4435,n4446);
and (n4435,n4436,n4442);
xor (n4436,n4437,n4438);
xor (n4437,n3926,n3927);
or (n4438,n4439,n1655);
and (n4439,n4021,n4440);
or (n4440,n4441,n2981);
and (n4441,n3942,n3943);
nand (n4442,n4443,n4445);
or (n4443,n4444,n4427);
not (n4444,n4015);
nand (n4445,n4444,n4427);
and (n4446,n4437,n4438);
nand (n4447,n4448,n4457);
not (n4448,n4449);
xor (n4449,n4450,n4454);
xor (n4450,n4451,n4452);
xor (n4451,n3887,n3888);
or (n4452,n4453,n1406);
and (n4453,n4009,n4431);
xor (n4454,n4003,n4455);
or (n4455,n4456,n2611);
and (n4456,n3912,n3913);
not (n4457,n4458);
or (n4458,n4459,n4460);
and (n4459,n4422,n4430);
and (n4460,n4423,n4424);
not (n4461,n4462);
nand (n4462,n4463,n4520);
or (n4463,n4464,n4503);
not (n4464,n4465);
or (n4465,n4466,n4502);
and (n4466,n4467,n4483);
xor (n4467,n4468,n4477);
or (n4468,n4469,n4476);
and (n4469,n4470,n4472);
xor (n4470,n4471,n1895);
xor (n4471,n1952,n3105);
nand (n4472,n4473,n4475);
or (n4473,n4474,n3949);
not (n4474,n3165);
nand (n4475,n4474,n3949);
and (n4476,n4471,n1895);
xor (n4477,n4478,n4481);
xor (n4478,n4479,n4480);
and (n4479,n1952,n3105);
xor (n4480,n3942,n3943);
xor (n4481,n4027,n4482);
and (n4482,n3949,n3165);
or (n4483,n4484,n4501);
and (n4484,n4485,n4500);
xor (n4485,n4486,n4488);
or (n4486,n4487,n2017);
and (n4487,n4039,n3983);
nand (n4488,n4489,n4499);
or (n4489,n4490,n4492);
nor (n4490,n4491,n3986);
xor (n4491,n4039,n3983);
nor (n4492,n4493,n4497);
nand (n4493,n4494,n4496);
or (n4494,n4495,n3986);
not (n4495,n2138);
not (n4496,n2137);
nor (n4497,n4498,n3986);
not (n4498,n2195);
nand (n4499,n4491,n3986);
xor (n4500,n4470,n4472);
and (n4501,n4486,n4488);
and (n4502,n4468,n4477);
not (n4503,n4504);
nor (n4504,n4505,n4515);
nor (n4505,n4506,n4507);
xor (n4506,n4436,n4442);
or (n4507,n4508,n4514);
and (n4508,n4509,n4513);
xor (n4509,n4510,n4511);
xor (n4510,n3934,n3935);
or (n4511,n4512,n1770);
and (n4512,n4027,n4482);
xor (n4513,n4021,n4440);
and (n4514,n4510,n4511);
nor (n4515,n4516,n4517);
xor (n4516,n4509,n4513);
or (n4517,n4518,n4519);
and (n4518,n4478,n4481);
and (n4519,n4479,n4480);
nor (n4520,n4521,n4525);
and (n4521,n4522,n4523);
not (n4522,n4505);
not (n4523,n4524);
nand (n4524,n4516,n4517);
and (n4525,n4506,n4507);
not (n4526,n4527);
nand (n4527,n4528,n4532);
or (n4528,n4529,n4531);
not (n4529,n4530);
and (n4530,n4421,n4434);
not (n4531,n4447);
nand (n4532,n4458,n4449);
and (n4533,n4534,n4565);
and (n4534,n4535,n4549);
nand (n4535,n4536,n4538);
not (n4536,n4537);
xor (n4537,n4377,n4384);
not (n4538,n4539);
or (n4539,n4540,n4548);
and (n4540,n4541,n4544);
xor (n4541,n4542,n4543);
xor (n4542,n2271,n3235);
xor (n4543,n1099,n4381);
or (n4544,n4545,n1198);
and (n4545,n3991,n4546);
or (n4546,n4547,n2383);
and (n4547,n3872,n3873);
and (n4548,n4542,n4543);
nand (n4549,n4550,n4552);
not (n4550,n4551);
xor (n4551,n4541,n4544);
not (n4552,n4553);
or (n4553,n4554,n4564);
and (n4554,n4555,n4558);
xor (n4555,n4556,n4557);
xor (n4556,n3851,n3852);
xor (n4557,n3991,n4546);
nand (n4558,n4559,n4563);
nand (n4559,n4560,n1208);
or (n4560,n1206,n4561);
or (n4561,n4562,n2503);
and (n4562,n3887,n3888);
nand (n4563,n4561,n1206);
and (n4564,n4556,n4557);
nor (n4565,n4566,n4579);
nor (n4566,n4567,n4568);
xor (n4567,n4555,n4558);
or (n4568,n4569,n4578);
and (n4569,n4570,n4576);
xor (n4570,n4571,n4572);
xor (n4571,n3872,n3873);
nand (n4572,n4573,n4575);
or (n4573,n4574,n4561);
not (n4574,n3997);
nand (n4575,n4561,n4574);
or (n4576,n4577,n1212);
and (n4577,n4003,n4455);
and (n4578,n4571,n4572);
nor (n4579,n4580,n4581);
xor (n4580,n4570,n4576);
or (n4581,n4582,n4583);
and (n4582,n4450,n4454);
and (n4583,n4451,n4452);
nand (n4584,n4344,n4585);
not (n4585,n4586);
nor (n4586,n4587,n4592);
and (n4587,n4534,n4588);
nand (n4588,n4589,n4591);
or (n4589,n4566,n4590);
nand (n4590,n4580,n4581);
nand (n4591,n4567,n4568);
nand (n4592,n4593,n4597);
or (n4593,n4594,n4596);
not (n4594,n4595);
nor (n4595,n4550,n4552);
not (n4596,n4535);
nand (n4597,n4537,n4539);
nor (n4598,n4599,n4607);
and (n4599,n4600,n4408);
not (n4600,n4601);
or (n4601,n4602,n4603);
not (n4602,n4390);
not (n4603,n4604);
nand (n4604,n4605,n4606);
nand (n4605,n4392,n4405);
nand (n4606,n4348,n4375);
and (n4607,n4410,n4412);
nand (n4608,n4243,n4342);
or (n4609,n4610,n4734,n4757);
and (n4610,n4611,n4720);
xor (n4611,n4612,n4713);
xor (n4612,n4613,n4629);
xor (n4613,n4322,n4614);
or (n4614,n4615,n4616,n4628);
and (n4615,n4328,n4335);
and (n4616,n4335,n4617);
or (n4617,n4618,n4619,n4627);
and (n4618,n4367,n4369);
and (n4619,n4369,n4620);
or (n4620,n4621,n4622,n4626);
and (n4621,n4354,n4361);
and (n4622,n4361,n4623);
or (n4623,n4383,n4624,n4625);
and (n4624,n1195,n1197);
and (n4625,n1100,n1197);
and (n4626,n4354,n4623);
and (n4627,n4367,n4620);
and (n4628,n4328,n4617);
nand (n4629,n4630,n4712);
or (n4630,n4631,n4637);
not (n4631,n4632);
nor (n4632,n4633,n4636);
not (n4633,n4634);
nand (n4634,n4635,n4323);
not (n4635,n4318);
nor (n4636,n4323,n4635);
nand (n4637,n4638,n4646,n4673);
not (n4638,n4639);
nand (n4639,n4640,n4645);
or (n4640,n4641,n4643);
not (n4641,n4642);
and (n4642,n4371,n4350);
not (n4643,n4644);
or (n4644,n4394,n4331);
nand (n4645,n4394,n4331);
nand (n4646,n4647,n4671);
not (n4647,n4648);
nor (n4648,n4649,n4665);
and (n4649,n4650,n4655);
and (n4650,n4651,n4652);
or (n4651,n4378,n4357);
nand (n4652,n4653,n4654);
not (n4653,n4542);
not (n4654,n4381);
not (n4655,n4656);
nor (n4656,n4657,n4664);
and (n4657,n4658,n4661);
nand (n4658,n4659,n4660);
not (n4659,n4546);
not (n4660,n4556);
nor (n4661,n4662,n4663);
not (n4662,n4561);
not (n4663,n4571);
nor (n4664,n4659,n4660);
nand (n4665,n4666,n4670);
or (n4666,n4667,n4669);
not (n4667,n4668);
nor (n4668,n4653,n4654);
not (n4669,n4651);
nand (n4670,n4378,n4357);
and (n4671,n4644,n4672);
or (n4672,n4350,n4371);
nand (n4673,n4674,n4678,n4671);
and (n4674,n4650,n4675);
nor (n4675,n4676,n4677);
not (n4676,n4658);
and (n4677,n4662,n4663);
nand (n4678,n4679,n4698);
nor (n4679,n4680,n4692);
and (n4680,n4681,n4686);
and (n4681,n4682,n4683);
or (n4682,n4451,n4455);
nand (n4683,n4684,n4685);
not (n4684,n4431);
not (n4685,n4423);
nor (n4686,n4687,n4690);
and (n4687,n4688,n4689);
nand (n4688,n4427,n4437);
nand (n4689,n4440,n4510);
not (n4690,n4691);
or (n4691,n4437,n4427);
nand (n4692,n4693,n4697);
or (n4693,n4694,n4696);
not (n4694,n4695);
nor (n4695,n4684,n4685);
not (n4696,n4682);
nand (n4697,n4451,n4455);
nand (n4698,n4681,n4699,n4701);
and (n4699,n4691,n4700);
or (n4700,n4440,n4510);
nand (n4701,n4702,n4708);
or (n4702,n4703,n4706);
not (n4703,n4704);
and (n4704,n4705,n3982);
or (n4705,n4472,n3105);
not (n4706,n4707);
or (n4707,n4480,n4482);
nor (n4708,n4709,n4711);
and (n4709,n4707,n4710);
and (n4710,n4472,n3105);
and (n4711,n4480,n4482);
nand (n4712,n4631,n4637);
or (n4713,n4714,n4716,n4733);
and (n4714,n4715,n4120);
xor (n4715,n4398,n4617);
and (n4716,n4120,n4717);
or (n4717,n4718,n4721,n4732);
and (n4718,n4719,n4720);
xor (n4719,n4366,n4620);
xor (n4720,n4235,n4237);
and (n4721,n4720,n4722);
or (n4722,n4723,n4726,n4731);
and (n4723,n4724,n4725);
xor (n4724,n4387,n4623);
xor (n4725,n4238,n4240);
and (n4726,n4725,n4727);
or (n4727,n4728,n4729,n4730);
and (n4728,n1098,n2267);
and (n4729,n2267,n3988);
and (n4730,n1098,n3988);
and (n4731,n4724,n4727);
and (n4732,n4719,n4722);
and (n4733,n4715,n4717);
and (n4734,n4720,n4735);
or (n4735,n4736,n4739,n4756);
and (n4736,n4737,n4725);
xor (n4737,n4738,n4717);
xor (n4738,n4715,n4120);
and (n4739,n4725,n4740);
or (n4740,n4741,n4744,n4755);
and (n4741,n4742,n2267);
xor (n4742,n4743,n4722);
xor (n4743,n4719,n4720);
and (n4744,n2267,n4745);
or (n4745,n4746,n4749,n4754);
and (n4746,n4747,n3992);
xor (n4747,n4748,n4727);
xor (n4748,n4724,n4725);
and (n4749,n3992,n4750);
or (n4750,n4751,n4752,n4753);
and (n4751,n1096,n3998);
and (n4752,n3998,n4053);
and (n4753,n1096,n4053);
and (n4754,n4747,n4750);
and (n4755,n4742,n4745);
and (n4756,n4737,n4740);
and (n4757,n4611,n4735);
and (n4758,n4759,n4761);
xor (n4759,n4760,n4735);
xor (n4760,n4611,n4720);
and (n4761,n4762,n4764);
xor (n4762,n4763,n4740);
xor (n4763,n4737,n4725);
and (n4764,n4765,n4767);
xor (n4765,n4766,n4745);
xor (n4766,n4742,n2267);
and (n4767,n4768,n4770);
xor (n4768,n4769,n4750);
xor (n4769,n4747,n3992);
and (n4770,n1094,n4098);
xor (n4771,n4118,n4772);
and (n4772,n4759,n4773);
and (n4773,n4762,n4774);
and (n4774,n4765,n4775);
and (n4775,n4768,n4776);
and (n4776,n1094,n4099);
wire s0n4777,s1n4777,notn4777;
or (n4777,s0n4777,s1n4777);
not(notn4777,n1102);
and (s0n4777,notn4777,n4778);
and (s1n4777,n1102,n4781);
wire s0n4778,s1n4778,notn4778;
or (n4778,s0n4778,s1n4778);
not(notn4778,n1102);
and (s0n4778,notn4778,n4779);
and (s1n4778,n1102,n4780);
xor (n4779,n4762,n4764);
xor (n4780,n4762,n4774);
wire s0n4781,s1n4781,notn4781;
or (n4781,s0n4781,s1n4781);
not(notn4781,n1102);
and (s0n4781,notn4781,n4782);
and (s1n4781,n1102,n4899);
xor (n4782,n4783,n4889);
xor (n4783,n4784,n4852);
nand (n4784,n4785,n4851);
or (n4785,n4786,n4811);
not (n4786,n4787);
xor (n4787,n4788,n4798);
xor (n4788,n4789,n4792);
or (n4789,n4790,n4791);
and (n4790,n4250,n4255);
and (n4791,n4251,n4253);
xor (n4792,n4793,n4255);
xor (n4793,n4794,n4796);
wire s0n4794,s1n4794,notn4794;
or (n4794,s0n4794,s1n4794);
not(notn4794,n1102);
and (s0n4794,notn4794,1'b0);
and (s1n4794,n1102,n4795);
wire s0n4796,s1n4796,notn4796;
or (n4796,s0n4796,s1n4796);
not(notn4796,n1102);
and (s0n4796,notn4796,1'b0);
and (s1n4796,n1102,n4797);
nand (n4798,n4799,n4803,n4804);
nand (n4799,n4647,n4800);
and (n4800,n4671,n4801);
and (n4801,n4802,n4634);
or (n4802,n4282,n4249);
nand (n4803,n4800,n4674,n4678);
nor (n4804,n4805,n4806);
and (n4805,n4639,n4801);
nand (n4806,n4807,n4810);
or (n4807,n4808,n4809);
not (n4808,n4802);
not (n4809,n4636);
nand (n4810,n4282,n4249);
nand (n4811,n4812,n4850);
or (n4812,n4813,n4832);
not (n4813,n4814);
xnor (n4814,n4815,n4820);
or (n4815,n4816,n4818);
and (n4816,n4817,n4282);
not (n4817,n4788);
and (n4818,n4792,n4819);
not (n4819,n4789);
nand (n4820,n4821,n4831);
or (n4821,n4819,n4822);
nand (n4822,n4823,n4830);
or (n4823,n4255,n4824);
not (n4824,n4825);
or (n4825,n4826,n4827);
and (n4826,n4793,n4255);
and (n4827,n4828,n4829);
not (n4828,n4794);
not (n4829,n4796);
or (n4830,n4825,n4256);
nand (n4831,n4822,n4819);
nand (n4832,n4833,n4847,n4849);
nand (n4833,n4834,n4835,n4586);
nand (n4834,n4415,n4533);
nand (n4835,n4836,n4845);
or (n4836,n4837,n4843);
nand (n4837,n4246,n4838);
nand (n4838,n4839,n4842);
or (n4839,n4840,n4841);
and (n4840,n4248,n4302);
and (n4841,n4249,n4281);
xor (n4842,n4817,n4282);
not (n4843,n4844);
nand (n4844,n4408,n4339);
nand (n4845,n4601,n4846);
nor (n4846,n4837,n4607);
nand (n4847,n4835,n4848);
nand (n4848,n4345,n4843);
or (n4849,n4839,n4842);
nand (n4850,n4813,n4832);
nand (n4851,n4811,n4786);
or (n4852,n4853,n4865,n4888);
and (n4853,n4811,n4854);
nand (n4854,n4855,n4864);
or (n4855,n4856,n4858);
not (n4856,n4857);
not (n4857,n4248);
nand (n4858,n4859,n4861,n4862);
nand (n4859,n4647,n4860);
and (n4860,n4671,n4634);
nand (n4861,n4860,n4674,n4678);
nor (n4862,n4863,n4636);
and (n4863,n4639,n4634);
nand (n4864,n4856,n4858);
and (n4865,n4854,n4866);
or (n4866,n4867,n4882,n4887);
and (n4867,n4629,n4868);
nand (n4868,n4869,n4881);
or (n4869,n4870,n4872);
not (n4870,n4871);
and (n4871,n4838,n4849);
nand (n4872,n4873,n4875,n4876);
nand (n4873,n4874,n4415,n4533);
not (n4874,n4848);
nand (n4875,n4874,n4585);
nor (n4876,n4877,n4878);
and (n4877,n4600,n4843);
nand (n4878,n4879,n4246);
or (n4879,n4880,n4338);
not (n4880,n4607);
nand (n4881,n4870,n4872);
and (n4882,n4629,n4883);
or (n4883,n4884,n4885,n4886);
and (n4884,n4120,n4241);
and (n4885,n4120,n4609);
and (n4886,n4241,n4609);
and (n4887,n4868,n4883);
and (n4888,n4811,n4866);
and (n4889,n4890,n4895);
xor (n4890,n4891,n4866);
nor (n4891,n4853,n4892);
and (n4892,n4893,n4894);
not (n4893,n4854);
not (n4894,n4811);
and (n4895,n4896,n4898);
xor (n4896,n4897,n4883);
xor (n4897,n4868,n4629);
and (n4898,n4118,n4758);
xor (n4899,n4783,n4900);
and (n4900,n4890,n4901);
and (n4901,n4896,n4902);
and (n4902,n4118,n4772);
wire s0n4903,s1n4903,notn4903;
or (n4903,s0n4903,s1n4903);
not(notn4903,n1102);
and (s0n4903,notn4903,n4904);
and (s1n4903,n1102,n4921);
xor (n4904,n4905,n4920);
xor (n4905,n4906,n4916);
nand (n4906,n4907,n4915);
or (n4907,n4908,n4811);
not (n4908,n4909);
nand (n4909,n4910,n4914);
or (n4910,n4911,n4822);
or (n4911,n4912,n4913);
and (n4912,n4788,n4798);
and (n4913,n4789,n4792);
nand (n4914,n4911,n4822);
nand (n4915,n4811,n4908);
or (n4916,n4917,n4918,n4919);
and (n4917,n4811,n4787);
and (n4918,n4787,n4852);
and (n4919,n4811,n4852);
and (n4920,n4783,n4889);
xor (n4921,n4905,n4922);
and (n4922,n4783,n4900);
and (n4923,n4924,n806);
not (n4924,n4925);
nor (n4925,n1184,n807,n800,n802);
and (n4926,n4927,n6);
wire s0n4927,s1n4927,notn4927;
or (n4927,s0n4927,s1n4927);
not(notn4927,n1194);
and (s0n4927,notn4927,1'b0);
and (s1n4927,n1194,n1089);
and (n4928,n1089,n4929);
not (n4929,n1229);
and (n4930,n4931,n7029);
wire s0n4931,s1n4931,notn4931;
or (n4931,s0n4931,s1n4931);
not(notn4931,n7024);
and (s0n4931,notn4931,n4932);
and (s1n4931,n7024,1'b0);
wire s0n4932,s1n4932,notn4932;
or (n4932,s0n4932,s1n4932);
not(notn4932,n6998);
and (s0n4932,notn4932,n4933);
and (s1n4932,n6998,1'b1);
wire s0n4933,s1n4933,notn4933;
or (n4933,s0n4933,s1n4933);
not(notn4933,n6991);
and (s0n4933,notn4933,1'b0);
and (s1n4933,n6991,n4934);
xor (n4934,n4935,n6974);
xor (n4935,n4936,n6930);
xor (n4936,n4937,n6865);
xor (n4937,n4938,n6426);
xor (n4938,n4939,n6394);
xnor (n4939,n4940,n5683);
or (n4940,n4941,n5096,n5682);
not (n4941,n4942);
or (n4942,n4943,n5053);
not (n4943,n4944);
nand (n4944,n4945,n5010);
nor (n4945,n4946,n4993);
nand (n4946,n4947,n4980,n4984,n4988);
nand (n4947,n4948,n4977);
not (n4948,n4949);
nand (n4949,n4950,n1331);
not (n4950,n4951);
nand (n4951,n4952,n4972);
nand (n4952,n4953,n4967);
not (n4953,n4954);
nand (n4954,n4955,n4961);
nand (n4955,n4956,n1183);
nand (n4956,n4957,n4958,n4960);
nand (n4957,n652,n1344,n1107);
not (n4958,n4959);
nor (n4959,n653,n726,n1106,n1107);
nand (n4960,n7,n653);
nor (n4961,n4962,n4966);
nor (n4962,n4963,n1236);
nand (n4963,n4964,n4965);
or (n4964,n726,n653);
not (n4965,n1230);
not (n4966,n1243);
and (n4967,n4968,n4969,n1231);
nand (n4968,n4956,n1187);
not (n4969,n4970);
and (n4970,n4971,n817);
not (n4971,n4963);
nand (n4972,n4973,n4955,n4974,n4975);
nand (n4973,n1186,n4956);
and (n4974,n4969,n1237);
nor (n4975,n4976,n4966);
and (n4976,n4971,n1183);
wire s0n4977,s1n4977,notn4977;
or (n4977,s0n4977,s1n4977);
not(notn4977,n4978);
and (s0n4977,notn4977,n2303);
and (s1n4977,n4978,n2367);
not (n4978,n4979);
nand (n4979,n7,n653,n726);
nand (n4980,n4981,n4983);
not (n4981,n4982);
nand (n4982,n4950,n1316);
wire s0n4983,s1n4983,notn4983;
or (n4983,s0n4983,s1n4983);
not(notn4983,n4978);
and (s0n4983,notn4983,n2291);
and (s1n4983,n4978,n2355);
nand (n4984,n4985,n4987);
not (n4985,n4986);
nand (n4986,n4950,n1265);
wire s0n4987,s1n4987,notn4987;
or (n4987,s0n4987,s1n4987);
not(notn4987,n4978);
and (s0n4987,notn4987,n2320);
and (s1n4987,n4978,n2374);
nand (n4988,n4989,n4992);
and (n4989,n4990,n1246);
and (n4990,n4952,n4991);
not (n4991,n4972);
wire s0n4992,s1n4992,notn4992;
or (n4992,s0n4992,s1n4992);
not(notn4992,n4978);
and (s0n4992,notn4992,n2308);
and (s1n4992,n4978,n2343);
nand (n4993,n4994,n4997,n5000,n5007);
nand (n4994,n4995,n4996);
and (n4995,n4990,n1316);
wire s0n4996,s1n4996,notn4996;
or (n4996,s0n4996,s1n4996);
not(notn4996,n4978);
and (s0n4996,notn4996,n2285);
and (s1n4996,n4978,n2349);
nand (n4997,n4998,n4999);
and (n4998,n4990,n1265);
wire s0n4999,s1n4999,notn4999;
or (n4999,s0n4999,s1n4999);
not(notn4999,n4978);
and (s0n4999,notn4999,n2315);
and (s1n4999,n4978,n2341);
nand (n5000,n5001,n5006);
not (n5001,n5002);
nand (n5002,n5003,n1246);
not (n5003,n5004);
nand (n5004,n4953,n4967,n5005);
nand (n5005,n4973,n4975,n1237);
wire s0n5006,s1n5006,notn5006;
or (n5006,s0n5006,s1n5006);
not(notn5006,n4978);
and (s0n5006,notn5006,n2313);
and (s1n5006,n4978,n2335);
nand (n5007,n5008,n5009);
and (n5008,n4990,n1331);
wire s0n5009,s1n5009,notn5009;
or (n5009,s0n5009,s1n5009);
not(notn5009,n4978);
and (s0n5009,notn5009,n2298);
and (s1n5009,n4978,n2362);
nor (n5010,n5011,n5022);
nand (n5011,n5012,n5015,n5018);
nand (n5012,n5013,n5014);
and (n5013,n5003,n1265);
wire s0n5014,s1n5014,notn5014;
or (n5014,s0n5014,s1n5014);
not(notn5014,n4978);
and (s0n5014,notn5014,n2311);
and (s1n5014,n4978,n2339);
nand (n5015,n5016,n5017);
and (n5016,n5003,n1331);
wire s0n5017,s1n5017,notn5017;
or (n5017,s0n5017,s1n5017);
not(notn5017,n4978);
and (s0n5017,notn5017,n2301);
and (s1n5017,n4978,n2365);
nand (n5018,n5019,n5021);
not (n5019,n5020);
nand (n5020,n5003,n1316);
wire s0n5021,s1n5021,notn5021;
or (n5021,s0n5021,s1n5021);
not(notn5021,n4978);
and (s0n5021,notn5021,n2289);
and (s1n5021,n4978,n2353);
nand (n5022,n5023,n5027);
or (n5023,n5024,n5026);
not (n5024,n5025);
wire s0n5025,s1n5025,notn5025;
or (n5025,s0n5025,s1n5025);
not(notn5025,n4978);
and (s0n5025,notn5025,n2325);
and (s1n5025,n4978,n2372);
nand (n5026,n4950,n1246);
nor (n5027,n5028,n5043);
nand (n5028,n5029,n5038);
or (n5029,n5030,n5036);
not (n5030,n5031);
and (n5031,n5032,n1316);
nand (n5032,n1259,n5033,n5035);
not (n5033,n5034);
and (n5034,n4971,n4925);
nand (n5035,n4956,n817);
not (n5036,n5037);
wire s0n5037,s1n5037,notn5037;
or (n5037,s0n5037,s1n5037);
not(notn5037,n4978);
and (s0n5037,notn5037,n2293);
and (s1n5037,n4978,n2357);
or (n5038,n5039,n5041);
not (n5039,n5040);
and (n5040,n5032,n1246);
not (n5041,n5042);
wire s0n5042,s1n5042,notn5042;
or (n5042,s0n5042,s1n5042);
not(notn5042,n4978);
and (s0n5042,notn5042,n2327);
and (s1n5042,n4978,n2377);
nand (n5043,n5044,n5048);
or (n5044,n5045,n5046);
nand (n5045,n5032,n1331);
not (n5046,n5047);
wire s0n5047,s1n5047,notn5047;
or (n5047,s0n5047,s1n5047);
not(notn5047,n4978);
and (s0n5047,notn5047,n2305);
and (s1n5047,n4978,n2369);
or (n5048,n5049,n5051);
not (n5049,n5050);
and (n5050,n5032,n1265);
not (n5051,n5052);
wire s0n5052,s1n5052,notn5052;
or (n5052,s0n5052,s1n5052);
not(notn5052,n4978);
and (s0n5052,notn5052,n2322);
and (s1n5052,n4978,n2379);
not (n5053,n5054);
nand (n5054,n5055,n5078,n5087);
nor (n5055,n5056,n5073);
nand (n5056,n5057,n5059,n5060);
nand (n5057,n5058,n5042);
not (n5058,n5026);
nand (n5059,n5019,n4983);
nor (n5060,n5061,n5066);
nand (n5061,n5062,n5064);
or (n5062,n5045,n5063);
not (n5063,n4996);
or (n5064,n5049,n5065);
not (n5065,n4992);
nand (n5066,n5067,n5070);
or (n5067,n5030,n5068);
not (n5068,n5069);
wire s0n5069,s1n5069,notn5069;
or (n5069,s0n5069,s1n5069);
not(notn5069,n4978);
and (s0n5069,notn5069,n2287);
and (s1n5069,n4978,n2351);
or (n5070,n5039,n5071);
not (n5071,n5072);
wire s0n5072,s1n5072,notn5072;
or (n5072,s0n5072,s1n5072);
not(notn5072,n4978);
and (s0n5072,notn5072,n2317);
and (s1n5072,n4978,n2337);
nand (n5073,n5074,n5077);
or (n5074,n5075,n5076);
not (n5075,n4987);
not (n5076,n5013);
nand (n5077,n5016,n4977);
nor (n5078,n5079,n5082);
nand (n5079,n5080,n5081);
or (n5080,n5051,n4986);
nand (n5081,n4948,n5047);
nand (n5082,n5083,n5086);
or (n5083,n5084,n5085);
not (n5084,n5017);
not (n5085,n5008);
nand (n5086,n4989,n5006);
nor (n5087,n5088,n5093);
nand (n5088,n5089,n5092);
or (n5089,n5090,n5091);
not (n5090,n5014);
not (n5091,n4998);
nand (n5092,n4995,n5021);
nand (n5093,n5094,n5095);
or (n5094,n5024,n5002);
nand (n5095,n4981,n5037);
and (n5096,n4944,n5097);
or (n5097,n5098,n5182,n5681);
and (n5098,n5099,n5153);
nand (n5099,n5100,n5126,n5139);
nor (n5100,n5101,n5120);
nand (n5101,n5102,n5104,n5106);
nand (n5102,n5058,n5103);
wire s0n5103,s1n5103,notn5103;
or (n5103,s0n5103,s1n5103);
not(notn5103,n4978);
and (s0n5103,notn5103,n2427);
and (s1n5103,n4978,n2493);
nand (n5104,n5016,n5105);
wire s0n5105,s1n5105,notn5105;
or (n5105,s0n5105,s1n5105);
not(notn5105,n4978);
and (s0n5105,notn5105,n2407);
and (s1n5105,n4978,n2454);
nor (n5106,n5107,n5114);
nand (n5107,n5108,n5111);
or (n5108,n5109,n5049);
not (n5109,n5110);
wire s0n5110,s1n5110,notn5110;
or (n5110,s0n5110,s1n5110);
not(notn5110,n4978);
and (s0n5110,notn5110,n2434);
and (s1n5110,n4978,n2482);
nand (n5111,n5112,n5113);
not (n5112,n5045);
wire s0n5113,s1n5113,notn5113;
or (n5113,s0n5113,s1n5113);
not(notn5113,n4978);
and (s0n5113,notn5113,n2411);
and (s1n5113,n4978,n2444);
nand (n5114,n5115,n5118);
or (n5115,n5116,n5039);
not (n5116,n5117);
wire s0n5117,s1n5117,notn5117;
or (n5117,s0n5117,s1n5117);
not(notn5117,n4978);
and (s0n5117,notn5117,n2432);
and (s1n5117,n4978,n2496);
nand (n5118,n5031,n5119);
wire s0n5119,s1n5119,notn5119;
or (n5119,s0n5119,s1n5119);
not(notn5119,n4978);
and (s0n5119,notn5119,n2399);
and (s1n5119,n4978,n2461);
nand (n5120,n5121,n5124);
or (n5121,n5122,n5076);
not (n5122,n5123);
wire s0n5123,s1n5123,notn5123;
or (n5123,s0n5123,s1n5123);
not(notn5123,n4978);
and (s0n5123,notn5123,n2424);
and (s1n5123,n4978,n2475);
nand (n5124,n5019,n5125);
wire s0n5125,s1n5125,notn5125;
or (n5125,s0n5125,s1n5125);
not(notn5125,n4978);
and (s0n5125,notn5125,n2395);
and (s1n5125,n4978,n2470);
nor (n5126,n5127,n5133);
nand (n5127,n5128,n5131);
or (n5128,n5129,n4986);
not (n5129,n5130);
wire s0n5130,s1n5130,notn5130;
or (n5130,s0n5130,s1n5130);
not(notn5130,n4978);
and (s0n5130,notn5130,n2429);
and (s1n5130,n4978,n2479);
nand (n5131,n4981,n5132);
wire s0n5132,s1n5132,notn5132;
or (n5132,s0n5132,s1n5132);
not(notn5132,n4978);
and (s0n5132,notn5132,n2397);
and (s1n5132,n4978,n2459);
nand (n5133,n5134,n5137);
or (n5134,n5135,n4949);
not (n5135,n5136);
wire s0n5136,s1n5136,notn5136;
or (n5136,s0n5136,s1n5136);
not(notn5136,n4978);
and (s0n5136,notn5136,n2409);
and (s1n5136,n4978,n2442);
nand (n5137,n4995,n5138);
wire s0n5138,s1n5138,notn5138;
or (n5138,s0n5138,s1n5138);
not(notn5138,n4978);
and (s0n5138,notn5138,n2391);
and (s1n5138,n4978,n2451);
nor (n5139,n5140,n5147);
nand (n5140,n5141,n5145);
or (n5141,n5142,n5144);
not (n5142,n5143);
wire s0n5143,s1n5143,notn5143;
or (n5143,s0n5143,s1n5143);
not(notn5143,n4978);
and (s0n5143,notn5143,n2414);
and (s1n5143,n4978,n2485);
not (n5144,n4989);
nand (n5145,n4998,n5146);
wire s0n5146,s1n5146,notn5146;
or (n5146,s0n5146,s1n5146);
not(notn5146,n4978);
and (s0n5146,notn5146,n2422);
and (s1n5146,n4978,n2476);
nand (n5147,n5148,n5151);
or (n5148,n5149,n5002);
not (n5149,n5150);
wire s0n5150,s1n5150,notn5150;
or (n5150,s0n5150,s1n5150);
not(notn5150,n4978);
and (s0n5150,notn5150,n2420);
and (s1n5150,n4978,n2490);
nand (n5151,n5008,n5152);
wire s0n5152,s1n5152,notn5152;
or (n5152,s0n5152,s1n5152);
not(notn5152,n4978);
and (s0n5152,notn5152,n2404);
and (s1n5152,n4978,n2449);
nand (n5153,n5154,n5165);
nor (n5154,n5155,n5160);
nand (n5155,n5156,n5157,n5158,n5159);
nand (n5156,n4948,n5113);
nand (n5157,n4981,n5119);
nand (n5158,n4985,n5110);
nand (n5159,n4989,n5150);
nand (n5160,n5161,n5162,n5163,n5164);
nand (n5161,n4995,n5125);
nand (n5162,n5001,n5103);
nand (n5163,n5008,n5105);
nand (n5164,n4998,n5123);
nor (n5165,n5166,n5179);
nand (n5166,n5167,n5168,n5169);
nand (n5167,n5058,n5117);
nand (n5168,n5016,n5136);
nor (n5169,n5170,n5173);
nand (n5170,n5171,n5172);
or (n5171,n5142,n5049);
nand (n5172,n5112,n5138);
nand (n5173,n5174,n5177);
or (n5174,n5175,n5030);
not (n5175,n5176);
wire s0n5176,s1n5176,notn5176;
or (n5176,s0n5176,s1n5176);
not(notn5176,n4978);
and (s0n5176,notn5176,n2393);
and (s1n5176,n4978,n2467);
nand (n5177,n5178,n5040);
wire s0n5178,s1n5178,notn5178;
or (n5178,s0n5178,s1n5178);
not(notn5178,n4978);
and (s0n5178,notn5178,n2418);
and (s1n5178,n4978,n2499);
nand (n5179,n5180,n5181);
or (n5180,n5129,n5076);
nand (n5181,n5019,n5132);
and (n5182,n5099,n5183);
or (n5183,n5184,n5261,n5680);
and (n5184,n5185,n5230);
nand (n5185,n5186,n5205);
nor (n5186,n5187,n5196);
nand (n5187,n5188,n5190,n5192,n5194);
nand (n5188,n4985,n5189);
wire s0n5189,s1n5189,notn5189;
or (n5189,s0n5189,s1n5189);
not(notn5189,n4978);
and (s0n5189,notn5189,n2550);
and (s1n5189,n4978,n2605);
nand (n5190,n4948,n5191);
wire s0n5191,s1n5191,notn5191;
or (n5191,s0n5191,s1n5191);
not(notn5191,n4978);
and (s0n5191,notn5191,n2537);
and (s1n5191,n4978,n2583);
nand (n5192,n4989,n5193);
wire s0n5193,s1n5193,notn5193;
or (n5193,s0n5193,s1n5193);
not(notn5193,n4978);
and (s0n5193,notn5193,n2508);
and (s1n5193,n4978,n2561);
nand (n5194,n4981,n5195);
wire s0n5195,s1n5195,notn5195;
or (n5195,s0n5195,s1n5195);
not(notn5195,n4978);
and (s0n5195,notn5195,n2524);
and (s1n5195,n4978,n2598);
nand (n5196,n5197,n5199,n5201,n5203);
nand (n5197,n4995,n5198);
wire s0n5198,s1n5198,notn5198;
or (n5198,s0n5198,s1n5198);
not(notn5198,n4978);
and (s0n5198,notn5198,n2529);
and (s1n5198,n4978,n2579);
nand (n5199,n5001,n5200);
wire s0n5200,s1n5200,notn5200;
or (n5200,s0n5200,s1n5200);
not(notn5200,n4978);
and (s0n5200,notn5200,n2512);
and (s1n5200,n4978,n2564);
nand (n5201,n4998,n5202);
wire s0n5202,s1n5202,notn5202;
or (n5202,s0n5202,s1n5202);
not(notn5202,n4978);
and (s0n5202,notn5202,n2517);
and (s1n5202,n4978,n2571);
nand (n5203,n5008,n5204);
wire s0n5204,s1n5204,notn5204;
or (n5204,s0n5204,s1n5204);
not(notn5204,n4978);
and (s0n5204,notn5204,n2542);
and (s1n5204,n4978,n2577);
nor (n5205,n5206,n5224);
nand (n5206,n5207,n5209,n5211);
nand (n5207,n5058,n5208);
wire s0n5208,s1n5208,notn5208;
or (n5208,s0n5208,s1n5208);
not(notn5208,n4978);
and (s0n5208,notn5208,n2548);
and (s1n5208,n4978,n2587);
nand (n5209,n5016,n5210);
wire s0n5210,s1n5210,notn5210;
or (n5210,s0n5210,s1n5210);
not(notn5210,n4978);
and (s0n5210,notn5210,n2545);
and (s1n5210,n4978,n2581);
nor (n5211,n5212,n5218);
nand (n5212,n5213,n5216);
or (n5213,n5214,n5045);
not (n5214,n5215);
wire s0n5215,s1n5215,notn5215;
or (n5215,s0n5215,s1n5215);
not(notn5215,n4978);
and (s0n5215,notn5215,n2539);
and (s1n5215,n4978,n2585);
nand (n5216,n5050,n5217);
wire s0n5217,s1n5217,notn5217;
or (n5217,s0n5217,s1n5217);
not(notn5217,n4978);
and (s0n5217,notn5217,n2555);
and (s1n5217,n4978,n2602);
nand (n5218,n5219,n5222);
or (n5219,n5220,n5039);
not (n5220,n5221);
wire s0n5221,s1n5221,notn5221;
or (n5221,s0n5221,s1n5221);
not(notn5221,n4978);
and (s0n5221,notn5221,n2553);
and (s1n5221,n4978,n2607);
nand (n5222,n5031,n5223);
wire s0n5223,s1n5223,notn5223;
or (n5223,s0n5223,s1n5223);
not(notn5223,n4978);
and (s0n5223,notn5223,n2526);
and (s1n5223,n4978,n2600);
nand (n5224,n5225,n5228);
or (n5225,n5226,n5076);
not (n5226,n5227);
wire s0n5227,s1n5227,notn5227;
or (n5227,s0n5227,s1n5227);
not(notn5227,n4978);
and (s0n5227,notn5227,n2519);
and (s1n5227,n4978,n2567);
nand (n5228,n5019,n5229);
wire s0n5229,s1n5229,notn5229;
or (n5229,s0n5229,s1n5229);
not(notn5229,n4978);
and (s0n5229,notn5229,n2533);
and (s1n5229,n4978,n2596);
nand (n5230,n5231,n5242);
nor (n5231,n5232,n5237);
nand (n5232,n5233,n5234,n5235,n5236);
nand (n5233,n4995,n5229);
nand (n5234,n4981,n5223);
nand (n5235,n4985,n5217);
nand (n5236,n4948,n5215);
nand (n5237,n5238,n5239,n5240,n5241);
nand (n5238,n5001,n5208);
nand (n5239,n4989,n5200);
nand (n5240,n4998,n5227);
nand (n5241,n5008,n5210);
nor (n5242,n5243,n5257);
nand (n5243,n5244,n5245,n5246);
nand (n5244,n5058,n5221);
nand (n5245,n5016,n5191);
nor (n5246,n5247,n5251);
nand (n5247,n5248,n5250);
or (n5248,n5249,n5049);
not (n5249,n5193);
nand (n5250,n5112,n5198);
nand (n5251,n5252,n5255);
or (n5252,n5253,n5030);
not (n5253,n5254);
wire s0n5254,s1n5254,notn5254;
or (n5254,s0n5254,s1n5254);
not(notn5254,n4978);
and (s0n5254,notn5254,n2531);
and (s1n5254,n4978,n2594);
nand (n5255,n5040,n5256);
wire s0n5256,s1n5256,notn5256;
or (n5256,s0n5256,s1n5256);
not(notn5256,n4978);
and (s0n5256,notn5256,n2515);
and (s1n5256,n4978,n2569);
nand (n5257,n5258,n5260);
or (n5258,n5259,n5020);
not (n5259,n5195);
nand (n5260,n5013,n5189);
and (n5261,n5185,n5262);
or (n5262,n5263,n5338,n5679);
and (n5263,n5264,n5308);
nand (n5264,n5265,n5284);
nor (n5265,n5266,n5275);
nand (n5266,n5267,n5269,n5271,n5273);
nand (n5267,n4995,n5268);
wire s0n5268,s1n5268,notn5268;
or (n5268,s0n5268,s1n5268);
not(notn5268,n4978);
and (s0n5268,notn5268,n2646);
and (s1n5268,n4978,n2706);
nand (n5269,n4985,n5270);
wire s0n5270,s1n5270,notn5270;
or (n5270,s0n5270,s1n5270);
not(notn5270,n4978);
and (s0n5270,notn5270,n2658);
and (s1n5270,n4978,n2718);
nand (n5271,n4948,n5272);
wire s0n5272,s1n5272,notn5272;
or (n5272,s0n5272,s1n5272);
not(notn5272,n4978);
and (s0n5272,notn5272,n2618);
and (s1n5272,n4978,n2691);
nand (n5273,n4981,n5274);
wire s0n5274,s1n5274,notn5274;
or (n5274,s0n5274,s1n5274);
not(notn5274,n4978);
and (s0n5274,notn5274,n2635);
and (s1n5274,n4978,n2698);
nand (n5275,n5276,n5278,n5280,n5282);
nand (n5276,n5001,n5277);
wire s0n5277,s1n5277,notn5277;
or (n5277,s0n5277,s1n5277);
not(notn5277,n4978);
and (s0n5277,notn5277,n2669);
and (s1n5277,n4978,n2729);
nand (n5278,n4989,n5279);
wire s0n5279,s1n5279,notn5279;
or (n5279,s0n5279,s1n5279);
not(notn5279,n4978);
and (s0n5279,notn5279,n2666);
and (s1n5279,n4978,n2726);
nand (n5280,n4998,n5281);
wire s0n5281,s1n5281,notn5281;
or (n5281,s0n5281,s1n5281);
not(notn5281,n4978);
and (s0n5281,notn5281,n2651);
and (s1n5281,n4978,n2711);
nand (n5282,n5008,n5283);
wire s0n5283,s1n5283,notn5283;
or (n5283,s0n5283,s1n5283);
not(notn5283,n4978);
and (s0n5283,notn5283,n2630);
and (s1n5283,n4978,n2687);
nor (n5284,n5285,n5292);
nand (n5285,n5286,n5288,n5290);
nand (n5286,n5019,n5287);
wire s0n5287,s1n5287,notn5287;
or (n5287,s0n5287,s1n5287);
not(notn5287,n4978);
and (s0n5287,notn5287,n2637);
and (s1n5287,n4978,n2696);
nand (n5288,n5013,n5289);
wire s0n5289,s1n5289,notn5289;
or (n5289,s0n5289,s1n5289);
not(notn5289,n4978);
and (s0n5289,notn5289,n2655);
and (s1n5289,n4978,n2715);
nand (n5290,n5016,n5291);
wire s0n5291,s1n5291,notn5291;
or (n5291,s0n5291,s1n5291);
not(notn5291,n4978);
and (s0n5291,notn5291,n2620);
and (s1n5291,n4978,n2689);
nand (n5292,n5293,n5296);
or (n5293,n5294,n5026);
not (n5294,n5295);
wire s0n5295,s1n5295,notn5295;
or (n5295,s0n5295,s1n5295);
not(notn5295,n4978);
and (s0n5295,notn5295,n2672);
and (s1n5295,n4978,n2732);
nor (n5296,n5297,n5303);
nand (n5297,n5298,n5301);
or (n5298,n5299,n5049);
not (n5299,n5300);
wire s0n5300,s1n5300,notn5300;
or (n5300,s0n5300,s1n5300);
not(notn5300,n4978);
and (s0n5300,notn5300,n2661);
and (s1n5300,n4978,n2721);
nand (n5301,n5112,n5302);
wire s0n5302,s1n5302,notn5302;
or (n5302,s0n5302,s1n5302);
not(notn5302,n4978);
and (s0n5302,notn5302,n2627);
and (s1n5302,n4978,n2685);
nand (n5303,n5304,n5306);
nand (n5304,n5031,n5305);
wire s0n5305,s1n5305,notn5305;
or (n5305,s0n5305,s1n5305);
not(notn5305,n4978);
and (s0n5305,notn5305,n2643);
and (s1n5305,n4978,n2704);
nand (n5306,n5040,n5307);
wire s0n5307,s1n5307,notn5307;
or (n5307,s0n5307,s1n5307);
not(notn5307,n4978);
and (s0n5307,notn5307,n2675);
and (s1n5307,n4978,n2735);
nand (n5308,n5309,n5322);
nor (n5309,n5310,n5315);
nand (n5310,n5311,n5312,n5313,n5314);
nand (n5311,n4985,n5289);
nand (n5312,n4948,n5291);
nand (n5313,n4995,n5302);
nand (n5314,n4981,n5287);
nand (n5315,n5316,n5317,n5318,n5320);
nand (n5316,n4989,n5300);
nand (n5317,n5001,n5279);
nand (n5318,n5008,n5319);
wire s0n5319,s1n5319,notn5319;
or (n5319,s0n5319,s1n5319);
not(notn5319,n4978);
and (s0n5319,notn5319,n2625);
and (s1n5319,n4978,n2683);
nand (n5320,n4998,n5321);
wire s0n5321,s1n5321,notn5321;
or (n5321,s0n5321,s1n5321);
not(notn5321,n4978);
and (s0n5321,notn5321,n2652);
and (s1n5321,n4978,n2712);
nor (n5322,n5323,n5334);
nand (n5323,n5324,n5325,n5326);
nand (n5324,n5058,n5277);
nand (n5325,n5016,n5283);
nor (n5326,n5327,n5331);
nand (n5327,n5328,n5330);
or (n5328,n5329,n5049);
not (n5329,n5270);
nand (n5330,n5112,n5272);
nand (n5331,n5332,n5333);
or (n5332,n5294,n5039);
nand (n5333,n5031,n5274);
nand (n5334,n5335,n5337);
or (n5335,n5336,n5076);
not (n5336,n5281);
nand (n5337,n5019,n5268);
and (n5338,n5308,n5339);
or (n5339,n5340,n5423,n5678);
and (n5340,n5341,n5386);
nand (n5341,n5342,n5361);
nor (n5342,n5343,n5352);
nand (n5343,n5344,n5346,n5348,n5350);
nand (n5344,n4989,n5345);
wire s0n5345,s1n5345,notn5345;
or (n5345,s0n5345,s1n5345);
not(notn5345,n4978);
and (s0n5345,notn5345,n2794);
and (s1n5345,n4978,n2851);
nand (n5346,n4985,n5347);
wire s0n5347,s1n5347,notn5347;
or (n5347,s0n5347,s1n5347);
not(notn5347,n4978);
and (s0n5347,notn5347,n2786);
and (s1n5347,n4978,n2843);
nand (n5348,n4948,n5349);
wire s0n5349,s1n5349,notn5349;
or (n5349,s0n5349,s1n5349);
not(notn5349,n4978);
and (s0n5349,notn5349,n2748);
and (s1n5349,n4978,n2812);
nand (n5350,n4981,n5351);
wire s0n5351,s1n5351,notn5351;
or (n5351,s0n5351,s1n5351);
not(notn5351,n4978);
and (s0n5351,notn5351,n2765);
and (s1n5351,n4978,n2825);
nand (n5352,n5353,n5355,n5357,n5359);
nand (n5353,n4995,n5354);
wire s0n5354,s1n5354,notn5354;
or (n5354,s0n5354,s1n5354);
not(notn5354,n4978);
and (s0n5354,notn5354,n2774);
and (s1n5354,n4978,n2831);
nand (n5355,n4998,n5356);
wire s0n5356,s1n5356,notn5356;
or (n5356,s0n5356,s1n5356);
not(notn5356,n4978);
and (s0n5356,notn5356,n2779);
and (s1n5356,n4978,n2836);
nand (n5357,n5001,n5358);
wire s0n5358,s1n5358,notn5358;
or (n5358,s0n5358,s1n5358);
not(notn5358,n4978);
and (s0n5358,notn5358,n2797);
and (s1n5358,n4978,n2854);
nand (n5359,n5008,n5360);
wire s0n5360,s1n5360,notn5360;
or (n5360,s0n5360,s1n5360);
not(notn5360,n4978);
and (s0n5360,notn5360,n2758);
and (s1n5360,n4978,n2819);
nor (n5361,n5362,n5380);
nand (n5362,n5363,n5365,n5367);
nand (n5363,n5364,n5016);
wire s0n5364,s1n5364,notn5364;
or (n5364,s0n5364,s1n5364);
not(notn5364,n4978);
and (s0n5364,notn5364,n2746);
and (s1n5364,n4978,n2810);
nand (n5365,n5058,n5366);
wire s0n5366,s1n5366,notn5366;
or (n5366,s0n5366,s1n5366);
not(notn5366,n4978);
and (s0n5366,notn5366,n2800);
and (s1n5366,n4978,n2857);
nor (n5367,n5368,n5374);
nand (n5368,n5369,n5372);
or (n5369,n5370,n5049);
not (n5370,n5371);
wire s0n5371,s1n5371,notn5371;
or (n5371,s0n5371,s1n5371);
not(notn5371,n4978);
and (s0n5371,notn5371,n2789);
and (s1n5371,n4978,n2846);
nand (n5372,n5112,n5373);
wire s0n5373,s1n5373,notn5373;
or (n5373,s0n5373,s1n5373);
not(notn5373,n4978);
and (s0n5373,notn5373,n2755);
and (s1n5373,n4978,n2817);
nand (n5374,n5375,n5378);
or (n5375,n5376,n5030);
not (n5376,n5377);
wire s0n5377,s1n5377,notn5377;
or (n5377,s0n5377,s1n5377);
not(notn5377,n4978);
and (s0n5377,notn5377,n2771);
and (s1n5377,n4978,n2829);
nand (n5378,n5040,n5379);
wire s0n5379,s1n5379,notn5379;
or (n5379,s0n5379,s1n5379);
not(notn5379,n4978);
and (s0n5379,notn5379,n2803);
and (s1n5379,n4978,n2860);
nand (n5380,n5381,n5384);
or (n5381,n5382,n5076);
not (n5382,n5383);
wire s0n5383,s1n5383,notn5383;
or (n5383,s0n5383,s1n5383);
not(notn5383,n4978);
and (s0n5383,notn5383,n2783);
and (s1n5383,n4978,n2840);
nand (n5384,n5019,n5385);
wire s0n5385,s1n5385,notn5385;
or (n5385,s0n5385,s1n5385);
not(notn5385,n4978);
and (s0n5385,notn5385,n2763);
and (s1n5385,n4978,n2823);
nand (n5386,n5387,n5404,n5413);
nor (n5387,n5388,n5392);
nand (n5388,n5389,n5390,n5391);
nand (n5389,n5016,n5360);
nand (n5390,n5019,n5354);
nand (n5391,n5013,n5356);
nand (n5392,n5393,n5395);
or (n5393,n5394,n5026);
not (n5394,n5358);
nor (n5395,n5396,n5400);
nand (n5396,n5397,n5399);
or (n5397,n5398,n5049);
not (n5398,n5347);
nand (n5399,n5112,n5349);
nand (n5400,n5401,n5403);
or (n5401,n5402,n5039);
not (n5402,n5366);
nand (n5403,n5031,n5351);
nor (n5404,n5405,n5410);
nand (n5405,n5406,n5409);
or (n5406,n5407,n5408);
not (n5407,n5373);
not (n5408,n4995);
nand (n5409,n4948,n5364);
nand (n5410,n5411,n5412);
or (n5411,n5382,n4986);
nand (n5412,n4981,n5385);
nor (n5413,n5414,n5418);
nand (n5414,n5415,n5416);
or (n5415,n5370,n5144);
nand (n5416,n4998,n5417);
wire s0n5417,s1n5417,notn5417;
or (n5417,s0n5417,s1n5417);
not(notn5417,n4978);
and (s0n5417,notn5417,n2780);
and (s1n5417,n4978,n2837);
nand (n5418,n5419,n5421);
or (n5419,n5420,n5002);
not (n5420,n5345);
nand (n5421,n5008,n5422);
wire s0n5422,s1n5422,notn5422;
or (n5422,s0n5422,s1n5422);
not(notn5422,n4978);
and (s0n5422,notn5422,n2753);
and (s1n5422,n4978,n2815);
and (n5423,n5386,n5424);
or (n5424,n5425,n5501,n5677);
and (n5425,n5426,n5471);
nand (n5426,n5427,n5446);
nor (n5427,n5428,n5437);
nand (n5428,n5429,n5431,n5433,n5435);
nand (n5429,n4948,n5430);
wire s0n5430,s1n5430,notn5430;
or (n5430,s0n5430,s1n5430);
not(notn5430,n4978);
and (s0n5430,notn5430,n2879);
and (s1n5430,n4978,n2936);
nand (n5431,n4981,n5432);
wire s0n5432,s1n5432,notn5432;
or (n5432,s0n5432,s1n5432);
not(notn5432,n4978);
and (s0n5432,notn5432,n2891);
and (s1n5432,n4978,n2948);
nand (n5433,n4985,n5434);
wire s0n5434,s1n5434,notn5434;
or (n5434,s0n5434,s1n5434);
not(notn5434,n4978);
and (s0n5434,notn5434,n2903);
and (s1n5434,n4978,n2960);
nand (n5435,n4989,n5436);
wire s0n5436,s1n5436,notn5436;
or (n5436,s0n5436,s1n5436);
not(notn5436,n4978);
and (s0n5436,notn5436,n2911);
and (s1n5436,n4978,n2968);
nand (n5437,n5438,n5440,n5442,n5444);
nand (n5438,n4995,n5439);
wire s0n5439,s1n5439,notn5439;
or (n5439,s0n5439,s1n5439);
not(notn5439,n4978);
and (s0n5439,notn5439,n2887);
and (s1n5439,n4978,n2944);
nand (n5440,n5008,n5441);
wire s0n5441,s1n5441,notn5441;
or (n5441,s0n5441,s1n5441);
not(notn5441,n4978);
and (s0n5441,notn5441,n2875);
and (s1n5441,n4978,n2932);
nand (n5442,n4998,n5443);
wire s0n5443,s1n5443,notn5443;
or (n5443,s0n5443,s1n5443);
not(notn5443,n4978);
and (s0n5443,notn5443,n2896);
and (s1n5443,n4978,n2953);
nand (n5444,n5001,n5445);
wire s0n5445,s1n5445,notn5445;
or (n5445,s0n5445,s1n5445);
not(notn5445,n4978);
and (s0n5445,notn5445,n2914);
and (s1n5445,n4978,n2971);
nor (n5446,n5447,n5454);
nand (n5447,n5448,n5450,n5452);
nand (n5448,n5019,n5449);
wire s0n5449,s1n5449,notn5449;
or (n5449,s0n5449,s1n5449);
not(notn5449,n4978);
and (s0n5449,notn5449,n2889);
and (s1n5449,n4978,n2946);
nand (n5450,n5013,n5451);
wire s0n5451,s1n5451,notn5451;
or (n5451,s0n5451,s1n5451);
not(notn5451,n4978);
and (s0n5451,notn5451,n2900);
and (s1n5451,n4978,n2957);
nand (n5452,n5016,n5453);
wire s0n5453,s1n5453,notn5453;
or (n5453,s0n5453,s1n5453);
not(notn5453,n4978);
and (s0n5453,notn5453,n2877);
and (s1n5453,n4978,n2934);
nand (n5454,n5455,n5458);
or (n5455,n5456,n5026);
not (n5456,n5457);
wire s0n5457,s1n5457,notn5457;
or (n5457,s0n5457,s1n5457);
not(notn5457,n4978);
and (s0n5457,notn5457,n2917);
and (s1n5457,n4978,n2974);
nor (n5458,n5459,n5465);
nand (n5459,n5460,n5463);
or (n5460,n5461,n5030);
not (n5461,n5462);
wire s0n5462,s1n5462,notn5462;
or (n5462,s0n5462,s1n5462);
not(notn5462,n4978);
and (s0n5462,notn5462,n2885);
and (s1n5462,n4978,n2941);
nand (n5463,n5040,n5464);
wire s0n5464,s1n5464,notn5464;
or (n5464,s0n5464,s1n5464);
not(notn5464,n4978);
and (s0n5464,notn5464,n2920);
and (s1n5464,n4978,n2977);
nand (n5465,n5466,n5469);
or (n5466,n5467,n5049);
not (n5467,n5468);
wire s0n5468,s1n5468,notn5468;
or (n5468,s0n5468,s1n5468);
not(notn5468,n4978);
and (s0n5468,notn5468,n2906);
and (s1n5468,n4978,n2963);
nand (n5469,n5112,n5470);
wire s0n5470,s1n5470,notn5470;
or (n5470,s0n5470,s1n5470);
not(notn5470,n4978);
and (s0n5470,notn5470,n2873);
and (s1n5470,n4978,n2930);
nand (n5471,n5472,n5485);
nor (n5472,n5473,n5478);
nand (n5473,n5474,n5475,n5476,n5477);
nand (n5474,n4995,n5470);
nand (n5475,n4981,n5449);
nand (n5476,n4948,n5453);
nand (n5477,n4985,n5451);
nand (n5478,n5479,n5481,n5482,n5483);
nand (n5479,n4998,n5480);
wire s0n5480,s1n5480,notn5480;
or (n5480,s0n5480,s1n5480);
not(notn5480,n4978);
and (s0n5480,notn5480,n2897);
and (s1n5480,n4978,n2954);
nand (n5481,n5468,n4989);
nand (n5482,n5001,n5436);
nand (n5483,n5008,n5484);
wire s0n5484,s1n5484,notn5484;
or (n5484,s0n5484,s1n5484);
not(notn5484,n4978);
and (s0n5484,notn5484,n2871);
and (s1n5484,n4978,n2928);
nor (n5485,n5486,n5497);
nand (n5486,n5487,n5488,n5489);
nand (n5487,n5016,n5441);
nand (n5488,n5058,n5445);
nor (n5489,n5490,n5493);
nand (n5490,n5491,n5492);
or (n5491,n5456,n5039);
nand (n5492,n5031,n5432);
nand (n5493,n5494,n5496);
or (n5494,n5495,n5049);
not (n5495,n5434);
nand (n5496,n5112,n5430);
nand (n5497,n5498,n5500);
or (n5498,n5499,n5076);
not (n5499,n5443);
nand (n5500,n5019,n5439);
and (n5501,n5471,n5502);
nand (n5502,n5503,n5592);
or (n5503,n5504,n5557);
not (n5504,n5505);
nand (n5505,n5506,n5531,n5544);
nor (n5506,n5507,n5514);
nand (n5507,n5508,n5510,n5512);
nand (n5508,n5016,n5509);
wire s0n5509,s1n5509,notn5509;
or (n5509,s0n5509,s1n5509);
not(notn5509,n4978);
and (s0n5509,notn5509,n2988);
and (s1n5509,n4978,n3055);
nand (n5510,n5019,n5511);
wire s0n5511,s1n5511,notn5511;
or (n5511,s0n5511,s1n5511);
not(notn5511,n4978);
and (s0n5511,notn5511,n3009);
and (s1n5511,n4978,n3068);
nand (n5512,n5013,n5513);
wire s0n5513,s1n5513,notn5513;
or (n5513,s0n5513,s1n5513);
not(notn5513,n4978);
and (s0n5513,notn5513,n3016);
and (s1n5513,n4978,n3077);
nand (n5514,n5515,n5518);
or (n5515,n5516,n5026);
not (n5516,n5517);
wire s0n5517,s1n5517,notn5517;
or (n5517,s0n5517,s1n5517);
not(notn5517,n4978);
and (s0n5517,notn5517,n3034);
and (s1n5517,n4978,n3095);
nor (n5518,n5519,n5525);
nand (n5519,n5520,n5523);
or (n5520,n5521,n5049);
not (n5521,n5522);
wire s0n5522,s1n5522,notn5522;
or (n5522,s0n5522,s1n5522);
not(notn5522,n4978);
and (s0n5522,notn5522,n3023);
and (s1n5522,n4978,n3084);
nand (n5523,n5112,n5524);
wire s0n5524,s1n5524,notn5524;
or (n5524,s0n5524,s1n5524);
not(notn5524,n4978);
and (s0n5524,notn5524,n2995);
and (s1n5524,n4978,n3059);
nand (n5525,n5526,n5529);
or (n5526,n5527,n5039);
not (n5527,n5528);
wire s0n5528,s1n5528,notn5528;
or (n5528,s0n5528,s1n5528);
not(notn5528,n4978);
and (s0n5528,notn5528,n3037);
and (s1n5528,n4978,n3098);
nand (n5529,n5031,n5530);
wire s0n5530,s1n5530,notn5530;
or (n5530,s0n5530,s1n5530);
not(notn5530,n4978);
and (s0n5530,notn5530,n3003);
and (s1n5530,n4978,n3072);
nor (n5531,n5532,n5538);
nand (n5532,n5533,n5536);
or (n5533,n5534,n4986);
not (n5534,n5535);
wire s0n5535,s1n5535,notn5535;
or (n5535,s0n5535,s1n5535);
not(notn5535,n4978);
and (s0n5535,notn5535,n3020);
and (s1n5535,n4978,n3081);
nand (n5536,n4981,n5537);
wire s0n5537,s1n5537,notn5537;
or (n5537,s0n5537,s1n5537);
not(notn5537,n4978);
and (s0n5537,notn5537,n3005);
and (s1n5537,n4978,n3070);
nand (n5538,n5539,n5542);
or (n5539,n5540,n4949);
not (n5540,n5541);
wire s0n5541,s1n5541,notn5541;
or (n5541,s0n5541,s1n5541);
not(notn5541,n4978);
and (s0n5541,notn5541,n2992);
and (s1n5541,n4978,n3057);
nand (n5542,n4995,n5543);
wire s0n5543,s1n5543,notn5543;
or (n5543,s0n5543,s1n5543);
not(notn5543,n4978);
and (s0n5543,notn5543,n2998);
and (s1n5543,n4978,n3053);
nor (n5544,n5545,n5551);
nand (n5545,n5546,n5549);
or (n5546,n5547,n5085);
not (n5547,n5548);
wire s0n5548,s1n5548,notn5548;
or (n5548,s0n5548,s1n5548);
not(notn5548,n4978);
and (s0n5548,notn5548,n2989);
and (s1n5548,n4978,n3051);
nand (n5549,n4998,n5550);
wire s0n5550,s1n5550,notn5550;
or (n5550,s0n5550,s1n5550);
not(notn5550,n4978);
and (s0n5550,notn5550,n3017);
and (s1n5550,n4978,n3078);
nand (n5551,n5552,n5555);
or (n5552,n5553,n5144);
not (n5553,n5554);
wire s0n5554,s1n5554,notn5554;
or (n5554,s0n5554,s1n5554);
not(notn5554,n4978);
and (s0n5554,notn5554,n3026);
and (s1n5554,n4978,n3087);
nand (n5555,n5001,n5556);
wire s0n5556,s1n5556,notn5556;
or (n5556,s0n5556,s1n5556);
not(notn5556,n4978);
and (s0n5556,notn5556,n3031);
and (s1n5556,n4978,n3092);
not (n5557,n5558);
nand (n5558,n5559,n5576,n5584);
nor (n5559,n5560,n5573);
nand (n5560,n5561,n5562,n5563);
nand (n5561,n5058,n5528);
nand (n5562,n5016,n5541);
nor (n5563,n5564,n5570);
nand (n5564,n5565,n5568);
or (n5565,n5566,n5030);
not (n5566,n5567);
wire s0n5567,s1n5567,notn5567;
or (n5567,s0n5567,s1n5567);
not(notn5567,n4978);
and (s0n5567,notn5567,n3011);
and (s1n5567,n4978,n3066);
nand (n5568,n5040,n5569);
wire s0n5569,s1n5569,notn5569;
or (n5569,s0n5569,s1n5569);
not(notn5569,n4978);
and (s0n5569,notn5569,n3040);
and (s1n5569,n4978,n3101);
nand (n5570,n5571,n5572);
or (n5571,n5553,n5049);
nand (n5572,n5112,n5543);
nand (n5573,n5574,n5575);
or (n5574,n5534,n5076);
nand (n5575,n5019,n5537);
nor (n5576,n5577,n5581);
nand (n5577,n5578,n5580);
or (n5578,n5579,n4949);
not (n5579,n5524);
nand (n5580,n4981,n5530);
nand (n5581,n5582,n5583);
or (n5582,n5521,n4986);
nand (n5583,n4989,n5556);
nor (n5584,n5585,n5589);
nand (n5585,n5586,n5588);
or (n5586,n5587,n5085);
not (n5587,n5509);
nand (n5588,n4995,n5511);
nand (n5589,n5590,n5591);
or (n5590,n5516,n5002);
nand (n5591,n4998,n5513);
or (n5592,n5593,n5676);
not (n5593,n5594);
and (n5594,n5595,n5646);
nand (n5595,n5596,n5620,n5633);
nor (n5596,n5597,n5604);
nand (n5597,n5598,n5600,n5602);
nand (n5598,n5016,n5599);
wire s0n5599,s1n5599,notn5599;
or (n5599,s0n5599,s1n5599);
not(notn5599,n4978);
and (s0n5599,notn5599,n3119);
and (s1n5599,n4978,n3176);
nand (n5600,n5013,n5601);
wire s0n5601,s1n5601,notn5601;
or (n5601,s0n5601,s1n5601);
not(notn5601,n4978);
and (s0n5601,notn5601,n3139);
and (s1n5601,n4978,n3202);
nand (n5602,n5019,n5603);
wire s0n5603,s1n5603,notn5603;
or (n5603,s0n5603,s1n5603);
not(notn5603,n4978);
and (s0n5603,notn5603,n3132);
and (s1n5603,n4978,n3192);
nand (n5604,n5605,n5608);
or (n5605,n5606,n5026);
not (n5606,n5607);
wire s0n5607,s1n5607,notn5607;
or (n5607,s0n5607,s1n5607);
not(notn5607,n4978);
and (s0n5607,notn5607,n3157);
and (s1n5607,n4978,n3220);
nor (n5608,n5609,n5614);
nand (n5609,n5610,n5612);
nand (n5610,n5050,n5611);
wire s0n5611,s1n5611,notn5611;
or (n5611,s0n5611,s1n5611);
not(notn5611,n4978);
and (s0n5611,notn5611,n3146);
and (s1n5611,n4978,n3209);
nand (n5612,n5112,n5613);
wire s0n5613,s1n5613,notn5613;
or (n5613,s0n5613,s1n5613);
not(notn5613,n4978);
and (s0n5613,notn5613,n3112);
and (s1n5613,n4978,n3173);
nand (n5614,n5615,n5618);
or (n5615,n5616,n5039);
not (n5616,n5617);
wire s0n5617,s1n5617,notn5617;
or (n5617,s0n5617,s1n5617);
not(notn5617,n4978);
and (s0n5617,notn5617,n3160);
and (s1n5617,n4978,n3223);
nand (n5618,n5031,n5619);
wire s0n5619,s1n5619,notn5619;
or (n5619,s0n5619,s1n5619);
not(notn5619,n4978);
and (s0n5619,notn5619,n3128);
and (s1n5619,n4978,n3189);
nor (n5620,n5621,n5627);
nand (n5621,n5622,n5625);
or (n5622,n5623,n4986);
not (n5623,n5624);
wire s0n5624,s1n5624,notn5624;
or (n5624,s0n5624,s1n5624);
not(notn5624,n4978);
and (s0n5624,notn5624,n3143);
and (s1n5624,n4978,n3206);
nand (n5625,n4981,n5626);
wire s0n5626,s1n5626,notn5626;
or (n5626,s0n5626,s1n5626);
not(notn5626,n4978);
and (s0n5626,notn5626,n3126);
and (s1n5626,n4978,n3187);
nand (n5627,n5628,n5631);
or (n5628,n5629,n5408);
not (n5629,n5630);
wire s0n5630,s1n5630,notn5630;
or (n5630,s0n5630,s1n5630);
not(notn5630,n4978);
and (s0n5630,notn5630,n3121);
and (s1n5630,n4978,n3182);
nand (n5631,n4948,n5632);
wire s0n5632,s1n5632,notn5632;
or (n5632,s0n5632,s1n5632);
not(notn5632,n4978);
and (s0n5632,notn5632,n3114);
and (s1n5632,n4978,n3171);
nor (n5633,n5634,n5640);
nand (n5634,n5635,n5638);
or (n5635,n5636,n5091);
not (n5636,n5637);
wire s0n5637,s1n5637,notn5637;
or (n5637,s0n5637,s1n5637);
not(notn5637,n4978);
and (s0n5637,notn5637,n3140);
and (s1n5637,n4978,n3203);
nand (n5638,n4989,n5639);
wire s0n5639,s1n5639,notn5639;
or (n5639,s0n5639,s1n5639);
not(notn5639,n4978);
and (s0n5639,notn5639,n3149);
and (s1n5639,n4978,n3212);
nand (n5640,n5641,n5644);
or (n5641,n5642,n5002);
not (n5642,n5643);
wire s0n5643,s1n5643,notn5643;
or (n5643,s0n5643,s1n5643);
not(notn5643,n4978);
and (s0n5643,notn5643,n3154);
and (s1n5643,n4978,n3217);
nand (n5644,n5008,n5645);
wire s0n5645,s1n5645,notn5645;
or (n5645,s0n5645,s1n5645);
not(notn5645,n4978);
and (s0n5645,notn5645,n3117);
and (s1n5645,n4978,n3180);
nand (n5646,n5647,n5658);
nor (n5647,n5648,n5653);
nand (n5648,n5649,n5650,n5651,n5652);
nand (n5649,n4981,n5619);
nand (n5650,n4985,n5611);
nand (n5651,n4948,n5613);
nand (n5652,n5008,n5599);
nand (n5653,n5654,n5655,n5656,n5657);
nand (n5654,n4989,n5643);
nand (n5655,n5001,n5607);
nand (n5656,n4995,n5603);
nand (n5657,n4998,n5601);
nor (n5658,n5659,n5663);
nand (n5659,n5660,n5661,n5662);
nand (n5660,n5013,n5624);
nand (n5661,n5016,n5632);
nand (n5662,n5019,n5626);
nand (n5663,n5664,n5665);
or (n5664,n5616,n5026);
nor (n5665,n5666,n5672);
nand (n5666,n5667,n5670);
or (n5667,n5668,n5030);
not (n5668,n5669);
wire s0n5669,s1n5669,notn5669;
or (n5669,s0n5669,s1n5669);
not(notn5669,n4978);
and (s0n5669,notn5669,n3134);
and (s1n5669,n4978,n3197);
nand (n5670,n5040,n5671);
wire s0n5671,s1n5671,notn5671;
or (n5671,s0n5671,s1n5671);
not(notn5671,n4978);
and (s0n5671,notn5671,n3163);
and (s1n5671,n4978,n3226);
nand (n5672,n5673,n5675);
or (n5673,n5674,n5049);
not (n5674,n5639);
nand (n5675,n5112,n5630);
and (n5676,n5504,n5557);
and (n5677,n5426,n5502);
and (n5678,n5341,n5424);
and (n5679,n5264,n5339);
and (n5680,n5230,n5262);
and (n5681,n5153,n5183);
and (n5682,n5054,n5097);
or (n5683,n5684,n5688);
xor (n5684,n5685,n5097);
not (n5685,n5686);
nand (n5686,n4942,n5687);
or (n5687,n5054,n4944);
or (n5688,n5689,n6310,n6393);
and (n5689,n5690,n5692);
xor (n5690,n5691,n5183);
xor (n5691,n5099,n5153);
nand (n5692,n5693,n6309);
or (n5693,n5694,n5770);
not (n5694,n5695);
nand (n5695,n5696,n5735);
nand (n5696,n5697,n5714,n5722);
nor (n5697,n5698,n5708);
and (n5698,n5699,n1265);
not (n5699,n5700);
nor (n5700,n5701,n5705);
nand (n5701,n5702,n5704);
or (n5702,n5075,n5703);
not (n5703,n4990);
nand (n5704,n4950,n4992);
nand (n5705,n5706,n5707);
or (n5706,n5051,n5004);
nand (n5707,n5032,n5006);
and (n5708,n5709,n1331);
nand (n5709,n5710,n5711,n5712,n5713);
nand (n5710,n5003,n5047);
nand (n5711,n4990,n4977);
nand (n5712,n4950,n4996);
nand (n5713,n5032,n5021);
nor (n5714,n5715,n5719);
nand (n5715,n5716,n5718);
or (n5716,n5717,n5408);
not (n5717,n4983);
nand (n5718,n5019,n5037);
nand (n5719,n5720,n5721);
or (n5720,n5024,n5144);
nand (n5721,n5058,n5072);
nor (n5722,n5723,n5734);
nand (n5723,n5724,n5725);
or (n5724,n5068,n4982);
nor (n5725,n5726,n5730);
and (n5726,n5031,n5727);
wire s0n5727,s1n5727,notn5727;
or (n5727,s0n5727,s1n5727);
not(notn5727,n4978);
and (s0n5727,notn5727,n5728);
and (s1n5727,n4978,n5729);
and (n5730,n5040,n5731);
wire s0n5731,s1n5731,notn5731;
or (n5731,s0n5731,s1n5731);
not(notn5731,n4978);
and (s0n5731,notn5731,n5732);
and (s1n5731,n4978,n5733);
and (n5734,n5001,n5042);
nand (n5735,n5736,n5754);
nor (n5736,n5737,n5748);
nand (n5737,n5738,n5742,n5746,n5747);
nand (n5738,n4998,n5739);
wire s0n5739,s1n5739,notn5739;
or (n5739,s0n5739,s1n5739);
not(notn5739,n4978);
and (s0n5739,notn5739,n5740);
and (s1n5739,n4978,n5741);
nand (n5742,n5008,n5743);
wire s0n5743,s1n5743,notn5743;
or (n5743,s0n5743,s1n5743);
not(notn5743,n4978);
and (s0n5743,notn5743,n5744);
and (s1n5743,n4978,n5745);
nand (n5746,n4985,n5014);
nand (n5747,n5016,n5009);
nand (n5748,n5749,n5750,n5751);
nand (n5749,n5013,n4999);
nand (n5750,n4948,n5017);
nor (n5751,n5752,n5753);
and (n5752,n5112,n4977);
and (n5753,n5050,n4987);
nor (n5754,n5755,n5764);
and (n5755,n5756,n1246);
nand (n5756,n5757,n5761);
not (n5757,n5758);
nand (n5758,n5759,n5760);
or (n5759,n5051,n5703);
nand (n5760,n4950,n5006);
nor (n5761,n5762,n5763);
and (n5762,n5032,n5025);
and (n5763,n5003,n4992);
and (n5764,n5765,n1316);
nand (n5765,n5766,n5767,n5768,n5769);
nand (n5766,n4990,n5047);
nand (n5767,n5003,n4996);
nand (n5768,n4950,n5021);
nand (n5769,n5032,n4983);
nand (n5770,n5771,n6308);
or (n5771,n5772,n5844);
not (n5772,n5773);
or (n5773,n5774,n5810);
nand (n5774,n5775,n5794);
nor (n5775,n5776,n5787);
nand (n5776,n5777,n5781,n5782,n5783);
nand (n5777,n4998,n5778);
wire s0n5778,s1n5778,notn5778;
or (n5778,s0n5778,s1n5778);
not(notn5778,n4978);
and (s0n5778,notn5778,n5779);
and (s1n5778,n4978,n5780);
nand (n5781,n4985,n5123);
nand (n5782,n5016,n5152);
nand (n5783,n5008,n5784);
wire s0n5784,s1n5784,notn5784;
or (n5784,s0n5784,s1n5784);
not(notn5784,n4978);
and (s0n5784,notn5784,n5785);
and (s1n5784,n4978,n5786);
nand (n5787,n5788,n5792,n5793);
not (n5788,n5789);
nand (n5789,n5790,n5791);
or (n5790,n5129,n5049);
nand (n5791,n5112,n5136);
nand (n5792,n5013,n5146);
nand (n5793,n4948,n5105);
nor (n5794,n5795,n5804);
and (n5795,n5796,n1246);
nand (n5796,n5797,n5801);
not (n5797,n5798);
nand (n5798,n5799,n5800);
or (n5799,n5109,n5703);
nand (n5800,n4950,n5150);
nor (n5801,n5802,n5803);
and (n5802,n5032,n5103);
and (n5803,n5003,n5143);
and (n5804,n5805,n1316);
nand (n5805,n5806,n5807,n5808,n5809);
nand (n5806,n5003,n5138);
nand (n5807,n4990,n5113);
nand (n5808,n4950,n5125);
nand (n5809,n5032,n5132);
nand (n5810,n5811,n5831);
nor (n5811,n5812,n5817);
nand (n5812,n5813,n5814,n5815,n5816);
nand (n5813,n5058,n5178);
nand (n5814,n4989,n5103);
nand (n5815,n4995,n5132);
nand (n5816,n5019,n5119);
nand (n5817,n5818,n5829,n5830);
not (n5818,n5819);
nand (n5819,n5820,n5825);
or (n5820,n5821,n5030);
not (n5821,n5822);
wire s0n5822,s1n5822,notn5822;
or (n5822,s0n5822,s1n5822);
not(notn5822,n4978);
and (s0n5822,notn5822,n5823);
and (s1n5822,n4978,n5824);
nand (n5825,n5040,n5826);
wire s0n5826,s1n5826,notn5826;
or (n5826,s0n5826,s1n5826);
not(notn5826,n4978);
and (s0n5826,notn5826,n5827);
and (s1n5826,n4978,n5828);
nand (n5829,n4981,n5176);
nand (n5830,n5001,n5117);
nor (n5831,n5832,n5838);
and (n5832,n5833,n1331);
nand (n5833,n5834,n5835,n5836,n5837);
nand (n5834,n5003,n5113);
nand (n5835,n4990,n5136);
nand (n5836,n4950,n5138);
nand (n5837,n5032,n5125);
and (n5838,n5839,n1265);
nand (n5839,n5840,n5841,n5842,n5843);
nand (n5840,n5003,n5110);
nand (n5841,n4990,n5130);
nand (n5842,n4950,n5143);
nand (n5843,n5032,n5150);
not (n5844,n5845);
nand (n5845,n5846,n6301);
or (n5846,n5847,n5993);
not (n5847,n5848);
nor (n5848,n5849,n5918);
nor (n5849,n5850,n5884);
nand (n5850,n5851,n5869);
nor (n5851,n5852,n5863);
nand (n5852,n5853,n5854,n5858,n5859);
nand (n5853,n4948,n5210);
nand (n5854,n5008,n5855);
wire s0n5855,s1n5855,notn5855;
or (n5855,s0n5855,s1n5855);
not(notn5855,n4978);
and (s0n5855,notn5855,n5856);
and (s1n5855,n4978,n5857);
nand (n5858,n5013,n5202);
nand (n5859,n4998,n5860);
wire s0n5860,s1n5860,notn5860;
or (n5860,s0n5860,s1n5860);
not(notn5860,n4978);
and (s0n5860,notn5860,n5861);
and (s1n5860,n4978,n5862);
nand (n5863,n5864,n5865,n5866);
nand (n5864,n4985,n5227);
nand (n5865,n5016,n5204);
nor (n5866,n5867,n5868);
and (n5867,n5050,n5189);
and (n5868,n5112,n5191);
nor (n5869,n5870,n5878);
and (n5870,n5871,n1246);
nand (n5871,n5872,n5875);
nor (n5872,n5873,n5874);
and (n5873,n4990,n5217);
and (n5874,n4950,n5200);
nor (n5875,n5876,n5877);
and (n5876,n5032,n5208);
and (n5877,n5003,n5193);
and (n5878,n5879,n1316);
nand (n5879,n5880,n5881,n5882,n5883);
nand (n5880,n5003,n5198);
nand (n5881,n4990,n5215);
nand (n5882,n4950,n5229);
nand (n5883,n5032,n5195);
nand (n5884,n5885,n5903);
nor (n5885,n5886,n5899);
nand (n5886,n5887,n5888,n5889,n5890);
nand (n5887,n4981,n5254);
nand (n5888,n5001,n5221);
nand (n5889,n5019,n5223);
nor (n5890,n5891,n5895);
and (n5891,n5040,n5892);
wire s0n5892,s1n5892,notn5892;
or (n5892,s0n5892,s1n5892);
not(notn5892,n4978);
and (s0n5892,notn5892,n5893);
and (s1n5892,n4978,n5894);
and (n5895,n5031,n5896);
wire s0n5896,s1n5896,notn5896;
or (n5896,s0n5896,s1n5896);
not(notn5896,n4978);
and (s0n5896,notn5896,n5897);
and (s1n5896,n4978,n5898);
nand (n5899,n5900,n5901,n5902);
nand (n5900,n4995,n5195);
nand (n5901,n4989,n5208);
nand (n5902,n5058,n5256);
nor (n5903,n5904,n5912);
and (n5904,n5905,n1331);
nand (n5905,n5906,n5909);
nor (n5906,n5907,n5908);
and (n5907,n4990,n5191);
and (n5908,n4950,n5198);
nor (n5909,n5910,n5911);
and (n5910,n5032,n5229);
and (n5911,n5003,n5215);
and (n5912,n5913,n1265);
nand (n5913,n5914,n5915,n5916,n5917);
nand (n5914,n4950,n5193);
nand (n5915,n4990,n5189);
nand (n5916,n5003,n5217);
nand (n5917,n5032,n5200);
nor (n5918,n5919,n5957);
nand (n5919,n5920,n5942);
nor (n5920,n5921,n5932);
nand (n5921,n5922,n5929);
not (n5922,n5923);
nand (n5923,n5924,n5926);
or (n5924,n5925,n5076);
not (n5925,n5321);
nor (n5926,n5927,n5928);
and (n5927,n5112,n5291);
and (n5928,n5050,n5289);
nor (n5929,n5930,n5931);
and (n5930,n5016,n5319);
and (n5931,n4948,n5283);
nand (n5932,n5933,n5937,n5938);
nand (n5933,n4998,n5934);
wire s0n5934,s1n5934,notn5934;
or (n5934,s0n5934,s1n5934);
not(notn5934,n4978);
and (s0n5934,notn5934,n5935);
and (s1n5934,n4978,n5936);
nand (n5937,n4985,n5281);
nand (n5938,n5008,n5939);
wire s0n5939,s1n5939,notn5939;
or (n5939,s0n5939,s1n5939);
not(notn5939,n4978);
and (s0n5939,notn5939,n5940);
and (s1n5939,n4978,n5941);
nor (n5942,n5943,n5951);
and (n5943,n5944,n1246);
nand (n5944,n5945,n5948);
nor (n5945,n5946,n5947);
and (n5946,n4950,n5279);
and (n5947,n4990,n5270);
nor (n5948,n5949,n5950);
and (n5949,n5032,n5277);
and (n5950,n5003,n5300);
and (n5951,n5952,n1316);
nand (n5952,n5953,n5954,n5955,n5956);
nand (n5953,n4950,n5268);
nand (n5954,n4990,n5272);
nand (n5955,n5003,n5302);
nand (n5956,n5032,n5287);
nand (n5957,n5958,n5975);
nor (n5958,n5959,n5967);
and (n5959,n5960,n1331);
nand (n5960,n5961,n5964);
nor (n5961,n5962,n5963);
and (n5962,n4950,n5302);
and (n5963,n4990,n5291);
nor (n5964,n5965,n5966);
and (n5965,n5032,n5268);
and (n5966,n5003,n5272);
and (n5967,n5968,n1265);
nand (n5968,n5969,n5972);
nor (n5969,n5970,n5971);
and (n5970,n4950,n5300);
and (n5971,n4990,n5289);
nor (n5972,n5973,n5974);
and (n5973,n5032,n5279);
and (n5974,n5003,n5270);
nor (n5975,n5976,n5989);
nand (n5976,n5977,n5978,n5979,n5980);
nand (n5977,n5001,n5295);
nand (n5978,n5019,n5274);
nand (n5979,n5058,n5307);
nor (n5980,n5981,n5985);
and (n5981,n5040,n5982);
wire s0n5982,s1n5982,notn5982;
or (n5982,s0n5982,s1n5982);
not(notn5982,n4978);
and (s0n5982,notn5982,n5983);
and (s1n5982,n4978,n5984);
and (n5985,n5031,n5986);
wire s0n5986,s1n5986,notn5986;
or (n5986,s0n5986,s1n5986);
not(notn5986,n4978);
and (s0n5986,notn5986,n5987);
and (s1n5986,n4978,n5988);
nand (n5989,n5990,n5991,n5992);
nand (n5990,n4989,n5277);
nand (n5991,n4995,n5287);
nand (n5992,n4981,n5305);
not (n5993,n5994);
nand (n5994,n5995,n6294);
or (n5995,n5996,n6146);
not (n5996,n5997);
nor (n5997,n5998,n6068);
nor (n5998,n5999,n6033);
nand (n5999,n6000,n6015);
nor (n6000,n6001,n6009);
and (n6001,n6002,n1246);
nand (n6002,n6003,n6006);
nor (n6003,n6004,n6005);
and (n6004,n4990,n5347);
and (n6005,n4950,n5345);
nor (n6006,n6007,n6008);
and (n6007,n5032,n5358);
and (n6008,n5003,n5371);
and (n6009,n6010,n1316);
nand (n6010,n6011,n6012,n6013,n6014);
nand (n6011,n5003,n5373);
nand (n6012,n4990,n5349);
nand (n6013,n4950,n5354);
nand (n6014,n5032,n5385);
nor (n6015,n6016,n6026);
nand (n6016,n6017,n6021,n6025);
nand (n6017,n4998,n6018);
wire s0n6018,s1n6018,notn6018;
or (n6018,s0n6018,s1n6018);
not(notn6018,n4978);
and (s0n6018,notn6018,n6019);
and (s1n6018,n4978,n6020);
nand (n6021,n5008,n6022);
wire s0n6022,s1n6022,notn6022;
or (n6022,s0n6022,s1n6022);
not(notn6022,n4978);
and (s0n6022,notn6022,n6023);
and (s1n6022,n4978,n6024);
nand (n6025,n4985,n5356);
nand (n6026,n6027,n6028,n6029,n6030);
nand (n6027,n4948,n5360);
nand (n6028,n5016,n5422);
nand (n6029,n5013,n5417);
nor (n6030,n6031,n6032);
and (n6031,n5112,n5364);
and (n6032,n5050,n5383);
nand (n6033,n6034,n6050);
not (n6034,n6035);
nand (n6035,n6036,n6044);
or (n6036,n6037,n6038);
not (n6037,n1265);
not (n6038,n6039);
nand (n6039,n6040,n6041,n6042,n6043);
nand (n6040,n4990,n5383);
nand (n6041,n5003,n5347);
nand (n6042,n4950,n5371);
nand (n6043,n5032,n5345);
nand (n6044,n6045,n1331);
nand (n6045,n6046,n6047,n6048,n6049);
nand (n6046,n4990,n5364);
nand (n6047,n5003,n5349);
nand (n6048,n4950,n5373);
nand (n6049,n5032,n5354);
nor (n6050,n6051,n6055);
nand (n6051,n6052,n6053,n6054);
nand (n6052,n4995,n5385);
nand (n6053,n5058,n5379);
nand (n6054,n4989,n5358);
nand (n6055,n6056,n6057,n6058,n6059);
nand (n6056,n5019,n5351);
nand (n6057,n4981,n5377);
nand (n6058,n5001,n5366);
nor (n6059,n6060,n6064);
and (n6060,n5040,n6061);
wire s0n6061,s1n6061,notn6061;
or (n6061,s0n6061,s1n6061);
not(notn6061,n4978);
and (s0n6061,notn6061,n6062);
and (s1n6061,n4978,n6063);
and (n6064,n5031,n6065);
wire s0n6065,s1n6065,notn6065;
or (n6065,s0n6065,s1n6065);
not(notn6065,n4978);
and (s0n6065,notn6065,n6066);
and (s1n6065,n4978,n6067);
nor (n6068,n6069,n6108);
nand (n6069,n6070,n6090);
nor (n6070,n6071,n6082);
and (n6071,n6072,n1331);
not (n6072,n6073);
nor (n6073,n6074,n6078);
nand (n6074,n6075,n6077);
or (n6075,n6076,n4951);
not (n6076,n5470);
nand (n6077,n4990,n5453);
nand (n6078,n6079,n6081);
or (n6079,n6080,n5004);
not (n6080,n5430);
nand (n6081,n5032,n5439);
and (n6082,n6083,n1265);
nand (n6083,n6084,n6087);
nor (n6084,n6085,n6086);
and (n6085,n4950,n5468);
and (n6086,n4990,n5451);
nor (n6087,n6088,n6089);
and (n6088,n5032,n5436);
and (n6089,n5003,n5434);
nor (n6090,n6091,n6104);
nand (n6091,n6092,n6093,n6094,n6095);
nand (n6092,n4981,n5462);
nand (n6093,n5001,n5457);
nand (n6094,n5019,n5432);
nor (n6095,n6096,n6100);
and (n6096,n5031,n6097);
wire s0n6097,s1n6097,notn6097;
or (n6097,s0n6097,s1n6097);
not(notn6097,n4978);
and (s0n6097,notn6097,n6098);
and (s1n6097,n4978,n6099);
and (n6100,n5040,n6101);
wire s0n6101,s1n6101,notn6101;
or (n6101,s0n6101,s1n6101);
not(notn6101,n4978);
and (s0n6101,notn6101,n6102);
and (s1n6101,n4978,n6103);
nand (n6104,n6105,n6106,n6107);
nand (n6105,n5058,n5464);
nand (n6106,n4989,n5445);
nand (n6107,n4995,n5449);
nand (n6108,n6109,n6128);
nor (n6109,n6110,n6120);
and (n6110,n6111,n1246);
not (n6111,n6112);
nor (n6112,n6113,n6117);
nand (n6113,n6114,n6116);
or (n6114,n6115,n4951);
not (n6115,n5436);
nand (n6116,n4990,n5434);
nand (n6117,n6118,n6119);
or (n6118,n5467,n5004);
nand (n6119,n5032,n5445);
and (n6120,n6121,n1316);
nand (n6121,n6122,n6125);
nor (n6122,n6123,n6124);
and (n6123,n4950,n5439);
and (n6124,n4990,n5430);
nor (n6125,n6126,n6127);
and (n6126,n5032,n5449);
and (n6127,n5003,n5470);
nor (n6128,n6129,n6136);
nand (n6129,n6130,n6131,n6132,n6133);
nand (n6130,n4985,n5443);
nand (n6131,n5013,n5480);
nand (n6132,n5016,n5484);
nor (n6133,n6134,n6135);
and (n6134,n5112,n5453);
and (n6135,n5050,n5451);
nand (n6136,n6137,n6138,n6142);
nand (n6137,n4948,n5441);
nand (n6138,n5008,n6139);
wire s0n6139,s1n6139,notn6139;
or (n6139,s0n6139,s1n6139);
not(notn6139,n4978);
and (s0n6139,notn6139,n6140);
and (s1n6139,n4978,n6141);
nand (n6142,n4998,n6143);
wire s0n6143,s1n6143,notn6143;
or (n6143,s0n6143,s1n6143);
not(notn6143,n4978);
and (s0n6143,notn6143,n6144);
and (s1n6143,n4978,n6145);
not (n6146,n6147);
nand (n6147,n6148,n6293);
or (n6148,n6149,n6221);
nor (n6149,n6150,n6186);
nand (n6150,n6151,n6159,n6174,n6180);
nor (n6151,n6152,n6157);
nand (n6152,n6153,n6154);
or (n6153,n5587,n4949);
nor (n6154,n6155,n6156);
and (n6155,n5112,n5541);
and (n6156,n5050,n5535);
nor (n6157,n6158,n5547);
not (n6158,n5016);
nor (n6159,n6160,n6167);
nand (n6160,n6161,n6163);
or (n6161,n6162,n4986);
not (n6162,n5513);
nand (n6163,n4998,n6164);
wire s0n6164,s1n6164,notn6164;
or (n6164,s0n6164,s1n6164);
not(notn6164,n4978);
and (s0n6164,notn6164,n6165);
and (s1n6164,n4978,n6166);
nand (n6167,n6168,n6173);
or (n6168,n6169,n5085);
not (n6169,n6170);
wire s0n6170,s1n6170,notn6170;
or (n6170,s0n6170,s1n6170);
not(notn6170,n4978);
and (s0n6170,notn6170,n6171);
and (s1n6170,n4978,n6172);
nand (n6173,n5013,n5550);
nand (n6174,n6175,n1316);
nand (n6175,n6176,n6177,n6178,n6179);
nand (n6176,n5003,n5543);
nand (n6177,n4990,n5524);
nand (n6178,n4950,n5511);
nand (n6179,n5032,n5537);
nand (n6180,n6181,n1246);
nand (n6181,n6182,n6183,n6184,n6185);
nand (n6182,n5003,n5554);
nand (n6183,n4990,n5522);
nand (n6184,n4950,n5556);
nand (n6185,n5032,n5517);
nand (n6186,n6187,n6195,n6209,n6215);
nor (n6187,n6188,n6191);
nand (n6188,n6189,n6190);
or (n6189,n5516,n5144);
nand (n6190,n5058,n5569);
nand (n6191,n6192,n6194);
or (n6192,n6193,n5408);
not (n6193,n5537);
nand (n6194,n5001,n5528);
nor (n6195,n6196,n6207);
nand (n6196,n6197,n6198);
or (n6197,n5566,n4982);
nor (n6198,n6199,n6203);
and (n6199,n5040,n6200);
wire s0n6200,s1n6200,notn6200;
or (n6200,s0n6200,s1n6200);
not(notn6200,n4978);
and (s0n6200,notn6200,n6201);
and (s1n6200,n4978,n6202);
and (n6203,n5031,n6204);
wire s0n6204,s1n6204,notn6204;
or (n6204,s0n6204,s1n6204);
not(notn6204,n4978);
and (s0n6204,notn6204,n6205);
and (s1n6204,n4978,n6206);
nor (n6207,n6208,n5020);
not (n6208,n5530);
nand (n6209,n6210,n1265);
nand (n6210,n6211,n6212,n6213,n6214);
nand (n6211,n5003,n5522);
nand (n6212,n4990,n5535);
nand (n6213,n4950,n5554);
nand (n6214,n5032,n5556);
nand (n6215,n6216,n1331);
nand (n6216,n6217,n6218,n6219,n6220);
nand (n6217,n5003,n5524);
nand (n6218,n4990,n5541);
nand (n6219,n4950,n5543);
nand (n6220,n5032,n5511);
nand (n6221,n6222,n6258);
nand (n6222,n6223,n6231,n6246,n6252);
nor (n6223,n6224,n6225);
and (n6224,n5016,n5645);
nand (n6225,n6226,n6228);
or (n6226,n6227,n4949);
not (n6227,n5599);
nor (n6228,n6229,n6230);
and (n6229,n5112,n5632);
and (n6230,n5050,n5624);
nor (n6231,n6232,n6239);
nand (n6232,n6233,n6235);
or (n6233,n6234,n4986);
not (n6234,n5601);
nand (n6235,n4998,n6236);
wire s0n6236,s1n6236,notn6236;
or (n6236,s0n6236,s1n6236);
not(notn6236,n4978);
and (s0n6236,notn6236,n6237);
and (s1n6236,n4978,n6238);
nand (n6239,n6240,n6245);
or (n6240,n6241,n5085);
not (n6241,n6242);
wire s0n6242,s1n6242,notn6242;
or (n6242,s0n6242,s1n6242);
not(notn6242,n4978);
and (s0n6242,notn6242,n6243);
and (s1n6242,n4978,n6244);
nand (n6245,n5013,n5637);
nand (n6246,n6247,n1316);
nand (n6247,n6248,n6249,n6250,n6251);
nand (n6248,n5003,n5630);
nand (n6249,n4990,n5613);
nand (n6250,n4950,n5603);
nand (n6251,n5032,n5626);
nand (n6252,n6253,n1246);
nand (n6253,n6254,n6255,n6256,n6257);
nand (n6254,n5003,n5639);
nand (n6255,n4990,n5611);
nand (n6256,n4950,n5643);
nand (n6257,n5032,n5607);
nand (n6258,n6259,n6266,n6281,n6287);
nor (n6259,n6260,n6263);
nand (n6260,n6261,n6262);
or (n6261,n5668,n4982);
nand (n6262,n4995,n5626);
nand (n6263,n6264,n6265);
or (n6264,n5606,n5144);
nand (n6265,n5001,n5617);
nor (n6266,n6267,n6279);
nand (n6267,n6268,n6270);
or (n6268,n6269,n5026);
not (n6269,n5671);
nor (n6270,n6271,n6275);
and (n6271,n5040,n6272);
wire s0n6272,s1n6272,notn6272;
or (n6272,s0n6272,s1n6272);
not(notn6272,n4978);
and (s0n6272,notn6272,n6273);
and (s1n6272,n4978,n6274);
and (n6275,n5031,n6276);
wire s0n6276,s1n6276,notn6276;
or (n6276,s0n6276,s1n6276);
not(notn6276,n4978);
and (s0n6276,notn6276,n6277);
and (s1n6276,n4978,n6278);
nor (n6279,n5020,n6280);
not (n6280,n5619);
nand (n6281,n6282,n1265);
nand (n6282,n6283,n6284,n6285,n6286);
nand (n6283,n5003,n5611);
nand (n6284,n4990,n5624);
nand (n6285,n4950,n5639);
nand (n6286,n5032,n5643);
nand (n6287,n6288,n1331);
nand (n6288,n6289,n6290,n6291,n6292);
nand (n6289,n5003,n5613);
nand (n6290,n4990,n5632);
nand (n6291,n4950,n5630);
nand (n6292,n5032,n5603);
nand (n6293,n6150,n6186);
nor (n6294,n6295,n6299);
and (n6295,n6296,n6297);
not (n6296,n5998);
not (n6297,n6298);
nand (n6298,n6069,n6108);
not (n6299,n6300);
nand (n6300,n5999,n6033);
nand (n6301,n6302,n6307);
or (n6302,n6303,n6305);
not (n6303,n6304);
nand (n6304,n5884,n5850);
not (n6305,n6306);
nand (n6306,n5957,n5919);
not (n6307,n5849);
nand (n6308,n5810,n5774);
or (n6309,n5696,n5735);
and (n6310,n5692,n6311);
or (n6311,n6312,n6321,n6392);
and (n6312,n6313,n6315);
xor (n6313,n6314,n5262);
xor (n6314,n5185,n5230);
nor (n6315,n6316,n6318);
and (n6316,n6317,n5770);
nand (n6317,n6309,n5695);
and (n6318,n6319,n6320);
not (n6319,n6317);
not (n6320,n5770);
and (n6321,n6315,n6322);
or (n6322,n6323,n6332,n6391);
and (n6323,n6324,n6327);
xor (n6324,n6325,n5339);
not (n6325,n6326);
xnor (n6326,n5308,n5264);
nor (n6327,n6328,n6330);
and (n6328,n5845,n6329);
nand (n6329,n5773,n6308);
and (n6330,n5844,n6331);
not (n6331,n6329);
and (n6332,n6327,n6333);
or (n6333,n6334,n6347,n6390);
and (n6334,n6335,n6339);
xor (n6335,n6336,n5424);
not (n6336,n6337);
xor (n6337,n5341,n6338);
not (n6338,n5386);
nor (n6339,n6340,n6344);
and (n6340,n6341,n6343);
nand (n6341,n6342,n6306);
or (n6342,n5918,n5993);
nand (n6343,n6307,n6304);
and (n6344,n6345,n6346);
not (n6345,n6341);
not (n6346,n6343);
and (n6347,n6339,n6348);
or (n6348,n6349,n6363,n6389);
and (n6349,n6350,n6357);
xor (n6350,n6351,n5502);
not (n6351,n6352);
nor (n6352,n6353,n6355);
and (n6353,n5471,n6354);
not (n6354,n5426);
and (n6355,n6356,n5426);
not (n6356,n5471);
nand (n6357,n6358,n6362);
or (n6358,n6359,n5994);
not (n6359,n6360);
nand (n6360,n6361,n6306);
not (n6361,n5918);
nand (n6362,n6359,n5994);
and (n6363,n6357,n6364);
or (n6364,n6365,n6379,n6388);
not (n6365,n6366);
nand (n6366,n6367,n6375);
nand (n6367,n6368,n6374);
or (n6368,n6369,n6371);
not (n6369,n6370);
nor (n6370,n5998,n6299);
not (n6371,n6372);
nand (n6372,n6373,n6298);
or (n6373,n6068,n6146);
or (n6374,n6372,n6370);
nand (n6375,n6376,n6378);
or (n6376,n6377,n5593);
xor (n6377,n5504,n5557);
nand (n6378,n5593,n6377);
and (n6379,n6367,n6380);
not (n6380,n6381);
nand (n6381,n6382,n6387);
nand (n6382,n6383,n6386);
or (n6383,n6384,n6146);
nand (n6384,n6385,n6298);
not (n6385,n6068);
nand (n6386,n6146,n6384);
xor (n6387,n5595,n5646);
and (n6388,n6375,n6380);
and (n6389,n6350,n6364);
and (n6390,n6335,n6348);
and (n6391,n6324,n6333);
and (n6392,n6313,n6322);
and (n6393,n5690,n6311);
and (n6394,n6395,n6396);
xnor (n6395,n5684,n5688);
and (n6396,n6397,n6399);
xor (n6397,n6398,n6311);
xor (n6398,n5690,n5692);
and (n6399,n6400,n6402);
xor (n6400,n6401,n6322);
xor (n6401,n6313,n6315);
and (n6402,n6403,n6405);
xor (n6403,n6404,n6333);
xor (n6404,n6324,n6327);
and (n6405,n6406,n6408);
xor (n6406,n6407,n6348);
xor (n6407,n6335,n6339);
and (n6408,n6409,n6411);
xor (n6409,n6410,n6364);
xor (n6410,n6350,n6357);
and (n6411,n6412,n6414);
xor (n6412,n6413,n6380);
xor (n6413,n6375,n6367);
and (n6414,n6415,n6416);
xor (n6415,n6387,n6382);
not (n6416,n6417);
nand (n6417,n6418,n6424);
not (n6418,n6419);
xor (n6419,n6420,n6423);
not (n6420,n6421);
nand (n6421,n6422,n6293);
not (n6422,n6149);
not (n6423,n6221);
not (n6424,n6425);
xor (n6425,n6222,n6258);
and (n6426,n6427,n6428);
xor (n6427,n6395,n6396);
or (n6428,n6429,n6866,n6929);
and (n6429,n6430,n6865);
or (n6430,n6431,n6490,n6864);
and (n6431,n6432,n6461);
nand (n6432,n6433,n6441,n6453,n6457);
nor (n6433,n6434,n6438);
and (n6434,n6435,n6437);
not (n6435,n6436);
nand (n6436,n4998,n4979);
and (n6438,n6439,n6440);
nor (n6439,n5091,n4979);
nor (n6441,n6442,n6449);
nand (n6442,n6443,n6444,n6445,n6446);
nand (n6443,n5709,n1316);
nand (n6444,n4948,n5009);
nand (n6445,n5016,n5743);
nor (n6446,n6447,n6448);
and (n6447,n5112,n5017);
and (n6448,n5050,n5014);
nand (n6449,n6450,n6451,n6452);
nand (n6450,n5699,n1246);
nand (n6451,n4985,n4999);
nand (n6452,n5013,n5739);
nand (n6453,n6454,n6456);
not (n6454,n6455);
nand (n6455,n5008,n4979);
nand (n6457,n6458,n6460);
not (n6458,n6459);
nand (n6459,n5008,n4978);
nand (n6461,n6462,n6471,n6482);
nor (n6462,n6463,n6468);
nand (n6463,n6464,n6465,n6466,n6467);
nand (n6464,n5058,n5731);
nand (n6465,n4981,n5727);
nand (n6466,n4989,n5042);
nand (n6467,n4995,n5037);
and (n6468,n6469,n6470);
and (n6469,n5040,n4978);
nor (n6471,n6472,n6476);
nand (n6472,n6473,n6474,n6475);
nand (n6473,n5756,n1265);
nand (n6474,n5001,n5072);
nand (n6475,n5019,n5069);
nand (n6476,n6477,n6479);
or (n6477,n3046,n6478);
not (n6478,n5765);
nand (n6479,n6480,n6481);
and (n6480,n5040,n4979);
nor (n6482,n6483,n6486);
and (n6483,n6484,n6485);
and (n6484,n5031,n4979);
and (n6486,n6487,n6489);
not (n6487,n6488);
nand (n6488,n5031,n4978);
and (n6490,n6432,n6491);
or (n6491,n6492,n6539,n6863);
and (n6492,n6493,n6517);
nand (n6493,n6494,n6502,n6512);
nor (n6494,n6495,n6500);
nand (n6495,n6496,n6497,n6498,n6499);
nand (n6496,n5058,n5826);
nand (n6497,n4981,n5822);
nand (n6498,n4989,n5117);
nand (n6499,n4995,n5119);
and (n6500,n6487,n6501);
nor (n6502,n6503,n6507);
nand (n6503,n6504,n6505,n6506);
nand (n6504,n5796,n1265);
nand (n6505,n5001,n5178);
nand (n6506,n5019,n5176);
nand (n6507,n6508,n6510);
or (n6508,n3046,n6509);
not (n6509,n5805);
nand (n6510,n6480,n6511);
nor (n6512,n6513,n6515);
and (n6513,n6484,n6514);
and (n6515,n6469,n6516);
nand (n6517,n6518,n6523,n6535,n6537);
nor (n6518,n6519,n6521);
and (n6519,n6435,n6520);
and (n6521,n6439,n6522);
nor (n6523,n6524,n6531);
nand (n6524,n6525,n6526,n6527,n6528);
nand (n6525,n5833,n1316);
nand (n6526,n4948,n5152);
nand (n6527,n5016,n5784);
nor (n6528,n6529,n6530);
and (n6529,n5112,n5105);
and (n6530,n5050,n5123);
nand (n6531,n6532,n6533,n6534);
nand (n6532,n5839,n1246);
nand (n6533,n4985,n5146);
nand (n6534,n5013,n5778);
nand (n6535,n6454,n6536);
nand (n6537,n6458,n6538);
and (n6539,n6517,n6540);
or (n6540,n6541,n6588,n6862);
and (n6541,n6542,n6566);
nand (n6542,n6543,n6551,n6561);
nor (n6543,n6544,n6549);
nand (n6544,n6545,n6546,n6547,n6548);
nand (n6545,n5892,n5058);
nand (n6546,n4981,n5896);
nand (n6547,n4989,n5221);
nand (n6548,n4995,n5223);
and (n6549,n6469,n6550);
nor (n6551,n6552,n6556);
nand (n6552,n6553,n6554,n6555);
nand (n6553,n5871,n1265);
nand (n6554,n5001,n5256);
nand (n6555,n5019,n5254);
nand (n6556,n6557,n6559);
or (n6557,n3046,n6558);
not (n6558,n5879);
nand (n6559,n6480,n6560);
nor (n6561,n6562,n6564);
and (n6562,n6487,n6563);
and (n6564,n6484,n6565);
nand (n6566,n6567,n6572,n6584,n6586);
nor (n6567,n6568,n6570);
and (n6568,n6435,n6569);
and (n6570,n6439,n6571);
nor (n6572,n6573,n6580);
nand (n6573,n6574,n6575,n6576,n6577);
nand (n6574,n5905,n1316);
nand (n6575,n4948,n5204);
nand (n6576,n5016,n5855);
nor (n6577,n6578,n6579);
and (n6578,n5112,n5210);
and (n6579,n5050,n5227);
nand (n6580,n6581,n6582,n6583);
nand (n6581,n5913,n1246);
nand (n6582,n4985,n5202);
nand (n6583,n5013,n5860);
nand (n6584,n6454,n6585);
nand (n6586,n6458,n6587);
and (n6588,n6566,n6589);
or (n6589,n6590,n6638,n6861);
and (n6590,n6591,n6615);
nand (n6591,n6592,n6602,n6610);
nor (n6592,n6593,n6597);
nand (n6593,n6594,n6595,n6596);
nand (n6594,n5944,n1265);
nand (n6595,n5001,n5307);
nand (n6596,n5019,n5305);
nand (n6597,n6598,n6600);
or (n6598,n3046,n6599);
not (n6599,n5952);
nand (n6600,n6480,n6601);
nor (n6602,n6603,n6608);
nand (n6603,n6604,n6605,n6606,n6607);
nand (n6604,n4995,n5274);
nand (n6605,n5982,n5058);
nand (n6606,n4981,n5986);
nand (n6607,n4989,n5295);
and (n6608,n6469,n6609);
nor (n6610,n6611,n6613);
and (n6611,n6487,n6612);
and (n6613,n6484,n6614);
nand (n6615,n6616,n6633);
and (n6616,n6617,n6629,n6631);
nor (n6617,n6618,n6625);
nand (n6618,n6619,n6620,n6621,n6622);
nand (n6619,n5968,n1246);
nand (n6620,n4948,n5319);
nand (n6621,n5016,n5939);
nor (n6622,n6623,n6624);
and (n6623,n5112,n5283);
and (n6624,n5050,n5281);
nand (n6625,n6626,n6627,n6628);
nand (n6626,n5960,n1316);
nand (n6627,n4985,n5321);
nand (n6628,n5013,n5934);
nand (n6629,n6454,n6630);
nand (n6631,n6435,n6632);
nor (n6633,n6634,n6636);
and (n6634,n6439,n6635);
and (n6636,n6458,n6637);
and (n6638,n6615,n6639);
or (n6639,n6640,n6694,n6860);
and (n6640,n6641,n6669);
nand (n6641,n6642,n6654,n6664);
nor (n6642,n6643,n6646,n6650);
nand (n6643,n6644,n6645);
or (n6644,n5402,n5144);
nand (n6645,n4995,n5351);
nand (n6646,n6647,n6649);
or (n6647,n6648,n4982);
not (n6648,n6065);
nand (n6649,n6061,n5058);
nor (n6650,n6651,n6653);
not (n6651,n6652);
not (n6653,n6469);
nor (n6654,n6655,n6659);
nand (n6655,n6656,n6657,n6658);
nand (n6656,n6002,n1265);
nand (n6657,n5001,n5379);
nand (n6658,n5019,n5377);
nand (n6659,n6660,n6662);
or (n6660,n3046,n6661);
not (n6661,n6010);
nand (n6662,n6480,n6663);
nor (n6664,n6665,n6667);
and (n6665,n6487,n6666);
and (n6667,n6484,n6668);
nand (n6669,n6670,n6687,n6692);
not (n6670,n6671);
nand (n6671,n6672,n6675);
or (n6672,n6673,n6455);
not (n6673,n6674);
nor (n6675,n6676,n6683);
nand (n6676,n6677,n6678,n6679,n6680);
nand (n6677,n6045,n1316);
nand (n6678,n4948,n5422);
nand (n6679,n5016,n6022);
nor (n6680,n6681,n6682);
and (n6681,n5112,n5360);
and (n6682,n5050,n5356);
nand (n6683,n6684,n6685,n6686);
nand (n6684,n6039,n1246);
nand (n6685,n5013,n6018);
nand (n6686,n4985,n5417);
nor (n6687,n6688,n6690);
and (n6688,n6435,n6689);
and (n6690,n6439,n6691);
nand (n6692,n6458,n6693);
and (n6694,n6669,n6695);
or (n6695,n6696,n6744,n6859);
and (n6696,n6697,n6721);
nand (n6697,n6698,n6706,n6716);
nor (n6698,n6699,n6704);
nand (n6699,n6700,n6701,n6702,n6703);
nand (n6700,n4995,n5432);
nand (n6701,n5058,n6101);
nand (n6702,n6097,n4981);
nand (n6703,n4989,n5457);
and (n6704,n6469,n6705);
nor (n6706,n6707,n6711);
nand (n6707,n6708,n6709,n6710);
nand (n6708,n5001,n5464);
nand (n6709,n6111,n1265);
nand (n6710,n5019,n5462);
nand (n6711,n6712,n6714);
or (n6712,n3046,n6713);
not (n6713,n6121);
nand (n6714,n6480,n6715);
nor (n6716,n6717,n6719);
and (n6717,n6487,n6718);
and (n6719,n6484,n6720);
nand (n6721,n6722,n6739);
and (n6722,n6723,n6735,n6737);
nor (n6723,n6724,n6731);
nand (n6724,n6725,n6726,n6727,n6728);
nand (n6725,n6072,n1316);
nand (n6726,n4948,n5484);
nand (n6727,n5016,n6139);
nor (n6728,n6729,n6730);
and (n6729,n5112,n5441);
and (n6730,n5050,n5443);
nand (n6731,n6732,n6733,n6734);
nand (n6732,n6083,n1246);
nand (n6733,n5013,n6143);
nand (n6734,n5480,n4985);
nand (n6735,n6454,n6736);
nand (n6737,n6458,n6738);
nor (n6739,n6740,n6742);
and (n6740,n6435,n6741);
and (n6742,n6439,n6743);
and (n6744,n6721,n6745);
or (n6745,n6746,n6799,n6858);
and (n6746,n6747,n6774);
nand (n6747,n6748,n6759,n6769);
nor (n6748,n6749,n6752,n6756);
nand (n6749,n6750,n6751);
or (n6750,n5527,n5144);
nand (n6751,n4995,n5530);
nand (n6752,n6753,n6755);
or (n6753,n6754,n4982);
not (n6754,n6204);
nand (n6755,n6200,n5058);
nor (n6756,n6757,n6653);
not (n6757,n6758);
nor (n6759,n6760,n6764);
nand (n6760,n6761,n6762,n6763);
nand (n6761,n6181,n1265);
nand (n6762,n5001,n5569);
nand (n6763,n5019,n5567);
nand (n6764,n6765,n6767);
or (n6765,n3046,n6766);
not (n6766,n6175);
nand (n6767,n6480,n6768);
nor (n6769,n6770,n6772);
and (n6770,n6487,n6771);
and (n6772,n6484,n6773);
nand (n6774,n6775,n6792,n6797);
not (n6775,n6776);
nand (n6776,n6777,n6780);
or (n6777,n6778,n6455);
not (n6778,n6779);
nor (n6780,n6781,n6788);
nand (n6781,n6782,n6783,n6784,n6785);
nand (n6782,n6216,n1316);
nand (n6783,n4948,n5548);
nand (n6784,n5016,n6170);
nor (n6785,n6786,n6787);
and (n6786,n5112,n5509);
and (n6787,n5050,n5513);
nand (n6788,n6789,n6790,n6791);
nand (n6789,n6210,n1246);
nand (n6790,n5013,n6164);
nand (n6791,n4985,n5550);
nor (n6792,n6793,n6795);
and (n6793,n6435,n6794);
and (n6795,n6439,n6796);
nand (n6797,n6458,n6798);
and (n6799,n6774,n6800);
and (n6800,n6801,n6833);
nand (n6801,n6802,n6820);
not (n6802,n6803);
nand (n6803,n6804,n6810,n6813,n6818);
not (n6804,n6805);
nand (n6805,n6806,n6808);
or (n6806,n4982,n6807);
not (n6807,n6276);
or (n6808,n5026,n6809);
not (n6809,n6272);
nor (n6810,n6811,n6812);
and (n6811,n4995,n5619);
and (n6812,n4989,n5617);
nor (n6813,n6814,n6816);
and (n6814,n6487,n6815);
and (n6816,n6484,n6817);
nand (n6818,n6469,n6819);
nor (n6820,n6821,n6826);
nand (n6821,n6822,n6824,n6825);
or (n6822,n6823,n6037);
not (n6823,n6253);
or (n6824,n5002,n6269);
or (n6825,n5020,n5668);
nand (n6826,n6827,n6831);
or (n6827,n6828,n6830);
not (n6828,n6829);
not (n6830,n6480);
or (n6831,n6832,n3046);
not (n6832,n6247);
nand (n6833,n6834,n6853);
and (n6834,n6835,n6849,n6851);
nor (n6835,n6836,n6843);
nand (n6836,n6837,n6838,n6839,n6840);
nand (n6837,n6288,n1316);
nand (n6838,n5013,n6236);
nand (n6839,n4985,n5637);
nor (n6840,n6841,n6842);
and (n6841,n5050,n5601);
and (n6842,n5112,n5599);
nand (n6843,n6844,n6846,n6848);
or (n6844,n6845,n1247);
not (n6845,n6282);
or (n6846,n4949,n6847);
not (n6847,n5645);
nand (n6848,n5016,n6242);
nand (n6849,n6454,n6850);
nand (n6851,n6458,n6852);
nor (n6853,n6854,n6856);
and (n6854,n6435,n6855);
and (n6856,n6439,n6857);
and (n6858,n6747,n6800);
and (n6859,n6697,n6745);
and (n6860,n6641,n6695);
and (n6861,n6591,n6639);
and (n6862,n6542,n6589);
and (n6863,n6493,n6540);
and (n6864,n6461,n6491);
xor (n6865,n6397,n6399);
and (n6866,n6865,n6867);
or (n6867,n6868,n6872,n6928);
and (n6868,n6869,n6871);
xor (n6869,n6870,n6491);
xor (n6870,n6432,n6461);
xor (n6871,n6400,n6402);
and (n6872,n6871,n6873);
or (n6873,n6874,n6878,n6927);
and (n6874,n6875,n6877);
xor (n6875,n6876,n6540);
xor (n6876,n6493,n6517);
xor (n6877,n6403,n6405);
and (n6878,n6877,n6879);
or (n6879,n6880,n6884,n6926);
and (n6880,n6881,n6883);
xor (n6881,n6882,n6589);
xor (n6882,n6542,n6566);
xor (n6883,n6406,n6408);
and (n6884,n6883,n6885);
or (n6885,n6886,n6901,n6925);
and (n6886,n6887,n6889);
xor (n6887,n6888,n6639);
xor (n6888,n6591,n6615);
xor (n6889,n6890,n6898);
xor (n6890,n5502,n6891);
nand (n6891,n6892,n6366);
or (n6892,n6893,n6897);
not (n6893,n6894);
nand (n6894,n6895,n6381);
or (n6895,n6896,n6417);
nor (n6896,n6382,n6387);
nor (n6897,n6367,n6375);
nand (n6898,n6899,n6900);
or (n6899,n6352,n6357);
nand (n6900,n6357,n6352);
and (n6901,n6889,n6902);
or (n6902,n6903,n6907,n6924);
and (n6903,n6904,n6906);
xor (n6904,n6905,n6695);
xor (n6905,n6641,n6669);
xor (n6906,n6412,n6414);
and (n6907,n6906,n6908);
or (n6908,n6909,n6913,n6923);
and (n6909,n6910,n6912);
xor (n6910,n6911,n6745);
xor (n6911,n6697,n6721);
xor (n6912,n6415,n6416);
and (n6913,n6912,n6914);
or (n6914,n6915,n6919,n6922);
and (n6915,n6916,n6918);
xor (n6916,n6917,n6800);
xor (n6917,n6747,n6774);
xor (n6918,n6418,n6424);
and (n6919,n6918,n6920);
and (n6920,n6921,n6425);
xor (n6921,n6801,n6833);
and (n6922,n6916,n6920);
and (n6923,n6910,n6914);
and (n6924,n6904,n6908);
and (n6925,n6887,n6902);
and (n6926,n6881,n6885);
and (n6927,n6875,n6879);
and (n6928,n6869,n6873);
and (n6929,n6430,n6867);
or (n6930,n6931,n6933,n6973);
and (n6931,n6932,n6871);
xor (n6932,n6427,n6428);
and (n6933,n6871,n6934);
or (n6934,n6935,n6938,n6972);
and (n6935,n6936,n6877);
xor (n6936,n6937,n6867);
xor (n6937,n6430,n6865);
and (n6938,n6877,n6939);
or (n6939,n6940,n6943,n6971);
and (n6940,n6941,n6883);
xor (n6941,n6942,n6873);
xor (n6942,n6869,n6871);
and (n6943,n6883,n6944);
or (n6944,n6945,n6948,n6970);
and (n6945,n6946,n6889);
xor (n6946,n6947,n6879);
xor (n6947,n6875,n6877);
and (n6948,n6889,n6949);
or (n6949,n6950,n6953,n6969);
and (n6950,n6951,n6906);
xor (n6951,n6952,n6885);
xor (n6952,n6881,n6883);
and (n6953,n6906,n6954);
or (n6954,n6955,n6958,n6968);
and (n6955,n6956,n6912);
xor (n6956,n6957,n6902);
xor (n6957,n6887,n6889);
and (n6958,n6912,n6959);
or (n6959,n6960,n6963,n6967);
and (n6960,n6961,n6918);
xor (n6961,n6962,n6908);
xor (n6962,n6904,n6906);
and (n6963,n6918,n6964);
and (n6964,n6965,n6425);
xor (n6965,n6966,n6914);
xor (n6966,n6910,n6912);
and (n6967,n6961,n6964);
and (n6968,n6956,n6959);
and (n6969,n6951,n6954);
and (n6970,n6946,n6949);
and (n6971,n6941,n6944);
and (n6972,n6936,n6939);
and (n6973,n6932,n6934);
and (n6974,n6975,n6977);
xor (n6975,n6976,n6934);
xor (n6976,n6932,n6871);
and (n6977,n6978,n6980);
xor (n6978,n6979,n6939);
xor (n6979,n6936,n6877);
and (n6980,n6981,n6983);
xor (n6981,n6982,n6944);
xor (n6982,n6941,n6883);
and (n6983,n6984,n6986);
xor (n6984,n6985,n6949);
xor (n6985,n6946,n6889);
and (n6986,n6987,n6989);
xor (n6987,n6988,n6954);
xor (n6988,n6951,n6906);
xor (n6989,n6990,n6959);
xor (n6990,n6956,n6912);
nor (n6991,n6992,n1105);
not (n6992,n6993);
nor (n6993,n6994,n6,n6997);
and (n6994,n6995,n6996);
nor (n6995,n7,n1107);
nand (n6996,n652,n726);
not (n6997,n806);
wire s0n6998,s1n6998,notn6998;
or (n6998,s0n6998,s1n6998);
not(notn6998,n6991);
and (s0n6998,notn6998,1'b0);
and (s1n6998,n6991,n6999);
xor (n6999,n7000,n7016);
xor (n7000,n7001,n7007);
and (n7001,n7002,n7006);
xor (n7002,n7003,n7005);
not (n7003,n7004);
or (n7004,n4940,n5683);
and (n7005,n4939,n6394);
and (n7006,n4938,n6426);
and (n7007,n4938,n7008);
or (n7008,n7009,n7010,n7015);
xor (n7009,n7002,n7006);
and (n7010,n6427,n7011);
or (n7011,n7012,n7013,n7014);
and (n7012,n4937,n6865);
and (n7013,n6865,n6930);
and (n7014,n4937,n6930);
and (n7015,n7009,n7011);
and (n7016,n7017,n7020);
xor (n7017,n7018,n7008);
xor (n7018,n7019,n4938);
xor (n7019,n7002,n7001);
and (n7020,n7021,n7023);
xor (n7021,n7022,n7011);
xor (n7022,n7009,n6427);
and (n7023,n4935,n6974);
wire s0n7024,s1n7024,notn7024;
or (n7024,s0n7024,s1n7024);
not(notn7024,n6991);
and (s0n7024,notn7024,1'b0);
and (s1n7024,n6991,n7025);
xor (n7025,n7026,n7028);
xor (n7026,n7001,n7027);
and (n7027,n7002,n7007);
and (n7028,n7000,n7016);
or (n7029,n4959,n7030);
and (n7030,n652,n1344,n7,n1107);
not (n7031,n7032);
or (n7032,1'b0,n7033,n7036,n7039,n7041);
and (n7033,n7034,n1189);
wire s0n7034,s1n7034,notn7034;
or (n7034,s0n7034,s1n7034);
not(notn7034,n4923);
and (s0n7034,notn7034,1'b0);
and (s1n7034,n4923,n7035);
and (n7036,n7037,n6);
wire s0n7037,s1n7037,notn7037;
or (n7037,s0n7037,s1n7037);
not(notn7037,n1194);
and (s0n7037,notn7037,1'b0);
and (s1n7037,n1194,n7038);
and (n7039,n4931,n7040);
not (n7040,n4960);
or (n7041,1'b0,n7042,n7065,n7085,n7105);
and (n7042,n7043,n1331);
or (n7043,1'b0,n7044,n7051,n7057);
and (n7044,n7045,n7050);
or (n7045,1'b0,n7046,n7047,n7048,n7049);
and (n7046,n2581,n1187);
and (n7047,n2583,n1186);
and (n7048,n2585,n1183);
and (n7049,n2579,n817);
nor (n7050,n652,n1344,n7,n1107);
and (n7051,n7052,n7030);
or (n7052,1'b0,n7053,n7054,n7055,n7056);
and (n7053,n2542,n1187);
and (n7054,n2545,n1186);
and (n7055,n2537,n1183);
and (n7056,n2539,n817);
and (n7057,n7058,n7063);
or (n7058,1'b0,n7059,n7060,n7061,n7062);
and (n7059,n2545,n1187);
and (n7060,n2537,n1186);
and (n7061,n2539,n1183);
and (n7062,n2529,n817);
or (n7063,n4959,n7064);
nor (n7064,n652,n726,n7,n1107);
and (n7065,n7066,n1316);
or (n7066,1'b0,n7067,n7073,n7079);
and (n7067,n7068,n7050);
or (n7068,1'b0,n7069,n7070,n7071,n7072);
and (n7069,n2596,n1187);
and (n7070,n2598,n1186);
and (n7071,n2600,n1183);
and (n7072,n2594,n817);
and (n7073,n7074,n7030);
or (n7074,1'b0,n7075,n7076,n7077,n7078);
and (n7075,n2529,n1187);
and (n7076,n2533,n1186);
and (n7077,n2524,n1183);
and (n7078,n2526,n817);
and (n7079,n7080,n7063);
or (n7080,1'b0,n7081,n7082,n7083,n7084);
and (n7081,n2533,n1187);
and (n7082,n2524,n1186);
and (n7083,n2526,n1183);
and (n7084,n2531,n817);
and (n7085,n7086,n1265);
or (n7086,1'b0,n7087,n7093,n7099);
and (n7087,n7088,n7050);
or (n7088,1'b0,n7089,n7090,n7091,n7092);
and (n7089,n2567,n1187);
and (n7090,n2605,n1186);
and (n7091,n2602,n1183);
and (n7092,n2561,n817);
and (n7093,n7094,n7030);
or (n7094,1'b0,n7095,n7096,n7097,n7098);
and (n7095,n2517,n1187);
and (n7096,n2519,n1186);
and (n7097,n2550,n1183);
and (n7098,n2555,n817);
and (n7099,n7100,n7063);
or (n7100,1'b0,n7101,n7102,n7103,n7104);
and (n7101,n2519,n1187);
and (n7102,n2550,n1186);
and (n7103,n2555,n1183);
and (n7104,n2508,n817);
and (n7105,n7106,n1246);
or (n7106,1'b0,n7107,n7113,n7119);
and (n7107,n7108,n7050);
or (n7108,1'b0,n7109,n7110,n7111,n7112);
and (n7109,n2564,n1187);
and (n7110,n2587,n1186);
and (n7111,n2607,n1183);
and (n7112,n2569,n817);
and (n7113,n7114,n7030);
or (n7114,1'b0,n7115,n7116,n7117,n7118);
and (n7115,n2508,n1187);
and (n7116,n2512,n1186);
and (n7117,n2548,n1183);
and (n7118,n2553,n817);
and (n7119,n7120,n7063);
or (n7120,1'b0,n7121,n7122,n7123,n7124);
and (n7121,n2512,n1187);
and (n7122,n2548,n1186);
and (n7123,n2553,n1183);
and (n7124,n2515,n817);
nand (n7125,n7126,n7147);
not (n7126,n7127);
or (n7127,1'b0,n7128,n7139,n7141,n7142);
and (n7128,n7129,n1189);
wire s0n7129,s1n7129,notn7129;
or (n7129,s0n7129,s1n7129);
not(notn7129,n4923);
and (s0n7129,notn7129,1'b0);
and (s1n7129,n4923,n7130);
wire s0n7130,s1n7130,notn7130;
or (n7130,s0n7130,s1n7130);
not(notn7130,n4903);
and (s0n7130,notn7130,n7131);
and (s1n7130,n4903,1'b0);
wire s0n7131,s1n7131,notn7131;
or (n7131,s0n7131,s1n7131);
not(notn7131,n4777);
and (s0n7131,notn7131,n7132);
and (s1n7131,n4777,1'b1);
wire s0n7132,s1n7132,notn7132;
or (n7132,s0n7132,s1n7132);
not(notn7132,n1102);
and (s0n7132,notn7132,n7133);
and (s1n7132,n1102,n7136);
wire s0n7133,s1n7133,notn7133;
or (n7133,s0n7133,s1n7133);
not(notn7133,n1102);
and (s0n7133,notn7133,n7134);
and (s1n7133,n1102,n7135);
xor (n7134,n4099,n4101);
not (n7135,n4099);
wire s0n7136,s1n7136,notn7136;
or (n7136,s0n7136,s1n7136);
not(notn7136,n1102);
and (s0n7136,notn7136,n7137);
and (s1n7136,n1102,n7138);
xor (n7137,n4759,n4761);
xor (n7138,n4759,n4773);
and (n7139,n7140,n6);
wire s0n7140,s1n7140,notn7140;
or (n7140,s0n7140,s1n7140);
not(notn7140,n1194);
and (s0n7140,notn7140,1'b0);
and (s1n7140,n1194,n7130);
and (n7141,n7130,n4929);
and (n7142,n7143,n7029);
wire s0n7143,s1n7143,notn7143;
or (n7143,s0n7143,s1n7143);
not(notn7143,n7024);
and (s0n7143,notn7143,n7144);
and (s1n7143,n7024,1'b0);
wire s0n7144,s1n7144,notn7144;
or (n7144,s0n7144,s1n7144);
not(notn7144,n6998);
and (s0n7144,notn7144,n7145);
and (s1n7144,n6998,1'b1);
wire s0n7145,s1n7145,notn7145;
or (n7145,s0n7145,s1n7145);
not(notn7145,n6991);
and (s0n7145,notn7145,1'b0);
and (s1n7145,n6991,n7146);
xor (n7146,n6975,n6977);
not (n7147,n7148);
or (n7148,1'b0,n7149,n7152,n7155,n7156);
and (n7149,n7150,n1189);
wire s0n7150,s1n7150,notn7150;
or (n7150,s0n7150,s1n7150);
not(notn7150,n4923);
and (s0n7150,notn7150,1'b0);
and (s1n7150,n4923,n7151);
and (n7152,n7153,n6);
wire s0n7153,s1n7153,notn7153;
or (n7153,s0n7153,s1n7153);
not(notn7153,n1194);
and (s0n7153,notn7153,1'b0);
and (s1n7153,n1194,n7154);
and (n7155,n7143,n7040);
or (n7156,1'b0,n7157,n7177,n7197,n7217);
and (n7157,n7158,n1331);
or (n7158,1'b0,n7159,n7165,n7171);
and (n7159,n7160,n7050);
or (n7160,1'b0,n7161,n7162,n7163,n7164);
and (n7161,n2687,n1187);
and (n7162,n2689,n1186);
and (n7163,n2691,n1183);
and (n7164,n2685,n817);
and (n7165,n7166,n7030);
or (n7166,1'b0,n7167,n7168,n7169,n7170);
and (n7167,n2625,n1187);
and (n7168,n2630,n1186);
and (n7169,n2620,n1183);
and (n7170,n2618,n817);
and (n7171,n7172,n7063);
or (n7172,1'b0,n7173,n7174,n7175,n7176);
and (n7173,n2630,n1187);
and (n7174,n2620,n1186);
and (n7175,n2618,n1183);
and (n7176,n2627,n817);
and (n7177,n7178,n1316);
or (n7178,1'b0,n7179,n7185,n7191);
and (n7179,n7180,n7050);
or (n7180,1'b0,n7181,n7182,n7183,n7184);
and (n7181,n2706,n1187);
and (n7182,n2696,n1186);
and (n7183,n2698,n1183);
and (n7184,n2704,n817);
and (n7185,n7186,n7030);
or (n7186,1'b0,n7187,n7188,n7189,n7190);
and (n7187,n2627,n1187);
and (n7188,n2646,n1186);
and (n7189,n2637,n1183);
and (n7190,n2635,n817);
and (n7191,n7192,n7063);
or (n7192,1'b0,n7193,n7194,n7195,n7196);
and (n7193,n2646,n1187);
and (n7194,n2637,n1186);
and (n7195,n2635,n1183);
and (n7196,n2643,n817);
and (n7197,n7198,n1265);
or (n7198,1'b0,n7199,n7205,n7211);
and (n7199,n7200,n7050);
or (n7200,1'b0,n7201,n7202,n7203,n7204);
and (n7201,n2711,n1187);
and (n7202,n2715,n1186);
and (n7203,n2718,n1183);
and (n7204,n2721,n817);
and (n7205,n7206,n7030);
or (n7206,1'b0,n7207,n7208,n7209,n7210);
and (n7207,n2652,n1187);
and (n7208,n2651,n1186);
and (n7209,n2655,n1183);
and (n7210,n2658,n817);
and (n7211,n7212,n7063);
or (n7212,1'b0,n7213,n7214,n7215,n7216);
and (n7213,n2651,n1187);
and (n7214,n2655,n1186);
and (n7215,n2658,n1183);
and (n7216,n2661,n817);
and (n7217,n7218,n1246);
or (n7218,1'b0,n7219,n7225,n7231);
and (n7219,n7220,n7050);
or (n7220,1'b0,n7221,n7222,n7223,n7224);
and (n7221,n2726,n1187);
and (n7222,n2729,n1186);
and (n7223,n2732,n1183);
and (n7224,n2735,n817);
and (n7225,n7226,n7030);
or (n7226,1'b0,n7227,n7228,n7229,n7230);
and (n7227,n2661,n1187);
and (n7228,n2666,n1186);
and (n7229,n2669,n1183);
and (n7230,n2672,n817);
and (n7231,n7232,n7063);
or (n7232,1'b0,n7233,n7234,n7235,n7236);
and (n7233,n2666,n1187);
and (n7234,n2669,n1186);
and (n7235,n2672,n1183);
and (n7236,n2675,n817);
nand (n7237,n7238,n7749);
or (n7238,n7239,n7347);
not (n7239,n7240);
not (n7240,n7241);
and (n7241,n7242,n7335);
or (n7242,1'b0,n7243,n7246,n7249,n7254);
and (n7243,n7244,n1189);
wire s0n7244,s1n7244,notn7244;
or (n7244,s0n7244,s1n7244);
not(notn7244,n4923);
and (s0n7244,notn7244,1'b0);
and (s1n7244,n4923,n7245);
and (n7246,n7247,n6);
wire s0n7247,s1n7247,notn7247;
or (n7247,s0n7247,s1n7247);
not(notn7247,n1194);
and (s0n7247,notn7247,1'b0);
and (s1n7247,n1194,n7248);
and (n7249,n7250,n7040);
wire s0n7250,s1n7250,notn7250;
or (n7250,s0n7250,s1n7250);
not(notn7250,n7024);
and (s0n7250,notn7250,n7251);
and (s1n7250,n7024,1'b0);
wire s0n7251,s1n7251,notn7251;
or (n7251,s0n7251,s1n7251);
not(notn7251,n6998);
and (s0n7251,notn7251,n7252);
and (s1n7251,n6998,1'b1);
wire s0n7252,s1n7252,notn7252;
or (n7252,s0n7252,s1n7252);
not(notn7252,n6991);
and (s0n7252,notn7252,1'b0);
and (s1n7252,n6991,n7253);
xor (n7253,n6978,n6980);
or (n7254,1'b0,n7255,n7275,n7295,n7315);
and (n7255,n7256,n1331);
or (n7256,1'b0,n7257,n7263,n7269);
and (n7257,n7258,n7050);
or (n7258,1'b0,n7259,n7260,n7261,n7262);
and (n7259,n2819,n1187);
and (n7260,n2810,n1186);
and (n7261,n2812,n1183);
and (n7262,n2817,n817);
and (n7263,n7264,n7030);
or (n7264,1'b0,n7265,n7266,n7267,n7268);
and (n7265,n2753,n1187);
and (n7266,n2758,n1186);
and (n7267,n2746,n1183);
and (n7268,n2748,n817);
and (n7269,n7270,n7063);
or (n7270,1'b0,n7271,n7272,n7273,n7274);
and (n7271,n2758,n1187);
and (n7272,n2746,n1186);
and (n7273,n2748,n1183);
and (n7274,n2755,n817);
and (n7275,n7276,n1316);
or (n7276,1'b0,n7277,n7283,n7289);
and (n7277,n7278,n7050);
or (n7278,1'b0,n7279,n7280,n7281,n7282);
and (n7279,n2831,n1187);
and (n7280,n2823,n1186);
and (n7281,n2825,n1183);
and (n7282,n2829,n817);
and (n7283,n7284,n7030);
or (n7284,1'b0,n7285,n7286,n7287,n7288);
and (n7285,n2755,n1187);
and (n7286,n2774,n1186);
and (n7287,n2763,n1183);
and (n7288,n2765,n817);
and (n7289,n7290,n7063);
or (n7290,1'b0,n7291,n7292,n7293,n7294);
and (n7291,n2774,n1187);
and (n7292,n2763,n1186);
and (n7293,n2765,n1183);
and (n7294,n2771,n817);
and (n7295,n7296,n1265);
or (n7296,1'b0,n7297,n7303,n7309);
and (n7297,n7298,n7050);
or (n7298,1'b0,n7299,n7300,n7301,n7302);
and (n7299,n2836,n1187);
and (n7300,n2840,n1186);
and (n7301,n2843,n1183);
and (n7302,n2846,n817);
and (n7303,n7304,n7030);
or (n7304,1'b0,n7305,n7306,n7307,n7308);
and (n7305,n2780,n1187);
and (n7306,n2779,n1186);
and (n7307,n2783,n1183);
and (n7308,n2786,n817);
and (n7309,n7310,n7063);
or (n7310,1'b0,n7311,n7312,n7313,n7314);
and (n7311,n2779,n1187);
and (n7312,n2783,n1186);
and (n7313,n2786,n1183);
and (n7314,n2789,n817);
and (n7315,n7316,n1246);
or (n7316,1'b0,n7317,n7323,n7329);
and (n7317,n7318,n7050);
or (n7318,1'b0,n7319,n7320,n7321,n7322);
and (n7319,n2851,n1187);
and (n7320,n2854,n1186);
and (n7321,n2857,n1183);
and (n7322,n2860,n817);
and (n7323,n7324,n7030);
or (n7324,1'b0,n7325,n7326,n7327,n7328);
and (n7325,n2789,n1187);
and (n7326,n2794,n1186);
and (n7327,n2797,n1183);
and (n7328,n2800,n817);
and (n7329,n7330,n7063);
or (n7330,1'b0,n7331,n7332,n7333,n7334);
and (n7331,n2794,n1187);
and (n7332,n2797,n1186);
and (n7333,n2800,n1183);
and (n7334,n2803,n817);
or (n7335,1'b0,n7336,n7343,n7345,n7346);
and (n7336,n7337,n1189);
wire s0n7337,s1n7337,notn7337;
or (n7337,s0n7337,s1n7337);
not(notn7337,n4923);
and (s0n7337,notn7337,1'b0);
and (s1n7337,n4923,n7338);
wire s0n7338,s1n7338,notn7338;
or (n7338,s0n7338,s1n7338);
not(notn7338,n4903);
and (s0n7338,notn7338,n7339);
and (s1n7338,n4903,1'b0);
wire s0n7339,s1n7339,notn7339;
or (n7339,s0n7339,s1n7339);
not(notn7339,n4777);
and (s0n7339,notn7339,n7340);
and (s1n7339,n4777,1'b1);
wire s0n7340,s1n7340,notn7340;
or (n7340,s0n7340,s1n7340);
not(notn7340,n1102);
and (s0n7340,notn7340,n7341);
and (s1n7340,n1102,n4778);
wire s0n7341,s1n7341,notn7341;
or (n7341,s0n7341,s1n7341);
not(notn7341,n1102);
and (s0n7341,notn7341,n7342);
and (s1n7341,n1102,n4102);
xor (n7342,n4102,n4104);
and (n7343,n7344,n6);
wire s0n7344,s1n7344,notn7344;
or (n7344,s0n7344,s1n7344);
not(notn7344,n1194);
and (s0n7344,notn7344,1'b0);
and (s1n7344,n1194,n7338);
and (n7345,n7338,n4929);
and (n7346,n7250,n7029);
not (n7347,n7348);
nor (n7348,n7349,n7748);
and (n7349,n7350,n7459);
or (n7350,n7351,n7370);
or (n7351,1'b0,n7352,n7362,n7364,n7365);
and (n7352,n7353,n1189);
wire s0n7353,s1n7353,notn7353;
or (n7353,s0n7353,s1n7353);
not(notn7353,n4923);
and (s0n7353,notn7353,1'b0);
and (s1n7353,n4923,n7354);
wire s0n7354,s1n7354,notn7354;
or (n7354,s0n7354,s1n7354);
not(notn7354,n4903);
and (s0n7354,notn7354,n7355);
and (s1n7354,n4903,1'b0);
wire s0n7355,s1n7355,notn7355;
or (n7355,s0n7355,s1n7355);
not(notn7355,n4777);
and (s0n7355,notn7355,n7356);
and (s1n7355,n4777,1'b1);
wire s0n7356,s1n7356,notn7356;
or (n7356,s0n7356,s1n7356);
not(notn7356,n1102);
and (s0n7356,notn7356,n7357);
and (s1n7356,n1102,n7359);
wire s0n7357,s1n7357,notn7357;
or (n7357,s0n7357,s1n7357);
not(notn7357,n1102);
and (s0n7357,notn7357,n7358);
and (s1n7357,n1102,n4105);
xor (n7358,n4105,n4107);
wire s0n7359,s1n7359,notn7359;
or (n7359,s0n7359,s1n7359);
not(notn7359,n1102);
and (s0n7359,notn7359,n7360);
and (s1n7359,n1102,n7361);
xor (n7360,n4765,n4767);
xor (n7361,n4765,n4775);
and (n7362,n7363,n6);
wire s0n7363,s1n7363,notn7363;
or (n7363,s0n7363,s1n7363);
not(notn7363,n1194);
and (s0n7363,notn7363,1'b0);
and (s1n7363,n1194,n7354);
and (n7364,n7354,n4929);
and (n7365,n7366,n7029);
wire s0n7366,s1n7366,notn7366;
or (n7366,s0n7366,s1n7366);
not(notn7366,n7024);
and (s0n7366,notn7366,n7367);
and (s1n7366,n7024,1'b0);
wire s0n7367,s1n7367,notn7367;
or (n7367,s0n7367,s1n7367);
not(notn7367,n6998);
and (s0n7367,notn7367,n7368);
and (s1n7367,n6998,1'b1);
wire s0n7368,s1n7368,notn7368;
or (n7368,s0n7368,s1n7368);
not(notn7368,n6991);
and (s0n7368,notn7368,1'b0);
and (s1n7368,n6991,n7369);
xor (n7369,n6981,n6983);
or (n7370,1'b0,n7371,n7374,n7377,n7378);
and (n7371,n7372,n1189);
wire s0n7372,s1n7372,notn7372;
or (n7372,s0n7372,s1n7372);
not(notn7372,n4923);
and (s0n7372,notn7372,1'b0);
and (s1n7372,n4923,n7373);
and (n7374,n7375,n6);
wire s0n7375,s1n7375,notn7375;
or (n7375,s0n7375,s1n7375);
not(notn7375,n1194);
and (s0n7375,notn7375,1'b0);
and (s1n7375,n1194,n7376);
and (n7377,n7366,n7040);
or (n7378,1'b0,n7379,n7399,n7419,n7439);
and (n7379,n7380,n1331);
or (n7380,1'b0,n7381,n7387,n7393);
and (n7381,n7382,n7050);
or (n7382,1'b0,n7383,n7384,n7385,n7386);
and (n7383,n2932,n1187);
and (n7384,n2934,n1186);
and (n7385,n2936,n1183);
and (n7386,n2930,n817);
and (n7387,n7388,n7030);
or (n7388,1'b0,n7389,n7390,n7391,n7392);
and (n7389,n2871,n1187);
and (n7390,n2875,n1186);
and (n7391,n2877,n1183);
and (n7392,n2879,n817);
and (n7393,n7394,n7063);
or (n7394,1'b0,n7395,n7396,n7397,n7398);
and (n7395,n2875,n1187);
and (n7396,n2877,n1186);
and (n7397,n2879,n1183);
and (n7398,n2873,n817);
and (n7399,n7400,n1316);
or (n7400,1'b0,n7401,n7407,n7413);
and (n7401,n7402,n7050);
or (n7402,1'b0,n7403,n7404,n7405,n7406);
and (n7403,n2944,n1187);
and (n7404,n2946,n1186);
and (n7405,n2948,n1183);
and (n7406,n2941,n817);
and (n7407,n7408,n7030);
or (n7408,1'b0,n7409,n7410,n7411,n7412);
and (n7409,n2873,n1187);
and (n7410,n2887,n1186);
and (n7411,n2889,n1183);
and (n7412,n2891,n817);
and (n7413,n7414,n7063);
or (n7414,1'b0,n7415,n7416,n7417,n7418);
and (n7415,n2887,n1187);
and (n7416,n2889,n1186);
and (n7417,n2891,n1183);
and (n7418,n2885,n817);
and (n7419,n7420,n1265);
or (n7420,1'b0,n7421,n7427,n7433);
and (n7421,n7422,n7050);
or (n7422,1'b0,n7423,n7424,n7425,n7426);
and (n7423,n2953,n1187);
and (n7424,n2957,n1186);
and (n7425,n2960,n1183);
and (n7426,n2963,n817);
and (n7427,n7428,n7030);
or (n7428,1'b0,n7429,n7430,n7431,n7432);
and (n7429,n2897,n1187);
and (n7430,n2896,n1186);
and (n7431,n2900,n1183);
and (n7432,n2903,n817);
and (n7433,n7434,n7063);
or (n7434,1'b0,n7435,n7436,n7437,n7438);
and (n7435,n2896,n1187);
and (n7436,n2900,n1186);
and (n7437,n2903,n1183);
and (n7438,n2906,n817);
and (n7439,n7440,n1246);
or (n7440,1'b0,n7441,n7447,n7453);
and (n7441,n7442,n7050);
or (n7442,1'b0,n7443,n7444,n7445,n7446);
and (n7443,n2968,n1187);
and (n7444,n2971,n1186);
and (n7445,n2974,n1183);
and (n7446,n2977,n817);
and (n7447,n7448,n7030);
or (n7448,1'b0,n7449,n7450,n7451,n7452);
and (n7449,n2906,n1187);
and (n7450,n2911,n1186);
and (n7451,n2914,n1183);
and (n7452,n2917,n817);
and (n7453,n7454,n7063);
or (n7454,1'b0,n7455,n7456,n7457,n7458);
and (n7455,n2911,n1187);
and (n7456,n2914,n1186);
and (n7457,n2917,n1183);
and (n7458,n2920,n817);
nand (n7459,n7460,n7740);
or (n7460,n7461,n7634);
not (n7461,n7462);
nand (n7462,n7463,n7476);
or (n7463,n7464,n7470);
not (n7464,n7465);
nand (n7465,n7466,n7467,n7468);
or (n7466,n1229,n6997);
not (n7467,n1193);
not (n7468,n7469);
and (n7469,n1189,n805,n4924);
not (n7470,n7471);
wire s0n7471,s1n7471,notn7471;
or (n7471,s0n7471,s1n7471);
not(notn7471,n4903);
and (s0n7471,notn7471,n7472);
and (s1n7471,n4903,1'b0);
wire s0n7472,s1n7472,notn7472;
or (n7472,s0n7472,s1n7472);
not(notn7472,n4777);
and (s0n7472,notn7472,n7473);
and (s1n7472,n4777,1'b1);
wire s0n7473,s1n7473,notn7473;
or (n7473,s0n7473,s1n7473);
not(notn7473,n1102);
and (s0n7473,notn7473,n7474);
and (s1n7473,n1102,n1092);
wire s0n7474,s1n7474,notn7474;
or (n7474,s0n7474,s1n7474);
not(notn7474,n1102);
and (s0n7474,notn7474,n7475);
and (s1n7474,n1102,n4111);
xor (n7475,n4111,n4113);
nor (n7476,n7477,n7544);
and (n7477,n7478,n7536);
wire s0n7478,s1n7478,notn7478;
or (n7478,s0n7478,s1n7478);
not(notn7478,n7024);
and (s0n7478,notn7478,n7479);
and (s1n7478,n7024,1'b0);
wire s0n7479,s1n7479,notn7479;
or (n7479,s0n7479,s1n7479);
not(notn7479,n6998);
and (s0n7479,notn7479,n7480);
and (s1n7479,n6998,1'b1);
wire s0n7480,s1n7480,notn7480;
or (n7480,s0n7480,s1n7480);
not(notn7480,n6991);
and (s0n7480,notn7480,1'b0);
and (s1n7480,n6991,n7481);
xor (n7481,n7482,n7505);
xor (n7482,n7483,n7488);
xor (n7483,n7484,n6883);
xor (n7484,n7485,n7487);
or (n7485,n7486,n6590);
and (n7486,n6888,n6912);
xor (n7487,n6882,n6906);
nand (n7488,n7489,n7504);
or (n7489,n7490,n7496);
or (n7490,n7491,n7495);
and (n7491,n7492,n6906);
xor (n7492,n7493,n7494);
and (n7493,n6721,n6425);
xor (n7494,n6905,n6918);
and (n7495,n7493,n7494);
not (n7496,n7497);
or (n7497,n7498,n7503);
and (n7498,n7499,n6889);
xor (n7499,n7500,n7502);
or (n7500,n7501,n6640);
and (n7501,n6905,n6918);
xor (n7502,n6888,n6912);
and (n7503,n7500,n7502);
nand (n7504,n7496,n7490);
or (n7505,n7506,n7535);
and (n7506,n7507,n7510);
xor (n7507,n7508,n7509);
xor (n7508,n7499,n6889);
not (n7509,n7490);
or (n7510,n7511,n7534);
and (n7511,n7512,n7519);
xor (n7512,n7513,n7518);
or (n7513,n7514,n7517);
and (n7514,n7515,n6912);
xor (n7515,n6697,n7516);
xor (n7516,n6721,n6425);
and (n7517,n6697,n7516);
xor (n7518,n7492,n6906);
or (n7519,n7520,n7533);
and (n7520,n7521,n7525);
xor (n7521,n7522,n7524);
or (n7522,n7523,n6746);
and (n7523,n6917,n6918);
xor (n7524,n7515,n6912);
or (n7525,n7526,n7532);
and (n7526,n7527,n7530);
xor (n7527,n7528,n7529);
and (n7528,n6833,n6425);
xor (n7529,n6917,n6918);
and (n7530,n7531,n6801);
xor (n7531,n6833,n6425);
and (n7532,n7528,n7529);
and (n7533,n7522,n7524);
and (n7534,n7513,n7518);
and (n7535,n7508,n7509);
nand (n7536,n7537,n7539);
not (n7537,n7538);
and (n7538,n7040,n806);
not (n7539,n7540);
and (n7540,n7541,n7542,n806);
and (n7541,n1344,n7);
nor (n7542,n7543,n653);
not (n7543,n651);
nand (n7544,n7545,n7627);
not (n7545,n7546);
or (n7546,1'b0,n7547,n7567,n7587,n7607);
and (n7547,n7548,n1331);
or (n7548,1'b0,n7549,n7555,n7561);
and (n7549,n7550,n7050);
or (n7550,1'b0,n7551,n7552,n7553,n7554);
and (n7551,n3176,n1187);
and (n7552,n3171,n1186);
and (n7553,n3173,n1183);
and (n7554,n3182,n817);
and (n7555,n7556,n7030);
or (n7556,1'b0,n7557,n7558,n7559,n7560);
and (n7557,n3117,n1187);
and (n7558,n3119,n1186);
and (n7559,n3114,n1183);
and (n7560,n3112,n817);
and (n7561,n7562,n7063);
or (n7562,1'b0,n7563,n7564,n7565,n7566);
and (n7563,n3119,n1187);
and (n7564,n3114,n1186);
and (n7565,n3112,n1183);
and (n7566,n3121,n817);
and (n7567,n7568,n1316);
or (n7568,1'b0,n7569,n7575,n7581);
and (n7569,n7570,n7050);
or (n7570,1'b0,n7571,n7572,n7573,n7574);
and (n7571,n3192,n1187);
and (n7572,n3187,n1186);
and (n7573,n3189,n1183);
and (n7574,n3197,n817);
and (n7575,n7576,n7030);
or (n7576,1'b0,n7577,n7578,n7579,n7580);
and (n7577,n3121,n1187);
and (n7578,n3132,n1186);
and (n7579,n3126,n1183);
and (n7580,n3128,n817);
and (n7581,n7582,n7063);
or (n7582,1'b0,n7583,n7584,n7585,n7586);
and (n7583,n3132,n1187);
and (n7584,n3126,n1186);
and (n7585,n3128,n1183);
and (n7586,n3134,n817);
and (n7587,n7588,n1265);
or (n7588,1'b0,n7589,n7595,n7601);
and (n7589,n7590,n7050);
or (n7590,1'b0,n7591,n7592,n7593,n7594);
and (n7591,n3202,n1187);
and (n7592,n3206,n1186);
and (n7593,n3209,n1183);
and (n7594,n3212,n817);
and (n7595,n7596,n7030);
or (n7596,1'b0,n7597,n7598,n7599,n7600);
and (n7597,n3140,n1187);
and (n7598,n3139,n1186);
and (n7599,n3143,n1183);
and (n7600,n3146,n817);
and (n7601,n7602,n7063);
or (n7602,1'b0,n7603,n7604,n7605,n7606);
and (n7603,n3139,n1187);
and (n7604,n3143,n1186);
and (n7605,n3146,n1183);
and (n7606,n3149,n817);
and (n7607,n7608,n1246);
or (n7608,1'b0,n7609,n7615,n7621);
and (n7609,n7610,n7050);
or (n7610,1'b0,n7611,n7612,n7613,n7614);
and (n7611,n3217,n1187);
and (n7612,n3220,n1186);
and (n7613,n3223,n1183);
and (n7614,n3226,n817);
and (n7615,n7616,n7030);
or (n7616,1'b0,n7617,n7618,n7619,n7620);
and (n7617,n3149,n1187);
and (n7618,n3154,n1186);
and (n7619,n3157,n1183);
and (n7620,n3160,n817);
and (n7621,n7622,n7063);
or (n7622,1'b0,n7623,n7624,n7625,n7626);
and (n7623,n3154,n1187);
and (n7624,n3157,n1186);
and (n7625,n3160,n1183);
and (n7626,n3163,n817);
nor (n7627,n7628,n7631);
and (n7628,n7629,n1189);
wire s0n7629,s1n7629,notn7629;
or (n7629,s0n7629,s1n7629);
not(notn7629,n4923);
and (s0n7629,notn7629,1'b0);
and (s1n7629,n4923,n7630);
and (n7631,n7632,n6);
wire s0n7632,s1n7632,notn7632;
or (n7632,s0n7632,s1n7632);
not(notn7632,n1194);
and (s0n7632,notn7632,1'b0);
and (s1n7632,n1194,n7633);
not (n7634,n7635);
nand (n7635,n7636,n7645);
nand (n7636,n7637,n7465);
wire s0n7637,s1n7637,notn7637;
or (n7637,s0n7637,s1n7637);
not(notn7637,n4903);
and (s0n7637,notn7637,n7638);
and (s1n7637,n4903,1'b0);
wire s0n7638,s1n7638,notn7638;
or (n7638,s0n7638,s1n7638);
not(notn7638,n4777);
and (s0n7638,notn7638,n7639);
and (s1n7638,n4777,1'b1);
wire s0n7639,s1n7639,notn7639;
or (n7639,s0n7639,s1n7639);
not(notn7639,n1102);
and (s0n7639,notn7639,n7640);
and (s1n7639,n1102,n7642);
wire s0n7640,s1n7640,notn7640;
or (n7640,s0n7640,s1n7640);
not(notn7640,n1102);
and (s0n7640,notn7640,n7641);
and (s1n7640,n1102,n4108);
xor (n7641,n4108,n4110);
wire s0n7642,s1n7642,notn7642;
or (n7642,s0n7642,s1n7642);
not(notn7642,n1102);
and (s0n7642,notn7642,n7643);
and (s1n7642,n1102,n7644);
xor (n7643,n4768,n4770);
xor (n7644,n4768,n4776);
nor (n7645,n7646,n7739);
or (n7646,1'b0,n7647,n7650,n7653,n7658);
and (n7647,n7648,n1189);
wire s0n7648,s1n7648,notn7648;
or (n7648,s0n7648,s1n7648);
not(notn7648,n4923);
and (s0n7648,notn7648,1'b0);
and (s1n7648,n4923,n7649);
and (n7650,n7651,n6);
wire s0n7651,s1n7651,notn7651;
or (n7651,s0n7651,s1n7651);
not(notn7651,n1194);
and (s0n7651,notn7651,1'b0);
and (s1n7651,n1194,n7652);
and (n7653,n7654,n7040);
wire s0n7654,s1n7654,notn7654;
or (n7654,s0n7654,s1n7654);
not(notn7654,n7024);
and (s0n7654,notn7654,n7655);
and (s1n7654,n7024,1'b0);
wire s0n7655,s1n7655,notn7655;
or (n7655,s0n7655,s1n7655);
not(notn7655,n6998);
and (s0n7655,notn7655,n7656);
and (s1n7655,n6998,1'b1);
wire s0n7656,s1n7656,notn7656;
or (n7656,s0n7656,s1n7656);
not(notn7656,n6991);
and (s0n7656,notn7656,1'b0);
and (s1n7656,n6991,n7657);
xor (n7657,n6984,n6986);
or (n7658,1'b0,n7659,n7679,n7699,n7719);
and (n7659,n7660,n1331);
or (n7660,1'b0,n7661,n7667,n7673);
and (n7661,n7662,n7050);
or (n7662,1'b0,n7663,n7664,n7665,n7666);
and (n7663,n3055,n1187);
and (n7664,n3057,n1186);
and (n7665,n3059,n1183);
and (n7666,n3053,n817);
and (n7667,n7668,n7030);
or (n7668,1'b0,n7669,n7670,n7671,n7672);
and (n7669,n2989,n1187);
and (n7670,n2988,n1186);
and (n7671,n2992,n1183);
and (n7672,n2995,n817);
and (n7673,n7674,n7063);
or (n7674,1'b0,n7675,n7676,n7677,n7678);
and (n7675,n2988,n1187);
and (n7676,n2992,n1186);
and (n7677,n2995,n1183);
and (n7678,n2998,n817);
and (n7679,n7680,n1316);
or (n7680,1'b0,n7681,n7687,n7693);
and (n7681,n7682,n7050);
or (n7682,1'b0,n7683,n7684,n7685,n7686);
and (n7683,n3068,n1187);
and (n7684,n3070,n1186);
and (n7685,n3072,n1183);
and (n7686,n3066,n817);
and (n7687,n7688,n7030);
or (n7688,1'b0,n7689,n7690,n7691,n7692);
and (n7689,n2998,n1187);
and (n7690,n3009,n1186);
and (n7691,n3005,n1183);
and (n7692,n3003,n817);
and (n7693,n7694,n7063);
or (n7694,1'b0,n7695,n7696,n7697,n7698);
and (n7695,n3009,n1187);
and (n7696,n3005,n1186);
and (n7697,n3003,n1183);
and (n7698,n3011,n817);
and (n7699,n7700,n1265);
or (n7700,1'b0,n7701,n7707,n7713);
and (n7701,n7702,n7050);
or (n7702,1'b0,n7703,n7704,n7705,n7706);
and (n7703,n3077,n1187);
and (n7704,n3081,n1186);
and (n7705,n3084,n1183);
and (n7706,n3087,n817);
and (n7707,n7708,n7030);
or (n7708,1'b0,n7709,n7710,n7711,n7712);
and (n7709,n3017,n1187);
and (n7710,n3016,n1186);
and (n7711,n3020,n1183);
and (n7712,n3023,n817);
and (n7713,n7714,n7063);
or (n7714,1'b0,n7715,n7716,n7717,n7718);
and (n7715,n3016,n1187);
and (n7716,n3020,n1186);
and (n7717,n3023,n1183);
and (n7718,n3026,n817);
and (n7719,n7720,n1246);
or (n7720,1'b0,n7721,n7727,n7733);
and (n7721,n7722,n7050);
or (n7722,1'b0,n7723,n7724,n7725,n7726);
and (n7723,n3092,n1187);
and (n7724,n3095,n1186);
and (n7725,n3098,n1183);
and (n7726,n3101,n817);
and (n7727,n7728,n7030);
or (n7728,1'b0,n7729,n7730,n7731,n7732);
and (n7729,n3026,n1187);
and (n7730,n3031,n1186);
and (n7731,n3034,n1183);
and (n7732,n3037,n817);
and (n7733,n7734,n7063);
or (n7734,1'b0,n7735,n7736,n7737,n7738);
and (n7735,n3031,n1187);
and (n7736,n3034,n1186);
and (n7737,n3037,n1183);
and (n7738,n3040,n817);
and (n7739,n7654,n7029);
not (n7740,n7741);
and (n7741,n7646,n7742);
or (n7742,1'b0,n7743,n7745,n7747,n7739);
and (n7743,n7744,n1189);
wire s0n7744,s1n7744,notn7744;
or (n7744,s0n7744,s1n7744);
not(notn7744,n4923);
and (s0n7744,notn7744,1'b0);
and (s1n7744,n4923,n7637);
and (n7745,n7746,n6);
wire s0n7746,s1n7746,notn7746;
or (n7746,s0n7746,s1n7746);
not(notn7746,n1194);
and (s0n7746,notn7746,1'b0);
and (s1n7746,n1194,n7637);
and (n7747,n7637,n4929);
and (n7748,n7370,n7351);
or (n7749,n7335,n7242);
not (n7750,n7751);
nand (n7751,n7752,n7756);
or (n7752,n7753,n7754);
not (n7753,n1084);
not (n7754,n7755);
and (n7755,n7148,n7127);
not (n7756,n7757);
and (n7757,n7032,n1086);
nor (n7758,n7759,n7869);
not (n7759,n7760);
nand (n7760,n7761,n7779);
not (n7761,n7762);
or (n7762,1'b0,n7763,n7771,n7773,n7774);
and (n7763,n7764,n1189);
wire s0n7764,s1n7764,notn7764;
or (n7764,s0n7764,s1n7764);
not(notn7764,n4923);
and (s0n7764,notn7764,1'b0);
and (s1n7764,n4923,n7765);
wire s0n7765,s1n7765,notn7765;
or (n7765,s0n7765,s1n7765);
not(notn7765,n4903);
and (s0n7765,notn7765,n7766);
and (s1n7765,n4903,1'b0);
wire s0n7766,s1n7766,notn7766;
or (n7766,s0n7766,s1n7766);
not(notn7766,n4777);
and (s0n7766,notn7766,n7767);
and (s1n7766,n4777,1'b1);
wire s0n7767,s1n7767,notn7767;
or (n7767,s0n7767,s1n7767);
not(notn7767,n1102);
and (s0n7767,notn7767,n7642);
and (s1n7767,n1102,n7768);
wire s0n7768,s1n7768,notn7768;
or (n7768,s0n7768,s1n7768);
not(notn7768,n1102);
and (s0n7768,notn7768,n7769);
and (s1n7768,n1102,n7770);
xor (n7769,n4896,n4898);
xor (n7770,n4896,n4902);
and (n7771,n7772,n6);
wire s0n7772,s1n7772,notn7772;
or (n7772,s0n7772,s1n7772);
not(notn7772,n1194);
and (s0n7772,notn7772,1'b0);
and (s1n7772,n1194,n7765);
and (n7773,n7765,n4929);
and (n7774,n7775,n7029);
wire s0n7775,s1n7775,notn7775;
or (n7775,s0n7775,s1n7775);
not(notn7775,n7024);
and (s0n7775,notn7775,n7776);
and (s1n7775,n7024,1'b0);
wire s0n7776,s1n7776,notn7776;
or (n7776,s0n7776,s1n7776);
not(notn7776,n6998);
and (s0n7776,notn7776,n7777);
and (s1n7776,n6998,1'b1);
wire s0n7777,s1n7777,notn7777;
or (n7777,s0n7777,s1n7777);
not(notn7777,n6991);
and (s0n7777,notn7777,1'b0);
and (s1n7777,n6991,n7778);
xor (n7778,n7021,n7023);
not (n7779,n7780);
or (n7780,1'b0,n7781,n7784,n7787,n7788);
and (n7781,n7782,n1189);
wire s0n7782,s1n7782,notn7782;
or (n7782,s0n7782,s1n7782);
not(notn7782,n4923);
and (s0n7782,notn7782,1'b0);
and (s1n7782,n4923,n7783);
and (n7784,n7785,n6);
wire s0n7785,s1n7785,notn7785;
or (n7785,s0n7785,s1n7785);
not(notn7785,n1194);
and (s0n7785,notn7785,1'b0);
and (s1n7785,n1194,n7786);
and (n7787,n7775,n7040);
or (n7788,1'b0,n7789,n7809,n7829,n7849);
and (n7789,n7790,n1331);
or (n7790,1'b0,n7791,n7797,n7803);
and (n7791,n7792,n7050);
or (n7792,1'b0,n7793,n7794,n7795,n7796);
and (n7793,n2454,n1187);
and (n7794,n2442,n1186);
and (n7795,n2444,n1183);
and (n7796,n2451,n817);
and (n7797,n7798,n7030);
or (n7798,1'b0,n7799,n7800,n7801,n7802);
and (n7799,n2404,n1187);
and (n7800,n2407,n1186);
and (n7801,n2409,n1183);
and (n7802,n2411,n817);
and (n7803,n7804,n7063);
or (n7804,1'b0,n7805,n7806,n7807,n7808);
and (n7805,n2407,n1187);
and (n7806,n2409,n1186);
and (n7807,n2411,n1183);
and (n7808,n2391,n817);
and (n7809,n7810,n1316);
or (n7810,1'b0,n7811,n7817,n7823);
and (n7811,n7812,n7050);
or (n7812,1'b0,n7813,n7814,n7815,n7816);
and (n7813,n2470,n1187);
and (n7814,n2459,n1186);
and (n7815,n2461,n1183);
and (n7816,n2467,n817);
and (n7817,n7818,n7030);
or (n7818,1'b0,n7819,n7820,n7821,n7822);
and (n7819,n2391,n1187);
and (n7820,n2395,n1186);
and (n7821,n2397,n1183);
and (n7822,n2399,n817);
and (n7823,n7824,n7063);
or (n7824,1'b0,n7825,n7826,n7827,n7828);
and (n7825,n2395,n1187);
and (n7826,n2397,n1186);
and (n7827,n2399,n1183);
and (n7828,n2393,n817);
and (n7829,n7830,n1265);
or (n7830,1'b0,n7831,n7837,n7843);
and (n7831,n7832,n7050);
or (n7832,1'b0,n7833,n7834,n7835,n7836);
and (n7833,n2475,n1187);
and (n7834,n2479,n1186);
and (n7835,n2482,n1183);
and (n7836,n2485,n817);
and (n7837,n7838,n7030);
or (n7838,1'b0,n7839,n7840,n7841,n7842);
and (n7839,n2422,n1187);
and (n7840,n2424,n1186);
and (n7841,n2429,n1183);
and (n7842,n2434,n817);
and (n7843,n7844,n7063);
or (n7844,1'b0,n7845,n7846,n7847,n7848);
and (n7845,n2424,n1187);
and (n7846,n2429,n1186);
and (n7847,n2434,n1183);
and (n7848,n2414,n817);
and (n7849,n7850,n1246);
or (n7850,1'b0,n7851,n7857,n7863);
and (n7851,n7852,n7050);
or (n7852,1'b0,n7853,n7854,n7855,n7856);
and (n7853,n2490,n1187);
and (n7854,n2493,n1186);
and (n7855,n2496,n1183);
and (n7856,n2499,n817);
and (n7857,n7858,n7030);
or (n7858,1'b0,n7859,n7860,n7861,n7862);
and (n7859,n2414,n1187);
and (n7860,n2420,n1186);
and (n7861,n2427,n1183);
and (n7862,n2432,n817);
and (n7863,n7864,n7063);
or (n7864,1'b0,n7865,n7866,n7867,n7868);
and (n7865,n2420,n1187);
and (n7866,n2427,n1186);
and (n7867,n2432,n1183);
and (n7868,n2418,n817);
and (n7869,n7870,n7888);
not (n7870,n7871);
or (n7871,1'b0,n7872,n7880,n7882,n7883);
and (n7872,n7873,n1189);
wire s0n7873,s1n7873,notn7873;
or (n7873,s0n7873,s1n7873);
not(notn7873,n4923);
and (s0n7873,notn7873,1'b0);
and (s1n7873,n4923,n7874);
wire s0n7874,s1n7874,notn7874;
or (n7874,s0n7874,s1n7874);
not(notn7874,n4903);
and (s0n7874,notn7874,n7875);
and (s1n7874,n4903,1'b0);
wire s0n7875,s1n7875,notn7875;
or (n7875,s0n7875,s1n7875);
not(notn7875,n4777);
and (s0n7875,notn7875,n7876);
and (s1n7875,n4777,1'b1);
wire s0n7876,s1n7876,notn7876;
or (n7876,s0n7876,s1n7876);
not(notn7876,n1102);
and (s0n7876,notn7876,n7359);
and (s1n7876,n1102,n7877);
wire s0n7877,s1n7877,notn7877;
or (n7877,s0n7877,s1n7877);
not(notn7877,n1102);
and (s0n7877,notn7877,n7878);
and (s1n7877,n1102,n7879);
xor (n7878,n4890,n4895);
xor (n7879,n4890,n4901);
and (n7880,n7881,n6);
wire s0n7881,s1n7881,notn7881;
or (n7881,s0n7881,s1n7881);
not(notn7881,n1194);
and (s0n7881,notn7881,1'b0);
and (s1n7881,n1194,n7874);
and (n7882,n7874,n4929);
and (n7883,n7884,n7029);
wire s0n7884,s1n7884,notn7884;
or (n7884,s0n7884,s1n7884);
not(notn7884,n7024);
and (s0n7884,notn7884,n7885);
and (s1n7884,n7024,1'b0);
wire s0n7885,s1n7885,notn7885;
or (n7885,s0n7885,s1n7885);
not(notn7885,n6998);
and (s0n7885,notn7885,n7886);
and (s1n7885,n6998,1'b1);
wire s0n7886,s1n7886,notn7886;
or (n7886,s0n7886,s1n7886);
not(notn7886,n6991);
and (s0n7886,notn7886,1'b0);
and (s1n7886,n6991,n7887);
xor (n7887,n7017,n7020);
not (n7888,n7889);
or (n7889,1'b0,n7890,n7893,n7896,n7897);
and (n7890,n7891,n1189);
wire s0n7891,s1n7891,notn7891;
or (n7891,s0n7891,s1n7891);
not(notn7891,n4923);
and (s0n7891,notn7891,1'b0);
and (s1n7891,n4923,n7892);
and (n7893,n7894,n6);
wire s0n7894,s1n7894,notn7894;
or (n7894,s0n7894,s1n7894);
not(notn7894,n1194);
and (s0n7894,notn7894,1'b0);
and (s1n7894,n1194,n7895);
and (n7896,n7884,n7040);
or (n7897,1'b0,n7898,n7918,n7938,n7958);
and (n7898,n7899,n1331);
or (n7899,1'b0,n7900,n7906,n7912);
and (n7900,n7901,n7050);
or (n7901,1'b0,n7902,n7903,n7904,n7905);
and (n7902,n2365,n1187);
and (n7903,n2367,n1186);
and (n7904,n2369,n1183);
and (n7905,n2349,n817);
and (n7906,n7907,n7030);
or (n7907,1'b0,n7908,n7909,n7910,n7911);
and (n7908,n2298,n1187);
and (n7909,n2301,n1186);
and (n7910,n2303,n1183);
and (n7911,n2305,n817);
and (n7912,n7913,n7063);
or (n7913,1'b0,n7914,n7915,n7916,n7917);
and (n7914,n2301,n1187);
and (n7915,n2303,n1186);
and (n7916,n2305,n1183);
and (n7917,n2285,n817);
and (n7918,n7919,n1316);
or (n7919,1'b0,n7920,n7926,n7932);
and (n7920,n7921,n7050);
or (n7921,1'b0,n7922,n7923,n7924,n7925);
and (n7922,n2353,n1187);
and (n7923,n2355,n1186);
and (n7924,n2357,n1183);
and (n7925,n2351,n817);
and (n7926,n7927,n7030);
or (n7927,1'b0,n7928,n7929,n7930,n7931);
and (n7928,n2285,n1187);
and (n7929,n2289,n1186);
and (n7930,n2291,n1183);
and (n7931,n2293,n817);
and (n7932,n7933,n7063);
or (n7933,1'b0,n7934,n7935,n7936,n7937);
and (n7934,n2289,n1187);
and (n7935,n2291,n1186);
and (n7936,n2293,n1183);
and (n7937,n2287,n817);
and (n7938,n7939,n1265);
or (n7939,1'b0,n7940,n7946,n7952);
and (n7940,n7941,n7050);
or (n7941,1'b0,n7942,n7943,n7944,n7945);
and (n7942,n2339,n1187);
and (n7943,n2374,n1186);
and (n7944,n2379,n1183);
and (n7945,n2343,n817);
and (n7946,n7947,n7030);
or (n7947,1'b0,n7948,n7949,n7950,n7951);
and (n7948,n2315,n1187);
and (n7949,n2311,n1186);
and (n7950,n2320,n1183);
and (n7951,n2322,n817);
and (n7952,n7953,n7063);
or (n7953,1'b0,n7954,n7955,n7956,n7957);
and (n7954,n2311,n1187);
and (n7955,n2320,n1186);
and (n7956,n2322,n1183);
and (n7957,n2308,n817);
and (n7958,n7959,n1246);
or (n7959,1'b0,n7960,n7966,n7972);
and (n7960,n7961,n7050);
or (n7961,1'b0,n7962,n7963,n7964,n7965);
and (n7962,n2335,n1187);
and (n7963,n2372,n1186);
and (n7964,n2377,n1183);
and (n7965,n2337,n817);
and (n7966,n7967,n7030);
or (n7967,1'b0,n7968,n7969,n7970,n7971);
and (n7968,n2308,n1187);
and (n7969,n2313,n1186);
and (n7970,n2325,n1183);
and (n7971,n2327,n817);
and (n7972,n7973,n7063);
or (n7973,1'b0,n7974,n7975,n7976,n7977);
and (n7974,n2313,n1187);
and (n7975,n2325,n1186);
and (n7976,n2327,n1183);
and (n7977,n2317,n817);
nand (n7978,n7979,n7982);
or (n7979,n7869,n7980);
not (n7980,n7981);
and (n7981,n7780,n7762);
not (n7982,n7983);
and (n7983,n7889,n7871);
and (n7984,n7467,n7985);
nand (n7985,n7986,n1180);
or (n7986,n7541,n653);
nor (n7987,n7988,n7995);
and (n7988,n7874,n7989);
and (n7989,n7990,n805);
nand (n7990,n7991,n7993);
or (n7991,n4925,n7992);
not (n7992,n1105);
not (n7993,n7994);
nor (n7994,n653,n1344,n7,n1107);
and (n7995,n7884,n7996);
nor (n7996,n653,n726,n7,n1191);
nor (n7997,n7998,n8114);
wire s0n7998,s1n7998,notn7998;
or (n7998,s0n7998,s1n7998);
not(notn7998,n8111);
and (s0n7998,notn7998,n7999);
and (s1n7998,n8111,n8106);
wire s0n7999,s1n7999,notn7999;
or (n7999,s0n7999,s1n7999);
not(notn7999,n8008);
and (s0n7999,notn7999,1'b0);
and (s1n7999,n8008,n8000);
wire s0n8000,s1n8000,notn8000;
or (n8000,s0n8000,s1n8000);
not(notn8000,n31);
and (s0n8000,notn8000,n8001);
and (s1n8000,n31,n8007);
or (n8001,1'b0,n8002,n8003,n8004,n8005);
and (n8002,n2317,n1187);
and (n8003,n6481,n1186);
and (n8004,n1262,n1183);
and (n8005,n8006,n817);
wire s0n8007,s1n8007,notn8007;
or (n8007,s0n8007,s1n8007);
not(notn8007,n806);
and (s0n8007,notn8007,1'b0);
and (s1n8007,n806,n8006);
and (n8008,n8009,n8058);
and (n8009,n601,n8010);
nor (n8010,n10,n1109,n8011);
wire s0n8011,s1n8011,notn8011;
or (n8011,s0n8011,s1n8011);
not(notn8011,n601);
and (s0n8011,notn8011,1'b0);
and (s1n8011,n601,n8012);
wire s0n8012,s1n8012,notn8012;
or (n8012,s0n8012,s1n8012);
not(notn8012,n600);
and (s0n8012,notn8012,n8013);
and (s1n8012,n600,n8049);
or (n8013,n8014,n8025,n8036,n8047);
and (n8014,n8015,n37);
wire s0n8015,s1n8015,notn8015;
or (n8015,s0n8015,s1n8015);
not(notn8015,n31);
and (s0n8015,notn8015,n8016);
and (s1n8015,n31,n8017);
or (n8017,n8018,n8020,n8022,n8024);
and (n8018,n8019,n19);
and (n8020,n8021,n24);
and (n8022,n8023,n28);
and (n8024,n8016,n30);
and (n8025,n8026,n42);
wire s0n8026,s1n8026,notn8026;
or (n8026,s0n8026,s1n8026);
not(notn8026,n31);
and (s0n8026,notn8026,n8027);
and (s1n8026,n31,n8028);
or (n8028,n8029,n8031,n8033,n8035);
and (n8029,n8030,n19);
and (n8031,n8032,n24);
and (n8033,n8034,n28);
and (n8035,n8027,n30);
and (n8036,n8037,n47);
wire s0n8037,s1n8037,notn8037;
or (n8037,s0n8037,s1n8037);
not(notn8037,n31);
and (s0n8037,notn8037,n8038);
and (s1n8037,n31,n8039);
or (n8039,n8040,n8042,n8044,n8046);
and (n8040,n8041,n19);
and (n8042,n8043,n24);
and (n8044,n8045,n28);
and (n8046,n8038,n30);
and (n8047,n8048,n50);
wire s0n8048,s1n8048,notn8048;
or (n8048,s0n8048,s1n8048);
not(notn8048,n31);
and (s0n8048,notn8048,n8049);
and (s1n8048,n31,n8050);
or (n8050,n8051,n8053,n8055,n8057);
and (n8051,n8052,n19);
and (n8053,n8054,n24);
and (n8055,n8056,n28);
and (n8057,n8049,n30);
nor (n8058,n655,n728,n8059);
wire s0n8059,s1n8059,notn8059;
or (n8059,s0n8059,s1n8059);
not(notn8059,n601);
and (s0n8059,notn8059,1'b0);
and (s1n8059,n601,n8060);
wire s0n8060,s1n8060,notn8060;
or (n8060,s0n8060,s1n8060);
not(notn8060,n600);
and (s0n8060,notn8060,n8061);
and (s1n8060,n600,n8097);
or (n8061,n8062,n8073,n8084,n8095);
and (n8062,n8063,n37);
wire s0n8063,s1n8063,notn8063;
or (n8063,s0n8063,s1n8063);
not(notn8063,n31);
and (s0n8063,notn8063,n8064);
and (s1n8063,n31,n8065);
or (n8065,n8066,n8068,n8070,n8072);
and (n8066,n8067,n19);
and (n8068,n8069,n24);
and (n8070,n8071,n28);
and (n8072,n8064,n30);
and (n8073,n8074,n42);
wire s0n8074,s1n8074,notn8074;
or (n8074,s0n8074,s1n8074);
not(notn8074,n31);
and (s0n8074,notn8074,n8075);
and (s1n8074,n31,n8076);
or (n8076,n8077,n8079,n8081,n8083);
and (n8077,n8078,n19);
and (n8079,n8080,n24);
and (n8081,n8082,n28);
and (n8083,n8075,n30);
and (n8084,n8085,n47);
wire s0n8085,s1n8085,notn8085;
or (n8085,s0n8085,s1n8085);
not(notn8085,n31);
and (s0n8085,notn8085,n8086);
and (s1n8085,n31,n8087);
or (n8087,n8088,n8090,n8092,n8094);
and (n8088,n8089,n19);
and (n8090,n8091,n24);
and (n8092,n8093,n28);
and (n8094,n8086,n30);
and (n8095,n8096,n50);
wire s0n8096,s1n8096,notn8096;
or (n8096,s0n8096,s1n8096);
not(notn8096,n31);
and (s0n8096,notn8096,n8097);
and (s1n8096,n31,n8098);
or (n8098,n8099,n8101,n8103,n8105);
and (n8099,n8100,n19);
and (n8101,n8102,n24);
and (n8103,n8104,n28);
and (n8105,n8097,n30);
or (n8106,1'b0,n8107,n8108,n8109,n8110);
and (n8107,n7913,n1331);
and (n8108,n7933,n1316);
and (n8109,n7953,n1265);
and (n8110,n7973,n1246);
and (n8111,n651,n8112);
not (n8112,n8113);
or (n8113,n653,n726,n7,n1107);
and (n8114,n8115,n9976);
nand (n8115,n8116,n9947);
not (n8116,n8117);
or (n8117,n8118,n9946);
and (n8118,n8119,n9471);
xor (n8119,n8120,n9398);
xor (n8120,n8121,n9335);
xor (n8121,n8122,n9304);
or (n8122,n8123,n9303);
and (n8123,n8124,n9109);
xor (n8124,n8125,n9064);
xor (n8125,n8126,n8918);
xor (n8126,n8127,n8511);
xor (n8127,n8128,n8505);
xor (n8128,n8129,n8323);
wire s0n8129,s1n8129,notn8129;
or (n8129,s0n8129,s1n8129);
not(notn8129,n8320);
and (s0n8129,notn8129,1'b0);
and (s1n8129,n8320,n8130);
xor (n8130,n8131,n8140);
wire s0n8131,s1n8131,notn8131;
or (n8131,s0n8131,s1n8131);
not(notn8131,n8010);
and (s0n8131,notn8131,1'b0);
and (s1n8131,n8010,n8132);
nand (n8132,n8133,n8138);
or (n8133,n8134,n8135);
not (n8134,n8006);
not (n8135,n8136);
and (n8136,n8137,n601);
nor (n8137,n1063,n1225);
nand (n8138,n8139,n8001);
and (n8139,n1063,n601);
or (n8140,n8141,n8261,n8319);
and (n8141,n8142,n8160);
xor (n8142,n8143,n8154);
wire s0n8143,s1n8143,notn8143;
or (n8143,s0n8143,s1n8143);
not(notn8143,n8010);
and (s0n8143,notn8143,1'b0);
and (s1n8143,n8010,n8144);
nand (n8144,n8145,n8148);
or (n8145,n8146,n8135);
not (n8146,n8147);
nand (n8148,n8139,n8149);
or (n8149,1'b0,n8150,n8151,n8152,n8153);
and (n8150,n2418,n1187);
and (n8151,n6511,n1186);
and (n8152,n1415,n1183);
and (n8153,n8147,n817);
wire s0n8154,s1n8154,notn8154;
or (n8154,s0n8154,s1n8154);
not(notn8154,n8155);
and (s0n8154,notn8154,1'b0);
and (s1n8154,n8155,n8132);
xor (n8155,n8156,n8157);
not (n8156,n8011);
and (n8157,n8158,n8159);
not (n8158,n1109);
not (n8159,n10);
and (n8160,n8161,n8163);
wire s0n8161,s1n8161,notn8161;
or (n8161,s0n8161,s1n8161);
not(notn8161,n8162);
and (s0n8161,notn8161,1'b0);
and (s1n8161,n8162,n8132);
xor (n8162,n8158,n8159);
or (n8163,n8164,n8167,n8260);
and (n8164,n8165,n8166);
wire s0n8165,s1n8165,notn8165;
or (n8165,s0n8165,s1n8165);
not(notn8165,n8162);
and (s0n8165,notn8165,1'b0);
and (s1n8165,n8162,n8144);
wire s0n8166,s1n8166,notn8166;
or (n8166,s0n8166,s1n8166);
not(notn8166,n10);
and (s0n8166,notn8166,1'b0);
and (s1n8166,n10,n8132);
and (n8167,n8166,n8168);
or (n8168,n8169,n8182,n8259);
and (n8169,n8170,n8181);
wire s0n8170,s1n8170,notn8170;
or (n8170,s0n8170,s1n8170);
not(notn8170,n8162);
and (s0n8170,notn8170,1'b0);
and (s1n8170,n8162,n8171);
nand (n8171,n8172,n8175);
or (n8172,n8173,n8135);
not (n8173,n8174);
nand (n8175,n8139,n8176);
or (n8176,1'b0,n8177,n8178,n8179,n8180);
and (n8177,n2515,n1187);
and (n8178,n6560,n1186);
and (n8179,n1587,n1183);
and (n8180,n8174,n817);
wire s0n8181,s1n8181,notn8181;
or (n8181,s0n8181,s1n8181);
not(notn8181,n10);
and (s0n8181,notn8181,1'b0);
and (s1n8181,n10,n8144);
and (n8182,n8181,n8183);
or (n8183,n8184,n8197,n8258);
and (n8184,n8185,n8196);
wire s0n8185,s1n8185,notn8185;
or (n8185,s0n8185,s1n8185);
not(notn8185,n8162);
and (s0n8185,notn8185,1'b0);
and (s1n8185,n8162,n8186);
nand (n8186,n8187,n8190);
or (n8187,n8188,n8135);
not (n8188,n8189);
nand (n8190,n8139,n8191);
or (n8191,1'b0,n8192,n8193,n8194,n8195);
and (n8192,n2675,n1187);
and (n8193,n6601,n1186);
and (n8194,n1664,n1183);
and (n8195,n8189,n817);
wire s0n8196,s1n8196,notn8196;
or (n8196,s0n8196,s1n8196);
not(notn8196,n10);
and (s0n8196,notn8196,1'b0);
and (s1n8196,n10,n8171);
and (n8197,n8196,n8198);
or (n8198,n8199,n8212,n8257);
and (n8199,n8200,n8211);
wire s0n8200,s1n8200,notn8200;
or (n8200,s0n8200,s1n8200);
not(notn8200,n8162);
and (s0n8200,notn8200,1'b0);
and (s1n8200,n8162,n8201);
nand (n8201,n8202,n8205);
or (n8202,n8203,n8135);
not (n8203,n8204);
nand (n8205,n8139,n8206);
or (n8206,1'b0,n8207,n8208,n8209,n8210);
and (n8207,n2803,n1187);
and (n8208,n6663,n1186);
and (n8209,n1826,n1183);
and (n8210,n8204,n817);
wire s0n8211,s1n8211,notn8211;
or (n8211,s0n8211,s1n8211);
not(notn8211,n10);
and (s0n8211,notn8211,1'b0);
and (s1n8211,n10,n8186);
and (n8212,n8211,n8213);
or (n8213,n8214,n8227,n8229);
and (n8214,n8215,n8226);
wire s0n8215,s1n8215,notn8215;
or (n8215,s0n8215,s1n8215);
not(notn8215,n8162);
and (s0n8215,notn8215,1'b0);
and (s1n8215,n8162,n8216);
nand (n8216,n8217,n8220);
or (n8217,n8218,n8135);
not (n8218,n8219);
nand (n8220,n8139,n8221);
or (n8221,1'b0,n8222,n8223,n8224,n8225);
and (n8222,n2920,n1187);
and (n8223,n6715,n1186);
and (n8224,n1950,n1183);
and (n8225,n8219,n817);
wire s0n8226,s1n8226,notn8226;
or (n8226,s0n8226,s1n8226);
not(notn8226,n10);
and (s0n8226,notn8226,1'b0);
and (s1n8226,n10,n8201);
and (n8227,n8226,n8228);
or (n8228,n8229,n8242,n8243);
and (n8229,n8230,n8241);
wire s0n8230,s1n8230,notn8230;
or (n8230,s0n8230,s1n8230);
not(notn8230,n8162);
and (s0n8230,notn8230,1'b0);
and (s1n8230,n8162,n8231);
nand (n8231,n8232,n8235);
or (n8232,n8233,n8135);
not (n8233,n8234);
nand (n8235,n8139,n8236);
or (n8236,1'b0,n8237,n8238,n8239,n8240);
and (n8237,n3040,n1187);
and (n8238,n6768,n1186);
and (n8239,n2073,n1183);
and (n8240,n8234,n817);
wire s0n8241,s1n8241,notn8241;
or (n8241,s0n8241,s1n8241);
not(notn8241,n10);
and (s0n8241,notn8241,1'b0);
and (s1n8241,n10,n8216);
and (n8242,n8241,n8243);
and (n8243,n8244,n8256);
wire s0n8244,s1n8244,notn8244;
or (n8244,s0n8244,s1n8244);
not(notn8244,n8162);
and (s0n8244,notn8244,1'b0);
and (s1n8244,n8162,n8245);
nand (n8245,n8246,n8255);
or (n8246,n8247,n8254);
not (n8247,n8248);
or (n8248,1'b0,n8249,n8250,n8251,n8252);
and (n8249,n3163,n1187);
and (n8250,n6829,n1186);
and (n8251,n2193,n1183);
and (n8252,n8253,n817);
not (n8254,n8139);
nand (n8255,n8136,n8253);
wire s0n8256,s1n8256,notn8256;
or (n8256,s0n8256,s1n8256);
not(notn8256,n10);
and (s0n8256,notn8256,1'b0);
and (s1n8256,n10,n8231);
and (n8257,n8200,n8213);
and (n8258,n8185,n8198);
and (n8259,n8170,n8183);
and (n8260,n8165,n8168);
and (n8261,n8160,n8262);
or (n8262,n8263,n8268,n8318);
and (n8263,n8264,n8267);
xor (n8264,n8265,n8266);
wire s0n8265,s1n8265,notn8265;
or (n8265,s0n8265,s1n8265);
not(notn8265,n8010);
and (s0n8265,notn8265,1'b0);
and (s1n8265,n8010,n8171);
wire s0n8266,s1n8266,notn8266;
or (n8266,s0n8266,s1n8266);
not(notn8266,n8155);
and (s0n8266,notn8266,1'b0);
and (s1n8266,n8155,n8144);
xor (n8267,n8161,n8163);
and (n8268,n8267,n8269);
or (n8269,n8270,n8276,n8317);
and (n8270,n8271,n8274);
xor (n8271,n8272,n8273);
wire s0n8272,s1n8272,notn8272;
or (n8272,s0n8272,s1n8272);
not(notn8272,n8010);
and (s0n8272,notn8272,1'b0);
and (s1n8272,n8010,n8186);
wire s0n8273,s1n8273,notn8273;
or (n8273,s0n8273,s1n8273);
not(notn8273,n8155);
and (s0n8273,notn8273,1'b0);
and (s1n8273,n8155,n8171);
xor (n8274,n8275,n8168);
xor (n8275,n8165,n8166);
and (n8276,n8274,n8277);
or (n8277,n8278,n8284,n8316);
and (n8278,n8279,n8282);
xor (n8279,n8280,n8281);
wire s0n8280,s1n8280,notn8280;
or (n8280,s0n8280,s1n8280);
not(notn8280,n8010);
and (s0n8280,notn8280,1'b0);
and (s1n8280,n8010,n8201);
wire s0n8281,s1n8281,notn8281;
or (n8281,s0n8281,s1n8281);
not(notn8281,n8155);
and (s0n8281,notn8281,1'b0);
and (s1n8281,n8155,n8186);
xor (n8282,n8283,n8183);
xor (n8283,n8170,n8181);
and (n8284,n8282,n8285);
or (n8285,n8286,n8292,n8315);
and (n8286,n8287,n8290);
xor (n8287,n8288,n8289);
wire s0n8288,s1n8288,notn8288;
or (n8288,s0n8288,s1n8288);
not(notn8288,n8010);
and (s0n8288,notn8288,1'b0);
and (s1n8288,n8010,n8216);
wire s0n8289,s1n8289,notn8289;
or (n8289,s0n8289,s1n8289);
not(notn8289,n8155);
and (s0n8289,notn8289,1'b0);
and (s1n8289,n8155,n8201);
xor (n8290,n8291,n8198);
xor (n8291,n8185,n8196);
and (n8292,n8290,n8293);
or (n8293,n8294,n8300,n8314);
and (n8294,n8295,n8298);
xor (n8295,n8296,n8297);
wire s0n8296,s1n8296,notn8296;
or (n8296,s0n8296,s1n8296);
not(notn8296,n8010);
and (s0n8296,notn8296,1'b0);
and (s1n8296,n8010,n8231);
wire s0n8297,s1n8297,notn8297;
or (n8297,s0n8297,s1n8297);
not(notn8297,n8155);
and (s0n8297,notn8297,1'b0);
and (s1n8297,n8155,n8216);
xor (n8298,n8299,n8213);
xor (n8299,n8200,n8211);
and (n8300,n8298,n8301);
or (n8301,n8302,n8308,n8313);
and (n8302,n8303,n8306);
xor (n8303,n8304,n8305);
wire s0n8304,s1n8304,notn8304;
or (n8304,s0n8304,s1n8304);
not(notn8304,n8010);
and (s0n8304,notn8304,1'b0);
and (s1n8304,n8010,n8245);
wire s0n8305,s1n8305,notn8305;
or (n8305,s0n8305,s1n8305);
not(notn8305,n8155);
and (s0n8305,notn8305,1'b0);
and (s1n8305,n8155,n8231);
xor (n8306,n8307,n8228);
xor (n8307,n8215,n8226);
and (n8308,n8306,n8309);
and (n8309,n8310,n8311);
wire s0n8310,s1n8310,notn8310;
or (n8310,s0n8310,s1n8310);
not(notn8310,n8155);
and (s0n8310,notn8310,1'b0);
and (s1n8310,n8155,n8245);
xor (n8311,n8312,n8243);
xor (n8312,n8230,n8241);
and (n8313,n8303,n8309);
and (n8314,n8295,n8301);
and (n8315,n8287,n8293);
and (n8316,n8279,n8285);
and (n8317,n8271,n8277);
and (n8318,n8264,n8269);
and (n8319,n8142,n8262);
xor (n8320,n8321,n8322);
not (n8321,n728);
not (n8322,n655);
wire s0n8323,s1n8323,notn8323;
or (n8323,s0n8323,s1n8323);
not(notn8323,n8059);
and (s0n8323,notn8323,1'b0);
and (s1n8323,n8059,n8324);
xor (n8324,n8325,n8448);
xor (n8325,n8326,n8349);
xor (n8326,n8327,n8338);
wire s0n8327,s1n8327,notn8327;
or (n8327,s0n8327,s1n8327);
not(notn8327,n8010);
and (s0n8327,notn8327,1'b0);
and (s1n8327,n8010,n8328);
nand (n8328,n8329,n8332);
or (n8329,n8330,n8135);
not (n8330,n8331);
nand (n8332,n8139,n8333);
or (n8333,1'b0,n8334,n8335,n8336,n8337);
and (n8334,n2499,n1187);
and (n8335,n6516,n1186);
and (n8336,n3287,n1183);
and (n8337,n8331,n817);
wire s0n8338,s1n8338,notn8338;
or (n8338,s0n8338,s1n8338);
not(notn8338,n8155);
and (s0n8338,notn8338,1'b0);
and (s1n8338,n8155,n8339);
nand (n8339,n8340,n8343);
or (n8340,n8341,n8135);
not (n8341,n8342);
nand (n8343,n8139,n8344);
or (n8344,1'b0,n8345,n8346,n8347,n8348);
and (n8345,n2337,n1187);
and (n8346,n6470,n1186);
and (n8347,n3355,n1183);
and (n8348,n8342,n817);
and (n8349,n8350,n8351);
wire s0n8350,s1n8350,notn8350;
or (n8350,s0n8350,s1n8350);
not(notn8350,n8162);
and (s0n8350,notn8350,1'b0);
and (s1n8350,n8162,n8339);
or (n8351,n8352,n8355,n8447);
and (n8352,n8353,n8354);
wire s0n8353,s1n8353,notn8353;
or (n8353,s0n8353,s1n8353);
not(notn8353,n8162);
and (s0n8353,notn8353,1'b0);
and (s1n8353,n8162,n8328);
wire s0n8354,s1n8354,notn8354;
or (n8354,s0n8354,s1n8354);
not(notn8354,n10);
and (s0n8354,notn8354,1'b0);
and (s1n8354,n10,n8339);
and (n8355,n8354,n8356);
or (n8356,n8357,n8370,n8446);
and (n8357,n8358,n8369);
wire s0n8358,s1n8358,notn8358;
or (n8358,s0n8358,s1n8358);
not(notn8358,n8162);
and (s0n8358,notn8358,1'b0);
and (s1n8358,n8162,n8359);
nand (n8359,n8360,n8363);
or (n8360,n8361,n8135);
not (n8361,n8362);
nand (n8363,n8139,n8364);
or (n8364,1'b0,n8365,n8366,n8367,n8368);
and (n8365,n2569,n1187);
and (n8366,n6550,n1186);
and (n8367,n3727,n1183);
and (n8368,n8362,n817);
wire s0n8369,s1n8369,notn8369;
or (n8369,s0n8369,s1n8369);
not(notn8369,n10);
and (s0n8369,notn8369,1'b0);
and (s1n8369,n10,n8328);
and (n8370,n8369,n8371);
or (n8371,n8372,n8385,n8445);
and (n8372,n8373,n8384);
wire s0n8373,s1n8373,notn8373;
or (n8373,s0n8373,s1n8373);
not(notn8373,n8162);
and (s0n8373,notn8373,1'b0);
and (s1n8373,n8162,n8374);
nand (n8374,n8375,n8378);
or (n8375,n8376,n8135);
not (n8376,n8377);
nand (n8378,n8139,n8379);
or (n8379,1'b0,n8380,n8381,n8382,n8383);
and (n8380,n2735,n1187);
and (n8381,n6609,n1186);
and (n8382,n3794,n1183);
and (n8383,n8377,n817);
wire s0n8384,s1n8384,notn8384;
or (n8384,s0n8384,s1n8384);
not(notn8384,n10);
and (s0n8384,notn8384,1'b0);
and (s1n8384,n10,n8359);
and (n8385,n8384,n8386);
or (n8386,n8387,n8400,n8444);
and (n8387,n8388,n8399);
wire s0n8388,s1n8388,notn8388;
or (n8388,s0n8388,s1n8388);
not(notn8388,n8162);
and (s0n8388,notn8388,1'b0);
and (s1n8388,n8162,n8389);
nand (n8389,n8390,n8393);
or (n8390,n8391,n8135);
not (n8391,n8392);
nand (n8393,n8139,n8394);
or (n8394,1'b0,n8395,n8396,n8397,n8398);
and (n8395,n2860,n1187);
and (n8396,n6652,n1186);
and (n8397,n3654,n1183);
and (n8398,n8392,n817);
wire s0n8399,s1n8399,notn8399;
or (n8399,s0n8399,s1n8399);
not(notn8399,n10);
and (s0n8399,notn8399,1'b0);
and (s1n8399,n10,n8374);
and (n8400,n8399,n8401);
or (n8401,n8402,n8415,n8417);
and (n8402,n8403,n8414);
wire s0n8403,s1n8403,notn8403;
or (n8403,s0n8403,s1n8403);
not(notn8403,n8162);
and (s0n8403,notn8403,1'b0);
and (s1n8403,n8162,n8404);
nand (n8404,n8405,n8413);
or (n8405,n8406,n8254);
not (n8406,n8407);
or (n8407,1'b0,n8408,n8409,n8410,n8411);
and (n8408,n2977,n1187);
and (n8409,n6705,n1186);
and (n8410,n3445,n1183);
and (n8411,n8412,n817);
nand (n8413,n8136,n8412);
wire s0n8414,s1n8414,notn8414;
or (n8414,s0n8414,s1n8414);
not(notn8414,n10);
and (s0n8414,notn8414,1'b0);
and (s1n8414,n10,n8389);
and (n8415,n8414,n8416);
or (n8416,n8417,n8430,n8431);
and (n8417,n8418,n8429);
wire s0n8418,s1n8418,notn8418;
or (n8418,s0n8418,s1n8418);
not(notn8418,n8162);
and (s0n8418,notn8418,1'b0);
and (s1n8418,n8162,n8419);
nand (n8419,n8420,n8428);
or (n8420,n8421,n8254);
not (n8421,n8422);
or (n8422,1'b0,n8423,n8424,n8425,n8426);
and (n8423,n3101,n1187);
and (n8424,n6758,n1186);
and (n8425,n3512,n1183);
and (n8426,n8427,n817);
nand (n8428,n8136,n8427);
wire s0n8429,s1n8429,notn8429;
or (n8429,s0n8429,s1n8429);
not(notn8429,n10);
and (s0n8429,notn8429,1'b0);
and (s1n8429,n10,n8404);
and (n8430,n8429,n8431);
and (n8431,n8432,n8443);
wire s0n8432,s1n8432,notn8432;
or (n8432,s0n8432,s1n8432);
not(notn8432,n8162);
and (s0n8432,notn8432,1'b0);
and (s1n8432,n8162,n8433);
nand (n8433,n8434,n8437);
or (n8434,n8435,n8135);
not (n8435,n8436);
nand (n8437,n8139,n8438);
or (n8438,1'b0,n8439,n8440,n8441,n8442);
and (n8439,n3226,n1187);
and (n8440,n6819,n1186);
and (n8441,n3581,n1183);
and (n8442,n8436,n817);
wire s0n8443,s1n8443,notn8443;
or (n8443,s0n8443,s1n8443);
not(notn8443,n10);
and (s0n8443,notn8443,1'b0);
and (s1n8443,n10,n8419);
and (n8444,n8388,n8401);
and (n8445,n8373,n8386);
and (n8446,n8358,n8371);
and (n8447,n8353,n8356);
or (n8448,n8449,n8454,n8504);
and (n8449,n8450,n8453);
xor (n8450,n8451,n8452);
wire s0n8451,s1n8451,notn8451;
or (n8451,s0n8451,s1n8451);
not(notn8451,n8010);
and (s0n8451,notn8451,1'b0);
and (s1n8451,n8010,n8359);
wire s0n8452,s1n8452,notn8452;
or (n8452,s0n8452,s1n8452);
not(notn8452,n8155);
and (s0n8452,notn8452,1'b0);
and (s1n8452,n8155,n8328);
xor (n8453,n8350,n8351);
and (n8454,n8453,n8455);
or (n8455,n8456,n8462,n8503);
and (n8456,n8457,n8460);
xor (n8457,n8458,n8459);
wire s0n8458,s1n8458,notn8458;
or (n8458,s0n8458,s1n8458);
not(notn8458,n8010);
and (s0n8458,notn8458,1'b0);
and (s1n8458,n8010,n8374);
wire s0n8459,s1n8459,notn8459;
or (n8459,s0n8459,s1n8459);
not(notn8459,n8155);
and (s0n8459,notn8459,1'b0);
and (s1n8459,n8155,n8359);
xor (n8460,n8461,n8356);
xor (n8461,n8353,n8354);
and (n8462,n8460,n8463);
or (n8463,n8464,n8470,n8502);
and (n8464,n8465,n8468);
xor (n8465,n8466,n8467);
wire s0n8466,s1n8466,notn8466;
or (n8466,s0n8466,s1n8466);
not(notn8466,n8010);
and (s0n8466,notn8466,1'b0);
and (s1n8466,n8010,n8389);
wire s0n8467,s1n8467,notn8467;
or (n8467,s0n8467,s1n8467);
not(notn8467,n8155);
and (s0n8467,notn8467,1'b0);
and (s1n8467,n8155,n8374);
xor (n8468,n8469,n8371);
xor (n8469,n8358,n8369);
and (n8470,n8468,n8471);
or (n8471,n8472,n8478,n8501);
and (n8472,n8473,n8476);
xor (n8473,n8474,n8475);
wire s0n8474,s1n8474,notn8474;
or (n8474,s0n8474,s1n8474);
not(notn8474,n8010);
and (s0n8474,notn8474,1'b0);
and (s1n8474,n8010,n8404);
wire s0n8475,s1n8475,notn8475;
or (n8475,s0n8475,s1n8475);
not(notn8475,n8155);
and (s0n8475,notn8475,1'b0);
and (s1n8475,n8155,n8389);
xor (n8476,n8477,n8386);
xor (n8477,n8373,n8384);
and (n8478,n8476,n8479);
or (n8479,n8480,n8486,n8500);
and (n8480,n8481,n8484);
xor (n8481,n8482,n8483);
wire s0n8482,s1n8482,notn8482;
or (n8482,s0n8482,s1n8482);
not(notn8482,n8010);
and (s0n8482,notn8482,1'b0);
and (s1n8482,n8010,n8419);
wire s0n8483,s1n8483,notn8483;
or (n8483,s0n8483,s1n8483);
not(notn8483,n8155);
and (s0n8483,notn8483,1'b0);
and (s1n8483,n8155,n8404);
xor (n8484,n8485,n8401);
xor (n8485,n8388,n8399);
and (n8486,n8484,n8487);
or (n8487,n8488,n8494,n8499);
and (n8488,n8489,n8492);
xor (n8489,n8490,n8491);
wire s0n8490,s1n8490,notn8490;
or (n8490,s0n8490,s1n8490);
not(notn8490,n8010);
and (s0n8490,notn8490,1'b0);
and (s1n8490,n8010,n8433);
wire s0n8491,s1n8491,notn8491;
or (n8491,s0n8491,s1n8491);
not(notn8491,n8155);
and (s0n8491,notn8491,1'b0);
and (s1n8491,n8155,n8419);
xor (n8492,n8493,n8416);
xor (n8493,n8403,n8414);
and (n8494,n8492,n8495);
and (n8495,n8496,n8497);
wire s0n8496,s1n8496,notn8496;
or (n8496,s0n8496,s1n8496);
not(notn8496,n8155);
and (s0n8496,notn8496,1'b0);
and (s1n8496,n8155,n8433);
xor (n8497,n8498,n8431);
xor (n8498,n8418,n8429);
and (n8499,n8489,n8495);
and (n8500,n8481,n8487);
and (n8501,n8473,n8479);
and (n8502,n8465,n8471);
and (n8503,n8457,n8463);
and (n8504,n8450,n8455);
wire s0n8505,s1n8505,notn8505;
or (n8505,s0n8505,s1n8505);
not(notn8505,n8508);
and (s0n8505,notn8505,1'b0);
and (s1n8505,n8508,n8506);
xor (n8506,n8507,n8262);
xor (n8507,n8142,n8160);
xor (n8508,n8509,n8510);
not (n8509,n8059);
and (n8510,n8321,n8322);
xor (n8511,n8512,n8907);
xor (n8512,n8513,n8891);
or (n8513,n8514,n8890);
and (n8514,n8515,n8758);
xor (n8515,n8516,n8746);
and (n8516,n8517,n8730);
xor (n8517,n8518,n8650);
wire s0n8518,s1n8518,notn8518;
or (n8518,s0n8518,s1n8518);
not(notn8518,n8058);
and (s0n8518,notn8518,1'b0);
and (s1n8518,n8058,n8519);
xor (n8519,n8520,n8622);
xor (n8520,n8521,n8533);
not (n8521,n8522);
nand (n8522,n8011,n8523);
nand (n8523,n8524,n8532);
or (n8524,n8525,n8254);
not (n8525,n8526);
or (n8526,1'b0,n8527,n8528,n8529,n8530);
and (n8527,n2672,n1187);
and (n8528,n5983,n1186);
and (n8529,n1704,n1183);
and (n8530,n8531,n817);
nand (n8532,n8136,n8531);
xor (n8533,n8534,n8557);
xor (n8534,n8535,n8546);
wire s0n8535,s1n8535,notn8535;
or (n8535,s0n8535,s1n8535);
not(notn8535,n1109);
and (s0n8535,notn8535,1'b0);
and (s1n8535,n1109,n8536);
nand (n8536,n8537,n8545);
or (n8537,n8538,n8254);
not (n8538,n8539);
or (n8539,1'b0,n8540,n8541,n8542,n8543);
and (n8540,n2553,n1187);
and (n8541,n5893,n1186);
and (n8542,n1584,n1183);
and (n8543,n8544,n817);
nand (n8545,n8136,n8544);
wire s0n8546,s1n8546,notn8546;
or (n8546,s0n8546,s1n8546);
not(notn8546,n10);
and (s0n8546,notn8546,1'b0);
and (s1n8546,n10,n8547);
nand (n8547,n8548,n8551);
or (n8548,n8549,n8135);
not (n8549,n8550);
nand (n8551,n8139,n8552);
or (n8552,1'b0,n8553,n8554,n8555,n8556);
and (n8553,n2432,n1187);
and (n8554,n5827,n1186);
and (n8555,n1456,n1183);
and (n8556,n8550,n817);
or (n8557,n8558,n8561,n8621);
and (n8558,n8559,n8560);
wire s0n8559,s1n8559,notn8559;
or (n8559,s0n8559,s1n8559);
not(notn8559,n1109);
and (s0n8559,notn8559,1'b0);
and (s1n8559,n1109,n8523);
wire s0n8560,s1n8560,notn8560;
or (n8560,s0n8560,s1n8560);
not(notn8560,n10);
and (s0n8560,notn8560,1'b0);
and (s1n8560,n10,n8536);
and (n8561,n8560,n8562);
or (n8562,n8563,n8576,n8620);
and (n8563,n8564,n8575);
wire s0n8564,s1n8564,notn8564;
or (n8564,s0n8564,s1n8564);
not(notn8564,n1109);
and (s0n8564,notn8564,1'b0);
and (s1n8564,n1109,n8565);
nand (n8565,n8566,n8569);
or (n8566,n8567,n8135);
not (n8567,n8568);
nand (n8569,n8139,n8570);
or (n8570,1'b0,n8571,n8572,n8573,n8574);
and (n8571,n2800,n1187);
and (n8572,n6062,n1186);
and (n8573,n1823,n1183);
and (n8574,n8568,n817);
wire s0n8575,s1n8575,notn8575;
or (n8575,s0n8575,s1n8575);
not(notn8575,n10);
and (s0n8575,notn8575,1'b0);
and (s1n8575,n10,n8523);
and (n8576,n8575,n8577);
or (n8577,n8578,n8591,n8593);
and (n8578,n8579,n8590);
wire s0n8579,s1n8579,notn8579;
or (n8579,s0n8579,s1n8579);
not(notn8579,n1109);
and (s0n8579,notn8579,1'b0);
and (s1n8579,n1109,n8580);
nand (n8580,n8581,n8589);
or (n8581,n8582,n8254);
not (n8582,n8583);
or (n8583,1'b0,n8584,n8585,n8586,n8587);
and (n8584,n2917,n1187);
and (n8585,n6102,n1186);
and (n8586,n1947,n1183);
and (n8587,n8588,n817);
nand (n8589,n8136,n8588);
wire s0n8590,s1n8590,notn8590;
or (n8590,s0n8590,s1n8590);
not(notn8590,n10);
and (s0n8590,notn8590,1'b0);
and (s1n8590,n10,n8565);
and (n8591,n8590,n8592);
or (n8592,n8593,n8606,n8607);
and (n8593,n8594,n8605);
wire s0n8594,s1n8594,notn8594;
or (n8594,s0n8594,s1n8594);
not(notn8594,n1109);
and (s0n8594,notn8594,1'b0);
and (s1n8594,n1109,n8595);
nand (n8595,n8596,n8599);
or (n8596,n8597,n8135);
not (n8597,n8598);
nand (n8599,n8139,n8600);
or (n8600,1'b0,n8601,n8602,n8603,n8604);
and (n8601,n3037,n1187);
and (n8602,n6201,n1186);
and (n8603,n2070,n1183);
and (n8604,n8598,n817);
wire s0n8605,s1n8605,notn8605;
or (n8605,s0n8605,s1n8605);
not(notn8605,n10);
and (s0n8605,notn8605,1'b0);
and (s1n8605,n10,n8580);
and (n8606,n8605,n8607);
and (n8607,n8608,n8619);
wire s0n8608,s1n8608,notn8608;
or (n8608,s0n8608,s1n8608);
not(notn8608,n1109);
and (s0n8608,notn8608,1'b0);
and (s1n8608,n1109,n8609);
nand (n8609,n8610,n8613);
or (n8610,n8611,n8135);
not (n8611,n8612);
nand (n8613,n8139,n8614);
or (n8614,1'b0,n8615,n8616,n8617,n8618);
and (n8615,n3160,n1187);
and (n8616,n6273,n1186);
and (n8617,n2190,n1183);
and (n8618,n8612,n817);
wire s0n8619,s1n8619,notn8619;
or (n8619,s0n8619,s1n8619);
not(notn8619,n10);
and (s0n8619,notn8619,1'b0);
and (s1n8619,n10,n8595);
and (n8620,n8564,n8577);
and (n8621,n8559,n8562);
or (n8622,n8623,n8628,n8649);
and (n8623,n8624,n8626);
not (n8624,n8625);
nand (n8625,n8011,n8565);
xor (n8626,n8627,n8562);
xor (n8627,n8559,n8560);
and (n8628,n8626,n8629);
or (n8629,n8630,n8635,n8648);
and (n8630,n8631,n8633);
not (n8631,n8632);
nand (n8632,n8011,n8580);
xor (n8633,n8634,n8577);
xor (n8634,n8564,n8575);
and (n8635,n8633,n8636);
or (n8636,n8637,n8642,n8647);
and (n8637,n8638,n8640);
not (n8638,n8639);
nand (n8639,n8011,n8595);
xor (n8640,n8641,n8592);
xor (n8641,n8579,n8590);
and (n8642,n8640,n8643);
and (n8643,n8644,n8645);
and (n8644,n8011,n8609);
xor (n8645,n8646,n8607);
xor (n8646,n8594,n8605);
and (n8647,n8638,n8643);
and (n8648,n8631,n8636);
and (n8649,n8624,n8629);
xor (n8650,n8651,n8692);
xor (n8651,n8652,n8680);
xor (n8652,n8653,n8678);
xor (n8653,n8654,n8666);
nor (n8654,n8655,n8322);
nand (n8655,n8011,n8656);
nand (n8656,n8657,n8665);
or (n8657,n8658,n8254);
not (n8658,n8659);
or (n8659,1'b0,n8660,n8661,n8662,n8663);
and (n8660,n2377,n1187);
and (n8661,n5733,n1186);
and (n8662,n3352,n1183);
and (n8663,n8664,n817);
nand (n8665,n8136,n8664);
and (n8666,n8667,n655);
and (n8667,n8011,n8668);
nand (n8668,n8669,n8672);
or (n8669,n8670,n8135);
not (n8670,n8671);
nand (n8672,n8139,n8673);
or (n8673,1'b0,n8674,n8675,n8676,n8677);
and (n8674,n2327,n1187);
and (n8675,n5732,n1186);
and (n8676,n1301,n1183);
and (n8677,n8671,n817);
and (n8678,n8666,n8679);
wire s0n8679,s1n8679,notn8679;
or (n8679,s0n8679,s1n8679);
not(notn8679,n1109);
and (s0n8679,notn8679,1'b0);
and (s1n8679,n1109,n8547);
and (n8680,n8654,n8681);
wire s0n8681,s1n8681,notn8681;
or (n8681,s0n8681,s1n8681);
not(notn8681,n1109);
and (s0n8681,notn8681,1'b0);
and (s1n8681,n1109,n8682);
nand (n8682,n8683,n8691);
or (n8683,n8684,n8254);
not (n8684,n8685);
or (n8685,1'b0,n8686,n8687,n8688,n8689);
and (n8686,n2496,n1187);
and (n8687,n5828,n1186);
and (n8688,n3284,n1183);
and (n8689,n8690,n817);
nand (n8691,n8136,n8690);
or (n8692,n8693,n8729);
and (n8693,n8694,n8708);
xor (n8694,n8695,n8700);
nor (n8695,n8696,n8322);
xnor (n8696,n8697,n8698);
nand (n8697,n8011,n8682);
not (n8698,n8699);
wire s0n8699,s1n8699,notn8699;
or (n8699,s0n8699,s1n8699);
not(notn8699,n1109);
and (s0n8699,notn8699,1'b0);
and (s1n8699,n1109,n8656);
and (n8700,n8701,n655);
nand (n8701,n8702,n8707);
or (n8702,n8703,n8705);
not (n8703,n8704);
wire s0n8704,s1n8704,notn8704;
or (n8704,s0n8704,s1n8704);
not(notn8704,n1109);
and (s0n8704,notn8704,1'b0);
and (s1n8704,n1109,n8668);
not (n8705,n8706);
nand (n8706,n8011,n8547);
or (n8707,n8706,n8704);
and (n8708,n8709,n655);
or (n8709,n8710,n8726);
nor (n8710,n8711,n8725);
and (n8711,n8712,n8723);
nand (n8712,n8011,n8713);
nand (n8713,n8714,n8722);
or (n8714,n8715,n8254);
not (n8715,n8716);
or (n8716,1'b0,n8717,n8718,n8719,n8720);
and (n8717,n2607,n1187);
and (n8718,n5894,n1186);
and (n8719,n3724,n1183);
and (n8720,n8721,n817);
nand (n8722,n8136,n8721);
not (n8723,n8724);
wire s0n8724,s1n8724,notn8724;
or (n8724,s0n8724,s1n8724);
not(notn8724,n10);
and (s0n8724,notn8724,1'b0);
and (s1n8724,n10,n8656);
not (n8725,n8681);
nor (n8726,n8727,n8655);
not (n8727,n8728);
wire s0n8728,s1n8728,notn8728;
or (n8728,s0n8728,s1n8728);
not(notn8728,n10);
and (s0n8728,notn8728,1'b0);
and (s1n8728,n10,n8713);
and (n8729,n8695,n8700);
wire s0n8730,s1n8730,notn8730;
or (n8730,s0n8730,s1n8730);
not(notn8730,n8508);
and (s0n8730,notn8730,1'b0);
and (s1n8730,n8508,n8731);
xor (n8731,n8732,n8742);
xor (n8732,n8733,n8735);
not (n8733,n8734);
nand (n8734,n8011,n8536);
xor (n8735,n8736,n8738);
xor (n8736,n8679,n8737);
wire s0n8737,s1n8737,notn8737;
or (n8737,s0n8737,s1n8737);
not(notn8737,n10);
and (s0n8737,notn8737,1'b0);
and (s1n8737,n10,n8668);
or (n8738,n8739,n8740,n8741);
and (n8739,n8535,n8546);
and (n8740,n8546,n8557);
and (n8741,n8535,n8557);
or (n8742,n8743,n8744,n8745);
and (n8743,n8521,n8533);
and (n8744,n8533,n8622);
and (n8745,n8521,n8622);
wire s0n8746,s1n8746,notn8746;
or (n8746,s0n8746,s1n8746);
not(notn8746,n8508);
and (s0n8746,notn8746,1'b0);
and (s1n8746,n8508,n8747);
xor (n8747,n8748,n8754);
xor (n8748,n8705,n8749);
xor (n8749,n8704,n8750);
or (n8750,n8751,n8752,n8753);
and (n8751,n8679,n8737);
and (n8752,n8737,n8738);
and (n8753,n8679,n8738);
or (n8754,n8755,n8756,n8757);
and (n8755,n8733,n8735);
and (n8756,n8735,n8742);
and (n8757,n8733,n8742);
wire s0n8758,s1n8758,notn8758;
or (n8758,s0n8758,s1n8758);
not(notn8758,n8059);
and (s0n8758,notn8758,1'b0);
and (s1n8758,n8059,n8759);
xor (n8759,n8760,n8847);
xor (n8760,n8761,n8762);
not (n8761,n8697);
xor (n8762,n8699,n8763);
or (n8763,n8764,n8765,n8846);
and (n8764,n8681,n8724);
and (n8765,n8724,n8766);
or (n8766,n8767,n8770,n8845);
and (n8767,n8768,n8769);
wire s0n8768,s1n8768,notn8768;
or (n8768,s0n8768,s1n8768);
not(notn8768,n1109);
and (s0n8768,notn8768,1'b0);
and (s1n8768,n1109,n8713);
wire s0n8769,s1n8769,notn8769;
or (n8769,s0n8769,s1n8769);
not(notn8769,n10);
and (s0n8769,notn8769,1'b0);
and (s1n8769,n10,n8682);
and (n8770,n8769,n8771);
or (n8771,n8772,n8784,n8844);
and (n8772,n8773,n8728);
wire s0n8773,s1n8773,notn8773;
or (n8773,s0n8773,s1n8773);
not(notn8773,n1109);
and (s0n8773,notn8773,1'b0);
and (s1n8773,n1109,n8774);
nand (n8774,n8775,n8783);
or (n8775,n8776,n8254);
not (n8776,n8777);
or (n8777,1'b0,n8778,n8779,n8780,n8781);
and (n8778,n2732,n1187);
and (n8779,n5984,n1186);
and (n8780,n3791,n1183);
and (n8781,n8782,n817);
nand (n8783,n8136,n8782);
and (n8784,n8728,n8785);
or (n8785,n8786,n8799,n8843);
and (n8786,n8787,n8798);
wire s0n8787,s1n8787,notn8787;
or (n8787,s0n8787,s1n8787);
not(notn8787,n1109);
and (s0n8787,notn8787,1'b0);
and (s1n8787,n1109,n8788);
nand (n8788,n8789,n8797);
or (n8789,n8790,n8254);
not (n8790,n8791);
or (n8791,1'b0,n8792,n8793,n8794,n8795);
and (n8792,n2857,n1187);
and (n8793,n6063,n1186);
and (n8794,n3651,n1183);
and (n8795,n8796,n817);
nand (n8797,n8136,n8796);
wire s0n8798,s1n8798,notn8798;
or (n8798,s0n8798,s1n8798);
not(notn8798,n10);
and (s0n8798,notn8798,1'b0);
and (s1n8798,n10,n8774);
and (n8799,n8798,n8800);
or (n8800,n8801,n8814,n8816);
and (n8801,n8802,n8813);
wire s0n8802,s1n8802,notn8802;
or (n8802,s0n8802,s1n8802);
not(notn8802,n1109);
and (s0n8802,notn8802,1'b0);
and (s1n8802,n1109,n8803);
nand (n8803,n8804,n8807);
or (n8804,n8805,n8135);
not (n8805,n8806);
nand (n8807,n8139,n8808);
or (n8808,1'b0,n8809,n8810,n8811,n8812);
and (n8809,n2974,n1187);
and (n8810,n6103,n1186);
and (n8811,n3442,n1183);
and (n8812,n8806,n817);
wire s0n8813,s1n8813,notn8813;
or (n8813,s0n8813,s1n8813);
not(notn8813,n10);
and (s0n8813,notn8813,1'b0);
and (s1n8813,n10,n8788);
and (n8814,n8813,n8815);
or (n8815,n8816,n8829,n8830);
and (n8816,n8817,n8828);
wire s0n8817,s1n8817,notn8817;
or (n8817,s0n8817,s1n8817);
not(notn8817,n1109);
and (s0n8817,notn8817,1'b0);
and (s1n8817,n1109,n8818);
nand (n8818,n8819,n8827);
or (n8819,n8820,n8254);
not (n8820,n8821);
or (n8821,1'b0,n8822,n8823,n8824,n8825);
and (n8822,n3098,n1187);
and (n8823,n6202,n1186);
and (n8824,n3509,n1183);
and (n8825,n8826,n817);
nand (n8827,n8136,n8826);
wire s0n8828,s1n8828,notn8828;
or (n8828,s0n8828,s1n8828);
not(notn8828,n10);
and (s0n8828,notn8828,1'b0);
and (s1n8828,n10,n8803);
and (n8829,n8828,n8830);
and (n8830,n8831,n8842);
wire s0n8831,s1n8831,notn8831;
or (n8831,s0n8831,s1n8831);
not(notn8831,n1109);
and (s0n8831,notn8831,1'b0);
and (s1n8831,n1109,n8832);
nand (n8832,n8833,n8841);
or (n8833,n8834,n8254);
not (n8834,n8835);
or (n8835,1'b0,n8836,n8837,n8838,n8839);
and (n8836,n3223,n1187);
and (n8837,n6274,n1186);
and (n8838,n3578,n1183);
and (n8839,n8840,n817);
nand (n8841,n8136,n8840);
wire s0n8842,s1n8842,notn8842;
or (n8842,s0n8842,s1n8842);
not(notn8842,n10);
and (s0n8842,notn8842,1'b0);
and (s1n8842,n10,n8818);
and (n8843,n8787,n8800);
and (n8844,n8773,n8785);
and (n8845,n8768,n8771);
and (n8846,n8681,n8766);
or (n8847,n8848,n8852,n8889);
and (n8848,n8849,n8850);
not (n8849,n8712);
xor (n8850,n8851,n8766);
xor (n8851,n8681,n8724);
and (n8852,n8850,n8853);
or (n8853,n8854,n8859,n8888);
and (n8854,n8855,n8857);
not (n8855,n8856);
nand (n8856,n8011,n8774);
xor (n8857,n8858,n8771);
xor (n8858,n8768,n8769);
and (n8859,n8857,n8860);
or (n8860,n8861,n8865,n8887);
and (n8861,n8862,n8863);
and (n8862,n8011,n8788);
xor (n8863,n8864,n8785);
xor (n8864,n8773,n8728);
and (n8865,n8863,n8866);
or (n8866,n8867,n8872,n8886);
and (n8867,n8868,n8870);
not (n8868,n8869);
nand (n8869,n8011,n8803);
xor (n8870,n8871,n8800);
xor (n8871,n8787,n8798);
and (n8872,n8870,n8873);
or (n8873,n8874,n8879,n8885);
and (n8874,n8875,n8877);
not (n8875,n8876);
nand (n8876,n8011,n8818);
xor (n8877,n8878,n8815);
xor (n8878,n8802,n8813);
and (n8879,n8877,n8880);
and (n8880,n8881,n8883);
not (n8881,n8882);
nand (n8882,n8011,n8832);
xor (n8883,n8884,n8830);
xor (n8884,n8817,n8828);
and (n8885,n8875,n8880);
and (n8886,n8868,n8873);
and (n8887,n8862,n8866);
and (n8888,n8855,n8860);
and (n8889,n8849,n8853);
and (n8890,n8516,n8746);
xor (n8891,n8892,n8904);
xor (n8892,n8893,n8903);
wire s0n8893,s1n8893,notn8893;
or (n8893,s0n8893,s1n8893);
not(notn8893,n8320);
and (s0n8893,notn8893,1'b0);
and (s1n8893,n8320,n8894);
or (n8894,n8895,n8897,n8902);
and (n8895,n8667,n8896);
and (n8896,n8704,n8750);
and (n8897,n8896,n8898);
or (n8898,n8899,n8900,n8901);
and (n8899,n8705,n8749);
and (n8900,n8749,n8754);
and (n8901,n8705,n8754);
and (n8902,n8667,n8898);
wire s0n8903,s1n8903,notn8903;
or (n8903,s0n8903,s1n8903);
not(notn8903,n8058);
and (s0n8903,notn8903,1'b0);
and (s1n8903,n8058,n8747);
wire s0n8904,s1n8904,notn8904;
or (n8904,s0n8904,s1n8904);
not(notn8904,n8508);
and (s0n8904,notn8904,1'b0);
and (s1n8904,n8508,n8905);
xor (n8905,n8906,n8898);
xor (n8906,n8667,n8896);
wire s0n8907,s1n8907,notn8907;
or (n8907,s0n8907,s1n8907);
not(notn8907,n728);
and (s0n8907,notn8907,1'b0);
and (s1n8907,n728,n8908);
or (n8908,n8909,n8912,n8917);
and (n8909,n8910,n8911);
not (n8910,n8655);
and (n8911,n8699,n8763);
and (n8912,n8911,n8913);
or (n8913,n8914,n8915,n8916);
and (n8914,n8761,n8762);
and (n8915,n8762,n8847);
and (n8916,n8761,n8847);
and (n8917,n8910,n8913);
or (n8918,n8919,n9063);
and (n8919,n8920,n8984);
xor (n8920,n8921,n8983);
or (n8921,n8922,n8982);
and (n8922,n8923,n8930);
xor (n8923,n8924,n8927);
wire s0n8924,s1n8924,notn8924;
or (n8924,s0n8924,s1n8924);
not(notn8924,n728);
and (s0n8924,notn8924,1'b0);
and (s1n8924,n728,n8925);
xor (n8925,n8926,n8455);
xor (n8926,n8450,n8453);
wire s0n8927,s1n8927,notn8927;
or (n8927,s0n8927,s1n8927);
not(notn8927,n8059);
and (s0n8927,notn8927,1'b0);
and (s1n8927,n8059,n8928);
xor (n8928,n8929,n8463);
xor (n8929,n8457,n8460);
and (n8930,n8931,n8508);
xor (n8931,n8932,n8944);
nor (n8932,n8933,n8943);
not (n8933,n8934);
or (n8934,n8935,n8938);
xor (n8935,n8936,n8169);
xor (n8936,n8273,n8937);
xor (n8937,n8275,n8272);
or (n8938,n8939,n8942);
and (n8939,n8940,n8184);
xor (n8940,n8281,n8941);
xor (n8941,n8283,n8280);
and (n8942,n8281,n8941);
and (n8943,n8935,n8938);
nand (n8944,n8945,n8981);
or (n8945,n8946,n8954);
not (n8946,n8947);
or (n8947,n8948,n8949);
xor (n8948,n8940,n8184);
or (n8949,n8950,n8953);
and (n8950,n8951,n8199);
xor (n8951,n8289,n8952);
xor (n8952,n8291,n8288);
and (n8953,n8289,n8952);
not (n8954,n8955);
nand (n8955,n8956,n8977,n8980);
nand (n8956,n8957,n8964,n8974);
or (n8957,n8958,n8959);
xor (n8958,n8951,n8199);
or (n8959,n8960,n8963);
and (n8960,n8961,n8962);
xor (n8961,n8297,n8214);
xor (n8962,n8299,n8296);
and (n8963,n8297,n8214);
or (n8964,n8965,n8973);
and (n8965,n8966,n8971);
xor (n8966,n8229,n8967);
or (n8967,n8968,n8970);
and (n8968,n8969,n8312);
xor (n8969,n8243,n8310);
and (n8970,n8243,n8310);
xor (n8971,n8972,n8305);
xor (n8972,n8304,n8307);
and (n8973,n8229,n8967);
or (n8974,n8975,n8976);
xor (n8975,n8961,n8962);
and (n8976,n8972,n8305);
nand (n8977,n8978,n8957);
not (n8978,n8979);
nand (n8979,n8975,n8976);
nand (n8980,n8958,n8959);
nand (n8981,n8948,n8949);
and (n8982,n8924,n8927);
xor (n8983,n8515,n8758);
and (n8984,n8985,n9060);
xor (n8985,n8986,n8989);
and (n8986,n8987,n8058);
xnor (n8987,n8955,n8988);
nand (n8988,n8947,n8981);
or (n8989,n8990,n9059);
and (n8990,n8991,n9027);
xor (n8991,n8992,n8995);
wire s0n8992,s1n8992,notn8992;
or (n8992,s0n8992,s1n8992);
not(notn8992,n8059);
and (s0n8992,notn8992,1'b0);
and (s1n8992,n8059,n8993);
xor (n8993,n8994,n8860);
xor (n8994,n8855,n8857);
and (n8995,n8996,n9021);
or (n8996,n8997,n9020);
and (n8997,n8998,n9012);
xor (n8998,n8999,n9006);
and (n8999,n9000,n655);
nand (n9000,n9001,n9003,n9005);
or (n9001,n9002,n8712);
not (n9002,n8813);
or (n9003,n8856,n9004);
not (n9004,n8787);
not (n9005,n8772);
nor (n9006,n8322,n9007);
nor (n9007,n8558,n9008);
nor (n9008,n9009,n8625);
and (n9009,n9010,n9011);
not (n9010,n8560);
not (n9011,n8559);
nor (n9012,n9013,n8322);
nor (n9013,n9014,n9018);
and (n9014,n9015,n8535);
not (n9015,n9016);
xor (n9016,n8522,n9017);
not (n9017,n8546);
and (n9018,n9016,n9019);
not (n9019,n8535);
and (n9020,n8999,n9006);
and (n9021,n9022,n655);
nor (n9022,n9023,n9025);
and (n9023,n9024,n8681);
xor (n9024,n8712,n8723);
and (n9025,n9026,n8725);
not (n9026,n9024);
or (n9027,n9028,n9058);
and (n9028,n9029,n9055);
xor (n9029,n9030,n9033);
wire s0n9030,s1n9030,notn9030;
or (n9030,s0n9030,s1n9030);
not(notn9030,n8508);
and (s0n9030,notn9030,1'b0);
and (s1n9030,n8508,n9031);
xor (n9031,n9032,n8629);
xor (n9032,n8624,n8626);
xor (n9033,n9034,n9047);
xor (n9034,n9035,n9040);
and (n9035,n9036,n655);
nand (n9036,n9037,n9038,n9039);
or (n9037,n8734,n9011);
not (n9038,n8739);
or (n9039,n8522,n9017);
and (n9040,n9041,n655);
nand (n9041,n9042,n9046);
or (n9042,n9043,n8856);
and (n9043,n9044,n9045);
not (n9044,n8768);
not (n9045,n8769);
not (n9046,n8767);
and (n9047,n9048,n655);
nor (n9048,n9049,n9052);
and (n9049,n9050,n8679);
xor (n9050,n9051,n8734);
not (n9051,n8737);
and (n9052,n9053,n9054);
not (n9053,n9050);
not (n9054,n8679);
wire s0n9055,s1n9055,notn9055;
or (n9055,s0n9055,s1n9055);
not(notn9055,n8059);
and (s0n9055,notn9055,1'b0);
and (s1n9055,n8059,n9056);
xor (n9056,n9057,n8866);
xor (n9057,n8862,n8863);
and (n9058,n9030,n9033);
and (n9059,n8992,n8995);
wire s0n9060,s1n9060,notn9060;
or (n9060,s0n9060,s1n9060);
not(notn9060,n8320);
and (s0n9060,notn9060,1'b0);
and (s1n9060,n8320,n9061);
xor (n9061,n9062,n8269);
xor (n9062,n8264,n8267);
and (n9063,n8921,n8983);
xor (n9064,n9065,n9096);
xor (n9065,n9066,n9079);
xor (n9066,n9067,n9076);
xor (n9067,n9068,n9069);
wire s0n9068,s1n9068,notn9068;
or (n9068,s0n9068,s1n9068);
not(notn9068,n8058);
and (s0n9068,notn9068,1'b0);
and (s1n9068,n8058,n9061);
and (n9069,n9070,n9073);
or (n9070,n9071,n9072);
and (n9071,n8651,n8692);
and (n9072,n8652,n8680);
or (n9073,n9074,n9075);
and (n9074,n8653,n8678);
and (n9075,n8654,n8666);
wire s0n9076,s1n9076,notn9076;
or (n9076,s0n9076,s1n9076);
not(notn9076,n8059);
and (s0n9076,notn9076,1'b0);
and (s1n9076,n8059,n9077);
xor (n9077,n9078,n8913);
xor (n9078,n8910,n8911);
or (n9079,n9080,n9095);
and (n9080,n9081,n9094);
xor (n9081,n9082,n9093);
or (n9082,n9083,n9092);
and (n9083,n9084,n9091);
xor (n9084,n9085,n9086);
xor (n9085,n8517,n8730);
and (n9086,n9087,n9090);
xor (n9087,n9088,n9089);
wire s0n9088,s1n9088,notn9088;
or (n9088,s0n9088,s1n9088);
not(notn9088,n8058);
and (s0n9088,notn9088,1'b0);
and (s1n9088,n8058,n9031);
wire s0n9089,s1n9089,notn9089;
or (n9089,s0n9089,s1n9089);
not(notn9089,n8508);
and (s0n9089,notn9089,1'b0);
and (s1n9089,n8508,n8519);
wire s0n9090,s1n9090,notn9090;
or (n9090,s0n9090,s1n9090);
not(notn9090,n8320);
and (s0n9090,notn9090,1'b0);
and (s1n9090,n8320,n8731);
wire s0n9091,s1n9091,notn9091;
or (n9091,s0n9091,s1n9091);
not(notn9091,n728);
and (s0n9091,notn9091,1'b0);
and (s1n9091,n728,n8759);
and (n9092,n9085,n9086);
wire s0n9093,s1n9093,notn9093;
or (n9093,s0n9093,s1n9093);
not(notn9093,n8059);
and (s0n9093,notn9093,1'b0);
and (s1n9093,n8059,n8925);
wire s0n9094,s1n9094,notn9094;
or (n9094,s0n9094,s1n9094);
not(notn9094,n8508);
and (s0n9094,notn9094,1'b0);
and (s1n9094,n8508,n9061);
and (n9095,n9082,n9093);
or (n9096,n9097,n9108);
and (n9097,n9098,n9107);
xor (n9098,n9099,n9100);
wire s0n9099,s1n9099,notn9099;
or (n9099,s0n9099,s1n9099);
not(notn9099,n655);
and (s0n9099,notn9099,1'b0);
and (s1n9099,n655,n8130);
wire s0n9100,s1n9100,notn9100;
or (n9100,s0n9100,s1n9100);
not(notn9100,n655);
and (s0n9100,notn9100,1'b0);
and (s1n9100,n655,n9101);
xor (n9101,n9102,n9103);
wire s0n9102,s1n9102,notn9102;
or (n9102,s0n9102,s1n9102);
not(notn9102,n8010);
and (s0n9102,notn9102,1'b0);
and (s1n9102,n8010,n8339);
or (n9103,n9104,n9105,n9106);
and (n9104,n8326,n8349);
and (n9105,n8349,n8448);
and (n9106,n8326,n8448);
wire s0n9107,s1n9107,notn9107;
or (n9107,s0n9107,s1n9107);
not(notn9107,n8320);
and (s0n9107,notn9107,1'b0);
and (s1n9107,n8320,n8506);
and (n9108,n9099,n9100);
or (n9109,n9110,n9302);
and (n9110,n9111,n9152);
xor (n9111,n9112,n9113);
xor (n9112,n8920,n8984);
or (n9113,n9114,n9151);
and (n9114,n9115,n9124);
xor (n9115,n9116,n9117);
xor (n9116,n8985,n9060);
or (n9117,n9118,n9123);
and (n9118,n9119,n9122);
xor (n9119,n9120,n9121);
and (n9120,n8987,n8508);
xor (n9121,n8991,n9027);
wire s0n9122,s1n9122,notn9122;
or (n9122,s0n9122,s1n9122);
not(notn9122,n655);
and (s0n9122,notn9122,1'b0);
and (s1n9122,n655,n8925);
and (n9123,n9120,n9121);
or (n9124,n9125,n9150);
and (n9125,n9126,n9149);
xor (n9126,n9127,n9128);
wire s0n9127,s1n9127,notn9127;
or (n9127,s0n9127,s1n9127);
not(notn9127,n728);
and (s0n9127,notn9127,1'b0);
and (s1n9127,n728,n8928);
or (n9128,n9129,n9148);
and (n9129,n9130,n9145);
xor (n9130,n9131,n9136);
xor (n9131,n9132,n9133);
xor (n9132,n8996,n9021);
wire s0n9133,s1n9133,notn9133;
or (n9133,s0n9133,s1n9133);
not(notn9133,n8058);
and (s0n9133,notn9133,1'b0);
and (s1n9133,n8058,n9134);
xor (n9134,n9135,n8636);
xor (n9135,n8631,n8633);
and (n9136,n9137,n9142);
xor (n9137,n9138,n9139);
xor (n9138,n8998,n9012);
wire s0n9139,s1n9139,notn9139;
or (n9139,s0n9139,s1n9139);
not(notn9139,n8058);
and (s0n9139,notn9139,1'b0);
and (s1n9139,n8058,n9140);
xor (n9140,n9141,n8643);
xor (n9141,n8638,n8640);
wire s0n9142,s1n9142,notn9142;
or (n9142,s0n9142,s1n9142);
not(notn9142,n8059);
and (s0n9142,notn9142,1'b0);
and (s1n9142,n8059,n9143);
xor (n9143,n9144,n8873);
xor (n9144,n8868,n8870);
wire s0n9145,s1n9145,notn9145;
or (n9145,s0n9145,s1n9145);
not(notn9145,n8058);
and (s0n9145,notn9145,1'b0);
and (s1n9145,n8058,n9146);
xor (n9146,n9147,n8301);
xor (n9147,n8295,n8298);
and (n9148,n9131,n9136);
and (n9149,n8931,n8320);
and (n9150,n9127,n9128);
and (n9151,n9116,n9117);
or (n9152,n9153,n9301);
and (n9153,n9154,n9277);
xor (n9154,n9155,n9276);
or (n9155,n9156,n9275);
and (n9156,n9157,n9274);
xor (n9157,n9158,n9191);
or (n9158,n9159,n9190);
and (n9159,n9160,n9187);
xor (n9160,n9161,n9162);
xor (n9161,n9029,n9055);
or (n9162,n9163,n9186);
and (n9163,n9164,n9185);
xor (n9164,n9165,n9166);
wire s0n9165,s1n9165,notn9165;
or (n9165,s0n9165,s1n9165);
not(notn9165,n8320);
and (s0n9165,notn9165,1'b0);
and (s1n9165,n8320,n9031);
or (n9166,n9167,n9184);
and (n9167,n9168,n9183);
xor (n9168,n9169,n9179);
and (n9169,n9170,n655);
nand (n9170,n9171,n9177);
or (n9171,n8773,n9172);
not (n9172,n9173);
nand (n9173,n9174,n9176);
or (n9174,n8728,n9175);
not (n9175,n8862);
or (n9176,n8862,n8727);
or (n9177,n9173,n9178);
not (n9178,n8773);
and (n9179,n9180,n655);
nand (n9180,n9181,n9182);
or (n9181,n8625,n8627);
nand (n9182,n8627,n8625);
wire s0n9183,s1n9183,notn9183;
or (n9183,s0n9183,s1n9183);
not(notn9183,n8508);
and (s0n9183,notn9183,1'b0);
and (s1n9183,n8508,n9140);
and (n9184,n9169,n9179);
wire s0n9185,s1n9185,notn9185;
or (n9185,s0n9185,s1n9185);
not(notn9185,n728);
and (s0n9185,notn9185,1'b0);
and (s1n9185,n728,n9056);
and (n9186,n9165,n9166);
wire s0n9187,s1n9187,notn9187;
or (n9187,s0n9187,s1n9187);
not(notn9187,n8059);
and (s0n9187,notn9187,1'b0);
and (s1n9187,n8059,n9188);
xor (n9188,n9189,n8479);
xor (n9189,n8473,n8476);
and (n9190,n9161,n9162);
or (n9191,n9192,n9273);
and (n9192,n9193,n9270);
xor (n9193,n9194,n9218);
xor (n9194,n9195,n9217);
xor (n9195,n9196,n9197);
wire s0n9196,s1n9196,notn9196;
or (n9196,s0n9196,s1n9196);
not(notn9196,n8320);
and (s0n9196,notn9196,1'b0);
and (s1n9196,n8320,n8519);
or (n9197,n9198,n9216);
and (n9198,n9199,n9215);
xor (n9199,n9200,n9213);
or (n9200,n9201,n9208);
and (n9201,n9202,n655);
nand (n9202,n9203,n9205,n9207);
or (n9203,n8522,n9204);
not (n9204,n8605);
or (n9205,n8625,n9206);
not (n9206,n8579);
not (n9207,n8563);
and (n9208,n9209,n655);
or (n9209,n9210,n8786);
nor (n9210,n9211,n8869);
and (n9211,n9212,n9004);
not (n9212,n8798);
nor (n9213,n9214,n8322);
xor (n9214,n8858,n8856);
wire s0n9215,s1n9215,notn9215;
or (n9215,s0n9215,s1n9215);
not(notn9215,n8508);
and (s0n9215,notn9215,1'b0);
and (s1n9215,n8508,n9134);
and (n9216,n9200,n9213);
wire s0n9217,s1n9217,notn9217;
or (n9217,s0n9217,s1n9217);
not(notn9217,n728);
and (s0n9217,notn9217,1'b0);
and (s1n9217,n728,n8993);
and (n9218,n9219,n9269);
xor (n9219,n9220,n9263);
or (n9220,n9221,n9262);
and (n9221,n9222,n9259);
xor (n9222,n9223,n9237);
and (n9223,n9224,n9235);
xor (n9224,n9225,n9233);
and (n9225,n9226,n9230);
nor (n9226,n9227,n8869);
not (n9227,n9228);
wire s0n9228,s1n9228,notn9228;
or (n9228,s0n9228,s1n9228);
not(notn9228,n655);
and (s0n9228,notn9228,1'b0);
and (s1n9228,n655,n9229);
wire s0n9229,s1n9229,notn9229;
or (n9229,s0n9229,s1n9229);
not(notn9229,n10);
and (s0n9229,notn9229,1'b0);
and (s1n9229,n10,n8832);
and (n9230,n9231,n655);
nor (n9231,n9232,n9204);
not (n9232,n8644);
wire s0n9233,s1n9233,notn9233;
or (n9233,s0n9233,s1n9233);
not(notn9233,n8058);
and (s0n9233,notn9233,1'b0);
and (s1n9233,n8058,n9234);
xor (n9234,n8608,n8619);
and (n9235,n9236,n655);
xnor (n9236,n8869,n8871);
or (n9237,n9238,n9258);
and (n9238,n9239,n9253);
xor (n9239,n9240,n9246);
and (n9240,n9241,n655);
nand (n9241,n9242,n9243,n9245);
or (n9242,n8639,n9206);
or (n9243,n8625,n9244);
not (n9244,n8619);
not (n9245,n8578);
and (n9246,n9247,n655);
not (n9247,n9248);
nor (n9248,n9249,n9250);
and (n9249,n8868,n8817);
nor (n9250,n9251,n9002);
and (n9251,n8876,n9252);
not (n9252,n8802);
and (n9253,n9254,n655);
xor (n9254,n9255,n9256);
not (n9255,n8564);
xnor (n9256,n8632,n9257);
not (n9257,n8575);
and (n9258,n9240,n9246);
wire s0n9259,s1n9259,notn9259;
or (n9259,s0n9259,s1n9259);
not(notn9259,n8059);
and (s0n9259,notn9259,1'b0);
and (s1n9259,n8059,n9260);
xor (n9260,n9261,n8880);
xor (n9261,n8875,n8877);
and (n9262,n9223,n9237);
and (n9263,n9264,n9268);
xor (n9264,n9265,n9266);
wire s0n9265,s1n9265,notn9265;
or (n9265,s0n9265,s1n9265);
not(notn9265,n728);
and (s0n9265,notn9265,1'b0);
and (s1n9265,n728,n9143);
wire s0n9266,s1n9266,notn9266;
or (n9266,s0n9266,s1n9266);
not(notn9266,n8058);
and (s0n9266,notn9266,1'b0);
and (s1n9266,n8058,n9267);
xor (n9267,n8644,n8645);
wire s0n9268,s1n9268,notn9268;
or (n9268,s0n9268,s1n9268);
not(notn9268,n8320);
and (s0n9268,notn9268,1'b0);
and (s1n9268,n8320,n9134);
xor (n9269,n9137,n9142);
wire s0n9270,s1n9270,notn9270;
or (n9270,s0n9270,s1n9270);
not(notn9270,n8508);
and (s0n9270,notn9270,1'b0);
and (s1n9270,n8508,n9271);
xor (n9271,n9272,n8293);
xor (n9272,n8287,n8290);
and (n9273,n9194,n9218);
wire s0n9274,s1n9274,notn9274;
or (n9274,s0n9274,s1n9274);
not(notn9274,n655);
and (s0n9274,notn9274,1'b0);
and (s1n9274,n655,n9061);
and (n9275,n9158,n9191);
xor (n9276,n8923,n8930);
xor (n9277,n9278,n9300);
xor (n9278,n9279,n9280);
wire s0n9279,s1n9279,notn9279;
or (n9279,s0n9279,s1n9279);
not(notn9279,n655);
and (s0n9279,notn9279,1'b0);
and (s1n9279,n655,n8324);
xor (n9280,n9281,n9297);
xor (n9281,n9282,n9283);
wire s0n9282,s1n9282,notn9282;
or (n9282,s0n9282,s1n9282);
not(notn9282,n8320);
and (s0n9282,notn9282,1'b0);
and (s1n9282,n8320,n8747);
or (n9283,n9284,n9296);
and (n9284,n9285,n9293);
xor (n9285,n9286,n9287);
xor (n9286,n8694,n8708);
and (n9287,n9288,n655);
nand (n9288,n9289,n9291);
or (n9289,n9290,n9054);
and (n9290,n9051,n8734);
or (n9291,n9010,n9292);
not (n9292,n8667);
or (n9293,n9294,n9295);
and (n9294,n9034,n9047);
and (n9295,n9035,n9040);
and (n9296,n9286,n9287);
wire s0n9297,s1n9297,notn9297;
or (n9297,s0n9297,s1n9297);
not(notn9297,n8059);
and (s0n9297,notn9297,1'b0);
and (s1n9297,n8059,n9298);
xor (n9298,n9299,n8853);
xor (n9299,n8849,n8850);
wire s0n9300,s1n9300,notn9300;
or (n9300,s0n9300,s1n9300);
not(notn9300,n655);
and (s0n9300,notn9300,1'b0);
and (s1n9300,n655,n8506);
and (n9301,n9155,n9276);
and (n9302,n9112,n9113);
and (n9303,n8125,n9064);
xor (n9304,n9305,n9328);
xor (n9305,n9306,n9309);
or (n9306,n9307,n9308);
and (n9307,n9065,n9096);
and (n9308,n9066,n9079);
and (n9309,n9310,n9321);
xor (n9310,n9311,n9320);
or (n9311,n9312,n9319);
and (n9312,n9313,n9318);
xor (n9313,n9314,n9315);
wire s0n9314,s1n9314,notn9314;
or (n9314,s0n9314,s1n9314);
not(notn9314,n8320);
and (s0n9314,notn9314,1'b0);
and (s1n9314,n8320,n8905);
xor (n9315,n9316,n9317);
xor (n9316,n9070,n9073);
wire s0n9317,s1n9317,notn9317;
or (n9317,s0n9317,s1n9317);
not(notn9317,n8058);
and (s0n9317,notn9317,1'b0);
and (s1n9317,n8058,n8731);
wire s0n9318,s1n9318,notn9318;
or (n9318,s0n9318,s1n9318);
not(notn9318,n728);
and (s0n9318,notn9318,1'b0);
and (s1n9318,n728,n8324);
and (n9319,n9314,n9315);
wire s0n9320,s1n9320,notn9320;
or (n9320,s0n9320,s1n9320);
not(notn9320,n728);
and (s0n9320,notn9320,1'b0);
and (s1n9320,n728,n9101);
and (n9321,n9322,n9327);
xor (n9322,n9323,n9324);
and (n9323,n8931,n8058);
or (n9324,n9325,n9326);
and (n9325,n9281,n9297);
and (n9326,n9282,n9283);
wire s0n9327,s1n9327,notn9327;
or (n9327,s0n9327,s1n9327);
not(notn9327,n728);
and (s0n9327,notn9327,1'b0);
and (s1n9327,n728,n9077);
xor (n9328,n9329,n9332);
xor (n9329,n9330,n9331);
and (n9330,n9067,n9076);
and (n9331,n8892,n8904);
or (n9332,n9333,n9334);
and (n9333,n8128,n8505);
and (n9334,n8129,n8323);
xor (n9335,n9336,n9355);
xor (n9336,n9337,n9340);
or (n9337,n9338,n9339);
and (n9338,n8126,n8918);
and (n9339,n8127,n8511);
xor (n9340,n9341,n9350);
xor (n9341,n9342,n9345);
or (n9342,n9343,n9344);
and (n9343,n8512,n8907);
and (n9344,n8513,n8891);
xor (n9345,n9346,n9349);
xor (n9346,n9347,n9348);
wire s0n9347,s1n9347,notn9347;
or (n9347,s0n9347,s1n9347);
not(notn9347,n8058);
and (s0n9347,notn9347,1'b0);
and (s1n9347,n8058,n8905);
wire s0n9348,s1n9348,notn9348;
or (n9348,s0n9348,s1n9348);
not(notn9348,n8508);
and (s0n9348,notn9348,1'b0);
and (s1n9348,n8508,n8894);
wire s0n9349,s1n9349,notn9349;
or (n9349,s0n9349,s1n9349);
not(notn9349,n8058);
and (s0n9349,notn9349,1'b0);
and (s1n9349,n8058,n8506);
xor (n9350,n9351,n9354);
xor (n9351,n9352,n9353);
wire s0n9352,s1n9352,notn9352;
or (n9352,s0n9352,s1n9352);
not(notn9352,n8059);
and (s0n9352,notn9352,1'b0);
and (s1n9352,n8059,n9101);
wire s0n9353,s1n9353,notn9353;
or (n9353,s0n9353,s1n9353);
not(notn9353,n8059);
and (s0n9353,notn9353,1'b0);
and (s1n9353,n8059,n8908);
wire s0n9354,s1n9354,notn9354;
or (n9354,s0n9354,s1n9354);
not(notn9354,n8508);
and (s0n9354,notn9354,1'b0);
and (s1n9354,n8508,n8130);
or (n9355,n9356,n9397);
and (n9356,n9357,n9368);
xor (n9357,n9358,n9367);
or (n9358,n9359,n9366);
and (n9359,n9360,n9363);
xor (n9360,n9361,n9362);
xor (n9361,n9081,n9094);
xor (n9362,n9313,n9318);
or (n9363,n9364,n9365);
and (n9364,n9278,n9300);
and (n9365,n9279,n9280);
and (n9366,n9361,n9362);
xor (n9367,n9310,n9321);
or (n9368,n9369,n9396);
and (n9369,n9370,n9395);
xor (n9370,n9371,n9372);
xor (n9371,n9322,n9327);
or (n9372,n9373,n9394);
and (n9373,n9374,n9385);
xor (n9374,n9375,n9376);
xor (n9375,n9084,n9091);
or (n9376,n9377,n9384);
and (n9377,n9378,n9383);
xor (n9378,n9379,n9382);
or (n9379,n9380,n9381);
and (n9380,n9195,n9217);
and (n9381,n9196,n9197);
xor (n9382,n9285,n9293);
wire s0n9383,s1n9383,notn9383;
or (n9383,s0n9383,s1n9383);
not(notn9383,n728);
and (s0n9383,notn9383,1'b0);
and (s1n9383,n728,n9298);
and (n9384,n9379,n9382);
or (n9385,n9386,n9393);
and (n9386,n9387,n9390);
xor (n9387,n9388,n9389);
wire s0n9388,s1n9388,notn9388;
or (n9388,s0n9388,s1n9388);
not(notn9388,n8058);
and (s0n9388,notn9388,1'b0);
and (s1n9388,n8058,n9271);
xor (n9389,n9087,n9090);
wire s0n9390,s1n9390,notn9390;
or (n9390,s0n9390,s1n9390);
not(notn9390,n8059);
and (s0n9390,notn9390,1'b0);
and (s1n9390,n8059,n9391);
xor (n9391,n9392,n8471);
xor (n9392,n8465,n8468);
and (n9393,n9388,n9389);
and (n9394,n9375,n9376);
xor (n9395,n9098,n9107);
and (n9396,n9371,n9372);
and (n9397,n9358,n9367);
or (n9398,n9399,n9470);
and (n9399,n9400,n9469);
xor (n9400,n9401,n9402);
xor (n9401,n9357,n9368);
or (n9402,n9403,n9468);
and (n9403,n9404,n9407);
xor (n9404,n9405,n9406);
xor (n9405,n9370,n9395);
xor (n9406,n9360,n9363);
or (n9407,n9408,n9467);
and (n9408,n9409,n9454);
xor (n9409,n9410,n9453);
or (n9410,n9411,n9452);
and (n9411,n9412,n9415);
xor (n9412,n9413,n9414);
xor (n9413,n9387,n9390);
xor (n9414,n9378,n9383);
or (n9415,n9416,n9451);
and (n9416,n9417,n9450);
xor (n9417,n9418,n9441);
or (n9418,n9419,n9440);
and (n9419,n9420,n9439);
xor (n9420,n9421,n9422);
xor (n9421,n9164,n9185);
or (n9422,n9423,n9438);
and (n9423,n9424,n9430);
xor (n9424,n9425,n9426);
xor (n9425,n9168,n9183);
nand (n9426,n9427,n9200);
or (n9427,n9428,n9429);
not (n9428,n9208);
not (n9429,n9201);
or (n9430,n9431,n9437);
and (n9431,n9432,n9436);
xor (n9432,n9433,n9434);
wire s0n9433,s1n9433,notn9433;
or (n9433,s0n9433,s1n9433);
not(notn9433,n8508);
and (s0n9433,notn9433,1'b0);
and (s1n9433,n8508,n9267);
wire s0n9434,s1n9434,notn9434;
or (n9434,s0n9434,s1n9434);
not(notn9434,n8059);
and (s0n9434,notn9434,1'b0);
and (s1n9434,n8059,n9435);
xor (n9435,n8881,n8883);
wire s0n9436,s1n9436,notn9436;
or (n9436,s0n9436,s1n9436);
not(notn9436,n8320);
and (s0n9436,notn9436,1'b0);
and (s1n9436,n8320,n9140);
and (n9437,n9433,n9434);
and (n9438,n9425,n9426);
wire s0n9439,s1n9439,notn9439;
or (n9439,s0n9439,s1n9439);
not(notn9439,n8508);
and (s0n9439,notn9439,1'b0);
and (s1n9439,n8508,n9146);
and (n9440,n9421,n9422);
and (n9441,n9442,n9447);
xor (n9442,n9443,n9446);
wire s0n9443,s1n9443,notn9443;
or (n9443,s0n9443,s1n9443);
not(notn9443,n8058);
and (s0n9443,notn9443,1'b0);
and (s1n9443,n8058,n9444);
xor (n9444,n9445,n8309);
xor (n9445,n8303,n8306);
xor (n9446,n9199,n9215);
wire s0n9447,s1n9447,notn9447;
or (n9447,s0n9447,s1n9447);
not(notn9447,n8059);
and (s0n9447,notn9447,1'b0);
and (s1n9447,n8059,n9448);
xor (n9448,n9449,n8487);
xor (n9449,n8481,n8484);
wire s0n9450,s1n9450,notn9450;
or (n9450,s0n9450,s1n9450);
not(notn9450,n655);
and (s0n9450,notn9450,1'b0);
and (s1n9450,n655,n8928);
and (n9451,n9418,n9441);
and (n9452,n9413,n9414);
xor (n9453,n9374,n9385);
or (n9454,n9455,n9466);
and (n9455,n9456,n9465);
xor (n9456,n9457,n9458);
xor (n9457,n9119,n9122);
or (n9458,n9459,n9464);
and (n9459,n9460,n9463);
xor (n9460,n9461,n9462);
and (n9461,n8987,n8320);
wire s0n9462,s1n9462,notn9462;
or (n9462,s0n9462,s1n9462);
not(notn9462,n728);
and (s0n9462,notn9462,1'b0);
and (s1n9462,n728,n9391);
and (n9463,n8931,n655);
and (n9464,n9461,n9462);
xor (n9465,n9126,n9149);
and (n9466,n9457,n9458);
and (n9467,n9410,n9453);
and (n9468,n9405,n9406);
xor (n9469,n8124,n9109);
and (n9470,n9401,n9402);
or (n9471,n9472,n9945);
and (n9472,n9473,n9550);
xor (n9473,n9474,n9475);
xor (n9474,n9400,n9469);
or (n9475,n9476,n9549);
and (n9476,n9477,n9548);
xor (n9477,n9478,n9479);
xor (n9478,n9111,n9152);
or (n9479,n9480,n9547);
and (n9480,n9481,n9484);
xor (n9481,n9482,n9483);
xor (n9482,n9115,n9124);
xor (n9483,n9154,n9277);
or (n9484,n9485,n9546);
and (n9485,n9486,n9525);
xor (n9486,n9487,n9488);
xor (n9487,n9157,n9274);
or (n9488,n9489,n9524);
and (n9489,n9490,n9493);
xor (n9490,n9491,n9492);
xor (n9491,n9160,n9187);
xor (n9492,n9130,n9145);
or (n9493,n9494,n9523);
and (n9494,n9495,n9522);
xor (n9495,n9496,n9521);
and (n9496,n9497,n9498);
xor (n9497,n9222,n9259);
or (n9498,n9499,n9520);
and (n9499,n9500,n9519);
xor (n9500,n9501,n9518);
or (n9501,n9502,n9517);
and (n9502,n9503,n9510);
xor (n9503,n9504,n9506);
wire s0n9504,s1n9504,notn9504;
or (n9504,s0n9504,s1n9504);
not(notn9504,n8059);
and (s0n9504,notn9504,1'b0);
and (s1n9504,n8059,n9505);
xor (n9505,n8831,n8842);
and (n9506,n9507,n9508);
wire s0n9507,s1n9507,notn9507;
or (n9507,s0n9507,s1n9507);
not(notn9507,n8059);
and (s0n9507,notn9507,1'b0);
and (s1n9507,n8059,n9229);
wire s0n9508,s1n9508,notn9508;
or (n9508,s0n9508,s1n9508);
not(notn9508,n8059);
and (s0n9508,notn9508,1'b0);
and (s1n9508,n8059,n9509);
wire s0n9509,s1n9509,notn9509;
or (n9509,s0n9509,s1n9509);
not(notn9509,n10);
and (s0n9509,notn9509,1'b0);
and (s1n9509,n10,n8433);
and (n9510,n9511,n655);
nand (n9511,n9512,n9516);
or (n9512,n9252,n9513);
nand (n9513,n9514,n9515);
or (n9514,n8813,n8876);
nand (n9515,n8813,n8876);
nand (n9516,n9513,n9252);
and (n9517,n9504,n9506);
xor (n9518,n9239,n9253);
wire s0n9519,s1n9519,notn9519;
or (n9519,s0n9519,s1n9519);
not(notn9519,n728);
and (s0n9519,notn9519,1'b0);
and (s1n9519,n728,n9260);
and (n9520,n9501,n9518);
wire s0n9521,s1n9521,notn9521;
or (n9521,s0n9521,s1n9521);
not(notn9521,n8320);
and (s0n9521,notn9521,1'b0);
and (s1n9521,n8320,n9271);
wire s0n9522,s1n9522,notn9522;
or (n9522,s0n9522,s1n9522);
not(notn9522,n728);
and (s0n9522,notn9522,1'b0);
and (s1n9522,n728,n9188);
and (n9523,n9496,n9521);
and (n9524,n9491,n9492);
or (n9525,n9526,n9545);
and (n9526,n9527,n9544);
xor (n9527,n9528,n9529);
xor (n9528,n9193,n9270);
or (n9529,n9530,n9543);
and (n9530,n9531,n9542);
xor (n9531,n9532,n9541);
or (n9532,n9533,n9540);
and (n9533,n9534,n9539);
xor (n9534,n9535,n9536);
xor (n9535,n9264,n9268);
wire s0n9536,s1n9536,notn9536;
or (n9536,s0n9536,s1n9536);
not(notn9536,n8059);
and (s0n9536,notn9536,1'b0);
and (s1n9536,n8059,n9537);
xor (n9537,n9538,n8495);
xor (n9538,n8489,n8492);
wire s0n9539,s1n9539,notn9539;
or (n9539,s0n9539,s1n9539);
not(notn9539,n8508);
and (s0n9539,notn9539,1'b0);
and (s1n9539,n8508,n9444);
and (n9540,n9535,n9536);
xor (n9541,n9219,n9269);
and (n9542,n8987,n655);
and (n9543,n9532,n9541);
xor (n9544,n9460,n9463);
and (n9545,n9528,n9529);
and (n9546,n9487,n9488);
and (n9547,n9482,n9483);
xor (n9548,n9404,n9407);
and (n9549,n9478,n9479);
or (n9550,n9551,n9944);
and (n9551,n9552,n9682);
xor (n9552,n9553,n9554);
xor (n9553,n9477,n9548);
or (n9554,n9555,n9681);
and (n9555,n9556,n9680);
xor (n9556,n9557,n9558);
xor (n9557,n9409,n9454);
or (n9558,n9559,n9679);
and (n9559,n9560,n9678);
xor (n9560,n9561,n9562);
xor (n9561,n9412,n9415);
or (n9562,n9563,n9677);
and (n9563,n9564,n9609);
xor (n9564,n9565,n9608);
or (n9565,n9566,n9607);
and (n9566,n9567,n9570);
xor (n9567,n9568,n9569);
xor (n9568,n9442,n9447);
wire s0n9569,s1n9569,notn9569;
or (n9569,s0n9569,s1n9569);
not(notn9569,n655);
and (s0n9569,notn9569,1'b0);
and (s1n9569,n655,n9391);
or (n9570,n9571,n9606);
and (n9571,n9572,n9605);
xor (n9572,n9573,n9587);
or (n9573,n9574,n9586);
and (n9574,n9575,n9584);
xor (n9575,n9576,n9578);
wire s0n9576,s1n9576,notn9576;
or (n9576,s0n9576,s1n9576);
not(notn9576,n8059);
and (s0n9576,notn9576,1'b0);
and (s1n9576,n8059,n9577);
xor (n9577,n8496,n8497);
and (n9578,n9579,n9583);
xor (n9579,n9580,n9581);
xor (n9580,n9226,n9230);
wire s0n9581,s1n9581,notn9581;
or (n9581,s0n9581,s1n9581);
not(notn9581,n8058);
and (s0n9581,notn9581,1'b0);
and (s1n9581,n8058,n9582);
wire s0n9582,s1n9582,notn9582;
or (n9582,s0n9582,s1n9582);
not(notn9582,n10);
and (s0n9582,notn9582,1'b0);
and (s1n9582,n10,n8609);
wire s0n9583,s1n9583,notn9583;
or (n9583,s0n9583,s1n9583);
not(notn9583,n728);
and (s0n9583,notn9583,1'b0);
and (s1n9583,n728,n9435);
wire s0n9584,s1n9584,notn9584;
or (n9584,s0n9584,s1n9584);
not(notn9584,n8508);
and (s0n9584,notn9584,1'b0);
and (s1n9584,n8508,n9585);
xor (n9585,n8310,n8311);
and (n9586,n9576,n9578);
or (n9587,n9588,n9604);
and (n9588,n9589,n9602);
xor (n9589,n9590,n9591);
xor (n9590,n9224,n9235);
and (n9591,n9592,n9601);
xor (n9592,n9593,n9599);
and (n9593,n9594,n655);
xnor (n9594,n9595,n9206);
nand (n9595,n9596,n9598);
or (n9596,n8638,n9597);
not (n9597,n8590);
nand (n9598,n8638,n9597);
wire s0n9599,s1n9599,notn9599;
or (n9599,s0n9599,s1n9599);
not(notn9599,n8058);
and (s0n9599,notn9599,1'b0);
and (s1n9599,n8058,n9600);
wire s0n9600,s1n9600,notn9600;
or (n9600,s0n9600,s1n9600);
not(notn9600,n10);
and (s0n9600,notn9600,1'b0);
and (s1n9600,n10,n8245);
wire s0n9601,s1n9601,notn9601;
or (n9601,s0n9601,s1n9601);
not(notn9601,n8508);
and (s0n9601,notn9601,1'b0);
and (s1n9601,n8508,n9234);
wire s0n9602,s1n9602,notn9602;
or (n9602,s0n9602,s1n9602);
not(notn9602,n8058);
and (s0n9602,notn9602,1'b0);
and (s1n9602,n8058,n9603);
xor (n9603,n8244,n8256);
and (n9604,n9590,n9591);
wire s0n9605,s1n9605,notn9605;
or (n9605,s0n9605,s1n9605);
not(notn9605,n8320);
and (s0n9605,notn9605,1'b0);
and (s1n9605,n8320,n9146);
and (n9606,n9573,n9587);
and (n9607,n9568,n9569);
xor (n9608,n9417,n9450);
or (n9609,n9610,n9676);
and (n9610,n9611,n9675);
xor (n9611,n9612,n9674);
or (n9612,n9613,n9673);
and (n9613,n9614,n9672);
xor (n9614,n9615,n9616);
xor (n9615,n9424,n9430);
or (n9616,n9617,n9671);
and (n9617,n9618,n9646);
xor (n9618,n9619,n9620);
xor (n9619,n9432,n9436);
or (n9620,n9621,n9645);
and (n9621,n9622,n9644);
xor (n9622,n9623,n9633);
or (n9623,n9624,n9632);
and (n9624,n9625,n9628);
xor (n9625,n9626,n9627);
wire s0n9626,s1n9626,notn9626;
or (n9626,s0n9626,s1n9626);
not(notn9626,n728);
and (s0n9626,notn9626,1'b0);
and (s1n9626,n728,n9505);
xor (n9627,n9507,n9508);
and (n9628,n9629,n655);
nand (n9629,n9630,n9631);
or (n9630,n8605,n9232);
or (n9631,n8644,n9204);
and (n9632,n9626,n9627);
or (n9633,n9634,n9643);
and (n9634,n9635,n9638);
xor (n9635,n9636,n9637);
and (n9636,n8594,n655);
and (n9637,n8817,n655);
and (n9638,n9639,n655);
nand (n9639,n9640,n9642);
or (n9640,n8881,n9641);
not (n9641,n8828);
nand (n9642,n8881,n9641);
and (n9643,n9636,n9637);
wire s0n9644,s1n9644,notn9644;
or (n9644,s0n9644,s1n9644);
not(notn9644,n8320);
and (s0n9644,notn9644,1'b0);
and (s1n9644,n8320,n9267);
and (n9645,n9623,n9633);
or (n9646,n9647,n9670);
and (n9647,n9648,n9668);
xor (n9648,n9649,n9650);
xor (n9649,n9503,n9510);
or (n9650,n9651,n9667);
and (n9651,n9652,n9666);
xor (n9652,n9653,n9661);
or (n9653,n9654,n9660);
and (n9654,n9655,n9658);
xor (n9655,n9656,n9657);
nor (n9656,n9244,n8322);
wire s0n9657,s1n9657,notn9657;
or (n9657,s0n9657,s1n9657);
not(notn9657,n728);
and (s0n9657,notn9657,1'b0);
and (s1n9657,n728,n9229);
nor (n9658,n9659,n8322);
not (n9659,n8842);
and (n9660,n9656,n9657);
and (n9661,n9662,n9664);
nor (n9662,n9663,n8322);
not (n9663,n8608);
nor (n9664,n9665,n8322);
not (n9665,n8831);
wire s0n9666,s1n9666,notn9666;
or (n9666,s0n9666,s1n9666);
not(notn9666,n8508);
and (s0n9666,notn9666,1'b0);
and (s1n9666,n8508,n9600);
and (n9667,n9653,n9661);
wire s0n9668,s1n9668,notn9668;
or (n9668,s0n9668,s1n9668);
not(notn9668,n8059);
and (s0n9668,notn9668,1'b0);
and (s1n9668,n8059,n9669);
xor (n9669,n8432,n8443);
and (n9670,n9649,n9650);
and (n9671,n9619,n9620);
wire s0n9672,s1n9672,notn9672;
or (n9672,s0n9672,s1n9672);
not(notn9672,n728);
and (s0n9672,notn9672,1'b0);
and (s1n9672,n728,n9448);
and (n9673,n9615,n9616);
xor (n9674,n9420,n9439);
xor (n9675,n9495,n9522);
and (n9676,n9612,n9674);
and (n9677,n9565,n9608);
xor (n9678,n9456,n9465);
and (n9679,n9561,n9562);
xor (n9680,n9481,n9484);
and (n9681,n9557,n9558);
or (n9682,n9683,n9943);
and (n9683,n9684,n9743);
xor (n9684,n9685,n9686);
xor (n9685,n9556,n9680);
or (n9686,n9687,n9742);
and (n9687,n9688,n9741);
xor (n9688,n9689,n9690);
xor (n9689,n9486,n9525);
or (n9690,n9691,n9740);
and (n9691,n9692,n9739);
xor (n9692,n9693,n9694);
xor (n9693,n9490,n9493);
or (n9694,n9695,n9738);
and (n9695,n9696,n9737);
xor (n9696,n9697,n9706);
or (n9697,n9698,n9705);
and (n9698,n9699,n9704);
xor (n9699,n9700,n9703);
xor (n9700,n9701,n9702);
xor (n9701,n9497,n9498);
wire s0n9702,s1n9702,notn9702;
or (n9702,s0n9702,s1n9702);
not(notn9702,n8058);
and (s0n9702,notn9702,1'b0);
and (s1n9702,n8058,n9585);
wire s0n9703,s1n9703,notn9703;
or (n9703,s0n9703,s1n9703);
not(notn9703,n655);
and (s0n9703,notn9703,1'b0);
and (s1n9703,n655,n9271);
wire s0n9704,s1n9704,notn9704;
or (n9704,s0n9704,s1n9704);
not(notn9704,n655);
and (s0n9704,notn9704,1'b0);
and (s1n9704,n655,n9188);
and (n9705,n9700,n9703);
or (n9706,n9707,n9736);
and (n9707,n9708,n9729);
xor (n9708,n9709,n9728);
or (n9709,n9710,n9727);
and (n9710,n9711,n9726);
xor (n9711,n9712,n9713);
xor (n9712,n9589,n9602);
or (n9713,n9714,n9725);
and (n9714,n9715,n9724);
xor (n9715,n9716,n9717);
wire s0n9716,s1n9716,notn9716;
or (n9716,s0n9716,s1n9716);
not(notn9716,n8508);
and (s0n9716,notn9716,1'b0);
and (s1n9716,n8508,n9603);
or (n9717,n9718,n9723);
and (n9718,n9719,n9722);
xor (n9719,n9720,n9721);
xor (n9720,n9635,n9638);
wire s0n9721,s1n9721,notn9721;
or (n9721,s0n9721,s1n9721);
not(notn9721,n8320);
and (s0n9721,notn9721,1'b0);
and (s1n9721,n8320,n9234);
wire s0n9722,s1n9722,notn9722;
or (n9722,s0n9722,s1n9722);
not(notn9722,n8508);
and (s0n9722,notn9722,1'b0);
and (s1n9722,n8508,n9582);
and (n9723,n9720,n9721);
xor (n9724,n9579,n9583);
and (n9725,n9716,n9717);
wire s0n9726,s1n9726,notn9726;
or (n9726,s0n9726,s1n9726);
not(notn9726,n8320);
and (s0n9726,notn9726,1'b0);
and (s1n9726,n8320,n9444);
and (n9727,n9712,n9713);
xor (n9728,n9534,n9539);
or (n9729,n9730,n9735);
and (n9730,n9731,n9734);
xor (n9731,n9732,n9733);
wire s0n9732,s1n9732,notn9732;
or (n9732,s0n9732,s1n9732);
not(notn9732,n728);
and (s0n9732,notn9732,1'b0);
and (s1n9732,n728,n9537);
xor (n9733,n9500,n9519);
wire s0n9734,s1n9734,notn9734;
or (n9734,s0n9734,s1n9734);
not(notn9734,n655);
and (s0n9734,notn9734,1'b0);
and (s1n9734,n655,n9146);
and (n9735,n9732,n9733);
and (n9736,n9709,n9728);
xor (n9737,n9531,n9542);
and (n9738,n9697,n9706);
xor (n9739,n9527,n9544);
and (n9740,n9693,n9694);
xor (n9741,n9560,n9678);
and (n9742,n9689,n9690);
or (n9743,n9744,n9942);
and (n9744,n9745,n9778);
xor (n9745,n9746,n9777);
or (n9746,n9747,n9776);
and (n9747,n9748,n9775);
xor (n9748,n9749,n9774);
or (n9749,n9750,n9773);
and (n9750,n9751,n9772);
xor (n9751,n9752,n9771);
or (n9752,n9753,n9770);
and (n9753,n9754,n9757);
xor (n9754,n9755,n9756);
xor (n9755,n9572,n9605);
xor (n9756,n9614,n9672);
or (n9757,n9758,n9769);
and (n9758,n9759,n9768);
xor (n9759,n9760,n9761);
xor (n9760,n9575,n9584);
or (n9761,n9762,n9767);
and (n9762,n9763,n9766);
xor (n9763,n9764,n9765);
xor (n9764,n9592,n9601);
wire s0n9765,s1n9765,notn9765;
or (n9765,s0n9765,s1n9765);
not(notn9765,n728);
and (s0n9765,notn9765,1'b0);
and (s1n9765,n728,n9577);
wire s0n9766,s1n9766,notn9766;
or (n9766,s0n9766,s1n9766);
not(notn9766,n8320);
and (s0n9766,notn9766,1'b0);
and (s1n9766,n8320,n9585);
and (n9767,n9764,n9765);
wire s0n9768,s1n9768,notn9768;
or (n9768,s0n9768,s1n9768);
not(notn9768,n655);
and (s0n9768,notn9768,1'b0);
and (s1n9768,n655,n9448);
and (n9769,n9760,n9761);
and (n9770,n9755,n9756);
xor (n9771,n9567,n9570);
xor (n9772,n9611,n9675);
and (n9773,n9752,n9771);
xor (n9774,n9564,n9609);
xor (n9775,n9692,n9739);
and (n9776,n9749,n9774);
xor (n9777,n9688,n9741);
or (n9778,n9779,n9941);
and (n9779,n9780,n9845);
xor (n9780,n9781,n9844);
or (n9781,n9782,n9843);
and (n9782,n9783,n9842);
xor (n9783,n9784,n9841);
or (n9784,n9785,n9840);
and (n9785,n9786,n9833);
xor (n9786,n9787,n9832);
or (n9787,n9788,n9831);
and (n9788,n9789,n9812);
xor (n9789,n9790,n9811);
or (n9790,n9791,n9810);
and (n9791,n9792,n9809);
xor (n9792,n9793,n9808);
or (n9793,n9794,n9807);
and (n9794,n9795,n9806);
xor (n9795,n9796,n9797);
xor (n9796,n9625,n9628);
or (n9797,n9798,n9805);
and (n9798,n9799,n9804);
xor (n9799,n9800,n9803);
and (n9800,n9801,n9802);
wire s0n9801,s1n9801,notn9801;
or (n9801,s0n9801,s1n9801);
not(notn9801,n655);
and (s0n9801,notn9801,1'b0);
and (s1n9801,n655,n9582);
wire s0n9802,s1n9802,notn9802;
or (n9802,s0n9802,s1n9802);
not(notn9802,n655);
and (s0n9802,notn9802,1'b0);
and (s1n9802,n655,n9509);
wire s0n9803,s1n9803,notn9803;
or (n9803,s0n9803,s1n9803);
not(notn9803,n728);
and (s0n9803,notn9803,1'b0);
and (s1n9803,n728,n9509);
xor (n9804,n9662,n9664);
and (n9805,n9800,n9803);
wire s0n9806,s1n9806,notn9806;
or (n9806,s0n9806,s1n9806);
not(notn9806,n8320);
and (s0n9806,notn9806,1'b0);
and (s1n9806,n8320,n9603);
and (n9807,n9796,n9797);
xor (n9808,n9622,n9644);
xor (n9809,n9648,n9668);
and (n9810,n9793,n9808);
xor (n9811,n9618,n9646);
or (n9812,n9813,n9830);
and (n9813,n9814,n9829);
xor (n9814,n9815,n9828);
or (n9815,n9816,n9827);
and (n9816,n9817,n9826);
xor (n9817,n9818,n9819);
wire s0n9818,s1n9818,notn9818;
or (n9818,s0n9818,s1n9818);
not(notn9818,n728);
and (s0n9818,notn9818,1'b0);
and (s1n9818,n728,n9669);
or (n9819,n9820,n9825);
and (n9820,n9821,n9824);
xor (n9821,n9822,n9823);
wire s0n9822,s1n9822,notn9822;
or (n9822,s0n9822,s1n9822);
not(notn9822,n8320);
and (s0n9822,notn9822,1'b0);
and (s1n9822,n8320,n9600);
xor (n9823,n9655,n9658);
wire s0n9824,s1n9824,notn9824;
or (n9824,s0n9824,s1n9824);
not(notn9824,n8320);
and (s0n9824,notn9824,1'b0);
and (s1n9824,n8320,n9582);
and (n9825,n9822,n9823);
xor (n9826,n9719,n9722);
and (n9827,n9818,n9819);
wire s0n9828,s1n9828,notn9828;
or (n9828,s0n9828,s1n9828);
not(notn9828,n655);
and (s0n9828,notn9828,1'b0);
and (s1n9828,n655,n9537);
wire s0n9829,s1n9829,notn9829;
or (n9829,s0n9829,s1n9829);
not(notn9829,n655);
and (s0n9829,notn9829,1'b0);
and (s1n9829,n655,n9444);
and (n9830,n9815,n9828);
and (n9831,n9790,n9811);
xor (n9832,n9699,n9704);
or (n9833,n9834,n9839);
and (n9834,n9835,n9838);
xor (n9835,n9836,n9837);
xor (n9836,n9711,n9726);
xor (n9837,n9731,n9734);
xor (n9838,n9759,n9768);
and (n9839,n9836,n9837);
and (n9840,n9787,n9832);
xor (n9841,n9696,n9737);
xor (n9842,n9751,n9772);
and (n9843,n9784,n9841);
xor (n9844,n9748,n9775);
or (n9845,n9846,n9940);
and (n9846,n9847,n9939);
xor (n9847,n9848,n9891);
or (n9848,n9849,n9890);
and (n9849,n9850,n9889);
xor (n9850,n9851,n9888);
or (n9851,n9852,n9887);
and (n9852,n9853,n9868);
xor (n9853,n9854,n9867);
or (n9854,n9855,n9866);
and (n9855,n9856,n9865);
xor (n9856,n9857,n9864);
or (n9857,n9858,n9863);
and (n9858,n9859,n9862);
xor (n9859,n9860,n9861);
wire s0n9860,s1n9860,notn9860;
or (n9860,s0n9860,s1n9860);
not(notn9860,n655);
and (s0n9860,notn9860,1'b0);
and (s1n9860,n655,n9577);
xor (n9861,n9652,n9666);
wire s0n9862,s1n9862,notn9862;
or (n9862,s0n9862,s1n9862);
not(notn9862,n655);
and (s0n9862,notn9862,1'b0);
and (s1n9862,n655,n9585);
and (n9863,n9860,n9861);
xor (n9864,n9715,n9724);
xor (n9865,n9763,n9766);
and (n9866,n9857,n9864);
xor (n9867,n9789,n9812);
or (n9868,n9869,n9886);
and (n9869,n9870,n9885);
xor (n9870,n9871,n9872);
xor (n9871,n9792,n9809);
or (n9872,n9873,n9884);
and (n9873,n9874,n9883);
xor (n9874,n9875,n9882);
or (n9875,n9876,n9881);
and (n9876,n9877,n9880);
xor (n9877,n9878,n9879);
wire s0n9878,s1n9878,notn9878;
or (n9878,s0n9878,s1n9878);
not(notn9878,n655);
and (s0n9878,notn9878,1'b0);
and (s1n9878,n655,n9603);
xor (n9879,n9799,n9804);
wire s0n9880,s1n9880,notn9880;
or (n9880,s0n9880,s1n9880);
not(notn9880,n655);
and (s0n9880,notn9880,1'b0);
and (s1n9880,n655,n9669);
and (n9881,n9878,n9879);
xor (n9882,n9795,n9806);
xor (n9883,n9817,n9826);
and (n9884,n9875,n9882);
xor (n9885,n9814,n9829);
and (n9886,n9871,n9872);
and (n9887,n9854,n9867);
xor (n9888,n9708,n9729);
xor (n9889,n9754,n9757);
and (n9890,n9851,n9888);
nand (n9891,n9892,n9935);
or (n9892,n9893,n9933);
not (n9893,n9894);
nand (n9894,n9895,n9897,n9932);
not (n9895,n9896);
xor (n9896,n9786,n9833);
nand (n9897,n9898,n9931);
or (n9898,n9899,n9900);
xor (n9899,n9853,n9868);
nand (n9900,n9901,n9928);
or (n9901,n9902,n9926);
not (n9902,n9903);
nand (n9903,n9904,n9923);
or (n9904,n9905,n9921);
not (n9905,n9906);
nand (n9906,n9907,n9918);
or (n9907,n9908,n9916);
not (n9908,n9909);
nand (n9909,n9910,n9913);
or (n9910,n9227,n9911);
not (n9911,n9912);
wire s0n9912,s1n9912,notn9912;
or (n9912,s0n9912,s1n9912);
not(notn9912,n655);
and (s0n9912,notn9912,1'b0);
and (s1n9912,n655,n9600);
nand (n9913,n9914,n9915);
or (n9914,n9912,n9228);
xor (n9915,n9801,n9802);
not (n9916,n9917);
xor (n9917,n9821,n9824);
nand (n9918,n9919,n9920);
or (n9919,n9917,n9909);
xor (n9920,n9877,n9880);
not (n9921,n9922);
xor (n9922,n9859,n9862);
nand (n9923,n9924,n9925);
or (n9924,n9922,n9906);
xor (n9925,n9874,n9883);
not (n9926,n9927);
xor (n9927,n9856,n9865);
nand (n9928,n9929,n9930);
or (n9929,n9927,n9903);
xor (n9930,n9870,n9885);
xor (n9931,n9835,n9838);
nand (n9932,n9899,n9900);
not (n9933,n9934);
xor (n9934,n9850,n9889);
nand (n9935,n9936,n9896);
or (n9936,n9937,n9938);
not (n9937,n9932);
not (n9938,n9897);
xor (n9939,n9783,n9842);
and (n9940,n9848,n9891);
and (n9941,n9781,n9844);
and (n9942,n9746,n9777);
and (n9943,n9685,n9686);
and (n9944,n9553,n9554);
and (n9945,n9474,n9475);
and (n9946,n8120,n9398);
nor (n9947,n9948,n9973);
not (n9948,n9949);
nor (n9949,n9950,n9970);
not (n9950,n9951);
nor (n9951,n9952,n9967);
not (n9952,n9953);
nor (n9953,n9954,n9964);
not (n9954,n9955);
nor (n9955,n9956,n9957);
and (n9956,n9351,n9354);
not (n9957,n9958);
nor (n9958,n9959,n9960);
and (n9959,n9346,n9349);
not (n9960,n9961);
xnor (n9961,n9962,n9963);
wire s0n9962,s1n9962,notn9962;
or (n9962,s0n9962,s1n9962);
not(notn9962,n8058);
and (s0n9962,notn9962,1'b0);
and (s1n9962,n8058,n8130);
wire s0n9963,s1n9963,notn9963;
or (n9963,s0n9963,s1n9963);
not(notn9963,n8058);
and (s0n9963,notn9963,1'b0);
and (s1n9963,n8058,n8894);
or (n9964,n9965,n9966);
and (n9965,n9341,n9350);
and (n9966,n9342,n9345);
or (n9967,n9968,n9969);
and (n9968,n9305,n9328);
and (n9969,n9306,n9309);
or (n9970,n9971,n9972);
and (n9971,n9336,n9355);
and (n9972,n9337,n9340);
or (n9973,n9974,n9975);
and (n9974,n8121,n9335);
and (n9975,n8122,n9304);
nor (n9976,n1065,n8008);
not (n9977,n9978);
wire s0n9978,s1n9978,notn9978;
or (n9978,s0n9978,s1n9978);
not(notn9978,n12915);
and (s0n9978,notn9978,n9979);
and (s1n9978,n12915,n9989);
wire s0n9979,s1n9979,notn9979;
or (n9979,s0n9979,s1n9979);
not(notn9979,n13472);
and (s0n9979,notn9979,n9980);
and (s1n9979,n13472,n13858);
wire s0n9980,s1n9980,notn9980;
or (n9980,s0n9980,s1n9980);
not(notn9980,n13854);
and (s0n9980,notn9980,n9981);
and (s1n9980,n13854,n13648);
wire s0n9981,s1n9981,notn9981;
or (n9981,s0n9981,s1n9981);
not(notn9981,n13645);
and (s0n9981,notn9981,n9982);
and (s1n9981,n13645,n13540);
wire s0n9982,s1n9982,notn9982;
or (n9982,s0n9982,s1n9982);
not(notn9982,n13539);
and (s0n9982,notn9982,n9983);
and (s1n9982,n13539,n13455);
xor (n9983,n9984,n13389);
xor (n9984,n9985,n13328);
xor (n9985,n9986,n12935);
wire s0n9986,s1n9986,notn9986;
or (n9986,s0n9986,s1n9986);
not(notn9986,n12915);
and (s0n9986,notn9986,n9987);
and (s1n9986,n12915,1'b0);
xor (n9987,n9988,n10531);
xor (n9988,n9989,n10397);
wire s0n9989,s1n9989,notn9989;
or (n9989,s0n9989,s1n9989);
not(notn9989,n10395);
and (s0n9989,notn9989,n9990);
and (s1n9989,n10395,n10276);
wire s0n9990,s1n9990,notn9990;
or (n9990,s0n9990,s1n9990);
not(notn9990,n1039);
and (s0n9990,notn9990,n9991);
and (s1n9990,n1039,n10262);
wire s0n9991,s1n9991,notn9991;
or (n9991,s0n9991,s1n9991);
not(notn9991,n10261);
and (s0n9991,notn9991,1'b0);
and (s1n9991,n10261,n9992);
or (n9992,n9993,n10022,n10127,n10235);
and (n9993,n9994,n10021);
wire s0n9994,s1n9994,notn9994;
or (n9994,s0n9994,s1n9994);
not(notn9994,n1057);
and (s0n9994,notn9994,1'b0);
and (s1n9994,n1057,n9995);
wire s0n9995,s1n9995,notn9995;
or (n9995,s0n9995,s1n9995);
not(notn9995,n10004);
and (s0n9995,notn9995,n9996);
and (s1n9995,n10004,n9997);
wire s0n9997,s1n9997,notn9997;
or (n9997,s0n9997,s1n9997);
not(notn9997,n10017);
and (s0n9997,notn9997,n9998);
and (s1n9997,n10017,n10006);
wire s0n9998,s1n9998,notn9998;
or (n9998,s0n9998,s1n9998);
not(notn9998,n10000);
and (s0n9998,notn9998,1'b0);
and (s1n9998,n10000,n9999);
and (n10000,n10001,n10004);
and (n10001,n10002,n1036);
nor (n10002,n10003,n1035);
not (n10003,n1037);
and (n10004,n10005,n44);
nor (n10005,n809,n810,n1051);
or (n10006,1'b0,n10007,n10010,n10013);
and (n10007,n10008,n10009);
or (n10009,n638,n621);
and (n10010,n10011,n10012);
or (n10012,n642,n626);
and (n10013,n9999,n10014);
or (n10014,n10015,n630);
or (n10015,n10016,n634);
or (n10016,n650,n646);
and (n10017,n10018,n619);
and (n10018,n10019,n10005);
and (n10019,n1040,n10020);
and (n10020,n1044,n1045);
and (n10021,n1036,n1037);
and (n10022,n10023,n10126);
or (n10023,1'b0,n10024,n10075,n10093,n10110);
and (n10024,n10025,n10073);
wire s0n10025,s1n10025,notn10025;
or (n10025,s0n10025,s1n10025);
not(notn10025,n65);
and (s0n10025,notn10025,1'b0);
and (s1n10025,n65,n10026);
wire s0n10026,s1n10026,notn10026;
or (n10026,s0n10026,s1n10026);
not(notn10026,n10068);
and (s0n10026,notn10026,n10027);
and (s1n10026,n10068,n10052);
wire s0n10027,s1n10027,notn10027;
or (n10027,s0n10027,s1n10027);
not(notn10027,n10047);
and (s0n10027,notn10027,1'b0);
and (s1n10027,n10047,n10028);
or (n10028,1'b0,n10029,n10038);
and (n10029,n10030,n10031);
or (n10031,n10032,n10037);
or (n10032,n10033,n10036);
or (n10033,n10034,n10035);
nor (n10034,n44,n39,n60,n56,n619);
nor (n10035,n44,n624,n60,n56,n619);
nor (n10036,n44,n39,n59,n56,n619);
nor (n10037,n44,n624,n59,n56,n619);
and (n10038,n10039,n10040);
or (n10040,n10041,n10046);
or (n10041,n10042,n10045);
or (n10042,n10043,n10044);
nor (n10043,n38,n39,n60,n56,n619);
nor (n10044,n38,n624,n60,n56,n619);
nor (n10045,n38,n39,n59,n56,n619);
nor (n10046,n38,n624,n59,n56,n619);
and (n10047,n10048,n1057);
and (n10048,n10049,n10051);
and (n10049,n51,n10050);
nand (n10050,n56,n51);
not (n10051,n1036);
or (n10052,1'b0,n10053,n10058,n10063,n10067);
and (n10053,n10054,n10055);
or (n10055,n10056,n618);
or (n10056,n10057,n623);
or (n10057,n640,n636);
and (n10058,n10059,n10060);
or (n10060,n10061,n621);
or (n10061,n10062,n626);
or (n10062,n642,n638);
and (n10063,n10030,n10064);
or (n10064,n10065,n628);
or (n10065,n10066,n632);
or (n10066,n648,n644);
and (n10067,n10039,n10014);
and (n10068,n10069,n10070);
and (n10069,n619,n1057);
or (n10070,n926,n10071);
and (n10071,n1041,n10072);
nor (n10072,n1044,n1045);
nor (n10073,n10074,n810,n811);
not (n10074,n809);
and (n10075,n10076,n10091);
wire s0n10076,s1n10076,notn10076;
or (n10076,s0n10076,s1n10076);
not(notn10076,n65);
and (s0n10076,notn10076,1'b0);
and (s1n10076,n65,n10077);
wire s0n10077,s1n10077,notn10077;
or (n10077,s0n10077,s1n10077);
not(notn10077,n10068);
and (s0n10077,notn10077,n10078);
and (s1n10077,n10068,n10084);
wire s0n10078,s1n10078,notn10078;
or (n10078,s0n10078,s1n10078);
not(notn10078,n10047);
and (s0n10078,notn10078,1'b0);
and (s1n10078,n10047,n10079);
or (n10079,1'b0,n10080,n10082);
and (n10080,n10081,n10031);
and (n10082,n10083,n10040);
or (n10084,1'b0,n10085,n10087,n10089,n10090);
and (n10085,n10086,n10055);
and (n10087,n10088,n10060);
and (n10089,n10081,n10064);
and (n10090,n10083,n10014);
nor (n10091,n809,n10092,n811);
not (n10092,n810);
and (n10093,n10094,n10109);
wire s0n10094,s1n10094,notn10094;
or (n10094,s0n10094,s1n10094);
not(notn10094,n65);
and (s0n10094,notn10094,1'b0);
and (s1n10094,n65,n10095);
wire s0n10095,s1n10095,notn10095;
or (n10095,s0n10095,s1n10095);
not(notn10095,n10068);
and (s0n10095,notn10095,n10096);
and (s1n10095,n10068,n10102);
wire s0n10096,s1n10096,notn10096;
or (n10096,s0n10096,s1n10096);
not(notn10096,n10047);
and (s0n10096,notn10096,1'b0);
and (s1n10096,n10047,n10097);
or (n10097,1'b0,n10098,n10100);
and (n10098,n10099,n10031);
and (n10100,n10101,n10040);
or (n10102,1'b0,n10103,n10105,n10107,n10108);
and (n10103,n10104,n10055);
and (n10105,n10106,n10060);
and (n10107,n10099,n10064);
and (n10108,n10101,n10014);
not (n10109,n1050);
and (n10110,n10111,n10005);
wire s0n10111,s1n10111,notn10111;
or (n10111,s0n10111,s1n10111);
not(notn10111,n65);
and (s0n10111,notn10111,1'b0);
and (s1n10111,n65,n10112);
wire s0n10112,s1n10112,notn10112;
or (n10112,s0n10112,s1n10112);
not(notn10112,n10068);
and (s0n10112,notn10112,n10113);
and (s1n10112,n10068,n10119);
wire s0n10113,s1n10113,notn10113;
or (n10113,s0n10113,s1n10113);
not(notn10113,n10047);
and (s0n10113,notn10113,1'b0);
and (s1n10113,n10047,n10114);
or (n10114,1'b0,n10115,n10117);
and (n10115,n10116,n10031);
and (n10117,n10118,n10040);
or (n10119,1'b0,n10120,n10122,n10124,n10125);
and (n10120,n10121,n10055);
and (n10122,n10123,n10060);
and (n10124,n10116,n10064);
and (n10125,n10118,n10014);
and (n10126,n10051,n1037);
and (n10127,n10128,n10215);
nand (n10128,n10129,n10195,n10208,n10226);
nor (n10129,n10130,n10185,n10190);
and (n10130,n10131,n10177);
nand (n10131,n10132,n10158);
or (n10132,n10133,n10135);
not (n10133,n10134);
not (n10135,n10136);
nor (n10136,n10137,n10157);
and (n10137,n10138,n10145);
nor (n10138,n926,n10139);
and (n10139,n10020,n10140);
or (n10140,n10141,n10142,n10143,n10144);
nand (n10145,n10146,n10156);
nand (n10146,n10147,n1045);
or (n10147,n1044,n10148);
not (n10148,n10149);
and (n10149,n65,n10150);
not (n10150,n10151);
nor (n10151,n10152,n10153,n10154,n10155);
nor (n10156,n10072,n808);
nand (n10157,n65,n619);
nor (n10158,n10159,n10172);
and (n10159,n10160,n10171);
not (n10160,n10161);
nand (n10161,n10162,n10168);
nand (n10162,n10163,n10165);
not (n10163,n10164);
and (n10164,n10021,n10140);
nand (n10165,n10166,n10167);
or (n10166,n1036,n10149);
nor (n10167,n808,n1037);
and (n10168,n65,n10169);
nor (n10169,n10170,n56);
nand (n10170,n51,n615);
and (n10172,n10173,n10176);
not (n10173,n10174);
nand (n10174,n10162,n10175);
and (n10175,n65,n10170,n51);
nor (n10177,n10178,n10184);
nand (n10178,n10179,n10182);
or (n10179,n926,n10180);
and (n10180,n1041,n10181);
nor (n10181,n1043,n1045);
not (n10182,n10183);
nand (n10183,n65,n1057,n619);
nand (n10184,n58,n39);
and (n10185,n10186,n10188);
and (n10186,n10136,n10187);
nor (n10188,n10178,n10189);
nand (n10189,n56,n624);
and (n10190,n10191,n10193);
and (n10191,n10136,n10192);
nor (n10193,n10178,n10194);
nand (n10194,n56,n39);
nand (n10195,n10196,n10205);
nand (n10196,n10197,n10200);
or (n10197,n10198,n10135);
not (n10198,n10199);
nor (n10200,n10201,n10203);
and (n10201,n10160,n10202);
and (n10203,n10173,n10204);
nor (n10205,n10178,n10206);
not (n10206,n10207);
nor (n10207,n39,n56);
nor (n10208,n10209,n10221);
and (n10209,n10210,n10176);
not (n10210,n10211);
nand (n10211,n10212,n10220);
nor (n10212,n10213,n10216);
nor (n10213,n10214,n10215);
nor (n10214,n10148,n1037);
nor (n10215,n10051,n1037);
nand (n10216,n10217,n59);
not (n10217,n10218);
nand (n10218,n65,n10219);
and (n10219,n51,n1057);
not (n10220,n10184);
and (n10221,n10222,n10202);
not (n10222,n10223);
nand (n10223,n10224,n10225);
nor (n10224,n10213,n10218);
nor (n10225,n10206,n59);
nor (n10226,n10227,n10230);
and (n10227,n10228,n10204);
not (n10228,n10229);
nand (n10229,n10212,n10207);
and (n10230,n10231,n10171);
not (n10231,n10232);
nand (n10232,n10224,n10233);
and (n10233,n10234,n58);
nor (n10234,n624,n59);
and (n10235,n10236,n10260);
or (n10236,n10237,n10251,n10255,n10258);
and (n10237,n10238,n10242);
wire s0n10238,s1n10238,notn10238;
or (n10238,s0n10238,s1n10238);
not(notn10238,n10005);
and (s0n10238,notn10238,n10239);
and (s1n10238,n10005,n10240);
wire s0n10239,s1n10239,notn10239;
or (n10239,s0n10239,s1n10239);
not(notn10239,n10109);
and (s0n10239,notn10239,1'b0);
and (s1n10239,n10109,n9996);
wire s0n10240,s1n10240,notn10240;
or (n10240,s0n10240,s1n10240);
not(notn10240,n10241);
and (s0n10240,notn10240,n10111);
and (s1n10240,n10241,1'b0);
or (n10241,n10044,n10046);
nor (n10242,n10243,n10148);
not (n10243,n10244);
and (n10244,n65,n10245);
not (n10245,n10246);
nor (n10246,n10247,n10248,n10249,n10250);
and (n10251,n10252,n10254);
wire s0n10252,s1n10252,notn10252;
or (n10252,s0n10252,s1n10252);
not(notn10252,n10109);
and (s0n10252,notn10252,1'b0);
and (s1n10252,n10109,n10253);
and (n10254,n10243,n10149);
and (n10255,n10256,n10257);
wire s0n10256,s1n10256,notn10256;
or (n10256,s0n10256,s1n10256);
not(notn10256,n10005);
and (s0n10256,notn10256,n10239);
and (s1n10256,n10005,n10111);
nor (n10257,n10243,n10149);
and (n10258,n10109,n10259);
and (n10259,n10243,n10148);
nor (n10260,n1036,n1037);
not (n10261,n1035);
or (n10262,n10263,n10264,n10274,n10275);
and (n10263,n9994,n10020);
and (n10264,n10265,n1042);
wire s0n10265,s1n10265,notn10265;
or (n10265,s0n10265,s1n10265);
not(notn10265,n650);
and (s0n10265,notn10265,1'b0);
and (s1n10265,n650,n10266);
or (n10266,1'b0,n10267,n10269,n10272);
and (n10267,n10268,n10073);
wire s0n10268,s1n10268,notn10268;
or (n10268,s0n10268,s1n10268);
not(notn10268,n10259);
and (s0n10268,notn10268,n9996);
and (s1n10268,n10259,1'b1);
and (n10269,n9996,n10270);
not (n10270,n10271);
nand (n10271,n1051,n810);
and (n10272,n10273,n10005);
wire s0n10273,s1n10273,notn10273;
or (n10273,s0n10273,s1n10273);
not(notn10273,n10148);
and (s0n10273,notn10273,n10196);
and (s1n10273,n10148,1'b0);
and (n10274,n10128,n10181);
and (n10275,n10023,n10072);
or (n10276,1'b0,n10277,n10288,n10297,n10349,n10354,n10360,n10368,n10391,n10393);
and (n10277,n10278,n10286);
or (n10278,1'b0,n10279,n10281,n10283);
and (n10279,n10280,n10073);
and (n10281,n10282,n10091);
and (n10283,n10128,n10284);
not (n10284,n10285);
nor (n10285,n10005,n10109);
nor (n10286,n826,n932,n966,n10287);
not (n10287,n1000);
and (n10288,n10289,n10296);
or (n10289,1'b0,n10290,n10292,n10294,n10110);
and (n10290,n10291,n10073);
and (n10292,n10293,n10091);
and (n10294,n10295,n10109);
and (n10296,n826,n932,n966,n10287);
and (n10297,n10298,n10340);
or (n10298,1'b0,n10299,n10300,n10283);
and (n10299,n10111,n10073);
and (n10300,n10301,n10091);
wire s0n10301,s1n10301,notn10301;
or (n10301,s0n10301,s1n10301);
not(notn10301,n10346);
and (s0n10301,notn10301,1'b0);
and (s1n10301,n10346,n10302);
wire s0n10302,s1n10302,notn10302;
or (n10302,s0n10302,s1n10302);
not(notn10302,n51);
and (s0n10302,notn10302,n10303);
and (s1n10302,n51,n10341);
wire s0n10303,s1n10303,notn10303;
or (n10303,s0n10303,s1n10303);
not(notn10303,n10335);
and (s0n10303,notn10303,n10304);
and (s1n10303,n10335,n10306);
wire s0n10304,s1n10304,notn10304;
or (n10304,s0n10304,s1n10304);
not(notn10304,n10020);
and (s0n10304,notn10304,1'b0);
and (s1n10304,n10020,n10305);
or (n10306,n10307,n10314,n10317,n10322,n10329,n10333);
and (n10307,n10308,n10309);
or (n10309,n10310,n10313);
or (n10310,n10311,n10312);
nor (n10311,n38,n39,n59,n56);
nor (n10312,n44,n624,n59,n56);
and (n10313,n44,n39,n60,n56);
and (n10314,n10315,n10316);
and (n10316,n44,n624,n60,n56);
and (n10317,n10318,n10319);
or (n10319,n10320,n10321);
and (n10320,n38,n624,n59,n56);
and (n10321,n38,n39,n60,n56);
and (n10322,n10323,n10324);
or (n10324,n10325,n10328);
or (n10325,n10326,n10327);
nor (n10326,n44,n39,n60,n56);
nor (n10327,n38,n624,n59,n56);
and (n10328,n38,n39,n59,n56);
and (n10329,n10330,n10331);
nor (n10331,n609,n10332,n44);
or (n10332,n10234,n1055);
and (n10333,n10305,n10334);
nor (n10334,n60,n38);
or (n10335,n10336,n10340);
or (n10336,n10337,n10339);
nor (n10337,n826,n932,n10338,n1000);
not (n10338,n966);
and (n10339,n826,n931,n966,n10287);
nor (n10340,n826,n931,n10338,n1000);
wire s0n10341,s1n10341,notn10341;
or (n10341,s0n10341,s1n10341);
not(notn10341,n10345);
and (s0n10341,notn10341,1'b0);
and (s1n10341,n10345,n10342);
wire s0n10342,s1n10342,notn10342;
or (n10342,s0n10342,s1n10342);
not(notn10342,n10170);
and (s0n10342,notn10342,n10343);
and (s1n10342,n10170,n10344);
and (n10345,n51,n10021);
not (n10346,n10347);
nand (n10347,n65,n10348);
or (n10348,n1057,n10140);
and (n10349,n10350,n10339);
or (n10350,1'b0,n10351,n10353);
and (n10351,n10076,n10352);
or (n10352,n10091,n10073);
and (n10353,n10111,n10284);
and (n10354,n10355,n10337);
or (n10355,1'b0,n10356,n10357,n10358);
and (n10356,n10094,n10073);
and (n10357,n10301,n10109);
and (n10358,n10111,n10359);
or (n10359,n10005,n10091);
and (n10360,n10361,n10366);
or (n10361,1'b0,n10362,n10364,n10365,n10110);
and (n10362,n10363,n10073);
and (n10364,n10295,n10091);
and (n10365,n10282,n10109);
nor (n10366,n10367,n931,n966,n1000);
not (n10367,n826);
and (n10368,n10369,n825);
or (n10369,1'b0,n10370,n10389);
and (n10370,n10371,n10109);
or (n10371,n10372,n10383,n10388);
and (n10372,n9996,n10373);
and (n10373,n10374,n10379);
not (n10374,n10375);
and (n10375,n825,n10376);
nor (n10376,n10377,n10150,n38);
not (n10377,n10378);
nor (n10378,n51,n60);
not (n10379,n10380);
and (n10380,n825,n10381);
nor (n10381,n10245,n10382);
nand (n10382,n10207,n619);
and (n10383,n10384,n10385);
wire s0n10384,s1n10384,notn10384;
or (n10384,s0n10384,s1n10384);
not(notn10384,n10379);
and (s0n10384,notn10384,1'b0);
and (s1n10384,n10379,n9996);
or (n10385,n10386,n10387);
and (n10386,n10374,n10380);
nor (n10387,n10374,n10380);
nor (n10388,n10374,n10379);
and (n10389,n10390,n10005);
wire s0n10390,s1n10390,notn10390;
or (n10390,s0n10390,s1n10390);
not(notn10390,n10379);
and (s0n10390,notn10390,1'b0);
and (s1n10390,n10379,n10111);
and (n10391,n10128,n10392);
nor (n10392,n10367,n932,n966,n1000);
and (n10393,n10023,n10394);
nor (n10394,n826,n932,n966,n1000);
and (n10395,n10396,n619);
and (n10396,n926,n65);
wire s0n10397,s1n10397,notn10397;
or (n10397,s0n10397,s1n10397);
not(notn10397,n10395);
and (s0n10397,notn10397,n10398);
and (s1n10397,n10395,n10438);
wire s0n10398,s1n10398,notn10398;
or (n10398,s0n10398,s1n10398);
not(notn10398,n1039);
and (s0n10398,notn10398,n10399);
and (s1n10398,n1039,n10413);
wire s0n10399,s1n10399,notn10399;
or (n10399,s0n10399,s1n10399);
not(notn10399,n10261);
and (s0n10399,notn10399,1'b0);
and (s1n10399,n10261,n10400);
or (n10400,n10401,1'b0,n10406);
and (n10401,n10402,n10021);
wire s0n10402,s1n10402,notn10402;
or (n10402,s0n10402,s1n10402);
not(notn10402,n1057);
and (s0n10402,notn10402,1'b0);
and (s1n10402,n1057,n10403);
wire s0n10403,s1n10403,notn10403;
or (n10403,s0n10403,s1n10403);
not(notn10403,n10004);
and (s0n10403,notn10403,n10404);
and (s1n10403,n10004,n10405);
and (n10406,n10407,n10260);
or (n10407,n10408,n10411,1'b0);
and (n10408,n10409,n10242);
wire s0n10409,s1n10409,notn10409;
or (n10409,s0n10409,s1n10409);
not(notn10409,n10005);
and (s0n10409,notn10409,n10252);
and (s1n10409,n10005,n10410);
wire s0n10410,s1n10410,notn10410;
or (n10410,s0n10410,s1n10410);
not(notn10410,n10241);
and (s0n10410,notn10410,n10094);
and (s1n10410,n10241,1'b0);
and (n10411,n10412,n10257);
wire s0n10412,s1n10412,notn10412;
or (n10412,s0n10412,s1n10412);
not(notn10412,n10005);
and (s0n10412,notn10412,1'b0);
and (s1n10412,n10005,n10094);
or (n10413,n10414,n10419,1'b0);
and (n10414,n10415,n10020);
wire s0n10415,s1n10415,notn10415;
or (n10415,s0n10415,s1n10415);
not(notn10415,n1057);
and (s0n10415,notn10415,1'b0);
and (s1n10415,n1057,n10416);
wire s0n10416,s1n10416,notn10416;
or (n10416,s0n10416,s1n10416);
not(notn10416,n10417);
and (s0n10416,notn10416,n10404);
and (s1n10416,n10417,n10405);
and (n10417,n10418,n44);
and (n10418,n10005,n59);
and (n10419,n10420,n1042);
wire s0n10420,s1n10420,notn10420;
or (n10420,s0n10420,s1n10420);
not(notn10420,n650);
and (s0n10420,notn10420,1'b0);
and (s1n10420,n650,n10421);
or (n10421,1'b0,n10422,n10423,n10425);
and (n10422,n10253,n10352);
and (n10423,n10424,n10109);
wire s0n10424,s1n10424,notn10424;
or (n10424,s0n10424,s1n10424);
not(notn10424,n10243);
and (s0n10424,notn10424,n10101);
and (s1n10424,n10243,1'b0);
and (n10425,n10426,n10005);
wire s0n10426,s1n10426,notn10426;
or (n10426,s0n10426,s1n10426);
not(notn10426,n10148);
and (s0n10426,notn10426,n10427);
and (s1n10426,n10148,1'b0);
nand (n10427,n10428,n10431);
or (n10428,n10429,n10135);
not (n10429,n10430);
nor (n10431,n10432,n10435);
nor (n10432,n10433,n10174);
not (n10433,n10434);
nor (n10435,n10436,n10161);
not (n10436,n10437);
or (n10438,n10439,n10507,n10508,n10514,n10517,n10523,n10525,1'b0);
and (n10439,n10440,n10286);
or (n10440,1'b0,n10441,n10477);
and (n10441,n10442,n10109);
nand (n10442,n10443,n10462);
and (n10443,n10444,n10454,n10458);
nand (n10444,n10445,n10205);
nand (n10445,n10446,n10449);
or (n10446,n10447,n10135);
not (n10447,n10448);
nor (n10449,n10450,n10452);
and (n10450,n10160,n10451);
and (n10452,n10173,n10453);
nor (n10454,n10455,n10457);
and (n10455,n10210,n10456);
and (n10457,n10222,n10451);
nor (n10458,n10459,n10460);
and (n10459,n10228,n10453);
and (n10460,n10231,n10461);
nor (n10462,n10463,n10471,n10474);
and (n10463,n10464,n10177);
nand (n10464,n10465,n10468);
or (n10465,n10466,n10135);
not (n10466,n10467);
nor (n10468,n10469,n10470);
and (n10469,n10160,n10461);
and (n10470,n10173,n10456);
and (n10471,n10472,n10188);
and (n10472,n10136,n10473);
and (n10474,n10475,n10193);
and (n10475,n10136,n10476);
and (n10477,n10478,n10005);
nand (n10478,n10479,n10493);
and (n10479,n10480,n10488,n10489);
nor (n10480,n10481,n10484);
and (n10481,n10482,n10188);
and (n10482,n10136,n10483);
and (n10484,n10485,n10193);
nor (n10485,n10135,n10486);
not (n10486,n10487);
nand (n10488,n10427,n10205);
nor (n10489,n10490,n10491);
and (n10490,n10228,n10434);
and (n10491,n10231,n10492);
nor (n10493,n10494,n10503);
and (n10494,n10495,n10177);
nand (n10495,n10496,n10499);
or (n10496,n10497,n10135);
not (n10497,n10498);
nor (n10499,n10500,n10501);
and (n10500,n10160,n10492);
and (n10501,n10173,n10502);
nand (n10503,n10504,n10505);
or (n10504,n10223,n10436);
or (n10505,n10211,n10506);
not (n10506,n10502);
and (n10507,n10412,n10296);
and (n10508,n10509,n10340);
or (n10509,1'b0,n10510,n10511,n10512,n10513);
and (n10510,n10076,n10073);
and (n10511,n10094,n10091);
and (n10512,n10111,n10109);
and (n10513,n10301,n10005);
and (n10514,n10515,n10339);
or (n10515,1'b0,n10024,n10516,n10513);
and (n10516,n10094,n10270);
and (n10517,n10518,n10337);
or (n10518,1'b0,n10024,n10075,n10093,n10519);
not (n10519,n10520);
or (n10520,n10521,n10522);
not (n10521,n10128);
not (n10522,n10005);
and (n10523,n10524,n10366);
wire s0n10524,s1n10524,notn10524;
or (n10524,s0n10524,s1n10524);
not(notn10524,n10005);
and (s0n10524,notn10524,1'b0);
and (s1n10524,n10005,n10076);
and (n10525,n10526,n825);
or (n10526,1'b0,n10527,n10529);
and (n10527,n10528,n10109);
wire s0n10528,s1n10528,notn10528;
or (n10528,s0n10528,s1n10528);
not(notn10528,n10374);
and (s0n10528,notn10528,1'b0);
and (s1n10528,n10374,n10253);
and (n10529,n10530,n10005);
wire s0n10530,s1n10530,notn10530;
or (n10530,s0n10530,s1n10530);
not(notn10530,n10379);
and (s0n10530,notn10530,1'b0);
and (s1n10530,n10379,n10094);
or (n10531,n10532,n10873,n12914);
and (n10532,n10533,n10740);
wire s0n10533,s1n10533,notn10533;
or (n10533,s0n10533,s1n10533);
not(notn10533,n10395);
and (s0n10533,notn10533,n10534);
and (s1n10533,n10395,n10676);
wire s0n10534,s1n10534,notn10534;
or (n10534,s0n10534,s1n10534);
not(notn10534,n1039);
and (s0n10534,notn10534,n10535);
and (s1n10534,n1039,n10664);
wire s0n10535,s1n10535,notn10535;
or (n10535,s0n10535,s1n10535);
not(notn10535,n10261);
and (s0n10535,notn10535,1'b0);
and (s1n10535,n10261,n10536);
or (n10536,n10537,n10550,n10616,n10653);
and (n10537,n10538,n10021);
wire s0n10538,s1n10538,notn10538;
or (n10538,s0n10538,s1n10538);
not(notn10538,n1057);
and (s0n10538,notn10538,1'b0);
and (s1n10538,n1057,n10539);
wire s0n10539,s1n10539,notn10539;
or (n10539,s0n10539,s1n10539);
not(notn10539,n10004);
and (s0n10539,notn10539,n10540);
and (s1n10539,n10004,n10541);
wire s0n10541,s1n10541,notn10541;
or (n10541,s0n10541,s1n10541);
not(notn10541,n10017);
and (s0n10541,notn10541,n10542);
and (s1n10541,n10017,n10544);
wire s0n10542,s1n10542,notn10542;
or (n10542,s0n10542,s1n10542);
not(notn10542,n10000);
and (s0n10542,notn10542,1'b0);
and (s1n10542,n10000,n10543);
or (n10544,1'b0,n10545,n10547,n10549);
and (n10545,n10546,n10009);
and (n10547,n10548,n10012);
and (n10549,n10543,n10014);
and (n10550,n10551,n10126);
or (n10551,1'b0,n10552,n10568,n10584,n10600);
and (n10552,n10553,n10073);
wire s0n10553,s1n10553,notn10553;
or (n10553,s0n10553,s1n10553);
not(notn10553,n65);
and (s0n10553,notn10553,1'b0);
and (s1n10553,n65,n10554);
wire s0n10554,s1n10554,notn10554;
or (n10554,s0n10554,s1n10554);
not(notn10554,n10068);
and (s0n10554,notn10554,n10555);
and (s1n10554,n10068,n10561);
wire s0n10555,s1n10555,notn10555;
or (n10555,s0n10555,s1n10555);
not(notn10555,n10047);
and (s0n10555,notn10555,1'b0);
and (s1n10555,n10047,n10556);
or (n10556,1'b0,n10557,n10559);
and (n10557,n10558,n10031);
and (n10559,n10560,n10040);
or (n10561,1'b0,n10562,n10564,n10566,n10567);
and (n10562,n10563,n10055);
and (n10564,n10565,n10060);
and (n10566,n10558,n10064);
and (n10567,n10560,n10014);
and (n10568,n10569,n10091);
wire s0n10569,s1n10569,notn10569;
or (n10569,s0n10569,s1n10569);
not(notn10569,n65);
and (s0n10569,notn10569,1'b0);
and (s1n10569,n65,n10570);
wire s0n10570,s1n10570,notn10570;
or (n10570,s0n10570,s1n10570);
not(notn10570,n10068);
and (s0n10570,notn10570,n10571);
and (s1n10570,n10068,n10577);
wire s0n10571,s1n10571,notn10571;
or (n10571,s0n10571,s1n10571);
not(notn10571,n10047);
and (s0n10571,notn10571,1'b0);
and (s1n10571,n10047,n10572);
or (n10572,1'b0,n10573,n10575);
and (n10573,n10574,n10031);
and (n10575,n10576,n10040);
or (n10577,1'b0,n10578,n10580,n10582,n10583);
and (n10578,n10579,n10055);
and (n10580,n10581,n10060);
and (n10582,n10574,n10064);
and (n10583,n10576,n10014);
and (n10584,n10585,n10109);
wire s0n10585,s1n10585,notn10585;
or (n10585,s0n10585,s1n10585);
not(notn10585,n65);
and (s0n10585,notn10585,1'b0);
and (s1n10585,n65,n10586);
wire s0n10586,s1n10586,notn10586;
or (n10586,s0n10586,s1n10586);
not(notn10586,n10068);
and (s0n10586,notn10586,n10587);
and (s1n10586,n10068,n10593);
wire s0n10587,s1n10587,notn10587;
or (n10587,s0n10587,s1n10587);
not(notn10587,n10047);
and (s0n10587,notn10587,1'b0);
and (s1n10587,n10047,n10588);
or (n10588,1'b0,n10589,n10591);
and (n10589,n10590,n10031);
and (n10591,n10592,n10040);
or (n10593,1'b0,n10594,n10596,n10598,n10599);
and (n10594,n10595,n10055);
and (n10596,n10597,n10060);
and (n10598,n10590,n10064);
and (n10599,n10592,n10014);
and (n10600,n10601,n10005);
wire s0n10601,s1n10601,notn10601;
or (n10601,s0n10601,s1n10601);
not(notn10601,n65);
and (s0n10601,notn10601,1'b0);
and (s1n10601,n65,n10602);
wire s0n10602,s1n10602,notn10602;
or (n10602,s0n10602,s1n10602);
not(notn10602,n10068);
and (s0n10602,notn10602,n10603);
and (s1n10602,n10068,n10609);
wire s0n10603,s1n10603,notn10603;
or (n10603,s0n10603,s1n10603);
not(notn10603,n10047);
and (s0n10603,notn10603,1'b0);
and (s1n10603,n10047,n10604);
or (n10604,1'b0,n10605,n10607);
and (n10605,n10606,n10031);
and (n10607,n10608,n10040);
or (n10609,1'b0,n10610,n10612,n10614,n10615);
and (n10610,n10611,n10055);
and (n10612,n10613,n10060);
and (n10614,n10606,n10064);
and (n10615,n10608,n10014);
and (n10616,n10617,n10215);
nand (n10617,n10618,n10638);
nor (n10618,n10619,n10629);
and (n10619,n10620,n10205);
nand (n10620,n10621,n10624);
or (n10621,n10622,n10135);
not (n10622,n10623);
nor (n10624,n10625,n10627);
and (n10625,n10160,n10626);
and (n10627,n10173,n10628);
nand (n10629,n10630,n10633);
nor (n10630,n10631,n10632);
and (n10631,n10228,n10628);
and (n10632,n10222,n10626);
nor (n10633,n10634,n10636);
and (n10634,n10210,n10635);
and (n10636,n10231,n10637);
nor (n10638,n10639,n10647,n10650);
and (n10639,n10640,n10177);
nand (n10640,n10641,n10644);
or (n10641,n10642,n10135);
not (n10642,n10643);
nor (n10644,n10645,n10646);
and (n10645,n10160,n10637);
and (n10646,n10173,n10635);
and (n10647,n10648,n10188);
and (n10648,n10136,n10649);
and (n10650,n10651,n10193);
and (n10651,n10136,n10652);
and (n10653,n10654,n10260);
or (n10654,n10655,n10659,n10662,1'b0);
and (n10655,n10656,n10242);
wire s0n10656,s1n10656,notn10656;
or (n10656,s0n10656,s1n10656);
not(notn10656,n10005);
and (s0n10656,notn10656,n10657);
and (s1n10656,n10005,n10658);
wire s0n10657,s1n10657,notn10657;
or (n10657,s0n10657,s1n10657);
not(notn10657,n10109);
and (s0n10657,notn10657,1'b0);
and (s1n10657,n10109,n10540);
wire s0n10658,s1n10658,notn10658;
or (n10658,s0n10658,s1n10658);
not(notn10658,n10241);
and (s0n10658,notn10658,n10601);
and (s1n10658,n10241,1'b0);
and (n10659,n10660,n10254);
wire s0n10660,s1n10660,notn10660;
or (n10660,s0n10660,s1n10660);
not(notn10660,n10109);
and (s0n10660,notn10660,1'b0);
and (s1n10660,n10109,n10661);
and (n10662,n10663,n10257);
wire s0n10663,s1n10663,notn10663;
or (n10663,s0n10663,s1n10663);
not(notn10663,n10005);
and (s0n10663,notn10663,n10657);
and (s1n10663,n10005,n10601);
or (n10664,n10665,n10666,n10674,n10675);
and (n10665,n10538,n10020);
and (n10666,n10667,n1042);
wire s0n10667,s1n10667,notn10667;
or (n10667,s0n10667,s1n10667);
not(notn10667,n650);
and (s0n10667,notn10667,1'b0);
and (s1n10667,n650,n10668);
or (n10668,1'b0,n10669,n10671,n10672);
and (n10669,n10670,n10073);
wire s0n10670,s1n10670,notn10670;
or (n10670,s0n10670,s1n10670);
not(notn10670,n10259);
and (s0n10670,notn10670,n10540);
and (s1n10670,n10259,1'b0);
and (n10671,n10540,n10270);
and (n10672,n10673,n10005);
wire s0n10673,s1n10673,notn10673;
or (n10673,s0n10673,s1n10673);
not(notn10673,n10148);
and (s0n10673,notn10673,n10620);
and (s1n10673,n10148,1'b0);
and (n10674,n10617,n10181);
and (n10675,n10551,n10072);
or (n10676,1'b0,n10677,n10684,n10692,n10717,n10721,n10726,n10732,n10738,n10739);
and (n10677,n10678,n10286);
or (n10678,1'b0,n10679,n10681,n10683);
and (n10679,n10680,n10073);
and (n10681,n10682,n10091);
and (n10683,n10617,n10284);
and (n10684,n10685,n10296);
or (n10685,1'b0,n10686,n10688,n10690,n10600);
and (n10686,n10687,n10073);
and (n10688,n10689,n10091);
and (n10690,n10691,n10109);
and (n10692,n10693,n10340);
or (n10693,1'b0,n10694,n10695,n10683);
and (n10694,n10601,n10073);
and (n10695,n10696,n10091);
wire s0n10696,s1n10696,notn10696;
or (n10696,s0n10696,s1n10696);
not(notn10696,n10346);
and (s0n10696,notn10696,1'b0);
and (s1n10696,n10346,n10697);
wire s0n10697,s1n10697,notn10697;
or (n10697,s0n10697,s1n10697);
not(notn10697,n51);
and (s0n10697,notn10697,n10698);
and (s1n10697,n51,n10713);
wire s0n10698,s1n10698,notn10698;
or (n10698,s0n10698,s1n10698);
not(notn10698,n10335);
and (s0n10698,notn10698,n10699);
and (s1n10698,n10335,n10701);
wire s0n10699,s1n10699,notn10699;
or (n10699,s0n10699,s1n10699);
not(notn10699,n10020);
and (s0n10699,notn10699,1'b0);
and (s1n10699,n10020,n10700);
or (n10701,n10702,n10704,n10706,n10708,n10710,n10712);
and (n10702,n10703,n10309);
and (n10704,n10705,n10316);
and (n10706,n10707,n10319);
and (n10708,n10709,n10324);
and (n10710,n10711,n10331);
and (n10712,n10700,n10334);
wire s0n10713,s1n10713,notn10713;
or (n10713,s0n10713,s1n10713);
not(notn10713,n10345);
and (s0n10713,notn10713,1'b0);
and (s1n10713,n10345,n10714);
wire s0n10714,s1n10714,notn10714;
or (n10714,s0n10714,s1n10714);
not(notn10714,n10170);
and (s0n10714,notn10714,n10715);
and (s1n10714,n10170,n10716);
and (n10717,n10718,n10339);
or (n10718,1'b0,n10719,n10720);
and (n10719,n10569,n10352);
and (n10720,n10601,n10284);
and (n10721,n10722,n10337);
or (n10722,1'b0,n10723,n10724,n10725);
and (n10723,n10585,n10073);
and (n10724,n10696,n10109);
and (n10725,n10601,n10359);
and (n10726,n10727,n10366);
or (n10727,1'b0,n10728,n10730,n10731,n10600);
and (n10728,n10729,n10073);
and (n10730,n10691,n10091);
and (n10731,n10682,n10109);
and (n10732,n10733,n825);
or (n10733,1'b0,n10734,n10736);
and (n10734,n10735,n10109);
wire s0n10735,s1n10735,notn10735;
or (n10735,s0n10735,s1n10735);
not(notn10735,n10379);
and (s0n10735,notn10735,1'b0);
and (s1n10735,n10379,n10540);
and (n10736,n10737,n10005);
wire s0n10737,s1n10737,notn10737;
or (n10737,s0n10737,s1n10737);
not(notn10737,n10379);
and (s0n10737,notn10737,1'b0);
and (s1n10737,n10379,n10601);
and (n10738,n10617,n10392);
and (n10739,n10551,n10394);
wire s0n10740,s1n10740,notn10740;
or (n10740,s0n10740,s1n10740);
not(notn10740,n10395);
and (s0n10740,notn10740,n10741);
and (s1n10740,n10395,n10779);
wire s0n10741,s1n10741,notn10741;
or (n10741,s0n10741,s1n10741);
not(notn10741,n1039);
and (s0n10741,notn10741,n10742);
and (s1n10741,n1039,n10756);
wire s0n10742,s1n10742,notn10742;
or (n10742,s0n10742,s1n10742);
not(notn10742,n10261);
and (s0n10742,notn10742,1'b0);
and (s1n10742,n10261,n10743);
or (n10743,n10744,1'b0,n10749);
and (n10744,n10745,n10021);
wire s0n10745,s1n10745,notn10745;
or (n10745,s0n10745,s1n10745);
not(notn10745,n1057);
and (s0n10745,notn10745,1'b0);
and (s1n10745,n1057,n10746);
wire s0n10746,s1n10746,notn10746;
or (n10746,s0n10746,s1n10746);
not(notn10746,n10004);
and (s0n10746,notn10746,n10747);
and (s1n10746,n10004,n10748);
and (n10749,n10750,n10260);
or (n10750,n10751,n10754,1'b0);
and (n10751,n10752,n10242);
wire s0n10752,s1n10752,notn10752;
or (n10752,s0n10752,s1n10752);
not(notn10752,n10005);
and (s0n10752,notn10752,n10660);
and (s1n10752,n10005,n10753);
wire s0n10753,s1n10753,notn10753;
or (n10753,s0n10753,s1n10753);
not(notn10753,n10241);
and (s0n10753,notn10753,n10585);
and (s1n10753,n10241,1'b0);
and (n10754,n10755,n10257);
wire s0n10755,s1n10755,notn10755;
or (n10755,s0n10755,s1n10755);
not(notn10755,n10005);
and (s0n10755,notn10755,1'b0);
and (s1n10755,n10005,n10585);
or (n10756,n10757,n10760,1'b0);
and (n10757,n10758,n10020);
wire s0n10758,s1n10758,notn10758;
or (n10758,s0n10758,s1n10758);
not(notn10758,n1057);
and (s0n10758,notn10758,1'b0);
and (s1n10758,n1057,n10759);
wire s0n10759,s1n10759,notn10759;
or (n10759,s0n10759,s1n10759);
not(notn10759,n10417);
and (s0n10759,notn10759,n10747);
and (s1n10759,n10417,n10748);
and (n10760,n10761,n1042);
wire s0n10761,s1n10761,notn10761;
or (n10761,s0n10761,s1n10761);
not(notn10761,n650);
and (s0n10761,notn10761,1'b0);
and (s1n10761,n650,n10762);
or (n10762,1'b0,n10763,n10764,n10766);
and (n10763,n10661,n10352);
and (n10764,n10765,n10109);
wire s0n10765,s1n10765,notn10765;
or (n10765,s0n10765,s1n10765);
not(notn10765,n10243);
and (s0n10765,notn10765,n10592);
and (s1n10765,n10243,1'b0);
and (n10766,n10767,n10005);
wire s0n10767,s1n10767,notn10767;
or (n10767,s0n10767,s1n10767);
not(notn10767,n10148);
and (s0n10767,notn10767,n10768);
and (s1n10767,n10148,1'b0);
nand (n10768,n10769,n10772);
or (n10769,n10770,n10135);
not (n10770,n10771);
nor (n10772,n10773,n10776);
nor (n10773,n10774,n10174);
not (n10774,n10775);
nor (n10776,n10777,n10161);
not (n10777,n10778);
or (n10779,n10780,n10850,n10851,n10857,n10860,n10865,n10867,1'b0);
and (n10780,n10781,n10286);
or (n10781,1'b0,n10782,n10822);
and (n10782,n10783,n10109);
nand (n10783,n10784,n10804);
nor (n10784,n10785,n10795);
and (n10785,n10786,n10205);
nand (n10786,n10787,n10790);
or (n10787,n10788,n10135);
not (n10788,n10789);
nor (n10790,n10791,n10793);
and (n10791,n10160,n10792);
and (n10793,n10173,n10794);
nand (n10795,n10796,n10800);
nor (n10796,n10797,n10798);
and (n10797,n10228,n10794);
and (n10798,n10231,n10799);
nor (n10800,n10801,n10803);
and (n10801,n10210,n10802);
and (n10803,n10222,n10792);
nor (n10804,n10805,n10813);
and (n10805,n10806,n10177);
nand (n10806,n10807,n10810);
or (n10807,n10808,n10135);
not (n10808,n10809);
nor (n10810,n10811,n10812);
and (n10811,n10160,n10799);
and (n10812,n10173,n10802);
not (n10813,n10814);
nor (n10814,n10815,n10818);
and (n10815,n10816,n10188);
and (n10816,n10136,n10817);
and (n10818,n10819,n10193);
nor (n10819,n10135,n10820);
not (n10820,n10821);
and (n10822,n10823,n10005);
nand (n10823,n10824,n10837);
and (n10824,n10825,n10832,n10833);
nor (n10825,n10826,n10829);
and (n10826,n10827,n10188);
and (n10827,n10136,n10828);
and (n10829,n10830,n10193);
and (n10830,n10136,n10831);
nand (n10832,n10768,n10205);
nor (n10833,n10834,n10835);
and (n10834,n10228,n10775);
and (n10835,n10231,n10836);
and (n10837,n10838,n10847);
nand (n10838,n10839,n10177);
nand (n10839,n10840,n10843);
or (n10840,n10841,n10135);
not (n10841,n10842);
nor (n10843,n10844,n10845);
and (n10844,n10160,n10836);
and (n10845,n10173,n10846);
nor (n10847,n10848,n10849);
and (n10848,n10210,n10846);
and (n10849,n10222,n10778);
and (n10850,n10755,n10296);
and (n10851,n10852,n10340);
or (n10852,1'b0,n10853,n10854,n10855,n10856);
and (n10853,n10569,n10073);
and (n10854,n10585,n10091);
and (n10855,n10601,n10109);
and (n10856,n10696,n10005);
and (n10857,n10858,n10339);
or (n10858,1'b0,n10552,n10859,n10856);
and (n10859,n10585,n10270);
and (n10860,n10861,n10337);
or (n10861,1'b0,n10552,n10568,n10584,n10862);
not (n10862,n10863);
or (n10863,n10522,n10864);
not (n10864,n10617);
and (n10865,n10866,n10366);
wire s0n10866,s1n10866,notn10866;
or (n10866,s0n10866,s1n10866);
not(notn10866,n10005);
and (s0n10866,notn10866,1'b0);
and (s1n10866,n10005,n10569);
and (n10867,n10868,n825);
or (n10868,1'b0,n10869,n10871);
and (n10869,n10870,n10109);
wire s0n10870,s1n10870,notn10870;
or (n10870,s0n10870,s1n10870);
not(notn10870,n10374);
and (s0n10870,notn10870,1'b0);
and (s1n10870,n10374,n10661);
and (n10871,n10872,n10005);
wire s0n10872,s1n10872,notn10872;
or (n10872,s0n10872,s1n10872);
not(notn10872,n10379);
and (s0n10872,notn10872,1'b0);
and (s1n10872,n10379,n10585);
and (n10873,n10740,n10874);
or (n10874,n10875,n11213,n12913);
and (n10875,n10876,n11083);
wire s0n10876,s1n10876,notn10876;
or (n10876,s0n10876,s1n10876);
not(notn10876,n10395);
and (s0n10876,notn10876,n10877);
and (s1n10876,n10395,n11019);
wire s0n10877,s1n10877,notn10877;
or (n10877,s0n10877,s1n10877);
not(notn10877,n1039);
and (s0n10877,notn10877,n10878);
and (s1n10877,n1039,n11007);
wire s0n10878,s1n10878,notn10878;
or (n10878,s0n10878,s1n10878);
not(notn10878,n10261);
and (s0n10878,notn10878,1'b0);
and (s1n10878,n10261,n10879);
or (n10879,n10880,n10893,n10959,n10996);
and (n10880,n10881,n10021);
wire s0n10881,s1n10881,notn10881;
or (n10881,s0n10881,s1n10881);
not(notn10881,n1057);
and (s0n10881,notn10881,1'b0);
and (s1n10881,n1057,n10882);
wire s0n10882,s1n10882,notn10882;
or (n10882,s0n10882,s1n10882);
not(notn10882,n10004);
and (s0n10882,notn10882,n10883);
and (s1n10882,n10004,n10884);
wire s0n10884,s1n10884,notn10884;
or (n10884,s0n10884,s1n10884);
not(notn10884,n10017);
and (s0n10884,notn10884,n10885);
and (s1n10884,n10017,n10887);
wire s0n10885,s1n10885,notn10885;
or (n10885,s0n10885,s1n10885);
not(notn10885,n10000);
and (s0n10885,notn10885,1'b0);
and (s1n10885,n10000,n10886);
or (n10887,1'b0,n10888,n10890,n10892);
and (n10888,n10889,n10009);
and (n10890,n10891,n10012);
and (n10892,n10886,n10014);
and (n10893,n10894,n10126);
or (n10894,1'b0,n10895,n10911,n10927,n10943);
and (n10895,n10896,n10073);
wire s0n10896,s1n10896,notn10896;
or (n10896,s0n10896,s1n10896);
not(notn10896,n65);
and (s0n10896,notn10896,1'b0);
and (s1n10896,n65,n10897);
wire s0n10897,s1n10897,notn10897;
or (n10897,s0n10897,s1n10897);
not(notn10897,n10068);
and (s0n10897,notn10897,n10898);
and (s1n10897,n10068,n10904);
wire s0n10898,s1n10898,notn10898;
or (n10898,s0n10898,s1n10898);
not(notn10898,n10047);
and (s0n10898,notn10898,1'b0);
and (s1n10898,n10047,n10899);
or (n10899,1'b0,n10900,n10902);
and (n10900,n10901,n10031);
and (n10902,n10903,n10040);
or (n10904,1'b0,n10905,n10907,n10909,n10910);
and (n10905,n10906,n10055);
and (n10907,n10908,n10060);
and (n10909,n10901,n10064);
and (n10910,n10903,n10014);
and (n10911,n10912,n10091);
wire s0n10912,s1n10912,notn10912;
or (n10912,s0n10912,s1n10912);
not(notn10912,n65);
and (s0n10912,notn10912,1'b0);
and (s1n10912,n65,n10913);
wire s0n10913,s1n10913,notn10913;
or (n10913,s0n10913,s1n10913);
not(notn10913,n10068);
and (s0n10913,notn10913,n10914);
and (s1n10913,n10068,n10920);
wire s0n10914,s1n10914,notn10914;
or (n10914,s0n10914,s1n10914);
not(notn10914,n10047);
and (s0n10914,notn10914,1'b0);
and (s1n10914,n10047,n10915);
or (n10915,1'b0,n10916,n10918);
and (n10916,n10917,n10031);
and (n10918,n10919,n10040);
or (n10920,1'b0,n10921,n10923,n10925,n10926);
and (n10921,n10922,n10055);
and (n10923,n10924,n10060);
and (n10925,n10917,n10064);
and (n10926,n10919,n10014);
and (n10927,n10928,n10109);
wire s0n10928,s1n10928,notn10928;
or (n10928,s0n10928,s1n10928);
not(notn10928,n65);
and (s0n10928,notn10928,1'b0);
and (s1n10928,n65,n10929);
wire s0n10929,s1n10929,notn10929;
or (n10929,s0n10929,s1n10929);
not(notn10929,n10068);
and (s0n10929,notn10929,n10930);
and (s1n10929,n10068,n10936);
wire s0n10930,s1n10930,notn10930;
or (n10930,s0n10930,s1n10930);
not(notn10930,n10047);
and (s0n10930,notn10930,1'b0);
and (s1n10930,n10047,n10931);
or (n10931,1'b0,n10932,n10934);
and (n10932,n10933,n10031);
and (n10934,n10935,n10040);
or (n10936,1'b0,n10937,n10939,n10941,n10942);
and (n10937,n10938,n10055);
and (n10939,n10940,n10060);
and (n10941,n10933,n10064);
and (n10942,n10935,n10014);
and (n10943,n10944,n10005);
wire s0n10944,s1n10944,notn10944;
or (n10944,s0n10944,s1n10944);
not(notn10944,n65);
and (s0n10944,notn10944,1'b0);
and (s1n10944,n65,n10945);
wire s0n10945,s1n10945,notn10945;
or (n10945,s0n10945,s1n10945);
not(notn10945,n10068);
and (s0n10945,notn10945,n10946);
and (s1n10945,n10068,n10952);
wire s0n10946,s1n10946,notn10946;
or (n10946,s0n10946,s1n10946);
not(notn10946,n10047);
and (s0n10946,notn10946,1'b0);
and (s1n10946,n10047,n10947);
or (n10947,1'b0,n10948,n10950);
and (n10948,n10949,n10031);
and (n10950,n10951,n10040);
or (n10952,1'b0,n10953,n10955,n10957,n10958);
and (n10953,n10954,n10055);
and (n10955,n10956,n10060);
and (n10957,n10949,n10064);
and (n10958,n10951,n10014);
and (n10959,n10960,n10215);
nand (n10960,n10961,n10981);
nor (n10961,n10962,n10972);
and (n10962,n10963,n10205);
nand (n10963,n10964,n10967);
or (n10964,n10965,n10135);
not (n10965,n10966);
nor (n10967,n10968,n10970);
and (n10968,n10160,n10969);
and (n10970,n10173,n10971);
nand (n10972,n10973,n10977);
nor (n10973,n10974,n10976);
and (n10974,n10210,n10975);
and (n10976,n10222,n10969);
nor (n10977,n10978,n10979);
and (n10978,n10228,n10971);
and (n10979,n10231,n10980);
nor (n10981,n10982,n10990,n10993);
and (n10982,n10983,n10177);
nand (n10983,n10984,n10987);
or (n10984,n10985,n10135);
not (n10985,n10986);
nor (n10987,n10988,n10989);
and (n10988,n10160,n10980);
and (n10989,n10173,n10975);
and (n10990,n10991,n10188);
and (n10991,n10136,n10992);
and (n10993,n10994,n10193);
and (n10994,n10136,n10995);
and (n10996,n10997,n10260);
or (n10997,n10998,n11002,n11005,1'b0);
and (n10998,n10999,n10242);
wire s0n10999,s1n10999,notn10999;
or (n10999,s0n10999,s1n10999);
not(notn10999,n10005);
and (s0n10999,notn10999,n11000);
and (s1n10999,n10005,n11001);
wire s0n11000,s1n11000,notn11000;
or (n11000,s0n11000,s1n11000);
not(notn11000,n10109);
and (s0n11000,notn11000,1'b0);
and (s1n11000,n10109,n10883);
wire s0n11001,s1n11001,notn11001;
or (n11001,s0n11001,s1n11001);
not(notn11001,n10241);
and (s0n11001,notn11001,n10944);
and (s1n11001,n10241,1'b0);
and (n11002,n11003,n10254);
wire s0n11003,s1n11003,notn11003;
or (n11003,s0n11003,s1n11003);
not(notn11003,n10109);
and (s0n11003,notn11003,1'b0);
and (s1n11003,n10109,n11004);
and (n11005,n11006,n10257);
wire s0n11006,s1n11006,notn11006;
or (n11006,s0n11006,s1n11006);
not(notn11006,n10005);
and (s0n11006,notn11006,n11000);
and (s1n11006,n10005,n10944);
or (n11007,n11008,n11009,n11017,n11018);
and (n11008,n10881,n10020);
and (n11009,n11010,n1042);
wire s0n11010,s1n11010,notn11010;
or (n11010,s0n11010,s1n11010);
not(notn11010,n650);
and (s0n11010,notn11010,1'b0);
and (s1n11010,n650,n11011);
or (n11011,1'b0,n11012,n11014,n11015);
and (n11012,n11013,n10073);
wire s0n11013,s1n11013,notn11013;
or (n11013,s0n11013,s1n11013);
not(notn11013,n10259);
and (s0n11013,notn11013,n10883);
and (s1n11013,n10259,1'b0);
and (n11014,n10883,n10270);
and (n11015,n11016,n10005);
wire s0n11016,s1n11016,notn11016;
or (n11016,s0n11016,s1n11016);
not(notn11016,n10148);
and (s0n11016,notn11016,n10963);
and (s1n11016,n10148,1'b0);
and (n11017,n10960,n10181);
and (n11018,n10894,n10072);
or (n11019,1'b0,n11020,n11027,n11035,n11060,n11064,n11069,n11075,n11081,n11082);
and (n11020,n11021,n10286);
or (n11021,1'b0,n11022,n11024,n11026);
and (n11022,n11023,n10073);
and (n11024,n11025,n10091);
and (n11026,n10960,n10284);
and (n11027,n11028,n10296);
or (n11028,1'b0,n11029,n11031,n11033,n10943);
and (n11029,n11030,n10073);
and (n11031,n11032,n10091);
and (n11033,n11034,n10109);
and (n11035,n11036,n10340);
or (n11036,1'b0,n11037,n11038,n11026);
and (n11037,n10944,n10073);
and (n11038,n11039,n10091);
wire s0n11039,s1n11039,notn11039;
or (n11039,s0n11039,s1n11039);
not(notn11039,n10346);
and (s0n11039,notn11039,1'b0);
and (s1n11039,n10346,n11040);
wire s0n11040,s1n11040,notn11040;
or (n11040,s0n11040,s1n11040);
not(notn11040,n51);
and (s0n11040,notn11040,n11041);
and (s1n11040,n51,n11056);
wire s0n11041,s1n11041,notn11041;
or (n11041,s0n11041,s1n11041);
not(notn11041,n10335);
and (s0n11041,notn11041,n11042);
and (s1n11041,n10335,n11044);
wire s0n11042,s1n11042,notn11042;
or (n11042,s0n11042,s1n11042);
not(notn11042,n10020);
and (s0n11042,notn11042,1'b0);
and (s1n11042,n10020,n11043);
or (n11044,n11045,n11047,n11049,n11051,n11053,n11055);
and (n11045,n11046,n10309);
and (n11047,n11048,n10316);
and (n11049,n11050,n10319);
and (n11051,n11052,n10324);
and (n11053,n11054,n10331);
and (n11055,n11043,n10334);
wire s0n11056,s1n11056,notn11056;
or (n11056,s0n11056,s1n11056);
not(notn11056,n10345);
and (s0n11056,notn11056,1'b0);
and (s1n11056,n10345,n11057);
wire s0n11057,s1n11057,notn11057;
or (n11057,s0n11057,s1n11057);
not(notn11057,n10170);
and (s0n11057,notn11057,n11058);
and (s1n11057,n10170,n11059);
and (n11060,n11061,n10339);
or (n11061,1'b0,n11062,n11063);
and (n11062,n10912,n10352);
and (n11063,n10944,n10284);
and (n11064,n11065,n10337);
or (n11065,1'b0,n11066,n11067,n11068);
and (n11066,n10928,n10073);
and (n11067,n11039,n10109);
and (n11068,n10944,n10359);
and (n11069,n11070,n10366);
or (n11070,1'b0,n11071,n11073,n11074,n10943);
and (n11071,n11072,n10073);
and (n11073,n11034,n10091);
and (n11074,n11025,n10109);
and (n11075,n11076,n825);
or (n11076,1'b0,n11077,n11079);
and (n11077,n11078,n10109);
wire s0n11078,s1n11078,notn11078;
or (n11078,s0n11078,s1n11078);
not(notn11078,n10379);
and (s0n11078,notn11078,1'b0);
and (s1n11078,n10379,n10883);
and (n11079,n11080,n10005);
wire s0n11080,s1n11080,notn11080;
or (n11080,s0n11080,s1n11080);
not(notn11080,n10379);
and (s0n11080,notn11080,1'b0);
and (s1n11080,n10379,n10944);
and (n11081,n10960,n10392);
and (n11082,n10894,n10394);
wire s0n11083,s1n11083,notn11083;
or (n11083,s0n11083,s1n11083);
not(notn11083,n10395);
and (s0n11083,notn11083,n11084);
and (s1n11083,n10395,n11120);
wire s0n11084,s1n11084,notn11084;
or (n11084,s0n11084,s1n11084);
not(notn11084,n1039);
and (s0n11084,notn11084,n11085);
and (s1n11084,n1039,n11099);
wire s0n11085,s1n11085,notn11085;
or (n11085,s0n11085,s1n11085);
not(notn11085,n10261);
and (s0n11085,notn11085,1'b0);
and (s1n11085,n10261,n11086);
or (n11086,n11087,1'b0,n11092);
and (n11087,n11088,n10021);
wire s0n11088,s1n11088,notn11088;
or (n11088,s0n11088,s1n11088);
not(notn11088,n1057);
and (s0n11088,notn11088,1'b0);
and (s1n11088,n1057,n11089);
wire s0n11089,s1n11089,notn11089;
or (n11089,s0n11089,s1n11089);
not(notn11089,n10004);
and (s0n11089,notn11089,n11090);
and (s1n11089,n10004,n11091);
and (n11092,n11093,n10260);
or (n11093,n11094,n11097,1'b0);
and (n11094,n11095,n10242);
wire s0n11095,s1n11095,notn11095;
or (n11095,s0n11095,s1n11095);
not(notn11095,n10005);
and (s0n11095,notn11095,n11003);
and (s1n11095,n10005,n11096);
wire s0n11096,s1n11096,notn11096;
or (n11096,s0n11096,s1n11096);
not(notn11096,n10241);
and (s0n11096,notn11096,n10928);
and (s1n11096,n10241,1'b0);
and (n11097,n11098,n10257);
wire s0n11098,s1n11098,notn11098;
or (n11098,s0n11098,s1n11098);
not(notn11098,n10005);
and (s0n11098,notn11098,1'b0);
and (s1n11098,n10005,n10928);
or (n11099,n11100,n11103,1'b0);
and (n11100,n11101,n10020);
wire s0n11101,s1n11101,notn11101;
or (n11101,s0n11101,s1n11101);
not(notn11101,n1057);
and (s0n11101,notn11101,1'b0);
and (s1n11101,n1057,n11102);
wire s0n11102,s1n11102,notn11102;
or (n11102,s0n11102,s1n11102);
not(notn11102,n10417);
and (s0n11102,notn11102,n11090);
and (s1n11102,n10417,n11091);
and (n11103,n11104,n1042);
wire s0n11104,s1n11104,notn11104;
or (n11104,s0n11104,s1n11104);
not(notn11104,n650);
and (s0n11104,notn11104,1'b0);
and (s1n11104,n650,n11105);
or (n11105,1'b0,n11106,n11107,n11109);
and (n11106,n11004,n10352);
and (n11107,n11108,n10109);
wire s0n11108,s1n11108,notn11108;
or (n11108,s0n11108,s1n11108);
not(notn11108,n10243);
and (s0n11108,notn11108,n10935);
and (s1n11108,n10243,1'b0);
and (n11109,n11110,n10005);
wire s0n11110,s1n11110,notn11110;
or (n11110,s0n11110,s1n11110);
not(notn11110,n10148);
and (s0n11110,notn11110,n11111);
and (s1n11110,n10148,1'b0);
nand (n11111,n11112,n11115);
or (n11112,n11113,n10135);
not (n11113,n11114);
nor (n11115,n11116,n11118);
and (n11116,n10160,n11117);
and (n11118,n10173,n11119);
or (n11120,n11121,n11190,n11191,n11197,n11200,n11205,n11207,1'b0);
and (n11121,n11122,n10286);
or (n11122,1'b0,n11123,n11159);
and (n11123,n11124,n10109);
nand (n11124,n11125,n11147);
and (n11125,n11126,n11136,n11143);
nand (n11126,n11127,n10205);
nand (n11127,n11128,n11131);
or (n11128,n11129,n10135);
not (n11129,n11130);
nor (n11131,n11132,n11134);
and (n11132,n10160,n11133);
and (n11134,n10173,n11135);
nor (n11136,n11137,n11140);
and (n11137,n11138,n10188);
and (n11138,n10136,n11139);
and (n11140,n11141,n10193);
and (n11141,n10136,n11142);
nor (n11143,n11144,n11145);
and (n11144,n10228,n11135);
and (n11145,n10231,n11146);
nor (n11147,n11148,n11157,n11158);
and (n11148,n11149,n10177);
nand (n11149,n11150,n11153);
or (n11150,n11151,n10135);
not (n11151,n11152);
nor (n11153,n11154,n11155);
and (n11154,n10160,n11146);
and (n11155,n10173,n11156);
and (n11157,n10210,n11156);
and (n11158,n10222,n11133);
and (n11159,n11160,n10005);
nand (n11160,n11161,n11176);
and (n11161,n11162,n11163,n11172);
nand (n11162,n11111,n10205);
nor (n11163,n11164,n11168);
and (n11164,n11165,n10188);
nor (n11165,n10135,n11166);
not (n11166,n11167);
and (n11168,n11169,n10193);
nor (n11169,n10135,n11170);
not (n11170,n11171);
nor (n11172,n11173,n11174);
and (n11173,n10228,n11119);
and (n11174,n10231,n11175);
nor (n11176,n11177,n11186);
and (n11177,n11178,n10177);
nand (n11178,n11179,n11182);
or (n11179,n11180,n10135);
not (n11180,n11181);
nor (n11182,n11183,n11184);
and (n11183,n10160,n11175);
and (n11184,n10173,n11185);
not (n11186,n11187);
nor (n11187,n11188,n11189);
and (n11188,n10210,n11185);
and (n11189,n10222,n11117);
and (n11190,n11098,n10296);
and (n11191,n11192,n10340);
or (n11192,1'b0,n11193,n11194,n11195,n11196);
and (n11193,n10912,n10073);
and (n11194,n10928,n10091);
and (n11195,n10944,n10109);
and (n11196,n11039,n10005);
and (n11197,n11198,n10339);
or (n11198,1'b0,n10895,n11199,n11196);
and (n11199,n10928,n10270);
and (n11200,n11201,n10337);
or (n11201,1'b0,n10895,n10911,n10927,n11202);
not (n11202,n11203);
or (n11203,n10522,n11204);
not (n11204,n10960);
and (n11205,n11206,n10366);
wire s0n11206,s1n11206,notn11206;
or (n11206,s0n11206,s1n11206);
not(notn11206,n10005);
and (s0n11206,notn11206,1'b0);
and (s1n11206,n10005,n10912);
and (n11207,n11208,n825);
or (n11208,1'b0,n11209,n11211);
and (n11209,n11210,n10109);
wire s0n11210,s1n11210,notn11210;
or (n11210,s0n11210,s1n11210);
not(notn11210,n10374);
and (s0n11210,notn11210,1'b0);
and (s1n11210,n10374,n11004);
and (n11211,n11212,n10005);
wire s0n11212,s1n11212,notn11212;
or (n11212,s0n11212,s1n11212);
not(notn11212,n10379);
and (s0n11212,notn11212,1'b0);
and (s1n11212,n10379,n10928);
and (n11213,n11083,n11214);
or (n11214,n11215,n11557,n12912);
and (n11215,n11216,n11425);
wire s0n11216,s1n11216,notn11216;
or (n11216,s0n11216,s1n11216);
not(notn11216,n10395);
and (s0n11216,notn11216,n11217);
and (s1n11216,n10395,n11361);
wire s0n11217,s1n11217,notn11217;
or (n11217,s0n11217,s1n11217);
not(notn11217,n1039);
and (s0n11217,notn11217,n11218);
and (s1n11217,n1039,n11349);
wire s0n11218,s1n11218,notn11218;
or (n11218,s0n11218,s1n11218);
not(notn11218,n10261);
and (s0n11218,notn11218,1'b0);
and (s1n11218,n10261,n11219);
or (n11219,n11220,n11233,n11299,n11338);
and (n11220,n11221,n10021);
wire s0n11221,s1n11221,notn11221;
or (n11221,s0n11221,s1n11221);
not(notn11221,n1057);
and (s0n11221,notn11221,1'b0);
and (s1n11221,n1057,n11222);
wire s0n11222,s1n11222,notn11222;
or (n11222,s0n11222,s1n11222);
not(notn11222,n10004);
and (s0n11222,notn11222,n11223);
and (s1n11222,n10004,n11224);
wire s0n11224,s1n11224,notn11224;
or (n11224,s0n11224,s1n11224);
not(notn11224,n10017);
and (s0n11224,notn11224,n11225);
and (s1n11224,n10017,n11227);
wire s0n11225,s1n11225,notn11225;
or (n11225,s0n11225,s1n11225);
not(notn11225,n10000);
and (s0n11225,notn11225,1'b0);
and (s1n11225,n10000,n11226);
or (n11227,1'b0,n11228,n11230,n11232);
and (n11228,n11229,n10009);
and (n11230,n11231,n10012);
and (n11232,n11226,n10014);
and (n11233,n11234,n10126);
or (n11234,1'b0,n11235,n11251,n11267,n11283);
and (n11235,n11236,n10073);
wire s0n11236,s1n11236,notn11236;
or (n11236,s0n11236,s1n11236);
not(notn11236,n65);
and (s0n11236,notn11236,1'b0);
and (s1n11236,n65,n11237);
wire s0n11237,s1n11237,notn11237;
or (n11237,s0n11237,s1n11237);
not(notn11237,n10068);
and (s0n11237,notn11237,n11238);
and (s1n11237,n10068,n11244);
wire s0n11238,s1n11238,notn11238;
or (n11238,s0n11238,s1n11238);
not(notn11238,n10047);
and (s0n11238,notn11238,1'b0);
and (s1n11238,n10047,n11239);
or (n11239,1'b0,n11240,n11242);
and (n11240,n11241,n10031);
and (n11242,n11243,n10040);
or (n11244,1'b0,n11245,n11247,n11249,n11250);
and (n11245,n11246,n10055);
and (n11247,n11248,n10060);
and (n11249,n11241,n10064);
and (n11250,n11243,n10014);
and (n11251,n11252,n10091);
wire s0n11252,s1n11252,notn11252;
or (n11252,s0n11252,s1n11252);
not(notn11252,n65);
and (s0n11252,notn11252,1'b0);
and (s1n11252,n65,n11253);
wire s0n11253,s1n11253,notn11253;
or (n11253,s0n11253,s1n11253);
not(notn11253,n10068);
and (s0n11253,notn11253,n11254);
and (s1n11253,n10068,n11260);
wire s0n11254,s1n11254,notn11254;
or (n11254,s0n11254,s1n11254);
not(notn11254,n10047);
and (s0n11254,notn11254,1'b0);
and (s1n11254,n10047,n11255);
or (n11255,1'b0,n11256,n11258);
and (n11256,n11257,n10031);
and (n11258,n11259,n10040);
or (n11260,1'b0,n11261,n11263,n11265,n11266);
and (n11261,n11262,n10055);
and (n11263,n11264,n10060);
and (n11265,n11257,n10064);
and (n11266,n11259,n10014);
and (n11267,n11268,n10109);
wire s0n11268,s1n11268,notn11268;
or (n11268,s0n11268,s1n11268);
not(notn11268,n65);
and (s0n11268,notn11268,1'b0);
and (s1n11268,n65,n11269);
wire s0n11269,s1n11269,notn11269;
or (n11269,s0n11269,s1n11269);
not(notn11269,n10068);
and (s0n11269,notn11269,n11270);
and (s1n11269,n10068,n11276);
wire s0n11270,s1n11270,notn11270;
or (n11270,s0n11270,s1n11270);
not(notn11270,n10047);
and (s0n11270,notn11270,1'b0);
and (s1n11270,n10047,n11271);
or (n11271,1'b0,n11272,n11274);
and (n11272,n11273,n10031);
and (n11274,n11275,n10040);
or (n11276,1'b0,n11277,n11279,n11281,n11282);
and (n11277,n11278,n10055);
and (n11279,n11280,n10060);
and (n11281,n11273,n10064);
and (n11282,n11275,n10014);
and (n11283,n11284,n10005);
wire s0n11284,s1n11284,notn11284;
or (n11284,s0n11284,s1n11284);
not(notn11284,n65);
and (s0n11284,notn11284,1'b0);
and (s1n11284,n65,n11285);
wire s0n11285,s1n11285,notn11285;
or (n11285,s0n11285,s1n11285);
not(notn11285,n10068);
and (s0n11285,notn11285,n11286);
and (s1n11285,n10068,n11292);
wire s0n11286,s1n11286,notn11286;
or (n11286,s0n11286,s1n11286);
not(notn11286,n10047);
and (s0n11286,notn11286,1'b0);
and (s1n11286,n10047,n11287);
or (n11287,1'b0,n11288,n11290);
and (n11288,n11289,n10031);
and (n11290,n11291,n10040);
or (n11292,1'b0,n11293,n11295,n11297,n11298);
and (n11293,n11294,n10055);
and (n11295,n11296,n10060);
and (n11297,n11289,n10064);
and (n11298,n11291,n10014);
and (n11299,n11300,n10215);
nand (n11300,n11301,n11320);
and (n11301,n11302,n11312,n11316);
nand (n11302,n11303,n10205);
nand (n11303,n11304,n11307);
or (n11304,n11305,n10135);
not (n11305,n11306);
nor (n11307,n11308,n11310);
and (n11308,n10160,n11309);
and (n11310,n10173,n11311);
nor (n11312,n11313,n11315);
and (n11313,n10210,n11314);
and (n11315,n10222,n11309);
nor (n11316,n11317,n11318);
and (n11317,n10228,n11311);
and (n11318,n10231,n11319);
nor (n11320,n11321,n11329);
and (n11321,n11322,n10177);
nand (n11322,n11323,n11326);
or (n11323,n11324,n10135);
not (n11324,n11325);
nor (n11326,n11327,n11328);
and (n11327,n10160,n11319);
and (n11328,n10173,n11314);
nand (n11329,n11330,n11335);
or (n11330,n11331,n11332);
not (n11331,n10193);
not (n11332,n11333);
and (n11333,n10136,n11334);
nand (n11335,n11336,n10188);
and (n11336,n10136,n11337);
and (n11338,n11339,n10260);
or (n11339,n11340,n11344,n11347,1'b0);
and (n11340,n11341,n10242);
wire s0n11341,s1n11341,notn11341;
or (n11341,s0n11341,s1n11341);
not(notn11341,n10005);
and (s0n11341,notn11341,n11342);
and (s1n11341,n10005,n11343);
wire s0n11342,s1n11342,notn11342;
or (n11342,s0n11342,s1n11342);
not(notn11342,n10109);
and (s0n11342,notn11342,1'b0);
and (s1n11342,n10109,n11223);
wire s0n11343,s1n11343,notn11343;
or (n11343,s0n11343,s1n11343);
not(notn11343,n10241);
and (s0n11343,notn11343,n11284);
and (s1n11343,n10241,1'b0);
and (n11344,n11345,n10254);
wire s0n11345,s1n11345,notn11345;
or (n11345,s0n11345,s1n11345);
not(notn11345,n10109);
and (s0n11345,notn11345,1'b0);
and (s1n11345,n10109,n11346);
and (n11347,n11348,n10257);
wire s0n11348,s1n11348,notn11348;
or (n11348,s0n11348,s1n11348);
not(notn11348,n10005);
and (s0n11348,notn11348,n11342);
and (s1n11348,n10005,n11284);
or (n11349,n11350,n11351,n11359,n11360);
and (n11350,n11221,n10020);
and (n11351,n11352,n1042);
wire s0n11352,s1n11352,notn11352;
or (n11352,s0n11352,s1n11352);
not(notn11352,n650);
and (s0n11352,notn11352,1'b0);
and (s1n11352,n650,n11353);
or (n11353,1'b0,n11354,n11356,n11357);
and (n11354,n11355,n10073);
wire s0n11355,s1n11355,notn11355;
or (n11355,s0n11355,s1n11355);
not(notn11355,n10259);
and (s0n11355,notn11355,n11223);
and (s1n11355,n10259,1'b0);
and (n11356,n11223,n10270);
and (n11357,n11358,n10005);
wire s0n11358,s1n11358,notn11358;
or (n11358,s0n11358,s1n11358);
not(notn11358,n10148);
and (s0n11358,notn11358,n11303);
and (s1n11358,n10148,1'b0);
and (n11359,n11300,n10181);
and (n11360,n11234,n10072);
or (n11361,1'b0,n11362,n11369,n11377,n11402,n11406,n11411,n11417,n11423,n11424);
and (n11362,n11363,n10286);
or (n11363,1'b0,n11364,n11366,n11368);
and (n11364,n11365,n10073);
and (n11366,n11367,n10091);
and (n11368,n11300,n10284);
and (n11369,n11370,n10296);
or (n11370,1'b0,n11371,n11373,n11375,n11283);
and (n11371,n11372,n10073);
and (n11373,n11374,n10091);
and (n11375,n11376,n10109);
and (n11377,n11378,n10340);
or (n11378,1'b0,n11379,n11380,n11368);
and (n11379,n11284,n10073);
and (n11380,n11381,n10091);
wire s0n11381,s1n11381,notn11381;
or (n11381,s0n11381,s1n11381);
not(notn11381,n10346);
and (s0n11381,notn11381,1'b0);
and (s1n11381,n10346,n11382);
wire s0n11382,s1n11382,notn11382;
or (n11382,s0n11382,s1n11382);
not(notn11382,n51);
and (s0n11382,notn11382,n11383);
and (s1n11382,n51,n11398);
wire s0n11383,s1n11383,notn11383;
or (n11383,s0n11383,s1n11383);
not(notn11383,n10335);
and (s0n11383,notn11383,n11384);
and (s1n11383,n10335,n11386);
wire s0n11384,s1n11384,notn11384;
or (n11384,s0n11384,s1n11384);
not(notn11384,n10020);
and (s0n11384,notn11384,1'b0);
and (s1n11384,n10020,n11385);
or (n11386,n11387,n11389,n11391,n11393,n11395,n11397);
and (n11387,n11388,n10309);
and (n11389,n11390,n10316);
and (n11391,n11392,n10319);
and (n11393,n11394,n10324);
and (n11395,n11396,n10331);
and (n11397,n11385,n10334);
wire s0n11398,s1n11398,notn11398;
or (n11398,s0n11398,s1n11398);
not(notn11398,n10345);
and (s0n11398,notn11398,1'b0);
and (s1n11398,n10345,n11399);
wire s0n11399,s1n11399,notn11399;
or (n11399,s0n11399,s1n11399);
not(notn11399,n10170);
and (s0n11399,notn11399,n11400);
and (s1n11399,n10170,n11401);
and (n11402,n11403,n10339);
or (n11403,1'b0,n11404,n11405);
and (n11404,n11252,n10352);
and (n11405,n11284,n10284);
and (n11406,n11407,n10337);
or (n11407,1'b0,n11408,n11409,n11410);
and (n11408,n11268,n10073);
and (n11409,n11381,n10109);
and (n11410,n11284,n10359);
and (n11411,n11412,n10366);
or (n11412,1'b0,n11413,n11415,n11416,n11283);
and (n11413,n11414,n10073);
and (n11415,n11376,n10091);
and (n11416,n11367,n10109);
and (n11417,n11418,n825);
or (n11418,1'b0,n11419,n11421);
and (n11419,n11420,n10109);
wire s0n11420,s1n11420,notn11420;
or (n11420,s0n11420,s1n11420);
not(notn11420,n10379);
and (s0n11420,notn11420,1'b0);
and (s1n11420,n10379,n11223);
and (n11421,n11422,n10005);
wire s0n11422,s1n11422,notn11422;
or (n11422,s0n11422,s1n11422);
not(notn11422,n10379);
and (s0n11422,notn11422,1'b0);
and (s1n11422,n10379,n11284);
and (n11423,n11300,n10392);
and (n11424,n11234,n10394);
wire s0n11425,s1n11425,notn11425;
or (n11425,s0n11425,s1n11425);
not(notn11425,n10395);
and (s0n11425,notn11425,n11426);
and (s1n11425,n10395,n11462);
wire s0n11426,s1n11426,notn11426;
or (n11426,s0n11426,s1n11426);
not(notn11426,n1039);
and (s0n11426,notn11426,n11427);
and (s1n11426,n1039,n11441);
wire s0n11427,s1n11427,notn11427;
or (n11427,s0n11427,s1n11427);
not(notn11427,n10261);
and (s0n11427,notn11427,1'b0);
and (s1n11427,n10261,n11428);
or (n11428,n11429,1'b0,n11434);
and (n11429,n11430,n10021);
wire s0n11430,s1n11430,notn11430;
or (n11430,s0n11430,s1n11430);
not(notn11430,n1057);
and (s0n11430,notn11430,1'b0);
and (s1n11430,n1057,n11431);
wire s0n11431,s1n11431,notn11431;
or (n11431,s0n11431,s1n11431);
not(notn11431,n10004);
and (s0n11431,notn11431,n11432);
and (s1n11431,n10004,n11433);
and (n11434,n11435,n10260);
or (n11435,n11436,n11439,1'b0);
and (n11436,n11437,n10242);
wire s0n11437,s1n11437,notn11437;
or (n11437,s0n11437,s1n11437);
not(notn11437,n10005);
and (s0n11437,notn11437,n11345);
and (s1n11437,n10005,n11438);
wire s0n11438,s1n11438,notn11438;
or (n11438,s0n11438,s1n11438);
not(notn11438,n10241);
and (s0n11438,notn11438,n11268);
and (s1n11438,n10241,1'b0);
and (n11439,n11440,n10257);
wire s0n11440,s1n11440,notn11440;
or (n11440,s0n11440,s1n11440);
not(notn11440,n10005);
and (s0n11440,notn11440,1'b0);
and (s1n11440,n10005,n11268);
or (n11441,n11442,n11445,1'b0);
and (n11442,n11443,n10020);
wire s0n11443,s1n11443,notn11443;
or (n11443,s0n11443,s1n11443);
not(notn11443,n1057);
and (s0n11443,notn11443,1'b0);
and (s1n11443,n1057,n11444);
wire s0n11444,s1n11444,notn11444;
or (n11444,s0n11444,s1n11444);
not(notn11444,n10417);
and (s0n11444,notn11444,n11432);
and (s1n11444,n10417,n11433);
and (n11445,n11446,n1042);
wire s0n11446,s1n11446,notn11446;
or (n11446,s0n11446,s1n11446);
not(notn11446,n650);
and (s0n11446,notn11446,1'b0);
and (s1n11446,n650,n11447);
or (n11447,1'b0,n11448,n11449,n11451);
and (n11448,n11346,n10352);
and (n11449,n11450,n10109);
wire s0n11450,s1n11450,notn11450;
or (n11450,s0n11450,s1n11450);
not(notn11450,n10243);
and (s0n11450,notn11450,n11275);
and (s1n11450,n10243,1'b0);
and (n11451,n11452,n10005);
wire s0n11452,s1n11452,notn11452;
or (n11452,s0n11452,s1n11452);
not(notn11452,n10148);
and (s0n11452,notn11452,n11453);
and (s1n11452,n10148,1'b0);
nand (n11453,n11454,n11457);
or (n11454,n11455,n10135);
not (n11455,n11456);
nor (n11457,n11458,n11460);
and (n11458,n10160,n11459);
and (n11460,n10173,n11461);
or (n11462,n11463,n11534,n11535,n11541,n11544,n11549,n11551,1'b0);
and (n11463,n11464,n10286);
or (n11464,1'b0,n11465,n11503);
and (n11465,n11466,n10109);
nand (n11466,n11467,n11489);
and (n11467,n11468,n11478,n11485);
nand (n11468,n11469,n10205);
nand (n11469,n11470,n11473);
or (n11470,n11471,n10135);
not (n11471,n11472);
nor (n11473,n11474,n11476);
and (n11474,n10160,n11475);
and (n11476,n10173,n11477);
nor (n11478,n11479,n11482);
and (n11479,n11480,n10188);
and (n11480,n10136,n11481);
and (n11482,n11483,n10193);
and (n11483,n10136,n11484);
nor (n11485,n11486,n11487);
and (n11486,n10228,n11477);
and (n11487,n10231,n11488);
nor (n11489,n11490,n11499);
and (n11490,n11491,n10177);
nand (n11491,n11492,n11495);
or (n11492,n11493,n10135);
not (n11493,n11494);
nor (n11495,n11496,n11497);
and (n11496,n10160,n11488);
and (n11497,n10173,n11498);
not (n11499,n11500);
nor (n11500,n11501,n11502);
and (n11501,n10210,n11498);
and (n11502,n10222,n11475);
and (n11503,n11504,n10005);
nand (n11504,n11505,n11520);
nor (n11505,n11506,n11507);
and (n11506,n11453,n10205);
nand (n11507,n11508,n11512,n11516);
nand (n11508,n11509,n10188);
nor (n11509,n10135,n11510);
not (n11510,n11511);
nand (n11512,n11513,n10193);
nor (n11513,n10135,n11514);
not (n11514,n11515);
nor (n11516,n11517,n11518);
and (n11517,n10228,n11461);
and (n11518,n10231,n11519);
nor (n11520,n11521,n11530);
and (n11521,n11522,n10177);
nand (n11522,n11523,n11526);
or (n11523,n11524,n10135);
not (n11524,n11525);
nor (n11526,n11527,n11528);
and (n11527,n10160,n11519);
and (n11528,n10173,n11529);
nand (n11530,n11531,n11533);
or (n11531,n11532,n10223);
not (n11532,n11459);
nand (n11533,n10210,n11529);
and (n11534,n11440,n10296);
and (n11535,n11536,n10340);
or (n11536,1'b0,n11537,n11538,n11539,n11540);
and (n11537,n11252,n10073);
and (n11538,n11268,n10091);
and (n11539,n11284,n10109);
and (n11540,n11381,n10005);
and (n11541,n11542,n10339);
or (n11542,1'b0,n11235,n11543,n11540);
and (n11543,n11268,n10270);
and (n11544,n11545,n10337);
or (n11545,1'b0,n11235,n11251,n11267,n11546);
not (n11546,n11547);
or (n11547,n10522,n11548);
not (n11548,n11300);
and (n11549,n11550,n10366);
wire s0n11550,s1n11550,notn11550;
or (n11550,s0n11550,s1n11550);
not(notn11550,n10005);
and (s0n11550,notn11550,1'b0);
and (s1n11550,n10005,n11252);
and (n11551,n11552,n825);
or (n11552,1'b0,n11553,n11555);
and (n11553,n11554,n10109);
wire s0n11554,s1n11554,notn11554;
or (n11554,s0n11554,s1n11554);
not(notn11554,n10374);
and (s0n11554,notn11554,1'b0);
and (s1n11554,n10374,n11346);
and (n11555,n11556,n10005);
wire s0n11556,s1n11556,notn11556;
or (n11556,s0n11556,s1n11556);
not(notn11556,n10379);
and (s0n11556,notn11556,1'b0);
and (s1n11556,n10379,n11268);
and (n11557,n11425,n11558);
or (n11558,n11559,n11891,n12911);
and (n11559,n11560,n11768);
wire s0n11560,s1n11560,notn11560;
or (n11560,s0n11560,s1n11560);
not(notn11560,n10395);
and (s0n11560,notn11560,n11561);
and (s1n11560,n10395,n11704);
wire s0n11561,s1n11561,notn11561;
or (n11561,s0n11561,s1n11561);
not(notn11561,n1039);
and (s0n11561,notn11561,n11562);
and (s1n11561,n1039,n11692);
wire s0n11562,s1n11562,notn11562;
or (n11562,s0n11562,s1n11562);
not(notn11562,n10261);
and (s0n11562,notn11562,1'b0);
and (s1n11562,n10261,n11563);
or (n11563,n11564,n11577,n11643,n11681);
and (n11564,n11565,n10021);
wire s0n11565,s1n11565,notn11565;
or (n11565,s0n11565,s1n11565);
not(notn11565,n1057);
and (s0n11565,notn11565,1'b0);
and (s1n11565,n1057,n11566);
wire s0n11566,s1n11566,notn11566;
or (n11566,s0n11566,s1n11566);
not(notn11566,n10004);
and (s0n11566,notn11566,n11567);
and (s1n11566,n10004,n11568);
wire s0n11568,s1n11568,notn11568;
or (n11568,s0n11568,s1n11568);
not(notn11568,n10017);
and (s0n11568,notn11568,n11569);
and (s1n11568,n10017,n11571);
wire s0n11569,s1n11569,notn11569;
or (n11569,s0n11569,s1n11569);
not(notn11569,n10000);
and (s0n11569,notn11569,1'b0);
and (s1n11569,n10000,n11570);
or (n11571,1'b0,n11572,n11574,n11576);
and (n11572,n11573,n10009);
and (n11574,n11575,n10012);
and (n11576,n11570,n10014);
and (n11577,n11578,n10126);
or (n11578,1'b0,n11579,n11595,n11611,n11627);
and (n11579,n11580,n10073);
wire s0n11580,s1n11580,notn11580;
or (n11580,s0n11580,s1n11580);
not(notn11580,n65);
and (s0n11580,notn11580,1'b0);
and (s1n11580,n65,n11581);
wire s0n11581,s1n11581,notn11581;
or (n11581,s0n11581,s1n11581);
not(notn11581,n10068);
and (s0n11581,notn11581,n11582);
and (s1n11581,n10068,n11588);
wire s0n11582,s1n11582,notn11582;
or (n11582,s0n11582,s1n11582);
not(notn11582,n10047);
and (s0n11582,notn11582,1'b0);
and (s1n11582,n10047,n11583);
or (n11583,1'b0,n11584,n11586);
and (n11584,n11585,n10031);
and (n11586,n11587,n10040);
or (n11588,1'b0,n11589,n11591,n11593,n11594);
and (n11589,n11590,n10055);
and (n11591,n11592,n10060);
and (n11593,n11585,n10064);
and (n11594,n11587,n10014);
and (n11595,n11596,n10091);
wire s0n11596,s1n11596,notn11596;
or (n11596,s0n11596,s1n11596);
not(notn11596,n65);
and (s0n11596,notn11596,1'b0);
and (s1n11596,n65,n11597);
wire s0n11597,s1n11597,notn11597;
or (n11597,s0n11597,s1n11597);
not(notn11597,n10068);
and (s0n11597,notn11597,n11598);
and (s1n11597,n10068,n11604);
wire s0n11598,s1n11598,notn11598;
or (n11598,s0n11598,s1n11598);
not(notn11598,n10047);
and (s0n11598,notn11598,1'b0);
and (s1n11598,n10047,n11599);
or (n11599,1'b0,n11600,n11602);
and (n11600,n11601,n10031);
and (n11602,n11603,n10040);
or (n11604,1'b0,n11605,n11607,n11609,n11610);
and (n11605,n11606,n10055);
and (n11607,n11608,n10060);
and (n11609,n11601,n10064);
and (n11610,n11603,n10014);
and (n11611,n11612,n10109);
wire s0n11612,s1n11612,notn11612;
or (n11612,s0n11612,s1n11612);
not(notn11612,n65);
and (s0n11612,notn11612,1'b0);
and (s1n11612,n65,n11613);
wire s0n11613,s1n11613,notn11613;
or (n11613,s0n11613,s1n11613);
not(notn11613,n10068);
and (s0n11613,notn11613,n11614);
and (s1n11613,n10068,n11620);
wire s0n11614,s1n11614,notn11614;
or (n11614,s0n11614,s1n11614);
not(notn11614,n10047);
and (s0n11614,notn11614,1'b0);
and (s1n11614,n10047,n11615);
or (n11615,1'b0,n11616,n11618);
and (n11616,n11617,n10031);
and (n11618,n11619,n10040);
or (n11620,1'b0,n11621,n11623,n11625,n11626);
and (n11621,n11622,n10055);
and (n11623,n11624,n10060);
and (n11625,n11617,n10064);
and (n11626,n11619,n10014);
and (n11627,n11628,n10005);
wire s0n11628,s1n11628,notn11628;
or (n11628,s0n11628,s1n11628);
not(notn11628,n65);
and (s0n11628,notn11628,1'b0);
and (s1n11628,n65,n11629);
wire s0n11629,s1n11629,notn11629;
or (n11629,s0n11629,s1n11629);
not(notn11629,n10068);
and (s0n11629,notn11629,n11630);
and (s1n11629,n10068,n11636);
wire s0n11630,s1n11630,notn11630;
or (n11630,s0n11630,s1n11630);
not(notn11630,n10047);
and (s0n11630,notn11630,1'b0);
and (s1n11630,n10047,n11631);
or (n11631,1'b0,n11632,n11634);
and (n11632,n11633,n10031);
and (n11634,n11635,n10040);
or (n11636,1'b0,n11637,n11639,n11641,n11642);
and (n11637,n11638,n10055);
and (n11639,n11640,n10060);
and (n11641,n11633,n10064);
and (n11642,n11635,n10014);
and (n11643,n11644,n10215);
nand (n11644,n11645,n11667);
nor (n11645,n11646,n11656);
and (n11646,n11647,n10205);
nand (n11647,n11648,n11651);
or (n11648,n11649,n10135);
not (n11649,n11650);
nor (n11651,n11652,n11654);
and (n11652,n10160,n11653);
and (n11654,n10173,n11655);
nand (n11656,n11657,n11660,n11663);
nand (n11657,n11658,n10188);
and (n11658,n10136,n11659);
nand (n11660,n11661,n10193);
and (n11661,n10136,n11662);
nor (n11663,n11664,n11665);
and (n11664,n10228,n11655);
and (n11665,n10231,n11666);
nor (n11667,n11668,n11677);
and (n11668,n11669,n10177);
nand (n11669,n11670,n11673);
or (n11670,n11671,n10135);
not (n11671,n11672);
nor (n11673,n11674,n11675);
and (n11674,n10160,n11666);
and (n11675,n10173,n11676);
not (n11677,n11678);
nor (n11678,n11679,n11680);
and (n11679,n10210,n11676);
and (n11680,n10222,n11653);
and (n11681,n11682,n10260);
or (n11682,n11683,n11687,n11690,1'b0);
and (n11683,n11684,n10242);
wire s0n11684,s1n11684,notn11684;
or (n11684,s0n11684,s1n11684);
not(notn11684,n10005);
and (s0n11684,notn11684,n11685);
and (s1n11684,n10005,n11686);
wire s0n11685,s1n11685,notn11685;
or (n11685,s0n11685,s1n11685);
not(notn11685,n10109);
and (s0n11685,notn11685,1'b0);
and (s1n11685,n10109,n11567);
wire s0n11686,s1n11686,notn11686;
or (n11686,s0n11686,s1n11686);
not(notn11686,n10241);
and (s0n11686,notn11686,n11628);
and (s1n11686,n10241,1'b0);
and (n11687,n11688,n10254);
wire s0n11688,s1n11688,notn11688;
or (n11688,s0n11688,s1n11688);
not(notn11688,n10109);
and (s0n11688,notn11688,1'b0);
and (s1n11688,n10109,n11689);
and (n11690,n11691,n10257);
wire s0n11691,s1n11691,notn11691;
or (n11691,s0n11691,s1n11691);
not(notn11691,n10005);
and (s0n11691,notn11691,n11685);
and (s1n11691,n10005,n11628);
or (n11692,n11693,n11694,n11702,n11703);
and (n11693,n11565,n10020);
and (n11694,n11695,n1042);
wire s0n11695,s1n11695,notn11695;
or (n11695,s0n11695,s1n11695);
not(notn11695,n650);
and (s0n11695,notn11695,1'b0);
and (s1n11695,n650,n11696);
or (n11696,1'b0,n11697,n11699,n11700);
and (n11697,n11698,n10073);
wire s0n11698,s1n11698,notn11698;
or (n11698,s0n11698,s1n11698);
not(notn11698,n10259);
and (s0n11698,notn11698,n11567);
and (s1n11698,n10259,1'b0);
and (n11699,n11567,n10270);
and (n11700,n11701,n10005);
wire s0n11701,s1n11701,notn11701;
or (n11701,s0n11701,s1n11701);
not(notn11701,n10148);
and (s0n11701,notn11701,n11647);
and (s1n11701,n10148,1'b0);
and (n11702,n11644,n10181);
and (n11703,n11578,n10072);
or (n11704,1'b0,n11705,n11712,n11720,n11745,n11749,n11754,n11760,n11766,n11767);
and (n11705,n11706,n10286);
or (n11706,1'b0,n11707,n11709,n11711);
and (n11707,n11708,n10073);
and (n11709,n11710,n10091);
and (n11711,n11644,n10284);
and (n11712,n11713,n10296);
or (n11713,1'b0,n11714,n11716,n11718,n11627);
and (n11714,n11715,n10073);
and (n11716,n11717,n10091);
and (n11718,n11719,n10109);
and (n11720,n11721,n10340);
or (n11721,1'b0,n11722,n11723,n11711);
and (n11722,n11628,n10073);
and (n11723,n11724,n10091);
wire s0n11724,s1n11724,notn11724;
or (n11724,s0n11724,s1n11724);
not(notn11724,n10346);
and (s0n11724,notn11724,1'b0);
and (s1n11724,n10346,n11725);
wire s0n11725,s1n11725,notn11725;
or (n11725,s0n11725,s1n11725);
not(notn11725,n51);
and (s0n11725,notn11725,n11726);
and (s1n11725,n51,n11741);
wire s0n11726,s1n11726,notn11726;
or (n11726,s0n11726,s1n11726);
not(notn11726,n10335);
and (s0n11726,notn11726,n11727);
and (s1n11726,n10335,n11729);
wire s0n11727,s1n11727,notn11727;
or (n11727,s0n11727,s1n11727);
not(notn11727,n10020);
and (s0n11727,notn11727,1'b0);
and (s1n11727,n10020,n11728);
or (n11729,n11730,n11732,n11734,n11736,n11738,n11740);
and (n11730,n11731,n10309);
and (n11732,n11733,n10316);
and (n11734,n11735,n10319);
and (n11736,n11737,n10324);
and (n11738,n11739,n10331);
and (n11740,n11728,n10334);
wire s0n11741,s1n11741,notn11741;
or (n11741,s0n11741,s1n11741);
not(notn11741,n10345);
and (s0n11741,notn11741,1'b0);
and (s1n11741,n10345,n11742);
wire s0n11742,s1n11742,notn11742;
or (n11742,s0n11742,s1n11742);
not(notn11742,n10170);
and (s0n11742,notn11742,n11743);
and (s1n11742,n10170,n11744);
and (n11745,n11746,n10339);
or (n11746,1'b0,n11747,n11748);
and (n11747,n11596,n10352);
and (n11748,n11628,n10284);
and (n11749,n11750,n10337);
or (n11750,1'b0,n11751,n11752,n11753);
and (n11751,n11612,n10073);
and (n11752,n11724,n10109);
and (n11753,n11628,n10359);
and (n11754,n11755,n10366);
or (n11755,1'b0,n11756,n11758,n11759,n11627);
and (n11756,n11757,n10073);
and (n11758,n11719,n10091);
and (n11759,n11710,n10109);
and (n11760,n11761,n825);
or (n11761,1'b0,n11762,n11764);
and (n11762,n11763,n10109);
wire s0n11763,s1n11763,notn11763;
or (n11763,s0n11763,s1n11763);
not(notn11763,n10379);
and (s0n11763,notn11763,1'b0);
and (s1n11763,n10379,n11567);
and (n11764,n11765,n10005);
wire s0n11765,s1n11765,notn11765;
or (n11765,s0n11765,s1n11765);
not(notn11765,n10379);
and (s0n11765,notn11765,1'b0);
and (s1n11765,n10379,n11628);
and (n11766,n11644,n10392);
and (n11767,n11578,n10394);
wire s0n11768,s1n11768,notn11768;
or (n11768,s0n11768,s1n11768);
not(notn11768,n10395);
and (s0n11768,notn11768,n11769);
and (s1n11768,n10395,n11803);
wire s0n11769,s1n11769,notn11769;
or (n11769,s0n11769,s1n11769);
not(notn11769,n1039);
and (s0n11769,notn11769,n11770);
and (s1n11769,n1039,n11784);
wire s0n11770,s1n11770,notn11770;
or (n11770,s0n11770,s1n11770);
not(notn11770,n10261);
and (s0n11770,notn11770,1'b0);
and (s1n11770,n10261,n11771);
or (n11771,n11772,1'b0,n11777);
and (n11772,n11773,n10021);
wire s0n11773,s1n11773,notn11773;
or (n11773,s0n11773,s1n11773);
not(notn11773,n1057);
and (s0n11773,notn11773,1'b0);
and (s1n11773,n1057,n11774);
wire s0n11774,s1n11774,notn11774;
or (n11774,s0n11774,s1n11774);
not(notn11774,n10004);
and (s0n11774,notn11774,n11775);
and (s1n11774,n10004,n11776);
and (n11777,n11778,n10260);
or (n11778,n11779,n11782,1'b0);
and (n11779,n11780,n10242);
wire s0n11780,s1n11780,notn11780;
or (n11780,s0n11780,s1n11780);
not(notn11780,n10005);
and (s0n11780,notn11780,n11688);
and (s1n11780,n10005,n11781);
wire s0n11781,s1n11781,notn11781;
or (n11781,s0n11781,s1n11781);
not(notn11781,n10241);
and (s0n11781,notn11781,n11612);
and (s1n11781,n10241,1'b0);
and (n11782,n11783,n10257);
wire s0n11783,s1n11783,notn11783;
or (n11783,s0n11783,s1n11783);
not(notn11783,n10005);
and (s0n11783,notn11783,1'b0);
and (s1n11783,n10005,n11612);
or (n11784,n11785,n11788,1'b0);
and (n11785,n11786,n10020);
wire s0n11786,s1n11786,notn11786;
or (n11786,s0n11786,s1n11786);
not(notn11786,n1057);
and (s0n11786,notn11786,1'b0);
and (s1n11786,n1057,n11787);
wire s0n11787,s1n11787,notn11787;
or (n11787,s0n11787,s1n11787);
not(notn11787,n10417);
and (s0n11787,notn11787,n11775);
and (s1n11787,n10417,n11776);
and (n11788,n11789,n1042);
wire s0n11789,s1n11789,notn11789;
or (n11789,s0n11789,s1n11789);
not(notn11789,n650);
and (s0n11789,notn11789,1'b0);
and (s1n11789,n650,n11790);
or (n11790,1'b0,n11791,n11792,n11794);
and (n11791,n11689,n10352);
and (n11792,n11793,n10109);
wire s0n11793,s1n11793,notn11793;
or (n11793,s0n11793,s1n11793);
not(notn11793,n10243);
and (s0n11793,notn11793,n11619);
and (s1n11793,n10243,1'b0);
and (n11794,n11795,n10005);
wire s0n11795,s1n11795,notn11795;
or (n11795,s0n11795,s1n11795);
not(notn11795,n10148);
and (s0n11795,notn11795,n11796);
and (s1n11795,n10148,1'b0);
nand (n11796,n11797,n11799,n11801);
nand (n11797,n10136,n11798);
nand (n11799,n10173,n11800);
nand (n11801,n10160,n11802);
or (n11803,n11804,n11870,n11871,n11877,n11880,n11883,n11885,1'b0);
and (n11804,n11805,n10286);
or (n11805,1'b0,n11806,n11843);
and (n11806,n11807,n10109);
nand (n11807,n11808,n11825,n11837);
nor (n11808,n11809,n11819);
and (n11809,n11810,n10177);
nand (n11810,n11811,n11814);
or (n11811,n11812,n10135);
not (n11812,n11813);
nor (n11814,n11815,n11817);
and (n11815,n10160,n11816);
and (n11817,n10173,n11818);
nand (n11819,n11820,n11823);
or (n11820,n10223,n11821);
not (n11821,n11822);
or (n11823,n10211,n11824);
not (n11824,n11818);
and (n11825,n11826,n11833);
nor (n11826,n11827,n11830);
and (n11827,n11828,n10188);
and (n11828,n10136,n11829);
and (n11830,n11831,n10193);
and (n11831,n10136,n11832);
nor (n11833,n11834,n11836);
and (n11834,n10228,n11835);
and (n11836,n10231,n11816);
nand (n11837,n11838,n10205);
nand (n11838,n11839,n11841,n11842);
nand (n11839,n10136,n11840);
nand (n11841,n10173,n11835);
nand (n11842,n10160,n11822);
and (n11843,n11844,n10005);
nand (n11844,n11845,n11858);
and (n11845,n11846,n11854,n11855);
nand (n11846,n11847,n10177);
nand (n11847,n11848,n11850,n11852);
nand (n11848,n10136,n11849);
nand (n11850,n10173,n11851);
nand (n11852,n10160,n11853);
nand (n11854,n11796,n10205);
nor (n11855,n11856,n11857);
and (n11856,n10231,n11853);
and (n11857,n10222,n11802);
and (n11858,n11859,n11863,n11867);
nand (n11859,n11860,n10188);
nor (n11860,n10135,n11861);
not (n11861,n11862);
nand (n11863,n11864,n10193);
nor (n11864,n10135,n11865);
not (n11865,n11866);
nor (n11867,n11868,n11869);
and (n11868,n10228,n11800);
and (n11869,n10210,n11851);
and (n11870,n11783,n10296);
and (n11871,n11872,n10340);
or (n11872,1'b0,n11873,n11874,n11875,n11876);
and (n11873,n11596,n10073);
and (n11874,n11612,n10091);
and (n11875,n11628,n10109);
and (n11876,n11724,n10005);
and (n11877,n11878,n10339);
or (n11878,1'b0,n11579,n11879,n11876);
and (n11879,n11612,n10270);
and (n11880,n11881,n10337);
or (n11881,1'b0,n11579,n11595,n11611,n11882);
and (n11882,n11644,n10005);
and (n11883,n11884,n10366);
wire s0n11884,s1n11884,notn11884;
or (n11884,s0n11884,s1n11884);
not(notn11884,n10005);
and (s0n11884,notn11884,1'b0);
and (s1n11884,n10005,n11596);
and (n11885,n11886,n825);
or (n11886,1'b0,n11887,n11889);
and (n11887,n11888,n10109);
wire s0n11888,s1n11888,notn11888;
or (n11888,s0n11888,s1n11888);
not(notn11888,n10374);
and (s0n11888,notn11888,1'b0);
and (s1n11888,n10374,n11689);
and (n11889,n11890,n10005);
wire s0n11890,s1n11890,notn11890;
or (n11890,s0n11890,s1n11890);
not(notn11890,n10379);
and (s0n11890,notn11890,1'b0);
and (s1n11890,n10379,n11612);
and (n11891,n11768,n11892);
or (n11892,n11893,n12238,n12910);
and (n11893,n11894,n12107);
wire s0n11894,s1n11894,notn11894;
or (n11894,s0n11894,s1n11894);
not(notn11894,n10395);
and (s0n11894,notn11894,n11895);
and (s1n11894,n10395,n12043);
wire s0n11895,s1n11895,notn11895;
or (n11895,s0n11895,s1n11895);
not(notn11895,n1039);
and (s0n11895,notn11895,n11896);
and (s1n11895,n1039,n12031);
wire s0n11896,s1n11896,notn11896;
or (n11896,s0n11896,s1n11896);
not(notn11896,n10261);
and (s0n11896,notn11896,1'b0);
and (s1n11896,n10261,n11897);
or (n11897,n11898,n11911,n11977,n12020);
and (n11898,n11899,n10021);
wire s0n11899,s1n11899,notn11899;
or (n11899,s0n11899,s1n11899);
not(notn11899,n1057);
and (s0n11899,notn11899,1'b0);
and (s1n11899,n1057,n11900);
wire s0n11900,s1n11900,notn11900;
or (n11900,s0n11900,s1n11900);
not(notn11900,n10004);
and (s0n11900,notn11900,n11901);
and (s1n11900,n10004,n11902);
wire s0n11902,s1n11902,notn11902;
or (n11902,s0n11902,s1n11902);
not(notn11902,n10017);
and (s0n11902,notn11902,n11903);
and (s1n11902,n10017,n11905);
wire s0n11903,s1n11903,notn11903;
or (n11903,s0n11903,s1n11903);
not(notn11903,n10000);
and (s0n11903,notn11903,1'b0);
and (s1n11903,n10000,n11904);
or (n11905,1'b0,n11906,n11908,n11910);
and (n11906,n11907,n10009);
and (n11908,n11909,n10012);
and (n11910,n11904,n10014);
and (n11911,n11912,n10126);
or (n11912,1'b0,n11913,n11929,n11945,n11961);
and (n11913,n11914,n10073);
wire s0n11914,s1n11914,notn11914;
or (n11914,s0n11914,s1n11914);
not(notn11914,n65);
and (s0n11914,notn11914,1'b0);
and (s1n11914,n65,n11915);
wire s0n11915,s1n11915,notn11915;
or (n11915,s0n11915,s1n11915);
not(notn11915,n10068);
and (s0n11915,notn11915,n11916);
and (s1n11915,n10068,n11922);
wire s0n11916,s1n11916,notn11916;
or (n11916,s0n11916,s1n11916);
not(notn11916,n10047);
and (s0n11916,notn11916,1'b0);
and (s1n11916,n10047,n11917);
or (n11917,1'b0,n11918,n11920);
and (n11918,n11919,n10031);
and (n11920,n11921,n10040);
or (n11922,1'b0,n11923,n11925,n11927,n11928);
and (n11923,n11924,n10055);
and (n11925,n11926,n10060);
and (n11927,n11919,n10064);
and (n11928,n11921,n10014);
and (n11929,n11930,n10091);
wire s0n11930,s1n11930,notn11930;
or (n11930,s0n11930,s1n11930);
not(notn11930,n65);
and (s0n11930,notn11930,1'b0);
and (s1n11930,n65,n11931);
wire s0n11931,s1n11931,notn11931;
or (n11931,s0n11931,s1n11931);
not(notn11931,n10068);
and (s0n11931,notn11931,n11932);
and (s1n11931,n10068,n11938);
wire s0n11932,s1n11932,notn11932;
or (n11932,s0n11932,s1n11932);
not(notn11932,n10047);
and (s0n11932,notn11932,1'b0);
and (s1n11932,n10047,n11933);
or (n11933,1'b0,n11934,n11936);
and (n11934,n11935,n10031);
and (n11936,n11937,n10040);
or (n11938,1'b0,n11939,n11941,n11943,n11944);
and (n11939,n11940,n10055);
and (n11941,n11942,n10060);
and (n11943,n11935,n10064);
and (n11944,n11937,n10014);
and (n11945,n11946,n10109);
wire s0n11946,s1n11946,notn11946;
or (n11946,s0n11946,s1n11946);
not(notn11946,n65);
and (s0n11946,notn11946,1'b0);
and (s1n11946,n65,n11947);
wire s0n11947,s1n11947,notn11947;
or (n11947,s0n11947,s1n11947);
not(notn11947,n10068);
and (s0n11947,notn11947,n11948);
and (s1n11947,n10068,n11954);
wire s0n11948,s1n11948,notn11948;
or (n11948,s0n11948,s1n11948);
not(notn11948,n10047);
and (s0n11948,notn11948,1'b0);
and (s1n11948,n10047,n11949);
or (n11949,1'b0,n11950,n11952);
and (n11950,n11951,n10031);
and (n11952,n11953,n10040);
or (n11954,1'b0,n11955,n11957,n11959,n11960);
and (n11955,n11956,n10055);
and (n11957,n11958,n10060);
and (n11959,n11951,n10064);
and (n11960,n11953,n10014);
and (n11961,n11962,n10005);
wire s0n11962,s1n11962,notn11962;
or (n11962,s0n11962,s1n11962);
not(notn11962,n65);
and (s0n11962,notn11962,1'b0);
and (s1n11962,n65,n11963);
wire s0n11963,s1n11963,notn11963;
or (n11963,s0n11963,s1n11963);
not(notn11963,n10068);
and (s0n11963,notn11963,n11964);
and (s1n11963,n10068,n11970);
wire s0n11964,s1n11964,notn11964;
or (n11964,s0n11964,s1n11964);
not(notn11964,n10047);
and (s0n11964,notn11964,1'b0);
and (s1n11964,n10047,n11965);
or (n11965,1'b0,n11966,n11968);
and (n11966,n11967,n10031);
and (n11968,n11969,n10040);
or (n11970,1'b0,n11971,n11973,n11975,n11976);
and (n11971,n11972,n10055);
and (n11973,n11974,n10060);
and (n11975,n11967,n10064);
and (n11976,n11969,n10014);
and (n11977,n11978,n10215);
nand (n11978,n11979,n12006);
nor (n11979,n11980,n11992);
and (n11980,n11981,n10205);
nand (n11981,n11982,n11985);
or (n11982,n11983,n10135);
not (n11983,n11984);
nor (n11985,n11986,n11989);
nor (n11986,n11987,n10174);
not (n11987,n11988);
nor (n11989,n11990,n10161);
not (n11990,n11991);
nand (n11992,n11993,n11997,n12001);
nand (n11993,n11994,n10188);
nor (n11994,n10135,n11995);
not (n11995,n11996);
nand (n11997,n11998,n10193);
nor (n11998,n10135,n11999);
not (n11999,n12000);
nor (n12001,n12002,n12004);
and (n12002,n10210,n12003);
and (n12004,n10231,n12005);
nor (n12006,n12007,n12017);
and (n12007,n12008,n10177);
nand (n12008,n12009,n12012);
or (n12009,n12010,n10135);
not (n12010,n12011);
nor (n12012,n12013,n12015);
nor (n12013,n12014,n10174);
not (n12014,n12003);
nor (n12015,n12016,n10161);
not (n12016,n12005);
nand (n12017,n12018,n12019);
or (n12018,n10223,n11990);
or (n12019,n10229,n11987);
and (n12020,n12021,n10260);
or (n12021,n12022,n12026,n12029,1'b0);
and (n12022,n12023,n10242);
wire s0n12023,s1n12023,notn12023;
or (n12023,s0n12023,s1n12023);
not(notn12023,n10005);
and (s0n12023,notn12023,n12024);
and (s1n12023,n10005,n12025);
wire s0n12024,s1n12024,notn12024;
or (n12024,s0n12024,s1n12024);
not(notn12024,n10109);
and (s0n12024,notn12024,1'b0);
and (s1n12024,n10109,n11901);
wire s0n12025,s1n12025,notn12025;
or (n12025,s0n12025,s1n12025);
not(notn12025,n10241);
and (s0n12025,notn12025,n11962);
and (s1n12025,n10241,1'b0);
and (n12026,n12027,n10254);
wire s0n12027,s1n12027,notn12027;
or (n12027,s0n12027,s1n12027);
not(notn12027,n10109);
and (s0n12027,notn12027,1'b0);
and (s1n12027,n10109,n12028);
and (n12029,n12030,n10257);
wire s0n12030,s1n12030,notn12030;
or (n12030,s0n12030,s1n12030);
not(notn12030,n10005);
and (s0n12030,notn12030,n12024);
and (s1n12030,n10005,n11962);
or (n12031,n12032,n12033,n12041,n12042);
and (n12032,n11899,n10020);
and (n12033,n12034,n1042);
wire s0n12034,s1n12034,notn12034;
or (n12034,s0n12034,s1n12034);
not(notn12034,n650);
and (s0n12034,notn12034,1'b0);
and (s1n12034,n650,n12035);
or (n12035,1'b0,n12036,n12038,n12039);
and (n12036,n12037,n10073);
wire s0n12037,s1n12037,notn12037;
or (n12037,s0n12037,s1n12037);
not(notn12037,n10259);
and (s0n12037,notn12037,n11901);
and (s1n12037,n10259,1'b0);
and (n12038,n11901,n10270);
and (n12039,n12040,n10005);
wire s0n12040,s1n12040,notn12040;
or (n12040,s0n12040,s1n12040);
not(notn12040,n10148);
and (s0n12040,notn12040,n11981);
and (s1n12040,n10148,1'b0);
and (n12041,n11978,n10181);
and (n12042,n11912,n10072);
or (n12043,1'b0,n12044,n12051,n12059,n12084,n12088,n12093,n12099,n12105,n12106);
and (n12044,n12045,n10286);
or (n12045,1'b0,n12046,n12048,n12050);
and (n12046,n12047,n10073);
and (n12048,n12049,n10091);
and (n12050,n11978,n10284);
and (n12051,n12052,n10296);
or (n12052,1'b0,n12053,n12055,n12057,n11961);
and (n12053,n12054,n10073);
and (n12055,n12056,n10091);
and (n12057,n12058,n10109);
and (n12059,n12060,n10340);
or (n12060,1'b0,n12061,n12062,n12050);
and (n12061,n11962,n10073);
and (n12062,n12063,n10091);
wire s0n12063,s1n12063,notn12063;
or (n12063,s0n12063,s1n12063);
not(notn12063,n10346);
and (s0n12063,notn12063,1'b0);
and (s1n12063,n10346,n12064);
wire s0n12064,s1n12064,notn12064;
or (n12064,s0n12064,s1n12064);
not(notn12064,n51);
and (s0n12064,notn12064,n12065);
and (s1n12064,n51,n12080);
wire s0n12065,s1n12065,notn12065;
or (n12065,s0n12065,s1n12065);
not(notn12065,n10335);
and (s0n12065,notn12065,n12066);
and (s1n12065,n10335,n12068);
wire s0n12066,s1n12066,notn12066;
or (n12066,s0n12066,s1n12066);
not(notn12066,n10020);
and (s0n12066,notn12066,1'b0);
and (s1n12066,n10020,n12067);
or (n12068,n12069,n12071,n12073,n12075,n12077,n12079);
and (n12069,n12070,n10309);
and (n12071,n12072,n10316);
and (n12073,n12074,n10319);
and (n12075,n12076,n10324);
and (n12077,n12078,n10331);
and (n12079,n12067,n10334);
wire s0n12080,s1n12080,notn12080;
or (n12080,s0n12080,s1n12080);
not(notn12080,n10345);
and (s0n12080,notn12080,1'b0);
and (s1n12080,n10345,n12081);
wire s0n12081,s1n12081,notn12081;
or (n12081,s0n12081,s1n12081);
not(notn12081,n10170);
and (s0n12081,notn12081,n12082);
and (s1n12081,n10170,n12083);
and (n12084,n12085,n10339);
or (n12085,1'b0,n12086,n12087);
and (n12086,n11930,n10352);
and (n12087,n11962,n10284);
and (n12088,n12089,n10337);
or (n12089,1'b0,n12090,n12091,n12092);
and (n12090,n11946,n10073);
and (n12091,n12063,n10109);
and (n12092,n11962,n10359);
and (n12093,n12094,n10366);
or (n12094,1'b0,n12095,n12097,n12098,n11961);
and (n12095,n12096,n10073);
and (n12097,n12058,n10091);
and (n12098,n12049,n10109);
and (n12099,n12100,n825);
or (n12100,1'b0,n12101,n12103);
and (n12101,n12102,n10109);
wire s0n12102,s1n12102,notn12102;
or (n12102,s0n12102,s1n12102);
not(notn12102,n10379);
and (s0n12102,notn12102,1'b0);
and (s1n12102,n10379,n11901);
and (n12103,n12104,n10005);
wire s0n12104,s1n12104,notn12104;
or (n12104,s0n12104,s1n12104);
not(notn12104,n10379);
and (s0n12104,notn12104,1'b0);
and (s1n12104,n10379,n11962);
and (n12105,n11978,n10392);
and (n12106,n11912,n10394);
wire s0n12107,s1n12107,notn12107;
or (n12107,s0n12107,s1n12107);
not(notn12107,n10395);
and (s0n12107,notn12107,n12108);
and (s1n12107,n10395,n12142);
wire s0n12108,s1n12108,notn12108;
or (n12108,s0n12108,s1n12108);
not(notn12108,n1039);
and (s0n12108,notn12108,n12109);
and (s1n12108,n1039,n12123);
wire s0n12109,s1n12109,notn12109;
or (n12109,s0n12109,s1n12109);
not(notn12109,n10261);
and (s0n12109,notn12109,1'b0);
and (s1n12109,n10261,n12110);
or (n12110,n12111,1'b0,n12116);
and (n12111,n12112,n10021);
wire s0n12112,s1n12112,notn12112;
or (n12112,s0n12112,s1n12112);
not(notn12112,n1057);
and (s0n12112,notn12112,1'b0);
and (s1n12112,n1057,n12113);
wire s0n12113,s1n12113,notn12113;
or (n12113,s0n12113,s1n12113);
not(notn12113,n10004);
and (s0n12113,notn12113,n12114);
and (s1n12113,n10004,n12115);
and (n12116,n12117,n10260);
or (n12117,n12118,n12121,1'b0);
and (n12118,n12119,n10242);
wire s0n12119,s1n12119,notn12119;
or (n12119,s0n12119,s1n12119);
not(notn12119,n10005);
and (s0n12119,notn12119,n12027);
and (s1n12119,n10005,n12120);
wire s0n12120,s1n12120,notn12120;
or (n12120,s0n12120,s1n12120);
not(notn12120,n10241);
and (s0n12120,notn12120,n11946);
and (s1n12120,n10241,1'b0);
and (n12121,n12122,n10257);
wire s0n12122,s1n12122,notn12122;
or (n12122,s0n12122,s1n12122);
not(notn12122,n10005);
and (s0n12122,notn12122,1'b0);
and (s1n12122,n10005,n11946);
or (n12123,n12124,n12127,1'b0);
and (n12124,n12125,n10020);
wire s0n12125,s1n12125,notn12125;
or (n12125,s0n12125,s1n12125);
not(notn12125,n1057);
and (s0n12125,notn12125,1'b0);
and (s1n12125,n1057,n12126);
wire s0n12126,s1n12126,notn12126;
or (n12126,s0n12126,s1n12126);
not(notn12126,n10417);
and (s0n12126,notn12126,n12114);
and (s1n12126,n10417,n12115);
and (n12127,n12128,n1042);
wire s0n12128,s1n12128,notn12128;
or (n12128,s0n12128,s1n12128);
not(notn12128,n650);
and (s0n12128,notn12128,1'b0);
and (s1n12128,n650,n12129);
or (n12129,1'b0,n12130,n12131,n12133);
and (n12130,n12028,n10352);
and (n12131,n12132,n10109);
wire s0n12132,s1n12132,notn12132;
or (n12132,s0n12132,s1n12132);
not(notn12132,n10243);
and (s0n12132,notn12132,n11953);
and (s1n12132,n10243,1'b0);
and (n12133,n12134,n10005);
wire s0n12134,s1n12134,notn12134;
or (n12134,s0n12134,s1n12134);
not(notn12134,n10148);
and (s0n12134,notn12134,n12135);
and (s1n12134,n10148,1'b0);
nand (n12135,n12136,n12138,n12140);
nand (n12136,n10136,n12137);
nand (n12138,n10173,n12139);
nand (n12140,n10160,n12141);
or (n12142,n12143,n12211,n12212,n12218,n12221,n12230,n12232,1'b0);
and (n12143,n12144,n10286);
or (n12144,1'b0,n12145,n12182);
and (n12145,n12146,n10109);
nand (n12146,n12147,n12166);
nor (n12147,n12148,n12158);
and (n12148,n12149,n10177);
nand (n12149,n12150,n12153);
or (n12150,n12151,n10135);
not (n12151,n12152);
nor (n12153,n12154,n12156);
and (n12154,n10160,n12155);
and (n12156,n10173,n12157);
nand (n12158,n12159,n12163);
or (n12159,n11331,n12160);
not (n12160,n12161);
and (n12161,n10136,n12162);
nand (n12163,n12164,n10188);
and (n12164,n10136,n12165);
nor (n12166,n12167,n12175);
and (n12167,n12168,n10205);
nand (n12168,n12169,n12171,n12173);
nand (n12169,n10136,n12170);
nand (n12171,n10173,n12172);
nand (n12173,n10160,n12174);
nand (n12175,n12176,n12179);
nor (n12176,n12177,n12178);
and (n12177,n10228,n12172);
and (n12178,n10231,n12155);
nor (n12179,n12180,n12181);
and (n12180,n10210,n12157);
and (n12181,n10222,n12174);
and (n12182,n12183,n10005);
nand (n12183,n12184,n12198);
not (n12184,n12185);
nand (n12185,n12186,n12194,n12195);
nand (n12186,n12187,n10177);
nand (n12187,n12188,n12190,n12192);
nand (n12188,n10136,n12189);
nand (n12190,n10173,n12191);
nand (n12192,n10160,n12193);
nand (n12194,n12135,n10205);
nor (n12195,n12196,n12197);
and (n12196,n10231,n12193);
and (n12197,n10222,n12141);
not (n12198,n12199);
nand (n12199,n12200,n12204,n12208);
nand (n12200,n12201,n10188);
nor (n12201,n10135,n12202);
not (n12202,n12203);
nand (n12204,n12205,n10193);
nor (n12205,n10135,n12206);
not (n12206,n12207);
nor (n12208,n12209,n12210);
and (n12209,n10228,n12139);
and (n12210,n10210,n12191);
and (n12211,n12122,n10296);
and (n12212,n12213,n10340);
or (n12213,1'b0,n12214,n12215,n12216,n12217);
and (n12214,n11930,n10073);
and (n12215,n11946,n10091);
and (n12216,n11962,n10109);
and (n12217,n12063,n10005);
and (n12218,n12219,n10339);
or (n12219,1'b0,n11913,n12220,n12217);
and (n12220,n11946,n10270);
not (n12221,n12222);
nand (n12222,n12223,n10337);
nand (n12223,n12224,n12226);
or (n12224,n10522,n12225);
not (n12225,n11978);
and (n12226,n12227,n12228,n12229);
not (n12227,n11913);
not (n12228,n11945);
not (n12229,n11929);
and (n12230,n12231,n10366);
wire s0n12231,s1n12231,notn12231;
or (n12231,s0n12231,s1n12231);
not(notn12231,n10005);
and (s0n12231,notn12231,1'b0);
and (s1n12231,n10005,n11930);
and (n12232,n12233,n825);
or (n12233,1'b0,n12234,n12236);
and (n12234,n12235,n10109);
wire s0n12235,s1n12235,notn12235;
or (n12235,s0n12235,s1n12235);
not(notn12235,n10374);
and (s0n12235,notn12235,1'b0);
and (s1n12235,n10374,n12028);
and (n12236,n12237,n10005);
wire s0n12237,s1n12237,notn12237;
or (n12237,s0n12237,s1n12237);
not(notn12237,n10379);
and (s0n12237,notn12237,1'b0);
and (s1n12237,n10379,n11946);
and (n12238,n12107,n12239);
or (n12239,n12240,n12573,n12909);
and (n12240,n12241,n12449);
wire s0n12241,s1n12241,notn12241;
or (n12241,s0n12241,s1n12241);
not(notn12241,n10395);
and (s0n12241,notn12241,n12242);
and (s1n12241,n10395,n12385);
wire s0n12242,s1n12242,notn12242;
or (n12242,s0n12242,s1n12242);
not(notn12242,n1039);
and (s0n12242,notn12242,n12243);
and (s1n12242,n1039,n12373);
wire s0n12243,s1n12243,notn12243;
or (n12243,s0n12243,s1n12243);
not(notn12243,n10261);
and (s0n12243,notn12243,1'b0);
and (s1n12243,n10261,n12244);
or (n12244,n12245,n12258,n12324,n12362);
and (n12245,n12246,n10021);
wire s0n12246,s1n12246,notn12246;
or (n12246,s0n12246,s1n12246);
not(notn12246,n1057);
and (s0n12246,notn12246,1'b0);
and (s1n12246,n1057,n12247);
wire s0n12247,s1n12247,notn12247;
or (n12247,s0n12247,s1n12247);
not(notn12247,n10004);
and (s0n12247,notn12247,n12248);
and (s1n12247,n10004,n12249);
wire s0n12249,s1n12249,notn12249;
or (n12249,s0n12249,s1n12249);
not(notn12249,n10017);
and (s0n12249,notn12249,n12250);
and (s1n12249,n10017,n12252);
wire s0n12250,s1n12250,notn12250;
or (n12250,s0n12250,s1n12250);
not(notn12250,n10000);
and (s0n12250,notn12250,1'b0);
and (s1n12250,n10000,n12251);
or (n12252,1'b0,n12253,n12255,n12257);
and (n12253,n12254,n10009);
and (n12255,n12256,n10012);
and (n12257,n12251,n10014);
and (n12258,n12259,n10126);
or (n12259,1'b0,n12260,n12276,n12292,n12308);
and (n12260,n12261,n10073);
wire s0n12261,s1n12261,notn12261;
or (n12261,s0n12261,s1n12261);
not(notn12261,n65);
and (s0n12261,notn12261,1'b0);
and (s1n12261,n65,n12262);
wire s0n12262,s1n12262,notn12262;
or (n12262,s0n12262,s1n12262);
not(notn12262,n10068);
and (s0n12262,notn12262,n12263);
and (s1n12262,n10068,n12269);
wire s0n12263,s1n12263,notn12263;
or (n12263,s0n12263,s1n12263);
not(notn12263,n10047);
and (s0n12263,notn12263,1'b0);
and (s1n12263,n10047,n12264);
or (n12264,1'b0,n12265,n12267);
and (n12265,n12266,n10031);
and (n12267,n12268,n10040);
or (n12269,1'b0,n12270,n12272,n12274,n12275);
and (n12270,n12271,n10055);
and (n12272,n12273,n10060);
and (n12274,n12266,n10064);
and (n12275,n12268,n10014);
and (n12276,n12277,n10091);
wire s0n12277,s1n12277,notn12277;
or (n12277,s0n12277,s1n12277);
not(notn12277,n65);
and (s0n12277,notn12277,1'b0);
and (s1n12277,n65,n12278);
wire s0n12278,s1n12278,notn12278;
or (n12278,s0n12278,s1n12278);
not(notn12278,n10068);
and (s0n12278,notn12278,n12279);
and (s1n12278,n10068,n12285);
wire s0n12279,s1n12279,notn12279;
or (n12279,s0n12279,s1n12279);
not(notn12279,n10047);
and (s0n12279,notn12279,1'b0);
and (s1n12279,n10047,n12280);
or (n12280,1'b0,n12281,n12283);
and (n12281,n12282,n10031);
and (n12283,n12284,n10040);
or (n12285,1'b0,n12286,n12288,n12290,n12291);
and (n12286,n12287,n10055);
and (n12288,n12289,n10060);
and (n12290,n12282,n10064);
and (n12291,n12284,n10014);
and (n12292,n12293,n10109);
wire s0n12293,s1n12293,notn12293;
or (n12293,s0n12293,s1n12293);
not(notn12293,n65);
and (s0n12293,notn12293,1'b0);
and (s1n12293,n65,n12294);
wire s0n12294,s1n12294,notn12294;
or (n12294,s0n12294,s1n12294);
not(notn12294,n10068);
and (s0n12294,notn12294,n12295);
and (s1n12294,n10068,n12301);
wire s0n12295,s1n12295,notn12295;
or (n12295,s0n12295,s1n12295);
not(notn12295,n10047);
and (s0n12295,notn12295,1'b0);
and (s1n12295,n10047,n12296);
or (n12296,1'b0,n12297,n12299);
and (n12297,n12298,n10031);
and (n12299,n12300,n10040);
or (n12301,1'b0,n12302,n12304,n12306,n12307);
and (n12302,n12303,n10055);
and (n12304,n12305,n10060);
and (n12306,n12298,n10064);
and (n12307,n12300,n10014);
and (n12308,n12309,n10005);
wire s0n12309,s1n12309,notn12309;
or (n12309,s0n12309,s1n12309);
not(notn12309,n65);
and (s0n12309,notn12309,1'b0);
and (s1n12309,n65,n12310);
wire s0n12310,s1n12310,notn12310;
or (n12310,s0n12310,s1n12310);
not(notn12310,n10068);
and (s0n12310,notn12310,n12311);
and (s1n12310,n10068,n12317);
wire s0n12311,s1n12311,notn12311;
or (n12311,s0n12311,s1n12311);
not(notn12311,n10047);
and (s0n12311,notn12311,1'b0);
and (s1n12311,n10047,n12312);
or (n12312,1'b0,n12313,n12315);
and (n12313,n12314,n10031);
and (n12315,n12316,n10040);
or (n12317,1'b0,n12318,n12320,n12322,n12323);
and (n12318,n12319,n10055);
and (n12320,n12321,n10060);
and (n12322,n12314,n10064);
and (n12323,n12316,n10014);
and (n12324,n12325,n10215);
nand (n12325,n12326,n12350);
nor (n12326,n12327,n12337);
and (n12327,n12328,n10205);
nand (n12328,n12329,n12332);
or (n12329,n12330,n10135);
not (n12330,n12331);
nor (n12332,n12333,n12335);
and (n12333,n10160,n12334);
and (n12335,n10173,n12336);
nand (n12337,n12338,n12342,n12346);
nand (n12338,n12339,n10188);
nor (n12339,n10135,n12340);
not (n12340,n12341);
nand (n12342,n12343,n10193);
nor (n12343,n10135,n12344);
not (n12344,n12345);
nor (n12346,n12347,n12348);
and (n12347,n10228,n12336);
and (n12348,n10231,n12349);
nor (n12350,n12351,n12358);
and (n12351,n12352,n10177);
nand (n12352,n12353,n12355,n12357);
nand (n12353,n10136,n12354);
nand (n12355,n10173,n12356);
nand (n12357,n10160,n12349);
nand (n12358,n12359,n12361);
or (n12359,n12360,n10223);
not (n12360,n12334);
nand (n12361,n10210,n12356);
and (n12362,n12363,n10260);
or (n12363,n12364,n12368,n12371,1'b0);
and (n12364,n12365,n10242);
wire s0n12365,s1n12365,notn12365;
or (n12365,s0n12365,s1n12365);
not(notn12365,n10005);
and (s0n12365,notn12365,n12366);
and (s1n12365,n10005,n12367);
wire s0n12366,s1n12366,notn12366;
or (n12366,s0n12366,s1n12366);
not(notn12366,n10109);
and (s0n12366,notn12366,1'b0);
and (s1n12366,n10109,n12248);
wire s0n12367,s1n12367,notn12367;
or (n12367,s0n12367,s1n12367);
not(notn12367,n10241);
and (s0n12367,notn12367,n12309);
and (s1n12367,n10241,1'b0);
and (n12368,n12369,n10254);
wire s0n12369,s1n12369,notn12369;
or (n12369,s0n12369,s1n12369);
not(notn12369,n10109);
and (s0n12369,notn12369,1'b0);
and (s1n12369,n10109,n12370);
and (n12371,n12372,n10257);
wire s0n12372,s1n12372,notn12372;
or (n12372,s0n12372,s1n12372);
not(notn12372,n10005);
and (s0n12372,notn12372,n12366);
and (s1n12372,n10005,n12309);
or (n12373,n12374,n12375,n12383,n12384);
and (n12374,n12246,n10020);
and (n12375,n12376,n1042);
wire s0n12376,s1n12376,notn12376;
or (n12376,s0n12376,s1n12376);
not(notn12376,n650);
and (s0n12376,notn12376,1'b0);
and (s1n12376,n650,n12377);
or (n12377,1'b0,n12378,n12380,n12381);
and (n12378,n12379,n10073);
wire s0n12379,s1n12379,notn12379;
or (n12379,s0n12379,s1n12379);
not(notn12379,n10259);
and (s0n12379,notn12379,n12248);
and (s1n12379,n10259,1'b0);
and (n12380,n12248,n10270);
and (n12381,n12382,n10005);
wire s0n12382,s1n12382,notn12382;
or (n12382,s0n12382,s1n12382);
not(notn12382,n10148);
and (s0n12382,notn12382,n12328);
and (s1n12382,n10148,1'b0);
and (n12383,n12325,n10181);
and (n12384,n12259,n10072);
or (n12385,1'b0,n12386,n12393,n12401,n12426,n12430,n12435,n12441,n12447,n12448);
and (n12386,n12387,n10286);
or (n12387,1'b0,n12388,n12390,n12392);
and (n12388,n12389,n10073);
and (n12390,n12391,n10091);
and (n12392,n12325,n10284);
and (n12393,n12394,n10296);
or (n12394,1'b0,n12395,n12397,n12399,n12308);
and (n12395,n12396,n10073);
and (n12397,n12398,n10091);
and (n12399,n12400,n10109);
and (n12401,n12402,n10340);
or (n12402,1'b0,n12403,n12404,n12392);
and (n12403,n12309,n10073);
and (n12404,n12405,n10091);
wire s0n12405,s1n12405,notn12405;
or (n12405,s0n12405,s1n12405);
not(notn12405,n10346);
and (s0n12405,notn12405,1'b0);
and (s1n12405,n10346,n12406);
wire s0n12406,s1n12406,notn12406;
or (n12406,s0n12406,s1n12406);
not(notn12406,n51);
and (s0n12406,notn12406,n12407);
and (s1n12406,n51,n12422);
wire s0n12407,s1n12407,notn12407;
or (n12407,s0n12407,s1n12407);
not(notn12407,n10335);
and (s0n12407,notn12407,n12408);
and (s1n12407,n10335,n12410);
wire s0n12408,s1n12408,notn12408;
or (n12408,s0n12408,s1n12408);
not(notn12408,n10020);
and (s0n12408,notn12408,1'b0);
and (s1n12408,n10020,n12409);
or (n12410,n12411,n12413,n12415,n12417,n12419,n12421);
and (n12411,n12412,n10309);
and (n12413,n12414,n10316);
and (n12415,n12416,n10319);
and (n12417,n12418,n10324);
and (n12419,n12420,n10331);
and (n12421,n12409,n10334);
wire s0n12422,s1n12422,notn12422;
or (n12422,s0n12422,s1n12422);
not(notn12422,n10345);
and (s0n12422,notn12422,1'b0);
and (s1n12422,n10345,n12423);
wire s0n12423,s1n12423,notn12423;
or (n12423,s0n12423,s1n12423);
not(notn12423,n10170);
and (s0n12423,notn12423,n12424);
and (s1n12423,n10170,n12425);
and (n12426,n12427,n10339);
or (n12427,1'b0,n12428,n12429);
and (n12428,n12277,n10352);
and (n12429,n12309,n10284);
and (n12430,n12431,n10337);
or (n12431,1'b0,n12432,n12433,n12434);
and (n12432,n12293,n10073);
and (n12433,n12405,n10109);
and (n12434,n12309,n10359);
and (n12435,n12436,n10366);
or (n12436,1'b0,n12437,n12439,n12440,n12308);
and (n12437,n12438,n10073);
and (n12439,n12400,n10091);
and (n12440,n12391,n10109);
and (n12441,n12442,n825);
or (n12442,1'b0,n12443,n12445);
and (n12443,n12444,n10109);
wire s0n12444,s1n12444,notn12444;
or (n12444,s0n12444,s1n12444);
not(notn12444,n10379);
and (s0n12444,notn12444,1'b0);
and (s1n12444,n10379,n12248);
and (n12445,n12446,n10005);
wire s0n12446,s1n12446,notn12446;
or (n12446,s0n12446,s1n12446);
not(notn12446,n10379);
and (s0n12446,notn12446,1'b0);
and (s1n12446,n10379,n12309);
and (n12447,n12325,n10392);
and (n12448,n12259,n10394);
wire s0n12449,s1n12449,notn12449;
or (n12449,s0n12449,s1n12449);
not(notn12449,n10395);
and (s0n12449,notn12449,n12450);
and (s1n12449,n10395,n12484);
wire s0n12450,s1n12450,notn12450;
or (n12450,s0n12450,s1n12450);
not(notn12450,n1039);
and (s0n12450,notn12450,n12451);
and (s1n12450,n1039,n12465);
wire s0n12451,s1n12451,notn12451;
or (n12451,s0n12451,s1n12451);
not(notn12451,n10261);
and (s0n12451,notn12451,1'b0);
and (s1n12451,n10261,n12452);
or (n12452,n12453,1'b0,n12458);
and (n12453,n12454,n10021);
wire s0n12454,s1n12454,notn12454;
or (n12454,s0n12454,s1n12454);
not(notn12454,n1057);
and (s0n12454,notn12454,1'b0);
and (s1n12454,n1057,n12455);
wire s0n12455,s1n12455,notn12455;
or (n12455,s0n12455,s1n12455);
not(notn12455,n10004);
and (s0n12455,notn12455,n12456);
and (s1n12455,n10004,n12457);
and (n12458,n12459,n10260);
or (n12459,n12460,n12463,1'b0);
and (n12460,n12461,n10242);
wire s0n12461,s1n12461,notn12461;
or (n12461,s0n12461,s1n12461);
not(notn12461,n10005);
and (s0n12461,notn12461,n12369);
and (s1n12461,n10005,n12462);
wire s0n12462,s1n12462,notn12462;
or (n12462,s0n12462,s1n12462);
not(notn12462,n10241);
and (s0n12462,notn12462,n12293);
and (s1n12462,n10241,1'b0);
and (n12463,n12464,n10257);
wire s0n12464,s1n12464,notn12464;
or (n12464,s0n12464,s1n12464);
not(notn12464,n10005);
and (s0n12464,notn12464,1'b0);
and (s1n12464,n10005,n12293);
or (n12465,n12466,n12469,1'b0);
and (n12466,n12467,n10020);
wire s0n12467,s1n12467,notn12467;
or (n12467,s0n12467,s1n12467);
not(notn12467,n1057);
and (s0n12467,notn12467,1'b0);
and (s1n12467,n1057,n12468);
wire s0n12468,s1n12468,notn12468;
or (n12468,s0n12468,s1n12468);
not(notn12468,n10417);
and (s0n12468,notn12468,n12456);
and (s1n12468,n10417,n12457);
and (n12469,n12470,n1042);
wire s0n12470,s1n12470,notn12470;
or (n12470,s0n12470,s1n12470);
not(notn12470,n650);
and (s0n12470,notn12470,1'b0);
and (s1n12470,n650,n12471);
or (n12471,1'b0,n12472,n12473,n12475);
and (n12472,n12370,n10352);
and (n12473,n12474,n10109);
wire s0n12474,s1n12474,notn12474;
or (n12474,s0n12474,s1n12474);
not(notn12474,n10243);
and (s0n12474,notn12474,n12300);
and (s1n12474,n10243,1'b0);
and (n12475,n12476,n10005);
wire s0n12476,s1n12476,notn12476;
or (n12476,s0n12476,s1n12476);
not(notn12476,n10148);
and (s0n12476,notn12476,n12477);
and (s1n12476,n10148,1'b0);
nand (n12477,n12478,n12480,n12482);
nand (n12478,n10136,n12479);
nand (n12480,n10173,n12481);
nand (n12482,n10160,n12483);
or (n12484,n12485,n12550,n12551,n12557,n12560,n12565,n12567,1'b0);
and (n12485,n12486,n10286);
or (n12486,1'b0,n12487,n12523);
and (n12487,n12488,n10109);
nand (n12488,n12489,n12511);
nor (n12489,n12490,n12498);
and (n12490,n12491,n10205);
nand (n12491,n12492,n12494,n12496);
nand (n12492,n10136,n12493);
nand (n12494,n10173,n12495);
nand (n12496,n10160,n12497);
nand (n12498,n12499,n12503,n12507);
nand (n12499,n12500,n10188);
nor (n12500,n10135,n12501);
not (n12501,n12502);
nand (n12503,n12504,n10193);
nor (n12504,n10135,n12505);
not (n12505,n12506);
nor (n12507,n12508,n12510);
and (n12508,n10231,n12509);
and (n12510,n10222,n12497);
nor (n12511,n12512,n12519);
and (n12512,n12513,n10177);
nand (n12513,n12514,n12516,n12518);
nand (n12514,n10136,n12515);
nand (n12516,n10173,n12517);
nand (n12518,n10160,n12509);
nand (n12519,n12520,n12522);
or (n12520,n12521,n10229);
not (n12521,n12495);
nand (n12522,n10210,n12517);
and (n12523,n12524,n10005);
nand (n12524,n12525,n12535,n12547);
and (n12525,n12526,n12534);
nand (n12526,n12527,n10177);
nand (n12527,n12528,n12530,n12532);
nand (n12528,n10136,n12529);
nand (n12530,n10173,n12531);
nand (n12532,n10160,n12533);
nand (n12534,n12477,n10205);
and (n12535,n12536,n12540,n12544);
nand (n12536,n12537,n10188);
nor (n12537,n10135,n12538);
not (n12538,n12539);
nand (n12540,n12541,n10193);
nor (n12541,n10135,n12542);
not (n12542,n12543);
nor (n12544,n12545,n12546);
and (n12545,n10228,n12481);
and (n12546,n10222,n12483);
nor (n12547,n12548,n12549);
and (n12548,n10210,n12531);
and (n12549,n10231,n12533);
and (n12550,n12464,n10296);
and (n12551,n12552,n10340);
or (n12552,1'b0,n12553,n12554,n12555,n12556);
and (n12553,n12277,n10073);
and (n12554,n12293,n10091);
and (n12555,n12309,n10109);
and (n12556,n12405,n10005);
and (n12557,n12558,n10339);
or (n12558,1'b0,n12260,n12559,n12556);
and (n12559,n12293,n10270);
and (n12560,n12561,n10337);
or (n12561,1'b0,n12260,n12276,n12292,n12562);
not (n12562,n12563);
or (n12563,n10522,n12564);
not (n12564,n12325);
and (n12565,n12566,n10366);
wire s0n12566,s1n12566,notn12566;
or (n12566,s0n12566,s1n12566);
not(notn12566,n10005);
and (s0n12566,notn12566,1'b0);
and (s1n12566,n10005,n12277);
and (n12567,n12568,n825);
or (n12568,1'b0,n12569,n12571);
and (n12569,n12570,n10109);
wire s0n12570,s1n12570,notn12570;
or (n12570,s0n12570,s1n12570);
not(notn12570,n10374);
and (s0n12570,notn12570,1'b0);
and (s1n12570,n10374,n12370);
and (n12571,n12572,n10005);
wire s0n12572,s1n12572,notn12572;
or (n12572,s0n12572,s1n12572);
not(notn12572,n10379);
and (s0n12572,notn12572,1'b0);
and (s1n12572,n10379,n12293);
and (n12573,n12449,n12574);
and (n12574,n12575,n12783);
wire s0n12575,s1n12575,notn12575;
or (n12575,s0n12575,s1n12575);
not(notn12575,n10395);
and (s0n12575,notn12575,n12576);
and (s1n12575,n10395,n12719);
wire s0n12576,s1n12576,notn12576;
or (n12576,s0n12576,s1n12576);
not(notn12576,n1039);
and (s0n12576,notn12576,n12577);
and (s1n12576,n1039,n12707);
wire s0n12577,s1n12577,notn12577;
or (n12577,s0n12577,s1n12577);
not(notn12577,n10261);
and (s0n12577,notn12577,1'b0);
and (s1n12577,n10261,n12578);
or (n12578,n12579,n12592,n12658,n12696);
and (n12579,n12580,n10021);
wire s0n12580,s1n12580,notn12580;
or (n12580,s0n12580,s1n12580);
not(notn12580,n1057);
and (s0n12580,notn12580,1'b0);
and (s1n12580,n1057,n12581);
wire s0n12581,s1n12581,notn12581;
or (n12581,s0n12581,s1n12581);
not(notn12581,n10004);
and (s0n12581,notn12581,n12582);
and (s1n12581,n10004,n12583);
wire s0n12583,s1n12583,notn12583;
or (n12583,s0n12583,s1n12583);
not(notn12583,n10017);
and (s0n12583,notn12583,n12584);
and (s1n12583,n10017,n12586);
wire s0n12584,s1n12584,notn12584;
or (n12584,s0n12584,s1n12584);
not(notn12584,n10000);
and (s0n12584,notn12584,1'b0);
and (s1n12584,n10000,n12585);
or (n12586,1'b0,n12587,n12589,n12591);
and (n12587,n12588,n10009);
and (n12589,n12590,n10012);
and (n12591,n12585,n10014);
and (n12592,n12593,n10126);
or (n12593,1'b0,n12594,n12610,n12626,n12642);
and (n12594,n12595,n10073);
wire s0n12595,s1n12595,notn12595;
or (n12595,s0n12595,s1n12595);
not(notn12595,n65);
and (s0n12595,notn12595,1'b0);
and (s1n12595,n65,n12596);
wire s0n12596,s1n12596,notn12596;
or (n12596,s0n12596,s1n12596);
not(notn12596,n10068);
and (s0n12596,notn12596,n12597);
and (s1n12596,n10068,n12603);
wire s0n12597,s1n12597,notn12597;
or (n12597,s0n12597,s1n12597);
not(notn12597,n10047);
and (s0n12597,notn12597,1'b0);
and (s1n12597,n10047,n12598);
or (n12598,1'b0,n12599,n12601);
and (n12599,n12600,n10031);
and (n12601,n12602,n10040);
or (n12603,1'b0,n12604,n12606,n12608,n12609);
and (n12604,n12605,n10055);
and (n12606,n12607,n10060);
and (n12608,n12600,n10064);
and (n12609,n12602,n10014);
and (n12610,n12611,n10091);
wire s0n12611,s1n12611,notn12611;
or (n12611,s0n12611,s1n12611);
not(notn12611,n65);
and (s0n12611,notn12611,1'b0);
and (s1n12611,n65,n12612);
wire s0n12612,s1n12612,notn12612;
or (n12612,s0n12612,s1n12612);
not(notn12612,n10068);
and (s0n12612,notn12612,n12613);
and (s1n12612,n10068,n12619);
wire s0n12613,s1n12613,notn12613;
or (n12613,s0n12613,s1n12613);
not(notn12613,n10047);
and (s0n12613,notn12613,1'b0);
and (s1n12613,n10047,n12614);
or (n12614,1'b0,n12615,n12617);
and (n12615,n12616,n10031);
and (n12617,n12618,n10040);
or (n12619,1'b0,n12620,n12622,n12624,n12625);
and (n12620,n12621,n10055);
and (n12622,n12623,n10060);
and (n12624,n12616,n10064);
and (n12625,n12618,n10014);
and (n12626,n12627,n10109);
wire s0n12627,s1n12627,notn12627;
or (n12627,s0n12627,s1n12627);
not(notn12627,n65);
and (s0n12627,notn12627,1'b0);
and (s1n12627,n65,n12628);
wire s0n12628,s1n12628,notn12628;
or (n12628,s0n12628,s1n12628);
not(notn12628,n10068);
and (s0n12628,notn12628,n12629);
and (s1n12628,n10068,n12635);
wire s0n12629,s1n12629,notn12629;
or (n12629,s0n12629,s1n12629);
not(notn12629,n10047);
and (s0n12629,notn12629,1'b0);
and (s1n12629,n10047,n12630);
or (n12630,1'b0,n12631,n12633);
and (n12631,n12632,n10031);
and (n12633,n12634,n10040);
or (n12635,1'b0,n12636,n12638,n12640,n12641);
and (n12636,n12637,n10055);
and (n12638,n12639,n10060);
and (n12640,n12632,n10064);
and (n12641,n12634,n10014);
and (n12642,n12643,n10005);
wire s0n12643,s1n12643,notn12643;
or (n12643,s0n12643,s1n12643);
not(notn12643,n65);
and (s0n12643,notn12643,1'b0);
and (s1n12643,n65,n12644);
wire s0n12644,s1n12644,notn12644;
or (n12644,s0n12644,s1n12644);
not(notn12644,n10068);
and (s0n12644,notn12644,n12645);
and (s1n12644,n10068,n12651);
wire s0n12645,s1n12645,notn12645;
or (n12645,s0n12645,s1n12645);
not(notn12645,n10047);
and (s0n12645,notn12645,1'b0);
and (s1n12645,n10047,n12646);
or (n12646,1'b0,n12647,n12649);
and (n12647,n12648,n10031);
and (n12649,n12650,n10040);
or (n12651,1'b0,n12652,n12654,n12656,n12657);
and (n12652,n12653,n10055);
and (n12654,n12655,n10060);
and (n12656,n12648,n10064);
and (n12657,n12650,n10014);
and (n12658,n12659,n10215);
nand (n12659,n12660,n12682);
nor (n12660,n12661,n12669);
and (n12661,n12662,n10205);
nand (n12662,n12663,n12665,n12667);
nand (n12663,n10136,n12664);
nand (n12665,n10173,n12666);
nand (n12667,n10160,n12668);
nand (n12669,n12670,n12674,n12678);
nand (n12670,n12671,n10188);
nor (n12671,n10135,n12672);
not (n12672,n12673);
nand (n12674,n12675,n10193);
nor (n12675,n10135,n12676);
not (n12676,n12677);
nor (n12678,n12679,n12680);
and (n12679,n10228,n12666);
and (n12680,n10231,n12681);
nor (n12682,n12683,n12692);
and (n12683,n12684,n10177);
nand (n12684,n12685,n12688);
or (n12685,n12686,n10135);
not (n12686,n12687);
nor (n12688,n12689,n12690);
and (n12689,n10160,n12681);
and (n12690,n10173,n12691);
nand (n12692,n12693,n12695);
or (n12693,n12694,n10223);
not (n12694,n12668);
nand (n12695,n10210,n12691);
and (n12696,n12697,n10260);
or (n12697,n12698,n12702,n12705,1'b0);
and (n12698,n12699,n10242);
wire s0n12699,s1n12699,notn12699;
or (n12699,s0n12699,s1n12699);
not(notn12699,n10005);
and (s0n12699,notn12699,n12700);
and (s1n12699,n10005,n12701);
wire s0n12700,s1n12700,notn12700;
or (n12700,s0n12700,s1n12700);
not(notn12700,n10109);
and (s0n12700,notn12700,1'b0);
and (s1n12700,n10109,n12582);
wire s0n12701,s1n12701,notn12701;
or (n12701,s0n12701,s1n12701);
not(notn12701,n10241);
and (s0n12701,notn12701,n12643);
and (s1n12701,n10241,1'b0);
and (n12702,n12703,n10254);
wire s0n12703,s1n12703,notn12703;
or (n12703,s0n12703,s1n12703);
not(notn12703,n10109);
and (s0n12703,notn12703,1'b0);
and (s1n12703,n10109,n12704);
and (n12705,n12706,n10257);
wire s0n12706,s1n12706,notn12706;
or (n12706,s0n12706,s1n12706);
not(notn12706,n10005);
and (s0n12706,notn12706,n12700);
and (s1n12706,n10005,n12643);
or (n12707,n12708,n12709,n12717,n12718);
and (n12708,n12580,n10020);
and (n12709,n12710,n1042);
wire s0n12710,s1n12710,notn12710;
or (n12710,s0n12710,s1n12710);
not(notn12710,n650);
and (s0n12710,notn12710,1'b0);
and (s1n12710,n650,n12711);
or (n12711,1'b0,n12712,n12714,n12715);
and (n12712,n12713,n10073);
wire s0n12713,s1n12713,notn12713;
or (n12713,s0n12713,s1n12713);
not(notn12713,n10259);
and (s0n12713,notn12713,n12582);
and (s1n12713,n10259,1'b0);
and (n12714,n12582,n10270);
and (n12715,n12716,n10005);
wire s0n12716,s1n12716,notn12716;
or (n12716,s0n12716,s1n12716);
not(notn12716,n10148);
and (s0n12716,notn12716,n12662);
and (s1n12716,n10148,1'b0);
and (n12717,n12659,n10181);
and (n12718,n12593,n10072);
or (n12719,1'b0,n12720,n12727,n12735,n12760,n12764,n12769,n12775,n12781,n12782);
and (n12720,n12721,n10286);
or (n12721,1'b0,n12722,n12724,n12726);
and (n12722,n12723,n10073);
and (n12724,n12725,n10091);
and (n12726,n12659,n10284);
and (n12727,n12728,n10296);
or (n12728,1'b0,n12729,n12731,n12733,n12642);
and (n12729,n12730,n10073);
and (n12731,n12732,n10091);
and (n12733,n12734,n10109);
and (n12735,n12736,n10340);
or (n12736,1'b0,n12737,n12738,n12726);
and (n12737,n12643,n10073);
and (n12738,n12739,n10091);
wire s0n12739,s1n12739,notn12739;
or (n12739,s0n12739,s1n12739);
not(notn12739,n10346);
and (s0n12739,notn12739,1'b0);
and (s1n12739,n10346,n12740);
wire s0n12740,s1n12740,notn12740;
or (n12740,s0n12740,s1n12740);
not(notn12740,n51);
and (s0n12740,notn12740,n12741);
and (s1n12740,n51,n12756);
wire s0n12741,s1n12741,notn12741;
or (n12741,s0n12741,s1n12741);
not(notn12741,n10335);
and (s0n12741,notn12741,n12742);
and (s1n12741,n10335,n12744);
wire s0n12742,s1n12742,notn12742;
or (n12742,s0n12742,s1n12742);
not(notn12742,n10020);
and (s0n12742,notn12742,1'b0);
and (s1n12742,n10020,n12743);
or (n12744,n12745,n12747,n12749,n12751,n12753,n12755);
and (n12745,n12746,n10309);
and (n12747,n12748,n10316);
and (n12749,n12750,n10319);
and (n12751,n12752,n10324);
and (n12753,n12754,n10331);
and (n12755,n12743,n10334);
wire s0n12756,s1n12756,notn12756;
or (n12756,s0n12756,s1n12756);
not(notn12756,n10345);
and (s0n12756,notn12756,1'b0);
and (s1n12756,n10345,n12757);
wire s0n12757,s1n12757,notn12757;
or (n12757,s0n12757,s1n12757);
not(notn12757,n10170);
and (s0n12757,notn12757,n12758);
and (s1n12757,n10170,n12759);
and (n12760,n12761,n10339);
or (n12761,1'b0,n12762,n12763);
and (n12762,n12611,n10352);
and (n12763,n12643,n10284);
and (n12764,n12765,n10337);
or (n12765,1'b0,n12766,n12767,n12768);
and (n12766,n12627,n10073);
and (n12767,n12739,n10109);
and (n12768,n12643,n10359);
and (n12769,n12770,n10366);
or (n12770,1'b0,n12771,n12773,n12774,n12642);
and (n12771,n12772,n10073);
and (n12773,n12734,n10091);
and (n12774,n12725,n10109);
and (n12775,n12776,n825);
or (n12776,1'b0,n12777,n12779);
and (n12777,n12778,n10109);
wire s0n12778,s1n12778,notn12778;
or (n12778,s0n12778,s1n12778);
not(notn12778,n10379);
and (s0n12778,notn12778,1'b0);
and (s1n12778,n10379,n12582);
and (n12779,n12780,n10005);
wire s0n12780,s1n12780,notn12780;
or (n12780,s0n12780,s1n12780);
not(notn12780,n10379);
and (s0n12780,notn12780,1'b0);
and (s1n12780,n10379,n12643);
and (n12781,n12659,n10392);
and (n12782,n12593,n10394);
wire s0n12783,s1n12783,notn12783;
or (n12783,s0n12783,s1n12783);
not(notn12783,n10395);
and (s0n12783,notn12783,n12784);
and (s1n12783,n10395,n12818);
wire s0n12784,s1n12784,notn12784;
or (n12784,s0n12784,s1n12784);
not(notn12784,n1039);
and (s0n12784,notn12784,n12785);
and (s1n12784,n1039,n12799);
wire s0n12785,s1n12785,notn12785;
or (n12785,s0n12785,s1n12785);
not(notn12785,n10261);
and (s0n12785,notn12785,1'b0);
and (s1n12785,n10261,n12786);
or (n12786,n12787,1'b0,n12792);
and (n12787,n12788,n10021);
wire s0n12788,s1n12788,notn12788;
or (n12788,s0n12788,s1n12788);
not(notn12788,n1057);
and (s0n12788,notn12788,1'b0);
and (s1n12788,n1057,n12789);
wire s0n12789,s1n12789,notn12789;
or (n12789,s0n12789,s1n12789);
not(notn12789,n10004);
and (s0n12789,notn12789,n12790);
and (s1n12789,n10004,n12791);
and (n12792,n12793,n10260);
or (n12793,n12794,n12797,1'b0);
and (n12794,n12795,n10242);
wire s0n12795,s1n12795,notn12795;
or (n12795,s0n12795,s1n12795);
not(notn12795,n10005);
and (s0n12795,notn12795,n12703);
and (s1n12795,n10005,n12796);
wire s0n12796,s1n12796,notn12796;
or (n12796,s0n12796,s1n12796);
not(notn12796,n10241);
and (s0n12796,notn12796,n12627);
and (s1n12796,n10241,1'b0);
and (n12797,n12798,n10257);
wire s0n12798,s1n12798,notn12798;
or (n12798,s0n12798,s1n12798);
not(notn12798,n10005);
and (s0n12798,notn12798,1'b0);
and (s1n12798,n10005,n12627);
or (n12799,n12800,n12803,1'b0);
and (n12800,n12801,n10020);
wire s0n12801,s1n12801,notn12801;
or (n12801,s0n12801,s1n12801);
not(notn12801,n1057);
and (s0n12801,notn12801,1'b0);
and (s1n12801,n1057,n12802);
wire s0n12802,s1n12802,notn12802;
or (n12802,s0n12802,s1n12802);
not(notn12802,n10417);
and (s0n12802,notn12802,n12790);
and (s1n12802,n10417,n12791);
and (n12803,n12804,n1042);
wire s0n12804,s1n12804,notn12804;
or (n12804,s0n12804,s1n12804);
not(notn12804,n650);
and (s0n12804,notn12804,1'b0);
and (s1n12804,n650,n12805);
or (n12805,1'b0,n12806,n12807,n12809);
and (n12806,n12704,n10352);
and (n12807,n12808,n10109);
wire s0n12808,s1n12808,notn12808;
or (n12808,s0n12808,s1n12808);
not(notn12808,n10243);
and (s0n12808,notn12808,n12634);
and (s1n12808,n10243,1'b0);
and (n12809,n12810,n10005);
wire s0n12810,s1n12810,notn12810;
or (n12810,s0n12810,s1n12810);
not(notn12810,n10148);
and (s0n12810,notn12810,n12811);
and (s1n12810,n10148,1'b0);
nand (n12811,n12812,n12814,n12816);
nand (n12812,n10136,n12813);
nand (n12814,n10173,n12815);
nand (n12816,n10160,n12817);
or (n12818,n12819,n12886,n12887,n12893,n12896,n12901,n12903,1'b0);
and (n12819,n12820,n10286);
or (n12820,1'b0,n12821,n12858);
and (n12821,n12822,n10109);
nand (n12822,n12823,n12838,n12850);
nor (n12823,n12824,n12832);
and (n12824,n12825,n10177);
nand (n12825,n12826,n12828,n12830);
nand (n12826,n10136,n12827);
nand (n12828,n10173,n12829);
nand (n12830,n10160,n12831);
nand (n12832,n12833,n12836);
or (n12833,n12834,n10229);
not (n12834,n12835);
nand (n12836,n10222,n12837);
and (n12838,n12839,n12843,n12847);
nand (n12839,n12840,n10188);
nor (n12840,n10135,n12841);
not (n12841,n12842);
nand (n12843,n12844,n10193);
nor (n12844,n10135,n12845);
not (n12845,n12846);
nor (n12847,n12848,n12849);
and (n12848,n10210,n12829);
and (n12849,n10231,n12831);
nand (n12850,n12851,n10205);
nand (n12851,n12852,n12855);
or (n12852,n12853,n10135);
not (n12853,n12854);
nor (n12855,n12856,n12857);
and (n12856,n10160,n12837);
and (n12857,n10173,n12835);
and (n12858,n12859,n10005);
nand (n12859,n12860,n12870,n12883);
and (n12860,n12861,n12862);
nand (n12861,n12811,n10205);
nand (n12862,n12863,n10177);
nand (n12863,n12864,n12866,n12868);
nand (n12864,n10136,n12865);
nand (n12866,n10173,n12867);
nand (n12868,n10160,n12869);
not (n12870,n12871);
nand (n12871,n12872,n12876,n12880);
nand (n12872,n12873,n10188);
nor (n12873,n10135,n12874);
not (n12874,n12875);
nand (n12876,n12877,n10193);
nor (n12877,n10135,n12878);
not (n12878,n12879);
nor (n12880,n12881,n12882);
and (n12881,n10228,n12815);
and (n12882,n10222,n12817);
nor (n12883,n12884,n12885);
and (n12884,n10210,n12867);
and (n12885,n10231,n12869);
and (n12886,n12798,n10296);
and (n12887,n12888,n10340);
or (n12888,1'b0,n12889,n12890,n12891,n12892);
and (n12889,n12611,n10073);
and (n12890,n12627,n10091);
and (n12891,n12643,n10109);
and (n12892,n12739,n10005);
and (n12893,n12894,n10339);
or (n12894,1'b0,n12594,n12895,n12892);
and (n12895,n12627,n10270);
and (n12896,n12897,n10337);
or (n12897,1'b0,n12594,n12610,n12626,n12898);
not (n12898,n12899);
or (n12899,n10522,n12900);
not (n12900,n12659);
and (n12901,n12902,n10366);
wire s0n12902,s1n12902,notn12902;
or (n12902,s0n12902,s1n12902);
not(notn12902,n10005);
and (s0n12902,notn12902,1'b0);
and (s1n12902,n10005,n12611);
and (n12903,n12904,n825);
or (n12904,1'b0,n12905,n12907);
and (n12905,n12906,n10109);
wire s0n12906,s1n12906,notn12906;
or (n12906,s0n12906,s1n12906);
not(notn12906,n10374);
and (s0n12906,notn12906,1'b0);
and (s1n12906,n10374,n12704);
and (n12907,n12908,n10005);
wire s0n12908,s1n12908,notn12908;
or (n12908,s0n12908,s1n12908);
not(notn12908,n10379);
and (s0n12908,notn12908,1'b0);
and (s1n12908,n10379,n12627);
and (n12909,n12241,n12574);
and (n12910,n11894,n12239);
and (n12911,n11560,n11892);
and (n12912,n11216,n11558);
and (n12913,n10876,n11214);
and (n12914,n10533,n10874);
wire s0n12915,s1n12915,notn12915;
or (n12915,s0n12915,s1n12915);
not(notn12915,n10395);
and (s0n12915,notn12915,n12916);
and (s1n12915,n10395,n12926);
wire s0n12916,s1n12916,notn12916;
or (n12916,s0n12916,s1n12916);
not(notn12916,n1039);
and (s0n12916,notn12916,n12917);
and (s1n12916,n1039,n12921);
and (n12917,n12918,n10261);
or (n12918,1'b0,n12919,n12920);
or (n12919,n10215,n10126);
and (n12920,n10258,n10260);
or (n12921,1'b0,n12922,n12925);
and (n12922,n12923,n1042);
and (n12923,n12924,n650);
and (n12924,n10259,n10073);
not (n12925,n1045);
or (n12926,n12927,1'b0,n12928,n12930,n12934);
and (n12927,n10285,n10286);
and (n12928,n10522,n12929);
or (n12929,n10366,n10296);
and (n12930,n12931,n825);
or (n12931,n10285,n12932,n12933);
and (n12932,n10388,n10109);
and (n12933,n10380,n10005);
or (n12934,n10394,n10392);
wire s0n12935,s1n12935,notn12935;
or (n12935,s0n12935,s1n12935);
not(notn12935,n13324);
and (s0n12935,notn12935,n12936);
and (s1n12935,n13324,n13008);
xor (n12936,n12937,n13005);
xor (n12937,n12938,n12970);
wire s0n12938,s1n12938,notn12938;
or (n12938,s0n12938,s1n12938);
not(notn12938,n10395);
and (s0n12938,notn12938,n12939);
and (s1n12938,n10395,n12956);
wire s0n12939,s1n12939,notn12939;
or (n12939,s0n12939,s1n12939);
not(notn12939,n1039);
and (s0n12939,notn12939,n12940);
and (s1n12939,n1039,n12947);
wire s0n12940,s1n12940,notn12940;
or (n12940,s0n12940,s1n12940);
not(notn12940,n10261);
and (s0n12940,notn12940,1'b0);
and (s1n12940,n10261,n12941);
and (n12941,n12942,n10260);
wire s0n12942,s1n12942,notn12942;
or (n12942,s0n12942,s1n12942);
not(notn12942,n12943);
and (s0n12942,notn12942,1'b0);
and (s1n12942,n12943,n10076);
and (n12943,n10244,n12944);
and (n12944,n10005,n12945);
not (n12945,n12946);
and (n12946,n10241,n10149);
and (n12947,n12948,n1042);
wire s0n12948,s1n12948,notn12948;
or (n12948,s0n12948,s1n12948);
not(notn12948,n650);
and (s0n12948,notn12948,1'b0);
and (s1n12948,n650,n12949);
or (n12949,1'b0,n12950,n12952,n12954);
and (n12950,n12951,n10091);
and (n12952,n12953,n10109);
wire s0n12953,s1n12953,notn12953;
or (n12953,s0n12953,s1n12953);
not(notn12953,n10243);
and (s0n12953,notn12953,n10083);
and (s1n12953,n10243,1'b0);
and (n12954,n12955,n10005);
wire s0n12955,s1n12955,notn12955;
or (n12955,s0n12955,s1n12955);
not(notn12955,n10148);
and (s0n12955,notn12955,n10445);
and (s1n12955,n10148,1'b0);
or (n12956,n12957,n12962,n12965,n12966,n12967,1'b0);
not (n12957,n12958);
or (n12958,n12959,n12960);
not (n12959,n10478);
not (n12960,n12961);
and (n12961,n10109,n10286);
and (n12962,n12963,n10340);
or (n12963,n10356,n12964,n10357,1'b0);
and (n12964,n10111,n10091);
and (n12965,n10509,n10337);
and (n12966,n10412,n10366);
and (n12967,n12968,n825);
and (n12968,n12969,n10005);
wire s0n12969,s1n12969,notn12969;
or (n12969,s0n12969,s1n12969);
not(notn12969,n10379);
and (s0n12969,notn12969,1'b0);
and (s1n12969,n10379,n10076);
nand (n12970,n12971,n12980);
or (n12971,n12972,n12979);
nand (n12972,n12973,n10005);
nand (n12973,n12974,n12976);
or (n12974,n12975,n10380);
not (n12975,n825);
or (n12976,n12977,n12978);
nand (n12977,n10244,n1034);
nor (n12978,n10148,n43,n56);
not (n12979,n10025);
nor (n12980,n12981,n12998,n13001);
and (n12981,n12982,n12991);
nand (n12982,n12983,n12986);
or (n12983,n12984,n10135);
not (n12984,n12985);
nor (n12986,n12987,n12989);
and (n12987,n10160,n12988);
and (n12989,n10173,n12990);
nor (n12991,n12992,n12997);
not (n12992,n12993);
nor (n12993,n12994,n12995);
not (n12994,n1039);
nand (n12995,n10207,n12996,n59,n1045);
nor (n12996,n38,n1044);
nand (n12997,n10149,n10005);
and (n12998,n12999,n10039);
nor (n12999,n13000,n10243);
nand (n13000,n12993,n10109);
and (n13001,n13002,n13004);
not (n13002,n13003);
nand (n13003,n12993,n10091);
or (n13005,n13006,n13323);
and (n13006,n13007,n13051);
xor (n13007,n13008,n13034);
wire s0n13008,s1n13008,notn13008;
or (n13008,s0n13008,s1n13008);
not(notn13008,n10395);
and (s0n13008,notn13008,n13009);
and (s1n13008,n10395,n13022);
wire s0n13009,s1n13009,notn13009;
or (n13009,s0n13009,s1n13009);
not(notn13009,n1039);
and (s0n13009,notn13009,n13010);
and (s1n13009,n1039,n13013);
wire s0n13010,s1n13010,notn13010;
or (n13010,s0n13010,s1n13010);
not(notn13010,n10261);
and (s0n13010,notn13010,1'b0);
and (s1n13010,n10261,n13011);
and (n13011,n13012,n10260);
wire s0n13012,s1n13012,notn13012;
or (n13012,s0n13012,s1n13012);
not(notn13012,n12943);
and (s0n13012,notn13012,1'b0);
and (s1n13012,n12943,n10569);
and (n13013,n13014,n1042);
wire s0n13014,s1n13014,notn13014;
or (n13014,s0n13014,s1n13014);
not(notn13014,n650);
and (s0n13014,notn13014,1'b0);
and (s1n13014,n650,n13015);
or (n13015,1'b0,n13016,n13018,n13020);
and (n13016,n13017,n10091);
and (n13018,n13019,n10109);
wire s0n13019,s1n13019,notn13019;
or (n13019,s0n13019,s1n13019);
not(notn13019,n10243);
and (s0n13019,notn13019,n10576);
and (s1n13019,n10243,1'b0);
and (n13020,n13021,n10005);
wire s0n13021,s1n13021,notn13021;
or (n13021,s0n13021,s1n13021);
not(notn13021,n10148);
and (s0n13021,notn13021,n10786);
and (s1n13021,n10148,1'b0);
or (n13022,n13023,n13026,n13029,n13030,n13031,1'b0);
not (n13023,n13024);
or (n13024,n13025,n12960);
not (n13025,n10823);
and (n13026,n13027,n10340);
or (n13027,n10723,n13028,n10724,1'b0);
and (n13028,n10601,n10091);
and (n13029,n10852,n10337);
and (n13030,n10755,n10366);
and (n13031,n13032,n825);
and (n13032,n13033,n10005);
wire s0n13033,s1n13033,notn13033;
or (n13033,s0n13033,s1n13033);
not(notn13033,n10379);
and (s0n13033,notn13033,1'b0);
and (s1n13033,n10379,n10569);
nand (n13034,n13035,n13037);
or (n13035,n12972,n13036);
not (n13036,n10553);
nor (n13037,n13038,n13048,n13049);
and (n13038,n13039,n12991);
nand (n13039,n13040,n13043);
or (n13040,n13041,n10135);
not (n13041,n13042);
nor (n13043,n13044,n13046);
and (n13044,n10160,n13045);
and (n13046,n10173,n13047);
and (n13048,n12999,n10560);
and (n13049,n13002,n13050);
or (n13051,n13052,n13322);
and (n13052,n13053,n13095);
xor (n13053,n13054,n13078);
wire s0n13054,s1n13054,notn13054;
or (n13054,s0n13054,s1n13054);
not(notn13054,n10395);
and (s0n13054,notn13054,n13055);
and (s1n13054,n10395,n13068);
wire s0n13055,s1n13055,notn13055;
or (n13055,s0n13055,s1n13055);
not(notn13055,n1039);
and (s0n13055,notn13055,n13056);
and (s1n13055,n1039,n13059);
wire s0n13056,s1n13056,notn13056;
or (n13056,s0n13056,s1n13056);
not(notn13056,n10261);
and (s0n13056,notn13056,1'b0);
and (s1n13056,n10261,n13057);
and (n13057,n13058,n10260);
wire s0n13058,s1n13058,notn13058;
or (n13058,s0n13058,s1n13058);
not(notn13058,n12943);
and (s0n13058,notn13058,1'b0);
and (s1n13058,n12943,n10912);
and (n13059,n13060,n1042);
wire s0n13060,s1n13060,notn13060;
or (n13060,s0n13060,s1n13060);
not(notn13060,n650);
and (s0n13060,notn13060,1'b0);
and (s1n13060,n650,n13061);
or (n13061,1'b0,n13062,n13064,n13066);
and (n13062,n13063,n10091);
and (n13064,n13065,n10109);
wire s0n13065,s1n13065,notn13065;
or (n13065,s0n13065,s1n13065);
not(notn13065,n10243);
and (s0n13065,notn13065,n10919);
and (s1n13065,n10243,1'b0);
and (n13066,n13067,n10005);
wire s0n13067,s1n13067,notn13067;
or (n13067,s0n13067,s1n13067);
not(notn13067,n10148);
and (s0n13067,notn13067,n11127);
and (s1n13067,n10148,1'b0);
or (n13068,n13069,n13070,n13073,n13074,n13075,1'b0);
and (n13069,n11160,n12961);
and (n13070,n13071,n10340);
or (n13071,n11066,n13072,n11067,1'b0);
and (n13072,n10944,n10091);
and (n13073,n11192,n10337);
and (n13074,n11098,n10366);
and (n13075,n13076,n825);
and (n13076,n13077,n10005);
wire s0n13077,s1n13077,notn13077;
or (n13077,s0n13077,s1n13077);
not(notn13077,n10379);
and (s0n13077,notn13077,1'b0);
and (s1n13077,n10379,n10912);
nand (n13078,n13079,n13081);
or (n13079,n13080,n12972);
not (n13080,n10896);
nor (n13081,n13082,n13092,n13093);
and (n13082,n13083,n12991);
nand (n13083,n13084,n13087);
or (n13084,n13085,n10135);
not (n13085,n13086);
nor (n13087,n13088,n13090);
and (n13088,n10160,n13089);
and (n13090,n10173,n13091);
and (n13092,n12999,n10903);
and (n13093,n13002,n13094);
or (n13095,n13096,n13321);
and (n13096,n13097,n13141);
xor (n13097,n13098,n13122);
wire s0n13098,s1n13098,notn13098;
or (n13098,s0n13098,s1n13098);
not(notn13098,n10395);
and (s0n13098,notn13098,n13099);
and (s1n13098,n10395,n13112);
wire s0n13099,s1n13099,notn13099;
or (n13099,s0n13099,s1n13099);
not(notn13099,n1039);
and (s0n13099,notn13099,n13100);
and (s1n13099,n1039,n13103);
wire s0n13100,s1n13100,notn13100;
or (n13100,s0n13100,s1n13100);
not(notn13100,n10261);
and (s0n13100,notn13100,1'b0);
and (s1n13100,n10261,n13101);
and (n13101,n13102,n10260);
wire s0n13102,s1n13102,notn13102;
or (n13102,s0n13102,s1n13102);
not(notn13102,n12943);
and (s0n13102,notn13102,1'b0);
and (s1n13102,n12943,n11252);
and (n13103,n13104,n1042);
wire s0n13104,s1n13104,notn13104;
or (n13104,s0n13104,s1n13104);
not(notn13104,n650);
and (s0n13104,notn13104,1'b0);
and (s1n13104,n650,n13105);
or (n13105,1'b0,n13106,n13108,n13110);
and (n13106,n13107,n10091);
and (n13108,n13109,n10109);
wire s0n13109,s1n13109,notn13109;
or (n13109,s0n13109,s1n13109);
not(notn13109,n10243);
and (s0n13109,notn13109,n11259);
and (s1n13109,n10243,1'b0);
and (n13110,n13111,n10005);
wire s0n13111,s1n13111,notn13111;
or (n13111,s0n13111,s1n13111);
not(notn13111,n10148);
and (s0n13111,notn13111,n11469);
and (s1n13111,n10148,1'b0);
or (n13112,n13113,n13114,n13117,n13118,n13119,1'b0);
and (n13113,n11504,n12961);
and (n13114,n13115,n10340);
or (n13115,n11408,n13116,n11409,1'b0);
and (n13116,n11284,n10091);
and (n13117,n11536,n10337);
and (n13118,n11440,n10366);
and (n13119,n13120,n825);
and (n13120,n13121,n10005);
wire s0n13121,s1n13121,notn13121;
or (n13121,s0n13121,s1n13121);
not(notn13121,n10379);
and (s0n13121,notn13121,1'b0);
and (s1n13121,n10379,n11252);
nand (n13122,n13123,n13125);
or (n13123,n12972,n13124);
not (n13124,n11236);
nor (n13125,n13126,n13136);
and (n13126,n13127,n12991);
nand (n13127,n13128,n13131);
or (n13128,n13129,n10135);
not (n13129,n13130);
nor (n13131,n13132,n13134);
and (n13132,n10160,n13133);
and (n13134,n10173,n13135);
not (n13136,n13137);
nor (n13137,n13138,n13139);
and (n13138,n12999,n11243);
and (n13139,n13002,n13140);
or (n13141,n13142,n13320);
and (n13142,n13143,n13186);
xor (n13143,n13144,n13168);
wire s0n13144,s1n13144,notn13144;
or (n13144,s0n13144,s1n13144);
not(notn13144,n10395);
and (s0n13144,notn13144,n13145);
and (s1n13144,n10395,n13158);
wire s0n13145,s1n13145,notn13145;
or (n13145,s0n13145,s1n13145);
not(notn13145,n1039);
and (s0n13145,notn13145,n13146);
and (s1n13145,n1039,n13149);
wire s0n13146,s1n13146,notn13146;
or (n13146,s0n13146,s1n13146);
not(notn13146,n10261);
and (s0n13146,notn13146,1'b0);
and (s1n13146,n10261,n13147);
and (n13147,n13148,n10260);
wire s0n13148,s1n13148,notn13148;
or (n13148,s0n13148,s1n13148);
not(notn13148,n12943);
and (s0n13148,notn13148,1'b0);
and (s1n13148,n12943,n11596);
and (n13149,n13150,n1042);
wire s0n13150,s1n13150,notn13150;
or (n13150,s0n13150,s1n13150);
not(notn13150,n650);
and (s0n13150,notn13150,1'b0);
and (s1n13150,n650,n13151);
or (n13151,1'b0,n13152,n13154,n13156);
and (n13152,n13153,n10091);
and (n13154,n13155,n10109);
wire s0n13155,s1n13155,notn13155;
or (n13155,s0n13155,s1n13155);
not(notn13155,n10243);
and (s0n13155,notn13155,n11603);
and (s1n13155,n10243,1'b0);
and (n13156,n13157,n10005);
wire s0n13157,s1n13157,notn13157;
or (n13157,s0n13157,s1n13157);
not(notn13157,n10148);
and (s0n13157,notn13157,n11838);
and (s1n13157,n10148,1'b0);
or (n13158,n13159,n13160,n13163,n13164,n13165,1'b0);
and (n13159,n11844,n12961);
and (n13160,n13161,n10340);
or (n13161,n11751,n13162,n11752,1'b0);
and (n13162,n11628,n10091);
and (n13163,n11872,n10337);
and (n13164,n11783,n10366);
and (n13165,n13166,n825);
and (n13166,n13167,n10005);
wire s0n13167,s1n13167,notn13167;
or (n13167,s0n13167,s1n13167);
not(notn13167,n10379);
and (s0n13167,notn13167,1'b0);
and (s1n13167,n10379,n11596);
nand (n13168,n13169,n13171);
or (n13169,n13170,n12972);
not (n13170,n11580);
and (n13171,n13172,n13182);
nand (n13172,n13173,n12991);
nand (n13173,n13174,n13177);
or (n13174,n13175,n10135);
not (n13175,n13176);
nor (n13177,n13178,n13180);
and (n13178,n10160,n13179);
and (n13180,n10173,n13181);
nor (n13182,n13183,n13184);
and (n13183,n12999,n11587);
and (n13184,n13002,n13185);
or (n13186,n13187,n13319);
and (n13187,n13188,n13231);
xor (n13188,n13189,n13213);
wire s0n13189,s1n13189,notn13189;
or (n13189,s0n13189,s1n13189);
not(notn13189,n10395);
and (s0n13189,notn13189,n13190);
and (s1n13189,n10395,n13203);
wire s0n13190,s1n13190,notn13190;
or (n13190,s0n13190,s1n13190);
not(notn13190,n1039);
and (s0n13190,notn13190,n13191);
and (s1n13190,n1039,n13194);
wire s0n13191,s1n13191,notn13191;
or (n13191,s0n13191,s1n13191);
not(notn13191,n10261);
and (s0n13191,notn13191,1'b0);
and (s1n13191,n10261,n13192);
and (n13192,n13193,n10260);
wire s0n13193,s1n13193,notn13193;
or (n13193,s0n13193,s1n13193);
not(notn13193,n12943);
and (s0n13193,notn13193,1'b0);
and (s1n13193,n12943,n11930);
and (n13194,n13195,n1042);
wire s0n13195,s1n13195,notn13195;
or (n13195,s0n13195,s1n13195);
not(notn13195,n650);
and (s0n13195,notn13195,1'b0);
and (s1n13195,n650,n13196);
or (n13196,1'b0,n13197,n13199,n13201);
and (n13197,n13198,n10091);
and (n13199,n13200,n10109);
wire s0n13200,s1n13200,notn13200;
or (n13200,s0n13200,s1n13200);
not(notn13200,n10243);
and (s0n13200,notn13200,n11937);
and (s1n13200,n10243,1'b0);
and (n13201,n13202,n10005);
wire s0n13202,s1n13202,notn13202;
or (n13202,s0n13202,s1n13202);
not(notn13202,n10148);
and (s0n13202,notn13202,n12168);
and (s1n13202,n10148,1'b0);
or (n13203,n13204,n13205,n13208,n13209,n13210,1'b0);
and (n13204,n12183,n12961);
and (n13205,n13206,n10340);
or (n13206,n12090,n13207,n12091,1'b0);
and (n13207,n11962,n10091);
and (n13208,n12213,n10337);
and (n13209,n12122,n10366);
and (n13210,n13211,n825);
and (n13211,n13212,n10005);
wire s0n13212,s1n13212,notn13212;
or (n13212,s0n13212,s1n13212);
not(notn13212,n10379);
and (s0n13212,notn13212,1'b0);
and (s1n13212,n10379,n11930);
nand (n13213,n13214,n13216);
or (n13214,n12972,n13215);
not (n13215,n11914);
nor (n13216,n13217,n13225);
and (n13217,n13218,n12991);
nand (n13218,n13219,n13221,n13223);
nand (n13219,n10136,n13220);
nand (n13221,n10173,n13222);
nand (n13223,n10160,n13224);
nand (n13225,n13226,n13229);
or (n13226,n13227,n13228);
not (n13227,n12999);
not (n13228,n11921);
nand (n13229,n13002,n13230);
nand (n13231,n13232,n13318);
or (n13232,n13233,n13283);
nand (n13233,n13234,n13267);
nand (n13234,n13235,n13239,n13246,n13262);
nand (n13235,n12739,n13236);
nand (n13236,n13237,n13238);
nand (n13237,n10340,n10109);
nand (n13238,n10337,n10005);
nand (n13239,n13240,n12627);
nand (n13240,n13241,n13245);
and (n13241,n13242,n13243);
nand (n13242,n10340,n10073);
not (n13243,n13244);
and (n13244,n10005,n10366);
nand (n13245,n10337,n10091);
nor (n13246,n13247,n13252);
and (n13247,n13248,n12611);
nand (n13248,n12972,n13249);
nand (n13249,n10336,n13250);
nor (n13250,n826,n13251);
not (n13251,n10073);
nand (n13252,n13253,n13255);
or (n13253,n12960,n13254);
not (n13254,n12859);
nor (n13255,n13256,n13257);
and (n13256,n12851,n12991);
nand (n13257,n13258,n13260);
or (n13258,n13259,n13227);
not (n13259,n12618);
nand (n13260,n13002,n13261);
nand (n13262,n13263,n12643);
nand (n13263,n13264,n13266);
or (n13264,n1050,n13265);
not (n13265,n10337);
nand (n13266,n10340,n10091);
nand (n13267,n13268,n13270);
or (n13268,n12972,n13269);
not (n13269,n12595);
and (n13270,n13271,n13279);
nand (n13271,n13272,n12991);
nand (n13272,n13273,n13275,n13277);
nand (n13273,n10136,n13274);
nand (n13275,n10173,n13276);
nand (n13277,n10160,n13278);
nor (n13279,n13280,n13281);
and (n13280,n12999,n12602);
and (n13281,n13002,n13282);
nor (n13283,n13284,n13300);
nand (n13284,n13285,n13286,n13287,n13299);
nand (n13285,n12405,n13236);
nand (n13286,n13240,n12293);
nor (n13287,n13288,n13289);
and (n13288,n13248,n12277);
nand (n13289,n13290,n13292);
or (n13290,n12960,n13291);
not (n13291,n12524);
nor (n13292,n13293,n13294);
and (n13293,n12491,n12991);
nand (n13294,n13295,n13297);
or (n13295,n13296,n13227);
not (n13296,n12284);
nand (n13297,n13002,n13298);
nand (n13299,n13263,n12309);
nand (n13300,n13301,n13303);
or (n13301,n12972,n13302);
not (n13302,n12261);
and (n13303,n13304,n13314);
nand (n13304,n13305,n12991);
nand (n13305,n13306,n13309);
or (n13306,n13307,n10135);
not (n13307,n13308);
nor (n13309,n13310,n13312);
and (n13310,n10160,n13311);
and (n13312,n10173,n13313);
nor (n13314,n13315,n13316);
and (n13315,n12999,n12268);
and (n13316,n13002,n13317);
nand (n13318,n13284,n13300);
and (n13319,n13189,n13213);
and (n13320,n13144,n13168);
and (n13321,n13098,n13122);
and (n13322,n13054,n13078);
and (n13323,n13008,n13034);
or (n13324,n12961,n13325,n13327,n13244,1'b0,1'b0);
and (n13325,n13326,n10340);
or (n13326,n10270,n10073);
and (n13327,n1057,n10337);
or (n13328,n13329,n13335,n13388);
and (n13329,n13330,n13333);
wire s0n13330,s1n13330,notn13330;
or (n13330,s0n13330,s1n13330);
not(notn13330,n12915);
and (s0n13330,notn13330,n13331);
and (s1n13330,n12915,1'b0);
xor (n13331,n13332,n10874);
xor (n13332,n10533,n10740);
wire s0n13333,s1n13333,notn13333;
or (n13333,s0n13333,s1n13333);
not(notn13333,n13324);
and (s0n13333,notn13333,n13334);
and (s1n13333,n13324,n13054);
xor (n13334,n13007,n13051);
and (n13335,n13333,n13336);
or (n13336,n13337,n13343,n13387);
and (n13337,n13338,n13341);
wire s0n13338,s1n13338,notn13338;
or (n13338,s0n13338,s1n13338);
not(notn13338,n12915);
and (s0n13338,notn13338,n13339);
and (s1n13338,n12915,1'b0);
xor (n13339,n13340,n11214);
xor (n13340,n10876,n11083);
wire s0n13341,s1n13341,notn13341;
or (n13341,s0n13341,s1n13341);
not(notn13341,n13324);
and (s0n13341,notn13341,n13342);
and (s1n13341,n13324,n13098);
xor (n13342,n13053,n13095);
and (n13343,n13341,n13344);
or (n13344,n13345,n13351,n13386);
and (n13345,n13346,n13349);
wire s0n13346,s1n13346,notn13346;
or (n13346,s0n13346,s1n13346);
not(notn13346,n12915);
and (s0n13346,notn13346,n13347);
and (s1n13346,n12915,1'b0);
xor (n13347,n13348,n11558);
xor (n13348,n11216,n11425);
wire s0n13349,s1n13349,notn13349;
or (n13349,s0n13349,s1n13349);
not(notn13349,n13324);
and (s0n13349,notn13349,n13350);
and (s1n13349,n13324,n13144);
xor (n13350,n13097,n13141);
and (n13351,n13349,n13352);
or (n13352,n13353,n13359,n13385);
and (n13353,n13354,n13357);
wire s0n13354,s1n13354,notn13354;
or (n13354,s0n13354,s1n13354);
not(notn13354,n12915);
and (s0n13354,notn13354,n13355);
and (s1n13354,n12915,1'b0);
xor (n13355,n13356,n11892);
xor (n13356,n11560,n11768);
wire s0n13357,s1n13357,notn13357;
or (n13357,s0n13357,s1n13357);
not(notn13357,n13324);
and (s0n13357,notn13357,n13358);
and (s1n13357,n13324,n13189);
xor (n13358,n13143,n13186);
and (n13359,n13357,n13360);
or (n13360,n13361,n13367,n13384);
and (n13361,n13362,n13365);
wire s0n13362,s1n13362,notn13362;
or (n13362,s0n13362,s1n13362);
not(notn13362,n12915);
and (s0n13362,notn13362,n13363);
and (s1n13362,n12915,1'b0);
xor (n13363,n13364,n12239);
xor (n13364,n11894,n12107);
wire s0n13365,s1n13365,notn13365;
or (n13365,s0n13365,s1n13365);
not(notn13365,n13324);
and (s0n13365,notn13365,n13366);
and (s1n13365,n13324,n13284);
xor (n13366,n13188,n13231);
and (n13367,n13365,n13368);
or (n13368,n13369,n13377,n13383);
and (n13369,n13370,n13373);
wire s0n13370,s1n13370,notn13370;
or (n13370,s0n13370,s1n13370);
not(notn13370,n12915);
and (s0n13370,notn13370,n13371);
and (s1n13370,n12915,1'b0);
xor (n13371,n13372,n12574);
xor (n13372,n12241,n12449);
wire s0n13373,s1n13373,notn13373;
or (n13373,s0n13373,s1n13373);
not(notn13373,n13324);
and (s0n13373,notn13373,n13374);
and (s1n13373,n13324,n13234);
xor (n13374,n13375,n13376);
xor (n13375,n13284,n13300);
not (n13376,n13233);
and (n13377,n13373,n13378);
and (n13378,n13379,n13381);
wire s0n13379,s1n13379,notn13379;
or (n13379,s0n13379,s1n13379);
not(notn13379,n12915);
and (s0n13379,notn13379,n13380);
and (s1n13379,n12915,1'b0);
xor (n13380,n12575,n12783);
wire s0n13381,s1n13381,notn13381;
or (n13381,s0n13381,s1n13381);
not(notn13381,n13324);
and (s0n13381,notn13381,n13382);
and (s1n13381,n13324,1'b0);
xor (n13382,n13267,n13234);
and (n13383,n13370,n13378);
and (n13384,n13362,n13368);
and (n13385,n13354,n13360);
and (n13386,n13346,n13352);
and (n13387,n13338,n13344);
and (n13388,n13330,n13336);
and (n13389,n13390,n13392);
xor (n13390,n13391,n13336);
xor (n13391,n13330,n13333);
and (n13392,n13393,n13395);
xor (n13393,n13394,n13344);
xor (n13394,n13338,n13341);
or (n13395,n13396,n13407,n13454);
and (n13396,n13397,n13399);
xor (n13397,n13398,n13352);
xor (n13398,n13346,n13349);
wire s0n13399,s1n13399,notn13399;
or (n13399,s0n13399,s1n13399);
not(notn13399,n1039);
and (s0n13399,notn13399,n13400);
and (s1n13399,n1039,n13402);
and (n13400,n13401,n10261);
and (n13401,n1057,n10021);
or (n13402,n13403,n13404,1'b0);
and (n13403,n1057,n10020);
and (n13404,n13405,n1042);
wire s0n13405,s1n13405,notn13405;
or (n13405,s0n13405,s1n13405);
not(notn13405,n650);
and (s0n13405,notn13405,1'b0);
and (s1n13405,n650,n13406);
and (n13406,n10242,n10073);
and (n13407,n13399,n13408);
or (n13408,n13409,n13417,n13453);
and (n13409,n13410,n13412);
xor (n13410,n13411,n13360);
xor (n13411,n13354,n13357);
wire s0n13412,s1n13412,notn13412;
or (n13412,s0n13412,s1n13412);
not(notn13412,n1039);
and (s0n13412,notn13412,1'b0);
and (s1n13412,n1039,n13413);
and (n13413,n13414,n1042);
wire s0n13414,s1n13414,notn13414;
or (n13414,s0n13414,s1n13414);
not(notn13414,n650);
and (s0n13414,notn13414,1'b0);
and (s1n13414,n650,n13415);
and (n13415,n13416,n10073);
not (n13416,n10242);
and (n13417,n13412,n13418);
or (n13418,n13419,n13430,n13452);
and (n13419,n13420,n13422);
xor (n13420,n13421,n13368);
xor (n13421,n13362,n13365);
nand (n13422,n13423,n13428);
or (n13423,n13424,n13426);
nand (n13424,n58,n10149,n13425,n43);
not (n13425,n47);
not (n13426,n13427);
nor (n13427,n12977,n1050);
or (n13428,n13429,n10380);
nand (n13429,n825,n10374,n10109);
and (n13430,n13422,n13431);
or (n13431,n13432,n13443,n13451);
and (n13432,n13433,n13435);
xor (n13433,n13434,n13378);
xor (n13434,n13370,n13373);
or (n13435,n13324,n13436);
nand (n13436,n13437,n13438);
or (n13437,n13429,n10379);
nor (n13438,n13439,n13440,n13441);
and (n13439,n13427,n13424);
nor (n13440,n12974,n10374,n1050);
and (n13441,n10243,n13442,n10149);
and (n13442,n1034,n10109);
and (n13443,n13435,n13444);
and (n13444,n13445,n13446);
xor (n13445,n13379,n13381);
or (n13446,n13447,n13448,n13449,n13450,1'b0,1'b0,1'b0,1'b0);
and (n13447,n10005,n10286);
and (n13448,n10005,n10296);
and (n13449,n10005,n10340);
and (n13450,n1057,n10339);
and (n13451,n13433,n13444);
and (n13452,n13420,n13431);
and (n13453,n13410,n13418);
and (n13454,n13397,n13408);
xor (n13455,n13456,n13538);
xor (n13456,n13457,n13534);
xor (n13457,n13458,n13518);
wire s0n13458,s1n13458,notn13458;
or (n13458,s0n13458,s1n13458);
not(notn13458,n12915);
and (s0n13458,notn13458,n13459);
and (s1n13458,n12915,1'b0);
xor (n13459,n13460,n13514);
xor (n13460,n13461,n13490);
nand (n13461,n13462,n13478);
or (n13462,n13463,n13465);
not (n13463,n13464);
not (n13465,n13466);
nand (n13466,n13467,n13469);
nand (n13467,n13468,n10109);
nand (n13468,n12974,n12977);
nor (n13469,n13470,n13473);
nor (n13470,n13471,n10004);
not (n13471,n13472);
wire s0n13472,s1n13472,notn13472;
or (n13472,s0n13472,s1n13472);
not(notn13472,n1039);
and (s0n13472,notn13472,n13400);
and (s1n13472,n1039,n13403);
nand (n13473,n13474,n13477);
or (n13474,n13475,n10259,n10005);
or (n13475,n12992,n13476);
nor (n13476,n10005,n13326);
or (n13477,n12992,n10271);
nor (n13478,n13479,n13481);
and (n13479,n13441,n13480);
wire s0n13481,s1n13481,notn13481;
or (n13481,s0n13481,s1n13481);
not(notn13481,n10017);
and (s0n13481,notn13481,n13482);
and (s1n13481,n10017,n13484);
wire s0n13482,s1n13482,notn13482;
or (n13482,s0n13482,s1n13482);
not(notn13482,n10000);
and (s0n13482,notn13482,1'b0);
and (s1n13482,n10000,n13483);
or (n13484,1'b0,n13485,n13487,n13489);
and (n13485,n13486,n10009);
and (n13487,n13488,n10012);
and (n13489,n13483,n10014);
nand (n13490,n13491,n13497,n13504);
nand (n13491,n13492,n13480);
nand (n13492,n13429,n13493);
nor (n13493,n13494,n13496);
and (n13494,n13495,n10285);
not (n13495,n13475);
and (n13496,n13427,n10149);
nand (n13497,n13498,n13503);
nand (n13498,n13499,n13500);
not (n13499,n13470);
nand (n13500,n13501,n1057,n60);
not (n13501,n13502);
nand (n13502,n1039,n10020);
nand (n13504,n13505,n13513);
and (n13505,n13506,n13510,n13511);
nand (n13506,n13507,n60);
nor (n13507,n926,n13508);
or (n13508,n13509,n51);
not (n13509,n10020);
or (n13510,n10345,n13507);
nor (n13511,n13512,n38);
nand (n13512,n65,n10005);
or (n13514,n13515,n13516,n13517);
and (n13515,n9989,n10397);
and (n13516,n10397,n10531);
and (n13517,n9989,n10531);
wire s0n13518,s1n13518,notn13518;
or (n13518,s0n13518,s1n13518);
not(notn13518,n13324);
and (s0n13518,notn13518,n13519);
and (s1n13518,n13324,n12938);
xor (n13519,n13520,n13531);
xor (n13520,n13521,n13526);
wire s0n13521,s1n13521,notn13521;
or (n13521,s0n13521,s1n13521);
not(notn13521,n1039);
and (s0n13521,notn13521,1'b0);
and (s1n13521,n1039,n13522);
and (n13522,n13523,n1042);
wire s0n13523,s1n13523,notn13523;
or (n13523,s0n13523,s1n13523);
not(notn13523,n650);
and (s0n13523,notn13523,1'b0);
and (s1n13523,n650,n13524);
and (n13524,n13525,n10091);
wire s0n13526,s1n13526,notn13526;
or (n13526,s0n13526,s1n13526);
not(notn13526,n1039);
and (s0n13526,notn13526,1'b0);
and (s1n13526,n1039,n13527);
and (n13527,n13528,n1042);
wire s0n13528,s1n13528,notn13528;
or (n13528,s0n13528,s1n13528);
not(notn13528,n650);
and (s0n13528,notn13528,1'b0);
and (s1n13528,n650,n13529);
and (n13529,n13530,n10091);
or (n13531,n13532,n13533);
and (n13532,n12937,n13005);
and (n13533,n12938,n12970);
or (n13534,n13535,n13536,n13537);
and (n13535,n9986,n12935);
and (n13536,n12935,n13328);
and (n13537,n9986,n13328);
and (n13538,n9984,n13389);
or (n13539,n13446,n13422,n13399);
wire s0n13540,s1n13540,notn13540;
or (n13540,s0n13540,s1n13540);
not(notn13540,n13539);
and (s0n13540,notn13540,n13541);
and (s1n13540,n13539,n13593);
xor (n13541,n13542,n13592);
xor (n13542,n13543,n13588);
xor (n13543,n13544,n13573);
wire s0n13544,s1n13544,notn13544;
or (n13544,s0n13544,s1n13544);
not(notn13544,n12915);
and (s0n13544,notn13544,n13545);
and (s1n13544,n12915,1'b0);
xor (n13545,n13546,n13569);
xor (n13546,n13547,n13563);
nand (n13547,n13548,n13551);
or (n13548,n13549,n13465);
not (n13549,n13550);
nor (n13551,n13552,n13554);
and (n13552,n13441,n13553);
wire s0n13554,s1n13554,notn13554;
or (n13554,s0n13554,s1n13554);
not(notn13554,n10017);
and (s0n13554,notn13554,n13555);
and (s1n13554,n10017,n13557);
wire s0n13555,s1n13555,notn13555;
or (n13555,s0n13555,s1n13555);
not(notn13555,n10000);
and (s0n13555,notn13555,1'b0);
and (s1n13555,n10000,n13556);
or (n13557,1'b0,n13558,n13560,n13562);
and (n13558,n13559,n10009);
and (n13560,n13561,n10012);
and (n13562,n13556,n10014);
nand (n13563,n13564,n13565,n13567);
nand (n13564,n13492,n13553);
nand (n13565,n13498,n13566);
nand (n13567,n13505,n13568);
or (n13569,n13570,n13571,n13572);
and (n13570,n13461,n13490);
and (n13571,n13490,n13514);
and (n13572,n13461,n13514);
xor (n13573,n13574,n13585);
xor (n13574,n13575,n13580);
wire s0n13575,s1n13575,notn13575;
or (n13575,s0n13575,s1n13575);
not(notn13575,n1039);
and (s0n13575,notn13575,1'b0);
and (s1n13575,n1039,n13576);
and (n13576,n13577,n1042);
wire s0n13577,s1n13577,notn13577;
or (n13577,s0n13577,s1n13577);
not(notn13577,n650);
and (s0n13577,notn13577,1'b0);
and (s1n13577,n650,n13578);
and (n13578,n13579,n10091);
wire s0n13580,s1n13580,notn13580;
or (n13580,s0n13580,s1n13580);
not(notn13580,n1039);
and (s0n13580,notn13580,1'b0);
and (s1n13580,n1039,n13581);
and (n13581,n13582,n1042);
wire s0n13582,s1n13582,notn13582;
or (n13582,s0n13582,s1n13582);
not(notn13582,n650);
and (s0n13582,notn13582,1'b0);
and (s1n13582,n650,n13583);
and (n13583,n13584,n10091);
or (n13585,n13586,n13587);
and (n13586,n13520,n13531);
and (n13587,n13521,n13526);
or (n13588,n13589,n13590,n13591);
and (n13589,n13458,n13518);
and (n13590,n13518,n13534);
and (n13591,n13458,n13534);
and (n13592,n13456,n13538);
xor (n13593,n13594,n13644);
xor (n13594,n13595,n13640);
xor (n13595,n13596,n13625);
wire s0n13596,s1n13596,notn13596;
or (n13596,s0n13596,s1n13596);
not(notn13596,n12915);
and (s0n13596,notn13596,n13597);
and (s1n13596,n12915,1'b0);
xor (n13597,n13598,n13621);
xor (n13598,n13599,n13615);
nand (n13599,n13600,n13603);
or (n13600,n13601,n13465);
not (n13601,n13602);
nor (n13603,n13604,n13606);
and (n13604,n13441,n13605);
wire s0n13606,s1n13606,notn13606;
or (n13606,s0n13606,s1n13606);
not(notn13606,n10017);
and (s0n13606,notn13606,n13607);
and (s1n13606,n10017,n13609);
wire s0n13607,s1n13607,notn13607;
or (n13607,s0n13607,s1n13607);
not(notn13607,n10000);
and (s0n13607,notn13607,1'b0);
and (s1n13607,n10000,n13608);
or (n13609,1'b0,n13610,n13612,n13614);
and (n13610,n13611,n10009);
and (n13612,n13613,n10012);
and (n13614,n13608,n10014);
nand (n13615,n13616,n13617,n13619);
nand (n13616,n13492,n13605);
nand (n13617,n13498,n13618);
nand (n13619,n13505,n13620);
or (n13621,n13622,n13623,n13624);
and (n13622,n13547,n13563);
and (n13623,n13563,n13569);
and (n13624,n13547,n13569);
xor (n13625,n13626,n13637);
xor (n13626,n13627,n13632);
wire s0n13627,s1n13627,notn13627;
or (n13627,s0n13627,s1n13627);
not(notn13627,n1039);
and (s0n13627,notn13627,1'b0);
and (s1n13627,n1039,n13628);
and (n13628,n13629,n1042);
wire s0n13629,s1n13629,notn13629;
or (n13629,s0n13629,s1n13629);
not(notn13629,n650);
and (s0n13629,notn13629,1'b0);
and (s1n13629,n650,n13630);
and (n13630,n13631,n10091);
wire s0n13632,s1n13632,notn13632;
or (n13632,s0n13632,s1n13632);
not(notn13632,n1039);
and (s0n13632,notn13632,1'b0);
and (s1n13632,n1039,n13633);
and (n13633,n13634,n1042);
wire s0n13634,s1n13634,notn13634;
or (n13634,s0n13634,s1n13634);
not(notn13634,n650);
and (s0n13634,notn13634,1'b0);
and (s1n13634,n650,n13635);
and (n13635,n13636,n10091);
or (n13637,n13638,n13639);
and (n13638,n13574,n13585);
and (n13639,n13575,n13580);
or (n13640,n13641,n13642,n13643);
and (n13641,n13544,n13573);
and (n13642,n13573,n13588);
and (n13643,n13544,n13588);
and (n13644,n13542,n13592);
or (n13645,n13324,n13646);
nand (n13646,n13467,n13429,n13647);
not (n13647,n13441);
wire s0n13648,s1n13648,notn13648;
or (n13648,s0n13648,s1n13648);
not(notn13648,n13645);
and (s0n13648,notn13648,n13649);
and (s1n13648,n13645,n13755);
wire s0n13649,s1n13649,notn13649;
or (n13649,s0n13649,s1n13649);
not(notn13649,n13539);
and (s0n13649,notn13649,n13650);
and (s1n13649,n13539,n13706);
xor (n13650,n13651,n13705);
xor (n13651,n13652,n13701);
xor (n13652,n13653,n13686);
wire s0n13653,s1n13653,notn13653;
or (n13653,s0n13653,s1n13653);
not(notn13653,n12915);
and (s0n13653,notn13653,n13654);
and (s1n13653,n12915,1'b0);
xor (n13654,n13655,n13682);
xor (n13655,n13656,n13672);
nand (n13656,n13657,n13660);
or (n13657,n13658,n13465);
not (n13658,n13659);
nor (n13660,n13661,n13663);
and (n13661,n13441,n13662);
wire s0n13663,s1n13663,notn13663;
or (n13663,s0n13663,s1n13663);
not(notn13663,n10017);
and (s0n13663,notn13663,n13664);
and (s1n13663,n10017,n13666);
wire s0n13664,s1n13664,notn13664;
or (n13664,s0n13664,s1n13664);
not(notn13664,n10000);
and (s0n13664,notn13664,1'b0);
and (s1n13664,n10000,n13665);
or (n13666,1'b0,n13667,n13669,n13671);
and (n13667,n13668,n10009);
and (n13669,n13670,n10012);
and (n13671,n13665,n10014);
nand (n13672,n13673,n13676);
or (n13673,n13674,n13675);
not (n13674,n13662);
not (n13675,n13492);
not (n13676,n13677);
nand (n13677,n13678,n13680);
nand (n13678,n13498,n13679);
nand (n13680,n13505,n13681);
or (n13682,n13683,n13684,n13685);
and (n13683,n13599,n13615);
and (n13684,n13615,n13621);
and (n13685,n13599,n13621);
xor (n13686,n13687,n13698);
xor (n13687,n13688,n13693);
wire s0n13688,s1n13688,notn13688;
or (n13688,s0n13688,s1n13688);
not(notn13688,n1039);
and (s0n13688,notn13688,1'b0);
and (s1n13688,n1039,n13689);
and (n13689,n13690,n1042);
wire s0n13690,s1n13690,notn13690;
or (n13690,s0n13690,s1n13690);
not(notn13690,n650);
and (s0n13690,notn13690,1'b0);
and (s1n13690,n650,n13691);
and (n13691,n13692,n10091);
wire s0n13693,s1n13693,notn13693;
or (n13693,s0n13693,s1n13693);
not(notn13693,n1039);
and (s0n13693,notn13693,1'b0);
and (s1n13693,n1039,n13694);
and (n13694,n13695,n1042);
wire s0n13695,s1n13695,notn13695;
or (n13695,s0n13695,s1n13695);
not(notn13695,n650);
and (s0n13695,notn13695,1'b0);
and (s1n13695,n650,n13696);
and (n13696,n13697,n10091);
or (n13698,n13699,n13700);
and (n13699,n13626,n13637);
and (n13700,n13627,n13632);
or (n13701,n13702,n13703,n13704);
and (n13702,n13596,n13625);
and (n13703,n13625,n13640);
and (n13704,n13596,n13640);
and (n13705,n13594,n13644);
xor (n13706,n13707,n13754);
xor (n13707,n13708,n13750);
xor (n13708,n13709,n13735);
wire s0n13709,s1n13709,notn13709;
or (n13709,s0n13709,s1n13709);
not(notn13709,n12915);
and (s0n13709,notn13709,n13710);
and (s1n13709,n12915,1'b0);
xor (n13710,n13711,n13731);
xor (n13711,n13712,n13728);
nand (n13712,n13713,n13716);
or (n13713,n13714,n13465);
not (n13714,n13715);
nor (n13716,n13717,n13719);
and (n13717,n13441,n13718);
wire s0n13719,s1n13719,notn13719;
or (n13719,s0n13719,s1n13719);
not(notn13719,n10017);
and (s0n13719,notn13719,n13720);
and (s1n13719,n10017,n13722);
wire s0n13720,s1n13720,notn13720;
or (n13720,s0n13720,s1n13720);
not(notn13720,n10000);
and (s0n13720,notn13720,1'b0);
and (s1n13720,n10000,n13721);
or (n13722,1'b0,n13723,n13725,n13727);
and (n13723,n13724,n10009);
and (n13725,n13726,n10012);
and (n13727,n13721,n10014);
nand (n13728,n13729,n13676);
or (n13729,n13730,n13675);
not (n13730,n13718);
or (n13731,n13732,n13733,n13734);
and (n13732,n13656,n13672);
and (n13733,n13672,n13682);
and (n13734,n13656,n13682);
xor (n13735,n13736,n13747);
xor (n13736,n13737,n13742);
wire s0n13737,s1n13737,notn13737;
or (n13737,s0n13737,s1n13737);
not(notn13737,n1039);
and (s0n13737,notn13737,1'b0);
and (s1n13737,n1039,n13738);
and (n13738,n13739,n1042);
wire s0n13739,s1n13739,notn13739;
or (n13739,s0n13739,s1n13739);
not(notn13739,n650);
and (s0n13739,notn13739,1'b0);
and (s1n13739,n650,n13740);
and (n13740,n13741,n10091);
wire s0n13742,s1n13742,notn13742;
or (n13742,s0n13742,s1n13742);
not(notn13742,n1039);
and (s0n13742,notn13742,1'b0);
and (s1n13742,n1039,n13743);
and (n13743,n13744,n1042);
wire s0n13744,s1n13744,notn13744;
or (n13744,s0n13744,s1n13744);
not(notn13744,n650);
and (s0n13744,notn13744,1'b0);
and (s1n13744,n650,n13745);
and (n13745,n13746,n10091);
or (n13747,n13748,n13749);
and (n13748,n13687,n13698);
and (n13749,n13688,n13693);
or (n13750,n13751,n13752,n13753);
and (n13751,n13653,n13686);
and (n13752,n13686,n13701);
and (n13753,n13653,n13701);
and (n13754,n13651,n13705);
wire s0n13755,s1n13755,notn13755;
or (n13755,s0n13755,s1n13755);
not(notn13755,n13539);
and (s0n13755,notn13755,n13756);
and (s1n13755,n13539,n13805);
xor (n13756,n13757,n13804);
xor (n13757,n13758,n13800);
xor (n13758,n13759,n13785);
wire s0n13759,s1n13759,notn13759;
or (n13759,s0n13759,s1n13759);
not(notn13759,n12915);
and (s0n13759,notn13759,n13760);
and (s1n13759,n12915,1'b0);
xor (n13760,n13761,n13781);
xor (n13761,n13762,n13778);
nand (n13762,n13763,n13766);
or (n13763,n13764,n13465);
not (n13764,n13765);
nor (n13766,n13767,n13769);
and (n13767,n13441,n13768);
wire s0n13769,s1n13769,notn13769;
or (n13769,s0n13769,s1n13769);
not(notn13769,n10017);
and (s0n13769,notn13769,n13770);
and (s1n13769,n10017,n13772);
wire s0n13770,s1n13770,notn13770;
or (n13770,s0n13770,s1n13770);
not(notn13770,n10000);
and (s0n13770,notn13770,1'b0);
and (s1n13770,n10000,n13771);
or (n13772,1'b0,n13773,n13775,n13777);
and (n13773,n13774,n10009);
and (n13775,n13776,n10012);
and (n13777,n13771,n10014);
nand (n13778,n13779,n13676);
or (n13779,n13780,n13675);
not (n13780,n13768);
or (n13781,n13782,n13783,n13784);
and (n13782,n13712,n13728);
and (n13783,n13728,n13731);
and (n13784,n13712,n13731);
xor (n13785,n13786,n13797);
xor (n13786,n13787,n13792);
wire s0n13787,s1n13787,notn13787;
or (n13787,s0n13787,s1n13787);
not(notn13787,n1039);
and (s0n13787,notn13787,1'b0);
and (s1n13787,n1039,n13788);
and (n13788,n13789,n1042);
wire s0n13789,s1n13789,notn13789;
or (n13789,s0n13789,s1n13789);
not(notn13789,n650);
and (s0n13789,notn13789,1'b0);
and (s1n13789,n650,n13790);
and (n13790,n13791,n10091);
wire s0n13792,s1n13792,notn13792;
or (n13792,s0n13792,s1n13792);
not(notn13792,n1039);
and (s0n13792,notn13792,1'b0);
and (s1n13792,n1039,n13793);
and (n13793,n13794,n1042);
wire s0n13794,s1n13794,notn13794;
or (n13794,s0n13794,s1n13794);
not(notn13794,n650);
and (s0n13794,notn13794,1'b0);
and (s1n13794,n650,n13795);
and (n13795,n13796,n10091);
or (n13797,n13798,n13799);
and (n13798,n13736,n13747);
and (n13799,n13737,n13742);
or (n13800,n13801,n13802,n13803);
and (n13801,n13709,n13735);
and (n13802,n13735,n13750);
and (n13803,n13709,n13750);
and (n13804,n13707,n13754);
xor (n13805,n13806,n13853);
xor (n13806,n13807,n13849);
xor (n13807,n13808,n13834);
wire s0n13808,s1n13808,notn13808;
or (n13808,s0n13808,s1n13808);
not(notn13808,n12915);
and (s0n13808,notn13808,n13809);
and (s1n13808,n12915,1'b0);
xor (n13809,n13810,n13830);
xor (n13810,n13811,n13827);
nand (n13811,n13812,n13815);
or (n13812,n13813,n13465);
not (n13813,n13814);
nor (n13815,n13816,n13818);
and (n13816,n13441,n13817);
wire s0n13818,s1n13818,notn13818;
or (n13818,s0n13818,s1n13818);
not(notn13818,n10017);
and (s0n13818,notn13818,n13819);
and (s1n13818,n10017,n13821);
wire s0n13819,s1n13819,notn13819;
or (n13819,s0n13819,s1n13819);
not(notn13819,n10000);
and (s0n13819,notn13819,1'b0);
and (s1n13819,n10000,n13820);
or (n13821,1'b0,n13822,n13824,n13826);
and (n13822,n13823,n10009);
and (n13824,n13825,n10012);
and (n13826,n13820,n10014);
nand (n13827,n13828,n13676);
or (n13828,n13829,n13675);
not (n13829,n13817);
or (n13830,n13831,n13832,n13833);
and (n13831,n13762,n13778);
and (n13832,n13778,n13781);
and (n13833,n13762,n13781);
xor (n13834,n13835,n13846);
xor (n13835,n13836,n13841);
wire s0n13836,s1n13836,notn13836;
or (n13836,s0n13836,s1n13836);
not(notn13836,n1039);
and (s0n13836,notn13836,1'b0);
and (s1n13836,n1039,n13837);
and (n13837,n13838,n1042);
wire s0n13838,s1n13838,notn13838;
or (n13838,s0n13838,s1n13838);
not(notn13838,n650);
and (s0n13838,notn13838,1'b0);
and (s1n13838,n650,n13839);
and (n13839,n13840,n10091);
wire s0n13841,s1n13841,notn13841;
or (n13841,s0n13841,s1n13841);
not(notn13841,n1039);
and (s0n13841,notn13841,1'b0);
and (s1n13841,n1039,n13842);
and (n13842,n13843,n1042);
wire s0n13843,s1n13843,notn13843;
or (n13843,s0n13843,s1n13843);
not(notn13843,n650);
and (s0n13843,notn13843,1'b0);
and (s1n13843,n650,n13844);
and (n13844,n13845,n10091);
or (n13846,n13847,n13848);
and (n13847,n13786,n13797);
and (n13848,n13787,n13792);
or (n13849,n13850,n13851,n13852);
and (n13850,n13759,n13785);
and (n13851,n13785,n13800);
and (n13852,n13759,n13800);
and (n13853,n13757,n13804);
wire s0n13854,s1n13854,notn13854;
or (n13854,s0n13854,s1n13854);
not(notn13854,n1039);
and (s0n13854,notn13854,n13400);
and (s1n13854,n1039,n13855);
or (n13855,n13403,n13856,1'b0);
and (n13856,n13857,n1042);
and (n13857,n650,n10073);
wire s0n13858,s1n13858,notn13858;
or (n13858,s0n13858,s1n13858);
not(notn13858,n13934);
and (s0n13858,notn13858,n13859);
and (s1n13858,n13934,1'b0);
wire s0n13859,s1n13859,notn13859;
or (n13859,s0n13859,s1n13859);
not(notn13859,n13860);
and (s0n13859,notn13859,1'b1);
and (s1n13859,n13860,n9980);
nor (n13860,n13861,n13919,n13924,n13928,n13930,n13932,n13933,n13934);
wire s0n13861,s1n13861,notn13861;
or (n13861,s0n13861,s1n13861);
not(notn13861,n13854);
and (s0n13861,notn13861,n13862);
and (s1n13861,n13854,n13865);
wire s0n13862,s1n13862,notn13862;
or (n13862,s0n13862,s1n13862);
not(notn13862,n13645);
and (s0n13862,notn13862,n13863);
and (s1n13862,n13645,n13864);
wire s0n13863,s1n13863,notn13863;
or (n13863,s0n13863,s1n13863);
not(notn13863,n13539);
and (s0n13863,notn13863,n13455);
and (s1n13863,n13539,n13541);
wire s0n13864,s1n13864,notn13864;
or (n13864,s0n13864,s1n13864);
not(notn13864,n13539);
and (s0n13864,notn13864,n13593);
and (s1n13864,n13539,n13650);
wire s0n13865,s1n13865,notn13865;
or (n13865,s0n13865,s1n13865);
not(notn13865,n13645);
and (s0n13865,notn13865,n13866);
and (s1n13865,n13645,n13867);
wire s0n13866,s1n13866,notn13866;
or (n13866,s0n13866,s1n13866);
not(notn13866,n13539);
and (s0n13866,notn13866,n13706);
and (s1n13866,n13539,n13756);
wire s0n13867,s1n13867,notn13867;
or (n13867,s0n13867,s1n13867);
not(notn13867,n13539);
and (s0n13867,notn13867,n13805);
and (s1n13867,n13539,n13868);
xor (n13868,n13869,n13918);
xor (n13869,n13870,n13914);
xor (n13870,n13871,n13897);
wire s0n13871,s1n13871,notn13871;
or (n13871,s0n13871,s1n13871);
not(notn13871,n12915);
and (s0n13871,notn13871,n13872);
and (s1n13871,n12915,1'b0);
xor (n13872,n13873,n13893);
xor (n13873,n13874,n13890);
nand (n13874,n13875,n13878);
or (n13875,n13876,n13465);
not (n13876,n13877);
nor (n13878,n13879,n13881);
and (n13879,n13441,n13880);
wire s0n13881,s1n13881,notn13881;
or (n13881,s0n13881,s1n13881);
not(notn13881,n10017);
and (s0n13881,notn13881,n13882);
and (s1n13881,n10017,n13884);
wire s0n13882,s1n13882,notn13882;
or (n13882,s0n13882,s1n13882);
not(notn13882,n10000);
and (s0n13882,notn13882,1'b0);
and (s1n13882,n10000,n13883);
or (n13884,1'b0,n13885,n13887,n13889);
and (n13885,n13886,n10009);
and (n13887,n13888,n10012);
and (n13889,n13883,n10014);
nand (n13890,n13891,n13676);
or (n13891,n13892,n13675);
not (n13892,n13880);
or (n13893,n13894,n13895,n13896);
and (n13894,n13811,n13827);
and (n13895,n13827,n13830);
and (n13896,n13811,n13830);
xor (n13897,n13898,n13910);
not (n13898,n13899);
xor (n13899,n13900,n13905);
wire s0n13900,s1n13900,notn13900;
or (n13900,s0n13900,s1n13900);
not(notn13900,n1039);
and (s0n13900,notn13900,1'b0);
and (s1n13900,n1039,n13901);
and (n13901,n13902,n1042);
wire s0n13902,s1n13902,notn13902;
or (n13902,s0n13902,s1n13902);
not(notn13902,n650);
and (s0n13902,notn13902,1'b0);
and (s1n13902,n650,n13903);
and (n13903,n13904,n10091);
wire s0n13905,s1n13905,notn13905;
or (n13905,s0n13905,s1n13905);
not(notn13905,n1039);
and (s0n13905,notn13905,1'b0);
and (s1n13905,n1039,n13906);
and (n13906,n13907,n1042);
wire s0n13907,s1n13907,notn13907;
or (n13907,s0n13907,s1n13907);
not(notn13907,n650);
and (s0n13907,notn13907,1'b0);
and (s1n13907,n650,n13908);
and (n13908,n13909,n10091);
nor (n13910,n13911,n13913);
and (n13911,n13846,n13912);
or (n13912,n13841,n13836);
and (n13913,n13836,n13841);
or (n13914,n13915,n13916,n13917);
and (n13915,n13808,n13834);
and (n13916,n13834,n13849);
and (n13917,n13808,n13849);
and (n13918,n13806,n13853);
wire s0n13919,s1n13919,notn13919;
or (n13919,s0n13919,s1n13919);
not(notn13919,n13854);
and (s0n13919,notn13919,n13920);
and (s1n13919,n13854,n13921);
wire s0n13920,s1n13920,notn13920;
or (n13920,s0n13920,s1n13920);
not(notn13920,n13645);
and (s0n13920,notn13920,n13540);
and (s1n13920,n13645,n13649);
wire s0n13921,s1n13921,notn13921;
or (n13921,s0n13921,s1n13921);
not(notn13921,n13645);
and (s0n13921,notn13921,n13755);
and (s1n13921,n13645,n13922);
wire s0n13922,s1n13922,notn13922;
or (n13922,s0n13922,s1n13922);
not(notn13922,n13539);
and (s0n13922,notn13922,n13868);
and (s1n13922,n13539,n13923);
and (n13923,n13869,n13918);
wire s0n13924,s1n13924,notn13924;
or (n13924,s0n13924,s1n13924);
not(notn13924,n13854);
and (s0n13924,notn13924,n13925);
and (s1n13924,n13854,n13926);
wire s0n13925,s1n13925,notn13925;
or (n13925,s0n13925,s1n13925);
not(notn13925,n13645);
and (s0n13925,notn13925,n13864);
and (s1n13925,n13645,n13866);
wire s0n13926,s1n13926,notn13926;
or (n13926,s0n13926,s1n13926);
not(notn13926,n13645);
and (s0n13926,notn13926,n13867);
and (s1n13926,n13645,n13927);
wire s0n13927,s1n13927,notn13927;
or (n13927,s0n13927,s1n13927);
not(notn13927,n13539);
and (s0n13927,notn13927,n13923);
and (s1n13927,n13539,1'b0);
wire s0n13928,s1n13928,notn13928;
or (n13928,s0n13928,s1n13928);
not(notn13928,n13854);
and (s0n13928,notn13928,n13648);
and (s1n13928,n13854,n13929);
wire s0n13929,s1n13929,notn13929;
or (n13929,s0n13929,s1n13929);
not(notn13929,n13645);
and (s0n13929,notn13929,n13922);
and (s1n13929,n13645,1'b0);
wire s0n13930,s1n13930,notn13930;
or (n13930,s0n13930,s1n13930);
not(notn13930,n13854);
and (s0n13930,notn13930,n13865);
and (s1n13930,n13854,n13931);
wire s0n13931,s1n13931,notn13931;
or (n13931,s0n13931,s1n13931);
not(notn13931,n13645);
and (s0n13931,notn13931,n13927);
and (s1n13931,n13645,1'b0);
wire s0n13932,s1n13932,notn13932;
or (n13932,s0n13932,s1n13932);
not(notn13932,n13854);
and (s0n13932,notn13932,n13921);
and (s1n13932,n13854,1'b0);
wire s0n13933,s1n13933,notn13933;
or (n13933,s0n13933,s1n13933);
not(notn13933,n13854);
and (s0n13933,notn13933,n13926);
and (s1n13933,n13854,1'b0);
wire s0n13934,s1n13934,notn13934;
or (n13934,s0n13934,s1n13934);
not(notn13934,n13854);
and (s0n13934,notn13934,n13929);
and (s1n13934,n13854,1'b0);
wire s0n13935,s1n13935,notn13935;
or (n13935,s0n13935,s1n13935);
not(notn13935,n1057);
and (s0n13935,notn13935,n13936);
and (s1n13935,n1057,n14701);
wire s0n13936,s1n13936,notn13936;
or (n13936,s0n13936,s1n13936);
not(notn13936,n805);
and (s0n13936,notn13936,n13937);
and (s1n13936,n805,n14695);
wire s0n13937,s1n13937,notn13937;
or (n13937,s0n13937,s1n13937);
not(notn13937,n1066);
and (s0n13937,notn13937,n1067);
and (s1n13937,n1066,n13938);
wire s0n13938,s1n13938,notn13938;
or (n13938,s0n13938,s1n13938);
not(notn13938,n31);
and (s0n13938,notn13938,n13939);
and (s1n13938,n31,n14691);
or (n13939,n13940,n14690);
and (n13940,n13941,n817);
wire s0n13941,s1n13941,notn13941;
or (n13941,s0n13941,s1n13941);
not(notn13941,n805);
and (s0n13941,notn13941,n13942);
and (s1n13941,n805,n14682);
wire s0n13942,s1n13942,notn13942;
or (n13942,s0n13942,s1n13942);
not(notn13942,n8008);
and (s0n13942,notn13942,n13943);
and (s1n13942,n8008,n7998);
xor (n13943,n13944,n14659);
xor (n13944,n13945,n14560);
xor (n13945,n13946,n14263);
xor (n13946,n13947,n14170);
xor (n13947,n13948,n14055);
xor (n13948,n9962,n13949);
or (n13949,n13950,n13988,n14054);
and (n13950,n13951,n13952);
xor (n13951,n9349,n9354);
and (n13952,n8129,n13953);
or (n13953,n13954,n13955,n13987);
and (n13954,n9107,n9099);
and (n13955,n9099,n13956);
or (n13956,n13957,n13958,n13986);
and (n13957,n9060,n9300);
and (n13958,n9300,n13959);
or (n13959,n13960,n13961,n13985);
and (n13960,n9149,n9274);
and (n13961,n9274,n13962);
or (n13962,n13963,n13964,n13984);
and (n13963,n9461,n9463);
and (n13964,n9463,n13965);
or (n13965,n13966,n13967,n13983);
and (n13966,n9521,n9542);
and (n13967,n9542,n13968);
or (n13968,n13969,n13970,n13982);
and (n13969,n9605,n9703);
and (n13970,n9703,n13971);
or (n13971,n13972,n13973,n13981);
and (n13972,n9726,n9734);
and (n13973,n9734,n13974);
or (n13974,n13975,n13976,n13978);
and (n13975,n9766,n9829);
and (n13976,n9829,n13977);
or (n13977,n13978,n13979,n13980);
and (n13978,n9806,n9862);
and (n13979,n9862,n13980);
and (n13980,n9822,n9878);
and (n13981,n9726,n13974);
and (n13982,n9605,n13971);
and (n13983,n9521,n13968);
and (n13984,n9461,n13965);
and (n13985,n9149,n13962);
and (n13986,n9060,n13959);
and (n13987,n9107,n13956);
and (n13988,n13952,n13989);
or (n13989,n13990,n13993,n14053);
and (n13990,n13991,n13992);
xor (n13991,n9068,n8505);
xor (n13992,n8129,n13953);
and (n13993,n13992,n13994);
or (n13994,n13995,n13999,n14052);
and (n13995,n13996,n13997);
xor (n13996,n9323,n9094);
xor (n13997,n13998,n13956);
xor (n13998,n9107,n9099);
and (n13999,n13997,n14000);
or (n14000,n14001,n14005,n14051);
and (n14001,n14002,n14003);
xor (n14002,n8986,n8930);
xor (n14003,n14004,n13959);
xor (n14004,n9060,n9300);
and (n14005,n14003,n14006);
or (n14006,n14007,n14011,n14050);
and (n14007,n14008,n14009);
xor (n14008,n9388,n9120);
xor (n14009,n14010,n13962);
xor (n14010,n9149,n9274);
and (n14011,n14009,n14012);
or (n14012,n14013,n14017,n14049);
and (n14013,n14014,n14015);
xor (n14014,n9145,n9270);
xor (n14015,n14016,n13965);
xor (n14016,n9461,n9463);
and (n14017,n14015,n14018);
or (n14018,n14019,n14023,n14048);
and (n14019,n14020,n14021);
xor (n14020,n9443,n9439);
xor (n14021,n14022,n13968);
xor (n14022,n9521,n9542);
and (n14023,n14021,n14024);
or (n14024,n14025,n14029,n14047);
and (n14025,n14026,n14027);
xor (n14026,n9702,n9539);
xor (n14027,n14028,n13971);
xor (n14028,n9605,n9703);
and (n14029,n14027,n14030);
or (n14030,n14031,n14035,n14046);
and (n14031,n14032,n14033);
xor (n14032,n9602,n9584);
xor (n14033,n14034,n13974);
xor (n14034,n9726,n9734);
and (n14035,n14033,n14036);
or (n14036,n14037,n14041,n14045);
and (n14037,n14038,n14039);
xor (n14038,n9599,n9716);
xor (n14039,n14040,n13977);
xor (n14040,n9766,n9829);
and (n14041,n14039,n14042);
and (n14042,n9666,n14043);
xor (n14043,n14044,n13980);
xor (n14044,n9806,n9862);
and (n14045,n14038,n14042);
and (n14046,n14032,n14036);
and (n14047,n14026,n14030);
and (n14048,n14020,n14024);
and (n14049,n14014,n14018);
and (n14050,n14008,n14012);
and (n14051,n14002,n14006);
and (n14052,n13996,n14000);
and (n14053,n13991,n13994);
and (n14054,n13951,n13989);
xor (n14055,n9963,n14056);
or (n14056,n14057,n14104,n14169);
and (n14057,n9346,n14058);
and (n14058,n8893,n14059);
or (n14059,n14060,n14062,n14103);
and (n14060,n9314,n14061);
wire s0n14061,s1n14061,notn14061;
or (n14061,s0n14061,s1n14061);
not(notn14061,n655);
and (s0n14061,notn14061,1'b0);
and (s1n14061,n655,n8894);
and (n14062,n14061,n14063);
or (n14063,n14064,n14066,n14102);
and (n14064,n9282,n14065);
wire s0n14065,s1n14065,notn14065;
or (n14065,s0n14065,s1n14065);
not(notn14065,n655);
and (s0n14065,notn14065,1'b0);
and (s1n14065,n655,n8905);
and (n14066,n14065,n14067);
or (n14067,n14068,n14070,n14101);
and (n14068,n9090,n14069);
wire s0n14069,s1n14069,notn14069;
or (n14069,s0n14069,s1n14069);
not(notn14069,n655);
and (s0n14069,notn14069,1'b0);
and (s1n14069,n655,n8747);
and (n14070,n14069,n14071);
or (n14071,n14072,n14074,n14100);
and (n14072,n9196,n14073);
wire s0n14073,s1n14073,notn14073;
or (n14073,s0n14073,s1n14073);
not(notn14073,n655);
and (s0n14073,notn14073,1'b0);
and (s1n14073,n655,n8731);
and (n14074,n14073,n14075);
or (n14075,n14076,n14078,n14099);
and (n14076,n9165,n14077);
wire s0n14077,s1n14077,notn14077;
or (n14077,s0n14077,s1n14077);
not(notn14077,n655);
and (s0n14077,notn14077,1'b0);
and (s1n14077,n655,n8519);
and (n14078,n14077,n14079);
or (n14079,n14080,n14082,n14098);
and (n14080,n9268,n14081);
wire s0n14081,s1n14081,notn14081;
or (n14081,s0n14081,s1n14081);
not(notn14081,n655);
and (s0n14081,notn14081,1'b0);
and (s1n14081,n655,n9031);
and (n14082,n14081,n14083);
or (n14083,n14084,n14086,n14097);
and (n14084,n9436,n14085);
wire s0n14085,s1n14085,notn14085;
or (n14085,s0n14085,s1n14085);
not(notn14085,n655);
and (s0n14085,notn14085,1'b0);
and (s1n14085,n655,n9134);
and (n14086,n14085,n14087);
or (n14087,n14088,n14090,n14092);
and (n14088,n9644,n14089);
wire s0n14089,s1n14089,notn14089;
or (n14089,s0n14089,s1n14089);
not(notn14089,n655);
and (s0n14089,notn14089,1'b0);
and (s1n14089,n655,n9140);
and (n14090,n14089,n14091);
or (n14091,n14092,n14094,n14095);
and (n14092,n9721,n14093);
wire s0n14093,s1n14093,notn14093;
or (n14093,s0n14093,s1n14093);
not(notn14093,n655);
and (s0n14093,notn14093,1'b0);
and (s1n14093,n655,n9267);
and (n14094,n14093,n14095);
and (n14095,n9824,n14096);
wire s0n14096,s1n14096,notn14096;
or (n14096,s0n14096,s1n14096);
not(notn14096,n655);
and (s0n14096,notn14096,1'b0);
and (s1n14096,n655,n9234);
and (n14097,n9436,n14087);
and (n14098,n9268,n14083);
and (n14099,n9165,n14079);
and (n14100,n9196,n14075);
and (n14101,n9090,n14071);
and (n14102,n9282,n14067);
and (n14103,n9314,n14063);
and (n14104,n14058,n14105);
or (n14105,n14106,n14109,n14168);
and (n14106,n14107,n14108);
xor (n14107,n8903,n8904);
xor (n14108,n8893,n14059);
and (n14109,n14108,n14110);
or (n14110,n14111,n14115,n14167);
and (n14111,n14112,n14113);
xor (n14112,n9317,n8746);
xor (n14113,n14114,n14063);
xor (n14114,n9314,n14061);
and (n14115,n14113,n14116);
or (n14116,n14117,n14121,n14166);
and (n14117,n14118,n14119);
xor (n14118,n8518,n8730);
xor (n14119,n14120,n14067);
xor (n14120,n9282,n14065);
and (n14121,n14119,n14122);
or (n14122,n14123,n14126,n14165);
and (n14123,n9087,n14124);
xor (n14124,n14125,n14071);
xor (n14125,n9090,n14069);
and (n14126,n14124,n14127);
or (n14127,n14128,n14132,n14164);
and (n14128,n14129,n14130);
xor (n14129,n9133,n9030);
xor (n14130,n14131,n14075);
xor (n14131,n9196,n14073);
and (n14132,n14130,n14133);
or (n14133,n14134,n14138,n14163);
and (n14134,n14135,n14136);
xor (n14135,n9139,n9215);
xor (n14136,n14137,n14079);
xor (n14137,n9165,n14077);
and (n14138,n14136,n14139);
or (n14139,n14140,n14144,n14162);
and (n14140,n14141,n14142);
xor (n14141,n9266,n9183);
xor (n14142,n14143,n14083);
xor (n14143,n9268,n14081);
and (n14144,n14142,n14145);
or (n14145,n14146,n14150,n14161);
and (n14146,n14147,n14148);
xor (n14147,n9233,n9433);
xor (n14148,n14149,n14087);
xor (n14149,n9436,n14085);
and (n14150,n14148,n14151);
or (n14151,n14152,n14156,n14160);
and (n14152,n14153,n14154);
xor (n14153,n9581,n9601);
xor (n14154,n14155,n14091);
xor (n14155,n9644,n14089);
and (n14156,n14154,n14157);
and (n14157,n9722,n14158);
xor (n14158,n14159,n14095);
xor (n14159,n9721,n14093);
and (n14160,n14153,n14157);
and (n14161,n14147,n14151);
and (n14162,n14141,n14145);
and (n14163,n14135,n14139);
and (n14164,n14129,n14133);
and (n14165,n9087,n14127);
and (n14166,n14118,n14122);
and (n14167,n14112,n14116);
and (n14168,n14107,n14110);
and (n14169,n9346,n14105);
or (n14170,n14171,n14176,n14262);
and (n14171,n14172,n14174);
xor (n14172,n14173,n13989);
xor (n14173,n13951,n13952);
xor (n14174,n14175,n14105);
xor (n14175,n9346,n14058);
and (n14176,n14174,n14177);
or (n14177,n14178,n14183,n14261);
and (n14178,n14179,n14181);
xor (n14179,n14180,n13994);
xor (n14180,n13991,n13992);
xor (n14181,n14182,n14110);
xor (n14182,n14107,n14108);
and (n14183,n14181,n14184);
or (n14184,n14185,n14190,n14260);
and (n14185,n14186,n14188);
xor (n14186,n14187,n14000);
xor (n14187,n13996,n13997);
xor (n14188,n14189,n14116);
xor (n14189,n14112,n14113);
and (n14190,n14188,n14191);
or (n14191,n14192,n14197,n14259);
and (n14192,n14193,n14195);
xor (n14193,n14194,n14006);
xor (n14194,n14002,n14003);
xor (n14195,n14196,n14122);
xor (n14196,n14118,n14119);
and (n14197,n14195,n14198);
or (n14198,n14199,n14204,n14258);
and (n14199,n14200,n14202);
xor (n14200,n14201,n14012);
xor (n14201,n14008,n14009);
xor (n14202,n14203,n14127);
xor (n14203,n9087,n14124);
and (n14204,n14202,n14205);
or (n14205,n14206,n14211,n14257);
and (n14206,n14207,n14209);
xor (n14207,n14208,n14018);
xor (n14208,n14014,n14015);
xor (n14209,n14210,n14133);
xor (n14210,n14129,n14130);
and (n14211,n14209,n14212);
or (n14212,n14213,n14218,n14256);
and (n14213,n14214,n14216);
xor (n14214,n14215,n14024);
xor (n14215,n14020,n14021);
xor (n14216,n14217,n14139);
xor (n14217,n14135,n14136);
and (n14218,n14216,n14219);
or (n14219,n14220,n14225,n14255);
and (n14220,n14221,n14223);
xor (n14221,n14222,n14030);
xor (n14222,n14026,n14027);
xor (n14223,n14224,n14145);
xor (n14224,n14141,n14142);
and (n14225,n14223,n14226);
or (n14226,n14227,n14232,n14254);
and (n14227,n14228,n14230);
xor (n14228,n14229,n14036);
xor (n14229,n14032,n14033);
xor (n14230,n14231,n14151);
xor (n14231,n14147,n14148);
and (n14232,n14230,n14233);
or (n14233,n14234,n14239,n14253);
and (n14234,n14235,n14237);
xor (n14235,n14236,n14042);
xor (n14236,n14038,n14039);
xor (n14237,n14238,n14157);
xor (n14238,n14153,n14154);
and (n14239,n14237,n14240);
or (n14240,n14241,n14244,n14252);
and (n14241,n14242,n14243);
xor (n14242,n9666,n14043);
xor (n14243,n9722,n14158);
and (n14244,n14243,n14245);
or (n14245,n14246,n14249,n14251);
and (n14246,n14247,n14248);
xor (n14247,n9822,n9878);
xor (n14248,n9824,n14096);
and (n14249,n14248,n14250);
and (n14250,n9912,n9801);
and (n14251,n14247,n14250);
and (n14252,n14242,n14245);
and (n14253,n14235,n14240);
and (n14254,n14228,n14233);
and (n14255,n14221,n14226);
and (n14256,n14214,n14219);
and (n14257,n14207,n14212);
and (n14258,n14200,n14205);
and (n14259,n14193,n14198);
and (n14260,n14186,n14191);
and (n14261,n14179,n14184);
and (n14262,n14172,n14177);
xor (n14263,n14264,n14467);
xor (n14264,n14265,n14361);
or (n14265,n14266,n14303,n14360);
and (n14266,n9352,n14267);
and (n14267,n9320,n14268);
or (n14268,n14269,n14270,n14302);
and (n14269,n9318,n9100);
and (n14270,n9100,n14271);
or (n14271,n14272,n14273,n14301);
and (n14272,n8924,n9279);
and (n14273,n9279,n14274);
or (n14274,n14275,n14276,n14300);
and (n14275,n9127,n9122);
and (n14276,n9122,n14277);
or (n14277,n14278,n14279,n14299);
and (n14278,n9462,n9450);
and (n14279,n9450,n14280);
or (n14280,n14281,n14282,n14298);
and (n14281,n9522,n9569);
and (n14282,n9569,n14283);
or (n14283,n14284,n14285,n14297);
and (n14284,n9672,n9704);
and (n14285,n9704,n14286);
or (n14286,n14287,n14288,n14296);
and (n14287,n9732,n9768);
and (n14288,n9768,n14289);
or (n14289,n14290,n14291,n14293);
and (n14290,n9765,n9828);
and (n14291,n9828,n14292);
or (n14292,n14293,n14294,n14295);
and (n14293,n9818,n9860);
and (n14294,n9860,n14295);
and (n14295,n9803,n9880);
and (n14296,n9732,n14289);
and (n14297,n9672,n14286);
and (n14298,n9522,n14283);
and (n14299,n9462,n14280);
and (n14300,n9127,n14277);
and (n14301,n8924,n14274);
and (n14302,n9318,n14271);
and (n14303,n14267,n14304);
or (n14304,n14305,n14307,n14359);
and (n14305,n8323,n14306);
xor (n14306,n9320,n14268);
and (n14307,n14306,n14308);
or (n14308,n14309,n14312,n14358);
and (n14309,n9093,n14310);
xor (n14310,n14311,n14271);
xor (n14311,n9318,n9100);
and (n14312,n14310,n14313);
or (n14313,n14314,n14317,n14357);
and (n14314,n8927,n14315);
xor (n14315,n14316,n14274);
xor (n14316,n8924,n9279);
and (n14317,n14315,n14318);
or (n14318,n14319,n14322,n14356);
and (n14319,n9390,n14320);
xor (n14320,n14321,n14277);
xor (n14321,n9127,n9122);
and (n14322,n14320,n14323);
or (n14323,n14324,n14327,n14355);
and (n14324,n9187,n14325);
xor (n14325,n14326,n14280);
xor (n14326,n9462,n9450);
and (n14327,n14325,n14328);
or (n14328,n14329,n14332,n14354);
and (n14329,n9447,n14330);
xor (n14330,n14331,n14283);
xor (n14331,n9522,n9569);
and (n14332,n14330,n14333);
or (n14333,n14334,n14337,n14353);
and (n14334,n9536,n14335);
xor (n14335,n14336,n14286);
xor (n14336,n9672,n9704);
and (n14337,n14335,n14338);
or (n14338,n14339,n14342,n14352);
and (n14339,n9576,n14340);
xor (n14340,n14341,n14289);
xor (n14341,n9732,n9768);
and (n14342,n14340,n14343);
or (n14343,n14344,n14347,n14351);
and (n14344,n9668,n14345);
xor (n14345,n14346,n14292);
xor (n14346,n9765,n9828);
and (n14347,n14345,n14348);
and (n14348,n9508,n14349);
xor (n14349,n14350,n14295);
xor (n14350,n9818,n9860);
and (n14351,n9668,n14348);
and (n14352,n9576,n14343);
and (n14353,n9536,n14338);
and (n14354,n9447,n14333);
and (n14355,n9187,n14328);
and (n14356,n9390,n14323);
and (n14357,n8927,n14318);
and (n14358,n9093,n14313);
and (n14359,n8323,n14308);
and (n14360,n9352,n14304);
or (n14361,n14362,n14409,n14466);
and (n14362,n9353,n14363);
and (n14363,n8907,n14364);
or (n14364,n14365,n14367,n14408);
and (n14365,n9327,n14366);
wire s0n14366,s1n14366,notn14366;
or (n14366,s0n14366,s1n14366);
not(notn14366,n655);
and (s0n14366,notn14366,1'b0);
and (s1n14366,n655,n8908);
and (n14367,n14366,n14368);
or (n14368,n14369,n14371,n14407);
and (n14369,n9091,n14370);
wire s0n14370,s1n14370,notn14370;
or (n14370,s0n14370,s1n14370);
not(notn14370,n655);
and (s0n14370,notn14370,1'b0);
and (s1n14370,n655,n9077);
and (n14371,n14370,n14372);
or (n14372,n14373,n14375,n14406);
and (n14373,n9383,n14374);
wire s0n14374,s1n14374,notn14374;
or (n14374,s0n14374,s1n14374);
not(notn14374,n655);
and (s0n14374,notn14374,1'b0);
and (s1n14374,n655,n8759);
and (n14375,n14374,n14376);
or (n14376,n14377,n14379,n14405);
and (n14377,n9217,n14378);
wire s0n14378,s1n14378,notn14378;
or (n14378,s0n14378,s1n14378);
not(notn14378,n655);
and (s0n14378,notn14378,1'b0);
and (s1n14378,n655,n9298);
and (n14379,n14378,n14380);
or (n14380,n14381,n14383,n14404);
and (n14381,n9185,n14382);
wire s0n14382,s1n14382,notn14382;
or (n14382,s0n14382,s1n14382);
not(notn14382,n655);
and (s0n14382,notn14382,1'b0);
and (s1n14382,n655,n8993);
and (n14383,n14382,n14384);
or (n14384,n14385,n14387,n14403);
and (n14385,n9265,n14386);
wire s0n14386,s1n14386,notn14386;
or (n14386,s0n14386,s1n14386);
not(notn14386,n655);
and (s0n14386,notn14386,1'b0);
and (s1n14386,n655,n9056);
and (n14387,n14386,n14388);
or (n14388,n14389,n14391,n14402);
and (n14389,n9519,n14390);
wire s0n14390,s1n14390,notn14390;
or (n14390,s0n14390,s1n14390);
not(notn14390,n655);
and (s0n14390,notn14390,1'b0);
and (s1n14390,n655,n9143);
and (n14391,n14390,n14392);
or (n14392,n14393,n14395,n14397);
and (n14393,n9583,n14394);
wire s0n14394,s1n14394,notn14394;
or (n14394,s0n14394,s1n14394);
not(notn14394,n655);
and (s0n14394,notn14394,1'b0);
and (s1n14394,n655,n9260);
and (n14395,n14394,n14396);
or (n14396,n14397,n14399,n14400);
and (n14397,n9626,n14398);
wire s0n14398,s1n14398,notn14398;
or (n14398,s0n14398,s1n14398);
not(notn14398,n655);
and (s0n14398,notn14398,1'b0);
and (s1n14398,n655,n9435);
and (n14399,n14398,n14400);
and (n14400,n9657,n14401);
wire s0n14401,s1n14401,notn14401;
or (n14401,s0n14401,s1n14401);
not(notn14401,n655);
and (s0n14401,notn14401,1'b0);
and (s1n14401,n655,n9505);
and (n14402,n9519,n14392);
and (n14403,n9265,n14388);
and (n14404,n9185,n14384);
and (n14405,n9217,n14380);
and (n14406,n9383,n14376);
and (n14407,n9091,n14372);
and (n14408,n9327,n14368);
and (n14409,n14363,n14410);
or (n14410,n14411,n14413,n14465);
and (n14411,n9076,n14412);
xor (n14412,n8907,n14364);
and (n14413,n14412,n14414);
or (n14414,n14415,n14418,n14464);
and (n14415,n8758,n14416);
xor (n14416,n14417,n14368);
xor (n14417,n9327,n14366);
and (n14418,n14416,n14419);
or (n14419,n14420,n14423,n14463);
and (n14420,n9297,n14421);
xor (n14421,n14422,n14372);
xor (n14422,n9091,n14370);
and (n14423,n14421,n14424);
or (n14424,n14425,n14428,n14462);
and (n14425,n8992,n14426);
xor (n14426,n14427,n14376);
xor (n14427,n9383,n14374);
and (n14428,n14426,n14429);
or (n14429,n14430,n14433,n14461);
and (n14430,n9055,n14431);
xor (n14431,n14432,n14380);
xor (n14432,n9217,n14378);
and (n14433,n14431,n14434);
or (n14434,n14435,n14438,n14460);
and (n14435,n9142,n14436);
xor (n14436,n14437,n14384);
xor (n14437,n9185,n14382);
and (n14438,n14436,n14439);
or (n14439,n14440,n14443,n14459);
and (n14440,n9259,n14441);
xor (n14441,n14442,n14388);
xor (n14442,n9265,n14386);
and (n14443,n14441,n14444);
or (n14444,n14445,n14448,n14458);
and (n14445,n9434,n14446);
xor (n14446,n14447,n14392);
xor (n14447,n9519,n14390);
and (n14448,n14446,n14449);
or (n14449,n14450,n14453,n14457);
and (n14450,n9504,n14451);
xor (n14451,n14452,n14396);
xor (n14452,n9583,n14394);
and (n14453,n14451,n14454);
and (n14454,n9507,n14455);
xor (n14455,n14456,n14400);
xor (n14456,n9626,n14398);
and (n14457,n9504,n14454);
and (n14458,n9434,n14449);
and (n14459,n9259,n14444);
and (n14460,n9142,n14439);
and (n14461,n9055,n14434);
and (n14462,n8992,n14429);
and (n14463,n9297,n14424);
and (n14464,n8758,n14419);
and (n14465,n9076,n14414);
and (n14466,n9353,n14410);
or (n14467,n14468,n14473,n14559);
and (n14468,n14469,n14471);
xor (n14469,n14470,n14304);
xor (n14470,n9352,n14267);
xor (n14471,n14472,n14410);
xor (n14472,n9353,n14363);
and (n14473,n14471,n14474);
or (n14474,n14475,n14480,n14558);
and (n14475,n14476,n14478);
xor (n14476,n14477,n14308);
xor (n14477,n8323,n14306);
xor (n14478,n14479,n14414);
xor (n14479,n9076,n14412);
and (n14480,n14478,n14481);
or (n14481,n14482,n14487,n14557);
and (n14482,n14483,n14485);
xor (n14483,n14484,n14313);
xor (n14484,n9093,n14310);
xor (n14485,n14486,n14419);
xor (n14486,n8758,n14416);
and (n14487,n14485,n14488);
or (n14488,n14489,n14494,n14556);
and (n14489,n14490,n14492);
xor (n14490,n14491,n14318);
xor (n14491,n8927,n14315);
xor (n14492,n14493,n14424);
xor (n14493,n9297,n14421);
and (n14494,n14492,n14495);
or (n14495,n14496,n14501,n14555);
and (n14496,n14497,n14499);
xor (n14497,n14498,n14323);
xor (n14498,n9390,n14320);
xor (n14499,n14500,n14429);
xor (n14500,n8992,n14426);
and (n14501,n14499,n14502);
or (n14502,n14503,n14508,n14554);
and (n14503,n14504,n14506);
xor (n14504,n14505,n14328);
xor (n14505,n9187,n14325);
xor (n14506,n14507,n14434);
xor (n14507,n9055,n14431);
and (n14508,n14506,n14509);
or (n14509,n14510,n14515,n14553);
and (n14510,n14511,n14513);
xor (n14511,n14512,n14333);
xor (n14512,n9447,n14330);
xor (n14513,n14514,n14439);
xor (n14514,n9142,n14436);
and (n14515,n14513,n14516);
or (n14516,n14517,n14522,n14552);
and (n14517,n14518,n14520);
xor (n14518,n14519,n14338);
xor (n14519,n9536,n14335);
xor (n14520,n14521,n14444);
xor (n14521,n9259,n14441);
and (n14522,n14520,n14523);
or (n14523,n14524,n14529,n14551);
and (n14524,n14525,n14527);
xor (n14525,n14526,n14343);
xor (n14526,n9576,n14340);
xor (n14527,n14528,n14449);
xor (n14528,n9434,n14446);
and (n14529,n14527,n14530);
or (n14530,n14531,n14536,n14550);
and (n14531,n14532,n14534);
xor (n14532,n14533,n14348);
xor (n14533,n9668,n14345);
xor (n14534,n14535,n14454);
xor (n14535,n9504,n14451);
and (n14536,n14534,n14537);
or (n14537,n14538,n14541,n14549);
and (n14538,n14539,n14540);
xor (n14539,n9508,n14349);
xor (n14540,n9507,n14455);
and (n14541,n14540,n14542);
or (n14542,n14543,n14546,n14548);
and (n14543,n14544,n14545);
xor (n14544,n9803,n9880);
xor (n14545,n9657,n14401);
and (n14546,n14545,n14547);
and (n14547,n9802,n9228);
and (n14548,n14544,n14547);
and (n14549,n14539,n14542);
and (n14550,n14532,n14537);
and (n14551,n14525,n14530);
and (n14552,n14518,n14523);
and (n14553,n14511,n14516);
and (n14554,n14504,n14509);
and (n14555,n14497,n14502);
and (n14556,n14490,n14495);
and (n14557,n14483,n14488);
and (n14558,n14476,n14481);
and (n14559,n14469,n14474);
or (n14560,n14561,n14566,n14658);
and (n14561,n14562,n14564);
xor (n14562,n14563,n14177);
xor (n14563,n14172,n14174);
xor (n14564,n14565,n14474);
xor (n14565,n14469,n14471);
and (n14566,n14564,n14567);
or (n14567,n14568,n14573,n14657);
and (n14568,n14569,n14571);
xor (n14569,n14570,n14184);
xor (n14570,n14179,n14181);
xor (n14571,n14572,n14481);
xor (n14572,n14476,n14478);
and (n14573,n14571,n14574);
or (n14574,n14575,n14580,n14656);
and (n14575,n14576,n14578);
xor (n14576,n14577,n14191);
xor (n14577,n14186,n14188);
xor (n14578,n14579,n14488);
xor (n14579,n14483,n14485);
and (n14580,n14578,n14581);
or (n14581,n14582,n14587,n14655);
and (n14582,n14583,n14585);
xor (n14583,n14584,n14198);
xor (n14584,n14193,n14195);
xor (n14585,n14586,n14495);
xor (n14586,n14490,n14492);
and (n14587,n14585,n14588);
or (n14588,n14589,n14594,n14654);
and (n14589,n14590,n14592);
xor (n14590,n14591,n14205);
xor (n14591,n14200,n14202);
xor (n14592,n14593,n14502);
xor (n14593,n14497,n14499);
and (n14594,n14592,n14595);
or (n14595,n14596,n14601,n14653);
and (n14596,n14597,n14599);
xor (n14597,n14598,n14212);
xor (n14598,n14207,n14209);
xor (n14599,n14600,n14509);
xor (n14600,n14504,n14506);
and (n14601,n14599,n14602);
or (n14602,n14603,n14608,n14652);
and (n14603,n14604,n14606);
xor (n14604,n14605,n14219);
xor (n14605,n14214,n14216);
xor (n14606,n14607,n14516);
xor (n14607,n14511,n14513);
and (n14608,n14606,n14609);
or (n14609,n14610,n14615,n14651);
and (n14610,n14611,n14613);
xor (n14611,n14612,n14226);
xor (n14612,n14221,n14223);
xor (n14613,n14614,n14523);
xor (n14614,n14518,n14520);
and (n14615,n14613,n14616);
or (n14616,n14617,n14622,n14650);
and (n14617,n14618,n14620);
xor (n14618,n14619,n14233);
xor (n14619,n14228,n14230);
xor (n14620,n14621,n14530);
xor (n14621,n14525,n14527);
and (n14622,n14620,n14623);
or (n14623,n14624,n14629,n14649);
and (n14624,n14625,n14627);
xor (n14625,n14626,n14240);
xor (n14626,n14235,n14237);
xor (n14627,n14628,n14537);
xor (n14628,n14532,n14534);
and (n14629,n14627,n14630);
or (n14630,n14631,n14636,n14648);
and (n14631,n14632,n14634);
xor (n14632,n14633,n14245);
xor (n14633,n14242,n14243);
xor (n14634,n14635,n14542);
xor (n14635,n14539,n14540);
and (n14636,n14634,n14637);
or (n14637,n14638,n14643,n14647);
and (n14638,n14639,n14641);
xor (n14639,n14640,n14250);
xor (n14640,n14247,n14248);
xor (n14641,n14642,n14547);
xor (n14642,n14544,n14545);
and (n14643,n14641,n14644);
and (n14644,n14645,n14646);
xor (n14645,n9912,n9801);
xor (n14646,n9802,n9228);
and (n14647,n14639,n14644);
and (n14648,n14632,n14637);
and (n14649,n14625,n14630);
and (n14650,n14618,n14623);
and (n14651,n14611,n14616);
and (n14652,n14604,n14609);
and (n14653,n14597,n14602);
and (n14654,n14590,n14595);
and (n14655,n14583,n14588);
and (n14656,n14576,n14581);
and (n14657,n14569,n14574);
and (n14658,n14562,n14567);
and (n14659,n14660,n14662);
xor (n14660,n14661,n14567);
xor (n14661,n14562,n14564);
and (n14662,n14663,n14665);
xor (n14663,n14664,n14574);
xor (n14664,n14569,n14571);
and (n14665,n14666,n14668);
xor (n14666,n14667,n14581);
xor (n14667,n14576,n14578);
and (n14668,n14669,n14671);
xor (n14669,n14670,n14588);
xor (n14670,n14583,n14585);
and (n14671,n14672,n14674);
xor (n14672,n14673,n14595);
xor (n14673,n14590,n14592);
and (n14674,n14675,n14677);
xor (n14675,n14676,n14602);
xor (n14676,n14597,n14599);
and (n14677,n14678,n14680);
xor (n14678,n14679,n14609);
xor (n14679,n14604,n14606);
xor (n14680,n14681,n14616);
xor (n14681,n14611,n14613);
or (n14682,n14683,n14688,n7998);
and (n14683,n14684,n14685);
wire s0n14684,s1n14684,notn14684;
or (n14684,s0n14684,s1n14684);
not(notn14684,n1180);
and (s0n14684,notn14684,1'b0);
and (s1n14684,n1180,n1077);
nor (n14685,n8112,n14686,n1346);
not (n14686,n14687);
nand (n14687,n652,n726,n7,n1191);
and (n14688,n14689,n6);
wire s0n14689,s1n14689,notn14689;
or (n14689,s0n14689,s1n14689);
not(notn14689,n1194);
and (s0n14689,notn14689,1'b0);
and (s1n14689,n1194,n1077);
and (n14690,n1067,n816);
or (n14691,n14692,n14693);
and (n14692,n13941,n30);
and (n14693,n1067,n14694);
not (n14694,n30);
wire s0n14695,s1n14695,notn14695;
or (n14695,s0n14695,s1n14695);
not(notn14695,n6);
and (s0n14695,notn14695,n13939);
and (s1n14695,n6,n14696);
or (n14696,n14697,n14699);
and (n14697,n13941,n14698);
and (n14698,n803,n807,n801,n1245);
and (n14699,n1067,n14700);
not (n14700,n14698);
wire s0n14701,s1n14701,notn14701;
or (n14701,s0n14701,s1n14701);
not(notn14701,n824);
and (s0n14701,notn14701,n14702);
and (s1n14701,n824,n14707);
wire s0n14702,s1n14702,notn14702;
or (n14702,s0n14702,s1n14702);
not(notn14702,n1038);
and (s0n14702,notn14702,n14703);
and (s1n14702,n1038,n14706);
or (n14703,n14704,n14705);
and (n14704,n9978,n10005);
and (n14705,n1067,n10522);
wire s0n14706,s1n14706,notn14706;
or (n14706,s0n14706,s1n14706);
not(notn14706,n13857);
and (s0n14706,notn14706,n1067);
and (s1n14706,n13857,n9978);
wire s0n14707,s1n14707,notn14707;
or (n14707,s0n14707,s1n14707);
not(notn14707,n10109);
and (s0n14707,notn14707,n1067);
and (s1n14707,n10109,n9978);
endmodule
