module top (out,n19,n21,n26,n32,n38,n46,n48,n56,n65
        ,n73,n74,n82,n88,n99,n106,n107,n118,n135,n139
        ,n146,n163,n191,n197,n255,n320,n392,n532,n540,n561
        ,n607,n627);
output out;
input n19;
input n21;
input n26;
input n32;
input n38;
input n46;
input n48;
input n56;
input n65;
input n73;
input n74;
input n82;
input n88;
input n99;
input n106;
input n107;
input n118;
input n135;
input n139;
input n146;
input n163;
input n191;
input n197;
input n255;
input n320;
input n392;
input n532;
input n540;
input n561;
input n607;
input n627;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n20;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
xor (out,n0,n1270);
nand (n0,n1,n1269);
or (n1,n2,n367);
not (n2,n3);
nand (n3,n4,n366);
not (n4,n5);
nor (n5,n6,n300);
xor (n6,n7,n240);
xor (n7,n8,n158);
xor (n8,n9,n121);
xor (n9,n10,n92);
or (n10,n11,n91);
and (n11,n12,n67);
xor (n12,n13,n41);
nand (n13,n14,n34);
or (n14,n15,n23);
not (n15,n16);
nor (n16,n17,n22);
and (n17,n18,n20);
not (n18,n19);
not (n20,n21);
and (n22,n21,n19);
nand (n23,n24,n28);
nand (n24,n25,n27);
or (n25,n26,n20);
nand (n27,n20,n26);
not (n28,n29);
nand (n29,n30,n33);
or (n30,n31,n26);
not (n31,n32);
nand (n33,n31,n26);
nand (n34,n35,n29);
not (n35,n36);
nor (n36,n37,n39);
and (n37,n20,n38);
and (n39,n21,n40);
not (n40,n38);
nand (n41,n42,n61);
or (n42,n43,n51);
not (n43,n44);
nand (n44,n45,n49);
or (n45,n46,n47);
not (n47,n48);
or (n49,n50,n48);
not (n50,n46);
not (n51,n52);
and (n52,n53,n58);
not (n53,n54);
nand (n54,n55,n57);
or (n55,n56,n20);
nand (n57,n56,n20);
nand (n58,n59,n60);
or (n59,n56,n50);
nand (n60,n50,n56);
or (n61,n53,n62);
nor (n62,n63,n66);
and (n63,n64,n46);
not (n64,n65);
and (n66,n65,n50);
nand (n67,n68,n85);
or (n68,n69,n80);
nand (n69,n70,n77);
nor (n70,n71,n75);
and (n71,n72,n74);
not (n72,n73);
and (n75,n73,n76);
not (n76,n74);
nand (n77,n78,n79);
or (n78,n74,n31);
nand (n79,n31,n74);
nor (n80,n81,n83);
and (n81,n31,n82);
and (n83,n32,n84);
not (n84,n82);
or (n85,n70,n86);
nor (n86,n87,n89);
and (n87,n31,n88);
and (n89,n32,n90);
not (n90,n88);
and (n91,n13,n41);
nand (n92,n93,n120);
not (n93,n94);
nand (n94,n95,n113);
or (n95,n96,n101);
nor (n96,n97,n100);
and (n97,n98,n73);
not (n98,n99);
and (n100,n99,n72);
not (n101,n102);
nor (n102,n103,n109);
nand (n103,n104,n108);
or (n104,n105,n107);
not (n105,n106);
nand (n108,n105,n107);
nor (n109,n110,n111);
and (n110,n72,n107);
and (n111,n73,n112);
not (n112,n107);
nand (n113,n114,n103);
not (n114,n115);
nor (n115,n116,n119);
and (n116,n117,n73);
not (n117,n118);
and (n119,n118,n72);
not (n120,n105);
xor (n121,n122,n154);
xor (n122,n123,n129);
nand (n123,n124,n125);
or (n124,n62,n51);
nand (n125,n54,n126);
nor (n126,n127,n128);
and (n127,n46,n19);
and (n128,n18,n50);
nand (n129,n130,n142);
or (n130,n131,n137);
not (n131,n132);
nor (n132,n133,n136);
and (n133,n47,n134);
not (n134,n135);
and (n136,n135,n48);
nor (n137,n138,n140);
and (n138,n50,n139);
and (n140,n46,n141);
not (n141,n139);
nand (n142,n143,n149);
not (n143,n144);
nor (n144,n145,n147);
and (n145,n146,n134);
and (n147,n148,n135);
not (n148,n146);
not (n149,n150);
nand (n150,n137,n151);
nand (n151,n152,n153);
or (n152,n141,n135);
nand (n153,n141,n135);
nand (n154,n155,n156);
or (n155,n101,n115);
or (n156,n157,n72);
not (n157,n103);
xor (n158,n159,n209);
xor (n159,n160,n180);
xor (n160,n161,n171);
xor (n161,n162,n164);
and (n162,n135,n163);
nand (n164,n165,n170);
or (n165,n166,n28);
not (n166,n167);
nor (n167,n168,n169);
and (n168,n21,n82);
and (n169,n84,n20);
or (n170,n23,n36);
nor (n171,n172,n175);
and (n172,n173,n174);
not (n173,n69);
not (n174,n86);
and (n175,n176,n177);
not (n176,n70);
nand (n177,n178,n179);
or (n178,n32,n98);
or (n179,n31,n99);
or (n180,n181,n208);
and (n181,n182,n192);
xor (n182,n183,n190);
nand (n183,n184,n189);
or (n184,n150,n185);
nor (n185,n186,n187);
and (n186,n134,n163);
and (n187,n135,n188);
not (n188,n163);
or (n189,n137,n144);
and (n190,n135,n191);
and (n192,n193,n202);
nand (n193,n194,n201);
or (n194,n195,n198);
nand (n195,n106,n196);
not (n196,n197);
nor (n198,n199,n200);
and (n199,n117,n106);
and (n200,n118,n105);
or (n201,n105,n196);
nand (n202,n203,n207);
or (n203,n101,n204);
nor (n204,n205,n206);
and (n205,n72,n88);
and (n206,n73,n90);
or (n207,n157,n96);
and (n208,n183,n190);
or (n209,n210,n239);
and (n210,n211,n238);
xor (n211,n212,n236);
or (n212,n213,n235);
and (n213,n214,n229);
xor (n214,n215,n222);
nand (n215,n216,n221);
or (n216,n217,n23);
not (n217,n218);
nor (n218,n219,n220);
and (n219,n64,n20);
and (n220,n21,n65);
nand (n221,n16,n29);
nand (n222,n223,n224);
or (n223,n43,n53);
nand (n224,n225,n52);
not (n225,n226);
nor (n226,n227,n228);
and (n227,n146,n50);
and (n228,n148,n46);
nand (n229,n230,n234);
or (n230,n69,n231);
nor (n231,n232,n233);
and (n232,n31,n38);
and (n233,n32,n40);
or (n234,n80,n70);
and (n235,n215,n222);
nand (n236,n237,n92);
or (n237,n120,n93);
xor (n238,n12,n67);
and (n239,n212,n236);
or (n240,n241,n299);
and (n241,n242,n258);
xor (n242,n243,n244);
xor (n243,n182,n192);
or (n244,n245,n257);
and (n245,n246,n256);
xor (n246,n247,n254);
nand (n247,n248,n253);
or (n248,n150,n249);
nor (n249,n250,n251);
and (n250,n134,n191);
and (n251,n135,n252);
not (n252,n191);
or (n253,n137,n185);
and (n254,n135,n255);
xor (n256,n193,n202);
and (n257,n247,n254);
or (n258,n259,n298);
and (n259,n260,n297);
xor (n260,n261,n274);
and (n261,n262,n268);
nand (n262,n263,n267);
or (n263,n195,n264);
nor (n264,n265,n266);
and (n265,n98,n106);
and (n266,n99,n105);
or (n267,n198,n196);
nand (n268,n269,n273);
or (n269,n101,n270);
nor (n270,n271,n272);
and (n271,n72,n82);
and (n272,n73,n84);
or (n273,n157,n204);
or (n274,n275,n296);
and (n275,n276,n290);
xor (n276,n277,n284);
nand (n277,n278,n283);
or (n278,n279,n23);
not (n279,n280);
nor (n280,n281,n282);
and (n281,n47,n20);
and (n282,n21,n48);
nand (n283,n29,n218);
nand (n284,n285,n289);
or (n285,n51,n286);
nor (n286,n287,n288);
and (n287,n188,n46);
and (n288,n163,n50);
or (n289,n53,n226);
nand (n290,n291,n295);
or (n291,n69,n292);
nor (n292,n293,n294);
and (n293,n31,n19);
and (n294,n32,n18);
or (n295,n70,n231);
and (n296,n277,n284);
xor (n297,n214,n229);
and (n298,n261,n274);
and (n299,n243,n244);
or (n300,n301,n365);
and (n301,n302,n305);
xor (n302,n303,n304);
xor (n303,n211,n238);
xor (n304,n242,n258);
or (n305,n306,n364);
and (n306,n307,n323);
xor (n307,n308,n309);
xor (n308,n246,n256);
or (n309,n310,n322);
and (n310,n311,n321);
xor (n311,n312,n319);
nand (n312,n313,n318);
or (n313,n150,n314);
nor (n314,n315,n316);
and (n315,n134,n255);
and (n316,n135,n317);
not (n317,n255);
or (n318,n137,n249);
and (n319,n135,n320);
xor (n321,n262,n268);
and (n322,n312,n319);
or (n323,n324,n363);
and (n324,n325,n362);
xor (n325,n326,n339);
and (n326,n327,n333);
nand (n327,n328,n332);
or (n328,n329,n195);
nor (n329,n330,n331);
and (n330,n105,n88);
and (n331,n106,n90);
or (n332,n264,n196);
nand (n333,n334,n338);
or (n334,n101,n335);
nor (n335,n336,n337);
and (n336,n72,n38);
and (n337,n73,n40);
or (n338,n157,n270);
or (n339,n340,n361);
and (n340,n341,n355);
xor (n341,n342,n349);
nand (n342,n343,n348);
or (n343,n344,n23);
not (n344,n345);
nand (n345,n346,n347);
or (n346,n21,n148);
or (n347,n20,n146);
nand (n348,n29,n280);
nand (n349,n350,n354);
or (n350,n51,n351);
nor (n351,n352,n353);
and (n352,n252,n46);
and (n353,n191,n50);
or (n354,n53,n286);
nand (n355,n356,n360);
or (n356,n69,n357);
nor (n357,n358,n359);
and (n358,n31,n65);
and (n359,n32,n64);
or (n360,n70,n292);
and (n361,n342,n349);
xor (n362,n276,n290);
and (n363,n326,n339);
and (n364,n308,n309);
and (n365,n303,n304);
nand (n366,n6,n300);
not (n367,n368);
nand (n368,n369,n1268);
or (n369,n370,n442);
nor (n370,n371,n372);
xor (n371,n302,n305);
or (n372,n373,n441);
and (n373,n374,n377);
xor (n374,n375,n376);
xor (n375,n260,n297);
xor (n376,n307,n323);
or (n377,n378,n440);
and (n378,n379,n395);
xor (n379,n380,n381);
xor (n380,n311,n321);
or (n381,n382,n394);
and (n382,n383,n393);
xor (n383,n384,n391);
nand (n384,n385,n390);
or (n385,n150,n386);
nor (n386,n387,n388);
and (n387,n134,n320);
and (n388,n135,n389);
not (n389,n320);
or (n390,n137,n314);
and (n391,n135,n392);
xor (n393,n327,n333);
and (n394,n384,n391);
or (n395,n396,n439);
and (n396,n397,n438);
xor (n397,n398,n414);
and (n398,n399,n406);
nand (n399,n400,n405);
or (n400,n401,n195);
not (n401,n402);
nor (n402,n403,n404);
and (n403,n84,n105);
and (n404,n106,n82);
or (n405,n329,n196);
nand (n406,n407,n412);
or (n407,n408,n101);
not (n408,n409);
nor (n409,n410,n411);
and (n410,n73,n19);
and (n411,n18,n72);
nand (n412,n413,n103);
not (n413,n335);
or (n414,n415,n437);
and (n415,n416,n431);
xor (n416,n417,n424);
nand (n417,n418,n423);
or (n418,n419,n23);
not (n419,n420);
nor (n420,n421,n422);
and (n421,n21,n163);
and (n422,n188,n20);
nand (n423,n29,n345);
nand (n424,n425,n430);
or (n425,n426,n51);
not (n426,n427);
nand (n427,n428,n429);
or (n428,n46,n317);
or (n429,n50,n255);
or (n430,n53,n351);
nand (n431,n432,n436);
or (n432,n69,n433);
nor (n433,n434,n435);
and (n434,n31,n48);
and (n435,n32,n47);
or (n436,n70,n357);
and (n437,n417,n424);
xor (n438,n341,n355);
and (n439,n398,n414);
and (n440,n380,n381);
and (n441,n375,n376);
not (n442,n443);
nand (n443,n444,n1253);
or (n444,n445,n1178);
not (n445,n446);
nand (n446,n447,n888);
nor (n447,n448,n883);
and (n448,n449,n771);
and (n449,n450,n735);
nand (n450,n451,n669);
not (n451,n452);
xor (n452,n453,n609);
xor (n453,n454,n524);
xor (n454,n455,n511);
xor (n455,n456,n477);
and (n456,n457,n467);
nand (n457,n458,n462);
or (n458,n459,n195);
nor (n459,n460,n461);
and (n460,n18,n106);
and (n461,n19,n105);
or (n462,n463,n196);
not (n463,n464);
nand (n464,n465,n466);
or (n465,n38,n105);
nand (n466,n105,n38);
nand (n467,n468,n473);
or (n468,n469,n101);
not (n469,n470);
nor (n470,n471,n472);
and (n471,n73,n48);
and (n472,n47,n72);
nand (n473,n103,n474);
nand (n474,n475,n476);
or (n475,n73,n64);
or (n476,n72,n65);
or (n477,n478,n510);
and (n478,n479,n500);
xor (n479,n480,n490);
nand (n480,n481,n486);
or (n481,n482,n23);
not (n482,n483);
nor (n483,n484,n485);
and (n484,n317,n20);
and (n485,n21,n255);
nand (n486,n487,n29);
nor (n487,n488,n489);
and (n488,n252,n20);
and (n489,n21,n191);
nand (n490,n491,n496);
or (n491,n51,n492);
nor (n492,n493,n494);
and (n493,n50,n392);
and (n494,n46,n495);
not (n495,n392);
nand (n496,n54,n497);
nand (n497,n498,n499);
or (n498,n46,n389);
or (n499,n50,n320);
nand (n500,n501,n506);
or (n501,n502,n69);
not (n502,n503);
nor (n503,n504,n505);
and (n504,n188,n31);
and (n505,n32,n163);
or (n506,n70,n507);
nor (n507,n508,n509);
and (n508,n31,n146);
and (n509,n32,n148);
and (n510,n480,n490);
xor (n511,n512,n521);
xor (n512,n513,n517);
nand (n513,n514,n516);
or (n514,n515,n23);
not (n515,n487);
nand (n516,n420,n29);
nand (n517,n518,n520);
or (n518,n519,n51);
not (n519,n497);
nand (n520,n54,n427);
nand (n521,n522,n523);
or (n522,n69,n507);
or (n523,n433,n70);
xor (n524,n525,n564);
xor (n525,n526,n550);
xor (n526,n527,n541);
xor (n527,n528,n539);
nand (n528,n529,n535);
or (n529,n150,n530);
nor (n530,n531,n533);
and (n531,n532,n134);
and (n533,n534,n135);
not (n534,n532);
or (n535,n137,n536);
nor (n536,n537,n538);
and (n537,n392,n134);
and (n538,n495,n135);
and (n539,n135,n540);
xor (n541,n542,n546);
nand (n542,n543,n544);
or (n543,n196,n401);
nand (n544,n464,n545);
not (n545,n195);
nand (n546,n547,n549);
or (n547,n548,n101);
not (n548,n474);
nand (n549,n103,n409);
or (n550,n551,n563);
and (n551,n552,n562);
xor (n552,n553,n560);
nand (n553,n554,n559);
or (n554,n555,n150);
nor (n555,n556,n557);
and (n556,n134,n540);
and (n557,n135,n558);
not (n558,n540);
or (n559,n137,n530);
and (n560,n135,n561);
xor (n562,n457,n467);
and (n563,n553,n560);
and (n564,n565,n589);
or (n565,n566,n588);
and (n566,n567,n582);
xor (n567,n568,n575);
nand (n568,n569,n574);
or (n569,n570,n101);
not (n570,n571);
nor (n571,n572,n573);
and (n572,n148,n72);
and (n573,n73,n146);
nand (n574,n103,n470);
nand (n575,n576,n581);
or (n576,n577,n23);
not (n577,n578);
nor (n578,n579,n580);
and (n579,n389,n20);
and (n580,n21,n320);
nand (n581,n29,n483);
nand (n582,n583,n587);
or (n583,n51,n584);
nor (n584,n585,n586);
and (n585,n50,n532);
and (n586,n46,n534);
or (n587,n53,n492);
and (n588,n568,n575);
or (n589,n590,n608);
and (n590,n591,n606);
xor (n591,n592,n599);
nand (n592,n593,n598);
or (n593,n594,n69);
not (n594,n595);
nand (n595,n596,n597);
or (n596,n32,n252);
or (n597,n31,n191);
nand (n598,n503,n176);
nand (n599,n600,n605);
or (n600,n150,n601);
nor (n601,n602,n603);
and (n602,n134,n561);
and (n603,n604,n135);
not (n604,n561);
or (n605,n137,n555);
and (n606,n135,n607);
and (n608,n592,n599);
or (n609,n610,n668);
and (n610,n611,n614);
xor (n611,n612,n613);
xor (n612,n479,n500);
xor (n613,n552,n562);
or (n614,n615,n667);
and (n615,n616,n642);
xor (n616,n617,n623);
nand (n617,n618,n622);
or (n618,n619,n195);
nor (n619,n620,n621);
and (n620,n64,n106);
and (n621,n65,n105);
or (n622,n459,n196);
or (n623,n624,n641);
and (n624,n625,n635);
xor (n625,n626,n628);
and (n626,n135,n627);
nand (n628,n629,n634);
or (n629,n630,n101);
not (n630,n631);
nand (n631,n632,n633);
or (n632,n73,n188);
or (n633,n72,n163);
nand (n634,n571,n103);
nand (n635,n636,n637);
or (n636,n577,n28);
or (n637,n23,n638);
nor (n638,n639,n640);
and (n639,n20,n392);
and (n640,n21,n495);
and (n641,n626,n628);
or (n642,n643,n666);
and (n643,n644,n657);
xor (n644,n645,n651);
nand (n645,n646,n650);
or (n646,n51,n647);
nor (n647,n648,n649);
and (n648,n50,n540);
and (n649,n46,n558);
or (n650,n53,n584);
nand (n651,n652,n656);
or (n652,n653,n195);
nor (n653,n654,n655);
and (n654,n47,n106);
and (n655,n48,n105);
or (n656,n619,n196);
nand (n657,n658,n663);
or (n658,n659,n150);
nor (n659,n660,n661);
and (n660,n607,n134);
and (n661,n662,n135);
not (n662,n607);
nand (n663,n664,n665);
not (n664,n601);
not (n665,n137);
and (n666,n645,n651);
and (n667,n617,n623);
and (n668,n612,n613);
not (n669,n670);
or (n670,n671,n734);
and (n671,n672,n678);
xor (n672,n673,n677);
nand (n673,n674,n676);
or (n674,n589,n675);
not (n675,n565);
nand (n676,n675,n589);
xor (n677,n611,n614);
or (n678,n679,n733);
and (n679,n680,n683);
xor (n680,n681,n682);
xor (n681,n591,n606);
xor (n682,n567,n582);
or (n683,n684,n732);
and (n684,n685,n707);
xor (n685,n686,n692);
nand (n686,n687,n691);
or (n687,n69,n688);
nor (n688,n689,n690);
and (n689,n31,n255);
and (n690,n32,n317);
or (n691,n70,n594);
nor (n692,n693,n701);
not (n693,n694);
nand (n694,n695,n700);
or (n695,n696,n101);
not (n696,n697);
nor (n697,n698,n699);
and (n698,n252,n72);
and (n699,n73,n191);
nand (n700,n103,n631);
nand (n701,n702,n135);
nand (n702,n703,n704);
or (n703,n46,n139);
nand (n704,n705,n706);
or (n705,n141,n50);
not (n706,n627);
or (n707,n708,n731);
and (n708,n709,n725);
xor (n709,n710,n718);
nand (n710,n711,n716);
or (n711,n712,n23);
not (n712,n713);
nand (n713,n714,n715);
or (n714,n21,n534);
or (n715,n20,n532);
nand (n716,n717,n29);
not (n717,n638);
nand (n718,n719,n724);
or (n719,n720,n51);
not (n720,n721);
nand (n721,n722,n723);
or (n722,n46,n604);
or (n723,n50,n561);
or (n724,n53,n647);
nand (n725,n726,n730);
or (n726,n727,n195);
nor (n727,n728,n729);
and (n728,n105,n146);
and (n729,n106,n148);
or (n730,n653,n196);
and (n731,n710,n718);
and (n732,n686,n692);
and (n733,n681,n682);
and (n734,n673,n677);
nand (n735,n736,n738);
not (n736,n737);
xor (n737,n672,n678);
not (n738,n739);
or (n739,n740,n770);
and (n740,n741,n769);
xor (n741,n742,n743);
xor (n742,n616,n642);
or (n743,n744,n768);
and (n744,n745,n748);
xor (n745,n746,n747);
xor (n746,n644,n657);
xor (n747,n625,n635);
or (n748,n749,n767);
and (n749,n750,n763);
xor (n750,n751,n757);
nand (n751,n752,n756);
or (n752,n150,n753);
nor (n753,n754,n755);
and (n754,n134,n627);
and (n755,n706,n135);
or (n756,n137,n659);
nand (n757,n758,n762);
or (n758,n69,n759);
nor (n759,n760,n761);
and (n760,n31,n320);
and (n761,n32,n389);
or (n762,n70,n688);
nand (n763,n764,n766);
or (n764,n765,n693);
not (n765,n701);
or (n766,n694,n701);
and (n767,n751,n757);
and (n768,n746,n747);
xor (n769,n680,n683);
and (n770,n742,n743);
not (n771,n772);
nand (n772,n773,n880);
or (n773,n774,n874);
not (n774,n775);
nand (n775,n776,n827);
xor (n776,n777,n826);
xor (n777,n778,n779);
xor (n778,n685,n707);
or (n779,n780,n825);
and (n780,n781,n824);
xor (n781,n782,n801);
or (n782,n783,n800);
and (n783,n784,n793);
xor (n784,n785,n786);
and (n785,n665,n627);
nand (n786,n787,n792);
or (n787,n788,n101);
not (n788,n789);
nand (n789,n790,n791);
or (n790,n73,n317);
or (n791,n72,n255);
nand (n792,n103,n697);
nand (n793,n794,n799);
or (n794,n795,n23);
not (n795,n796);
nor (n796,n797,n798);
and (n797,n558,n20);
and (n798,n21,n540);
nand (n799,n29,n713);
and (n800,n785,n786);
or (n801,n802,n823);
and (n802,n803,n817);
xor (n803,n804,n811);
nand (n804,n805,n810);
or (n805,n806,n51);
not (n806,n807);
nand (n807,n808,n809);
or (n808,n46,n662);
or (n809,n50,n607);
nand (n810,n54,n721);
nand (n811,n812,n816);
or (n812,n813,n195);
nor (n813,n814,n815);
and (n814,n105,n163);
and (n815,n106,n188);
or (n816,n727,n196);
nand (n817,n818,n822);
or (n818,n69,n819);
nor (n819,n820,n821);
and (n820,n31,n392);
and (n821,n32,n495);
or (n822,n759,n70);
and (n823,n804,n811);
xor (n824,n709,n725);
and (n825,n782,n801);
xor (n826,n745,n748);
or (n827,n828,n873);
and (n828,n829,n832);
xor (n829,n830,n831);
xor (n830,n750,n763);
xor (n831,n781,n824);
or (n832,n833,n872);
and (n833,n834,n871);
xor (n834,n835,n849);
and (n835,n836,n842);
and (n836,n837,n46);
nand (n837,n838,n839);
or (n838,n21,n56);
nand (n839,n840,n706);
or (n840,n841,n20);
not (n841,n56);
nand (n842,n843,n844);
or (n843,n157,n788);
nand (n844,n845,n102);
not (n845,n846);
nor (n846,n847,n848);
and (n847,n72,n320);
and (n848,n73,n389);
or (n849,n850,n870);
and (n850,n851,n864);
xor (n851,n852,n858);
nand (n852,n853,n857);
or (n853,n23,n854);
nor (n854,n855,n856);
and (n855,n604,n21);
and (n856,n561,n20);
nand (n857,n796,n29);
nand (n858,n859,n860);
or (n859,n53,n806);
nand (n860,n52,n861);
nand (n861,n862,n863);
or (n862,n46,n706);
or (n863,n50,n627);
nand (n864,n865,n869);
or (n865,n195,n866);
nor (n866,n867,n868);
and (n867,n105,n191);
and (n868,n106,n252);
or (n869,n813,n196);
and (n870,n852,n858);
xor (n871,n784,n793);
and (n872,n835,n849);
and (n873,n830,n831);
not (n874,n875);
nand (n875,n876,n877);
xor (n876,n741,n769);
or (n877,n878,n879);
and (n878,n777,n826);
and (n879,n778,n779);
nand (n880,n881,n882);
not (n881,n876);
not (n882,n877);
nand (n883,n884,n887);
or (n884,n885,n886);
not (n885,n450);
nand (n886,n737,n739);
nand (n887,n452,n670);
nand (n888,n889,n1176,n449);
nand (n889,n890,n1166,n1175);
nand (n890,n891,n1026,n1033);
nor (n891,n892,n965);
not (n892,n893);
nand (n893,n894,n928);
not (n894,n895);
xor (n895,n896,n927);
xor (n896,n897,n898);
xor (n897,n803,n817);
or (n898,n899,n926);
and (n899,n900,n908);
xor (n900,n901,n907);
nand (n901,n902,n906);
or (n902,n69,n903);
nor (n903,n904,n905);
and (n904,n532,n31);
and (n905,n32,n534);
or (n906,n819,n70);
xor (n907,n836,n842);
or (n908,n909,n925);
and (n909,n910,n918);
xor (n910,n911,n912);
and (n911,n54,n627);
nand (n912,n913,n917);
or (n913,n914,n195);
nor (n914,n915,n916);
and (n915,n317,n106);
and (n916,n255,n105);
or (n917,n866,n196);
nand (n918,n919,n924);
or (n919,n23,n920);
not (n920,n921);
nor (n921,n922,n923);
and (n922,n662,n20);
and (n923,n21,n607);
or (n924,n28,n854);
and (n925,n911,n912);
and (n926,n901,n907);
xor (n927,n834,n871);
not (n928,n929);
or (n929,n930,n964);
and (n930,n931,n963);
xor (n931,n932,n933);
xor (n932,n851,n864);
or (n933,n934,n962);
and (n934,n935,n948);
xor (n935,n936,n942);
nand (n936,n937,n941);
or (n937,n101,n938);
nor (n938,n939,n940);
and (n939,n495,n73);
and (n940,n392,n72);
or (n941,n157,n846);
nand (n942,n943,n947);
or (n943,n69,n944);
nor (n944,n945,n946);
and (n945,n540,n31);
and (n946,n32,n558);
or (n947,n70,n903);
and (n948,n949,n955);
nor (n949,n950,n20);
nor (n950,n951,n953);
and (n951,n952,n706);
nand (n952,n32,n26);
and (n953,n31,n954);
not (n954,n26);
nand (n955,n956,n961);
or (n956,n195,n957);
not (n957,n958);
nor (n958,n959,n960);
and (n959,n106,n320);
and (n960,n389,n105);
or (n961,n914,n196);
and (n962,n936,n942);
xor (n963,n900,n908);
and (n964,n932,n933);
nand (n965,n966,n1000);
not (n966,n967);
nor (n967,n968,n969);
xor (n968,n931,n963);
or (n969,n970,n999);
and (n970,n971,n998);
xor (n971,n972,n997);
or (n972,n973,n996);
and (n973,n974,n990);
xor (n974,n975,n982);
nand (n975,n976,n981);
or (n976,n977,n23);
not (n977,n978);
nand (n978,n979,n980);
or (n979,n21,n706);
or (n980,n20,n627);
nand (n981,n921,n29);
nand (n982,n983,n988);
or (n983,n984,n101);
not (n984,n985);
nand (n985,n986,n987);
or (n986,n73,n534);
or (n987,n72,n532);
nand (n988,n989,n103);
not (n989,n938);
nand (n990,n991,n995);
or (n991,n69,n992);
nor (n992,n993,n994);
and (n993,n31,n561);
and (n994,n32,n604);
or (n995,n70,n944);
and (n996,n975,n982);
xor (n997,n910,n918);
xor (n998,n935,n948);
and (n999,n972,n997);
or (n1000,n1001,n1002);
xor (n1001,n971,n998);
or (n1002,n1003,n1025);
and (n1003,n1004,n1024);
xor (n1004,n1005,n1006);
xor (n1005,n949,n955);
or (n1006,n1007,n1023);
and (n1007,n1008,n1016);
xor (n1008,n1009,n1010);
and (n1009,n29,n627);
nand (n1010,n1011,n1012);
or (n1011,n196,n957);
or (n1012,n195,n1013);
nor (n1013,n1014,n1015);
and (n1014,n105,n392);
and (n1015,n106,n495);
nand (n1016,n1017,n1022);
or (n1017,n1018,n101);
not (n1018,n1019);
nor (n1019,n1020,n1021);
and (n1020,n73,n540);
and (n1021,n558,n72);
nand (n1022,n103,n985);
and (n1023,n1009,n1010);
xor (n1024,n974,n990);
and (n1025,n1005,n1006);
nand (n1026,n1027,n1029);
not (n1027,n1028);
xor (n1028,n829,n832);
not (n1029,n1030);
or (n1030,n1031,n1032);
and (n1031,n896,n927);
and (n1032,n897,n898);
or (n1033,n1034,n1165);
and (n1034,n1035,n1060);
xor (n1035,n1036,n1059);
or (n1036,n1037,n1058);
and (n1037,n1038,n1057);
xor (n1038,n1039,n1045);
nand (n1039,n1040,n1044);
or (n1040,n69,n1041);
nor (n1041,n1042,n1043);
and (n1042,n31,n607);
and (n1043,n32,n662);
or (n1044,n70,n992);
and (n1045,n1046,n1051);
and (n1046,n1047,n32);
nand (n1047,n1048,n1049);
or (n1048,n73,n74);
nand (n1049,n1050,n706);
or (n1050,n76,n72);
nand (n1051,n1052,n1056);
or (n1052,n1053,n195);
nor (n1053,n1054,n1055);
and (n1054,n105,n532);
and (n1055,n106,n534);
or (n1056,n1013,n196);
xor (n1057,n1008,n1016);
and (n1058,n1039,n1045);
xor (n1059,n1004,n1024);
or (n1060,n1061,n1164);
and (n1061,n1062,n1083);
xor (n1062,n1063,n1082);
or (n1063,n1064,n1081);
and (n1064,n1065,n1080);
xor (n1065,n1066,n1073);
nand (n1066,n1067,n1072);
or (n1067,n1068,n101);
not (n1068,n1069);
nor (n1069,n1070,n1071);
and (n1070,n604,n72);
and (n1071,n73,n561);
nand (n1072,n103,n1019);
nand (n1073,n1074,n1079);
or (n1074,n1075,n69);
not (n1075,n1076);
nand (n1076,n1077,n1078);
or (n1077,n706,n32);
or (n1078,n31,n627);
or (n1079,n70,n1041);
xor (n1080,n1046,n1051);
and (n1081,n1066,n1073);
xor (n1082,n1038,n1057);
or (n1083,n1084,n1163);
and (n1084,n1085,n1105);
xor (n1085,n1086,n1104);
or (n1086,n1087,n1103);
and (n1087,n1088,n1096);
xor (n1088,n1089,n1090);
nor (n1089,n70,n706);
nand (n1090,n1091,n1095);
or (n1091,n1092,n101);
nor (n1092,n1093,n1094);
and (n1093,n607,n72);
and (n1094,n662,n73);
nand (n1095,n1069,n103);
nand (n1096,n1097,n1102);
or (n1097,n195,n1098);
not (n1098,n1099);
nand (n1099,n1100,n1101);
or (n1100,n540,n105);
nand (n1101,n105,n540);
or (n1102,n1053,n196);
and (n1103,n1089,n1090);
xor (n1104,n1065,n1080);
or (n1105,n1106,n1162);
and (n1106,n1107,n1161);
xor (n1107,n1108,n1123);
nor (n1108,n1109,n1117);
not (n1109,n1110);
nand (n1110,n1111,n1116);
or (n1111,n195,n1112);
not (n1112,n1113);
nand (n1113,n1114,n1115);
or (n1114,n561,n105);
nand (n1115,n105,n561);
nand (n1116,n1099,n197);
nand (n1117,n1118,n73);
nand (n1118,n1119,n1122);
nand (n1119,n1120,n706);
not (n1120,n1121);
and (n1121,n106,n107);
or (n1122,n107,n106);
nand (n1123,n1124,n1160);
nand (n1124,n1125,n1138);
or (n1125,n1126,n1133);
not (n1126,n1127);
nor (n1127,n1128,n1132);
and (n1128,n102,n1129);
nand (n1129,n1130,n1131);
or (n1130,n73,n706);
or (n1131,n72,n627);
nor (n1132,n157,n1092);
not (n1133,n1134);
nor (n1134,n1135,n1136);
and (n1135,n1117,n1110);
and (n1136,n1137,n1109);
not (n1137,n1117);
nand (n1138,n1139,n1159);
or (n1139,n1140,n1149);
nor (n1140,n1141,n1143);
not (n1141,n1142);
nand (n1142,n103,n627);
nand (n1143,n1144,n1145);
or (n1144,n196,n1112);
nand (n1145,n1146,n545);
nand (n1146,n1147,n1148);
or (n1147,n662,n106);
nand (n1148,n106,n662);
nand (n1149,n1150,n1157);
nand (n1150,n1151,n1155);
or (n1151,n1152,n195);
nor (n1152,n1153,n1154);
and (n1153,n706,n106);
and (n1154,n627,n105);
or (n1155,n1156,n196);
not (n1156,n1146);
nor (n1157,n1158,n105);
and (n1158,n627,n197);
nand (n1159,n1141,n1143);
or (n1160,n1134,n1127);
xor (n1161,n1088,n1096);
and (n1162,n1108,n1123);
and (n1163,n1086,n1104);
and (n1164,n1063,n1082);
and (n1165,n1036,n1059);
nand (n1166,n1167,n1026);
nand (n1167,n1168,n1174);
or (n1168,n1169,n892);
not (n1169,n1170);
nand (n1170,n1171,n1173);
or (n1171,n967,n1172);
nand (n1172,n1001,n1002);
nand (n1173,n968,n969);
nand (n1174,n895,n929);
nand (n1175,n1028,n1030);
and (n1176,n880,n1177);
or (n1177,n776,n827);
not (n1178,n1179);
and (n1179,n1180,n1213,n1247);
not (n1180,n1181);
nor (n1181,n1182,n1183);
xor (n1182,n374,n377);
or (n1183,n1184,n1212);
and (n1184,n1185,n1188);
xor (n1185,n1186,n1187);
xor (n1186,n325,n362);
xor (n1187,n379,n395);
or (n1188,n1189,n1211);
and (n1189,n1190,n1202);
xor (n1190,n1191,n1192);
xor (n1191,n383,n393);
or (n1192,n1193,n1201);
and (n1193,n1194,n1200);
xor (n1194,n1195,n1199);
nand (n1195,n1196,n1197);
or (n1196,n536,n150);
nand (n1197,n1198,n665);
not (n1198,n386);
and (n1199,n135,n532);
xor (n1200,n399,n406);
and (n1201,n1195,n1199);
or (n1202,n1203,n1210);
and (n1203,n1204,n1209);
xor (n1204,n1205,n1206);
and (n1205,n542,n546);
or (n1206,n1207,n1208);
and (n1207,n512,n521);
and (n1208,n513,n517);
xor (n1209,n416,n431);
and (n1210,n1205,n1206);
and (n1211,n1191,n1192);
and (n1212,n1186,n1187);
nor (n1213,n1214,n1242);
not (n1214,n1215);
nand (n1215,n1216,n1232);
not (n1216,n1217);
xor (n1217,n1218,n1221);
xor (n1218,n1219,n1220);
xor (n1219,n397,n438);
xor (n1220,n1190,n1202);
or (n1221,n1222,n1231);
and (n1222,n1223,n1228);
xor (n1223,n1224,n1225);
xor (n1224,n1194,n1200);
or (n1225,n1226,n1227);
and (n1226,n527,n541);
and (n1227,n528,n539);
or (n1228,n1229,n1230);
and (n1229,n455,n511);
and (n1230,n456,n477);
and (n1231,n1224,n1225);
not (n1232,n1233);
or (n1233,n1234,n1241);
and (n1234,n1235,n1240);
xor (n1235,n1236,n1237);
xor (n1236,n1204,n1209);
or (n1237,n1238,n1239);
and (n1238,n525,n564);
and (n1239,n526,n550);
xor (n1240,n1223,n1228);
and (n1241,n1236,n1237);
nor (n1242,n1243,n1244);
xor (n1243,n1235,n1240);
or (n1244,n1245,n1246);
and (n1245,n453,n609);
and (n1246,n454,n524);
not (n1247,n1248);
nor (n1248,n1249,n1250);
xor (n1249,n1185,n1188);
or (n1250,n1251,n1252);
and (n1251,n1218,n1221);
and (n1252,n1219,n1220);
not (n1253,n1254);
nand (n1254,n1255,n1264);
or (n1255,n1256,n1258);
not (n1256,n1257);
nor (n1257,n1181,n1248);
nand (n1258,n1259,n1215);
or (n1259,n1260,n1262);
not (n1260,n1261);
nand (n1261,n1243,n1244);
not (n1262,n1263);
nand (n1263,n1217,n1233);
nor (n1264,n1265,n1267);
and (n1265,n1180,n1266);
and (n1266,n1249,n1250);
and (n1267,n1182,n1183);
nand (n1268,n371,n372);
or (n1269,n368,n3);
xor (n1270,n1271,n2214);
xor (n1271,n1272,n2213);
xor (n1272,n1273,n2192);
xor (n1273,n1274,n2191);
xor (n1274,n1275,n2164);
xor (n1275,n1276,n2163);
xor (n1276,n1277,n2131);
xor (n1277,n1278,n2130);
xor (n1278,n1279,n2091);
xor (n1279,n1280,n2090);
xor (n1280,n1281,n2047);
xor (n1281,n1282,n2046);
xor (n1282,n1283,n1996);
xor (n1283,n1284,n1995);
xor (n1284,n1285,n1940);
xor (n1285,n1286,n1939);
xor (n1286,n1287,n1877);
xor (n1287,n1288,n1876);
or (n1288,n1289,n1813);
and (n1289,n1290,n162);
or (n1290,n1291,n1750);
and (n1291,n1292,n190);
or (n1292,n1293,n1686);
and (n1293,n1294,n254);
or (n1294,n1295,n1623);
and (n1295,n1296,n319);
or (n1296,n1297,n1558);
and (n1297,n1298,n391);
or (n1298,n1299,n1493);
and (n1299,n1300,n1199);
or (n1300,n1301,n1430);
and (n1301,n1302,n539);
or (n1302,n1303,n1366);
and (n1303,n1304,n560);
and (n1304,n606,n1305);
or (n1305,n1306,n1308);
and (n1306,n626,n1307);
and (n1307,n139,n607);
and (n1308,n1309,n1310);
xor (n1309,n626,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
and (n1312,n139,n627);
and (n1313,n46,n607);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
and (n1318,n46,n627);
and (n1319,n56,n607);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1325);
and (n1323,n1324,n923);
and (n1324,n56,n627);
and (n1325,n1326,n1327);
xor (n1326,n1324,n923);
or (n1327,n1328,n1331);
and (n1328,n1329,n1330);
and (n1329,n21,n627);
and (n1330,n26,n607);
and (n1331,n1332,n1333);
xor (n1332,n1329,n1330);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
and (n1335,n26,n627);
and (n1336,n32,n607);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
and (n1341,n32,n627);
and (n1342,n74,n607);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
and (n1347,n74,n627);
and (n1348,n73,n607);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
and (n1353,n73,n627);
and (n1354,n107,n607);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
and (n1359,n107,n627);
and (n1360,n106,n607);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
and (n1363,n1364,n1365);
and (n1364,n106,n627);
and (n1365,n197,n607);
and (n1366,n1367,n1368);
xor (n1367,n1304,n560);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n606,n1305);
and (n1371,n139,n561);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1309,n1310);
and (n1377,n46,n561);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1315,n1316);
and (n1383,n56,n561);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1321,n1322);
and (n1389,n21,n561);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
or (n1392,n1393,n1396);
and (n1393,n1394,n1395);
xor (n1394,n1326,n1327);
and (n1395,n26,n561);
and (n1396,n1397,n1398);
xor (n1397,n1394,n1395);
or (n1398,n1399,n1402);
and (n1399,n1400,n1401);
xor (n1400,n1332,n1333);
and (n1401,n32,n561);
and (n1402,n1403,n1404);
xor (n1403,n1400,n1401);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1338,n1339);
and (n1407,n74,n561);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1413);
and (n1411,n1412,n1071);
xor (n1412,n1344,n1345);
and (n1413,n1414,n1415);
xor (n1414,n1412,n1071);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1350,n1351);
and (n1418,n107,n561);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1356,n1357);
and (n1424,n106,n561);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
and (n1427,n1428,n1429);
xor (n1428,n1362,n1363);
and (n1429,n197,n561);
and (n1430,n1431,n1432);
xor (n1431,n1302,n539);
or (n1432,n1433,n1436);
and (n1433,n1434,n1435);
xor (n1434,n1367,n1368);
and (n1435,n139,n540);
and (n1436,n1437,n1438);
xor (n1437,n1434,n1435);
or (n1438,n1439,n1442);
and (n1439,n1440,n1441);
xor (n1440,n1373,n1374);
and (n1441,n46,n540);
and (n1442,n1443,n1444);
xor (n1443,n1440,n1441);
or (n1444,n1445,n1448);
and (n1445,n1446,n1447);
xor (n1446,n1379,n1380);
and (n1447,n56,n540);
and (n1448,n1449,n1450);
xor (n1449,n1446,n1447);
or (n1450,n1451,n1453);
and (n1451,n1452,n798);
xor (n1452,n1385,n1386);
and (n1453,n1454,n1455);
xor (n1454,n1452,n798);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1391,n1392);
and (n1458,n26,n540);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1397,n1398);
and (n1464,n32,n540);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1403,n1404);
and (n1470,n74,n540);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
or (n1473,n1474,n1476);
and (n1474,n1475,n1020);
xor (n1475,n1409,n1410);
and (n1476,n1477,n1478);
xor (n1477,n1475,n1020);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1414,n1415);
and (n1481,n107,n540);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1420,n1421);
and (n1487,n106,n540);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
and (n1490,n1491,n1492);
xor (n1491,n1426,n1427);
and (n1492,n197,n540);
and (n1493,n1494,n1495);
xor (n1494,n1300,n1199);
or (n1495,n1496,n1499);
and (n1496,n1497,n1498);
xor (n1497,n1431,n1432);
and (n1498,n139,n532);
and (n1499,n1500,n1501);
xor (n1500,n1497,n1498);
or (n1501,n1502,n1505);
and (n1502,n1503,n1504);
xor (n1503,n1437,n1438);
and (n1504,n46,n532);
and (n1505,n1506,n1507);
xor (n1506,n1503,n1504);
or (n1507,n1508,n1511);
and (n1508,n1509,n1510);
xor (n1509,n1443,n1444);
and (n1510,n56,n532);
and (n1511,n1512,n1513);
xor (n1512,n1509,n1510);
or (n1513,n1514,n1517);
and (n1514,n1515,n1516);
xor (n1515,n1449,n1450);
and (n1516,n21,n532);
and (n1517,n1518,n1519);
xor (n1518,n1515,n1516);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1454,n1455);
and (n1522,n26,n532);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1460,n1461);
and (n1528,n32,n532);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1466,n1467);
and (n1534,n74,n532);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1472,n1473);
and (n1540,n73,n532);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1477,n1478);
and (n1546,n107,n532);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1483,n1484);
and (n1552,n106,n532);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
and (n1555,n1556,n1557);
xor (n1556,n1489,n1490);
and (n1557,n197,n532);
and (n1558,n1559,n1560);
xor (n1559,n1298,n391);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1494,n1495);
and (n1563,n139,n392);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
or (n1566,n1567,n1570);
and (n1567,n1568,n1569);
xor (n1568,n1500,n1501);
and (n1569,n46,n392);
and (n1570,n1571,n1572);
xor (n1571,n1568,n1569);
or (n1572,n1573,n1576);
and (n1573,n1574,n1575);
xor (n1574,n1506,n1507);
and (n1575,n56,n392);
and (n1576,n1577,n1578);
xor (n1577,n1574,n1575);
or (n1578,n1579,n1582);
and (n1579,n1580,n1581);
xor (n1580,n1512,n1513);
and (n1581,n21,n392);
and (n1582,n1583,n1584);
xor (n1583,n1580,n1581);
or (n1584,n1585,n1588);
and (n1585,n1586,n1587);
xor (n1586,n1518,n1519);
and (n1587,n26,n392);
and (n1588,n1589,n1590);
xor (n1589,n1586,n1587);
or (n1590,n1591,n1594);
and (n1591,n1592,n1593);
xor (n1592,n1524,n1525);
and (n1593,n32,n392);
and (n1594,n1595,n1596);
xor (n1595,n1592,n1593);
or (n1596,n1597,n1600);
and (n1597,n1598,n1599);
xor (n1598,n1530,n1531);
and (n1599,n74,n392);
and (n1600,n1601,n1602);
xor (n1601,n1598,n1599);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1536,n1537);
and (n1605,n73,n392);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1542,n1543);
and (n1611,n107,n392);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1548,n1549);
and (n1617,n106,n392);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
and (n1620,n1621,n1622);
xor (n1621,n1554,n1555);
and (n1622,n197,n392);
and (n1623,n1624,n1625);
xor (n1624,n1296,n319);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1559,n1560);
and (n1628,n139,n320);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1565,n1566);
and (n1634,n46,n320);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1571,n1572);
and (n1640,n56,n320);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1646);
and (n1644,n1645,n580);
xor (n1645,n1577,n1578);
and (n1646,n1647,n1648);
xor (n1647,n1645,n580);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1583,n1584);
and (n1651,n26,n320);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1589,n1590);
and (n1657,n32,n320);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1595,n1596);
and (n1663,n74,n320);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1601,n1602);
and (n1669,n73,n320);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1607,n1608);
and (n1675,n107,n320);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1681);
and (n1679,n1680,n959);
xor (n1680,n1613,n1614);
and (n1681,n1682,n1683);
xor (n1682,n1680,n959);
and (n1683,n1684,n1685);
xor (n1684,n1619,n1620);
and (n1685,n197,n320);
and (n1686,n1687,n1688);
xor (n1687,n1294,n254);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1624,n1625);
and (n1691,n139,n255);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1630,n1631);
and (n1697,n46,n255);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1636,n1637);
and (n1703,n56,n255);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1709);
and (n1707,n1708,n485);
xor (n1708,n1642,n1643);
and (n1709,n1710,n1711);
xor (n1710,n1708,n485);
or (n1711,n1712,n1715);
and (n1712,n1713,n1714);
xor (n1713,n1647,n1648);
and (n1714,n26,n255);
and (n1715,n1716,n1717);
xor (n1716,n1713,n1714);
or (n1717,n1718,n1721);
and (n1718,n1719,n1720);
xor (n1719,n1653,n1654);
and (n1720,n32,n255);
and (n1721,n1722,n1723);
xor (n1722,n1719,n1720);
or (n1723,n1724,n1727);
and (n1724,n1725,n1726);
xor (n1725,n1659,n1660);
and (n1726,n74,n255);
and (n1727,n1728,n1729);
xor (n1728,n1725,n1726);
or (n1729,n1730,n1733);
and (n1730,n1731,n1732);
xor (n1731,n1665,n1666);
and (n1732,n73,n255);
and (n1733,n1734,n1735);
xor (n1734,n1731,n1732);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1671,n1672);
and (n1738,n107,n255);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
or (n1741,n1742,n1745);
and (n1742,n1743,n1744);
xor (n1743,n1677,n1678);
and (n1744,n106,n255);
and (n1745,n1746,n1747);
xor (n1746,n1743,n1744);
and (n1747,n1748,n1749);
xor (n1748,n1682,n1683);
and (n1749,n197,n255);
and (n1750,n1751,n1752);
xor (n1751,n1292,n190);
or (n1752,n1753,n1756);
and (n1753,n1754,n1755);
xor (n1754,n1687,n1688);
and (n1755,n139,n191);
and (n1756,n1757,n1758);
xor (n1757,n1754,n1755);
or (n1758,n1759,n1762);
and (n1759,n1760,n1761);
xor (n1760,n1693,n1694);
and (n1761,n46,n191);
and (n1762,n1763,n1764);
xor (n1763,n1760,n1761);
or (n1764,n1765,n1768);
and (n1765,n1766,n1767);
xor (n1766,n1699,n1700);
and (n1767,n56,n191);
and (n1768,n1769,n1770);
xor (n1769,n1766,n1767);
or (n1770,n1771,n1773);
and (n1771,n1772,n489);
xor (n1772,n1705,n1706);
and (n1773,n1774,n1775);
xor (n1774,n1772,n489);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1710,n1711);
and (n1778,n26,n191);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1716,n1717);
and (n1784,n32,n191);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1722,n1723);
and (n1790,n74,n191);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1796);
and (n1794,n1795,n699);
xor (n1795,n1728,n1729);
and (n1796,n1797,n1798);
xor (n1797,n1795,n699);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1734,n1735);
and (n1801,n107,n191);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1740,n1741);
and (n1807,n106,n191);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
and (n1810,n1811,n1812);
xor (n1811,n1746,n1747);
and (n1812,n197,n191);
and (n1813,n1814,n1815);
xor (n1814,n1290,n162);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1751,n1752);
and (n1818,n139,n163);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1825);
and (n1822,n1823,n1824);
xor (n1823,n1757,n1758);
and (n1824,n46,n163);
and (n1825,n1826,n1827);
xor (n1826,n1823,n1824);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1763,n1764);
and (n1830,n56,n163);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
or (n1833,n1834,n1836);
and (n1834,n1835,n421);
xor (n1835,n1769,n1770);
and (n1836,n1837,n1838);
xor (n1837,n1835,n421);
or (n1838,n1839,n1842);
and (n1839,n1840,n1841);
xor (n1840,n1774,n1775);
and (n1841,n26,n163);
and (n1842,n1843,n1844);
xor (n1843,n1840,n1841);
or (n1844,n1845,n1847);
and (n1845,n1846,n505);
xor (n1846,n1780,n1781);
and (n1847,n1848,n1849);
xor (n1848,n1846,n505);
or (n1849,n1850,n1853);
and (n1850,n1851,n1852);
xor (n1851,n1786,n1787);
and (n1852,n74,n163);
and (n1853,n1854,n1855);
xor (n1854,n1851,n1852);
or (n1855,n1856,n1859);
and (n1856,n1857,n1858);
xor (n1857,n1792,n1793);
and (n1858,n73,n163);
and (n1859,n1860,n1861);
xor (n1860,n1857,n1858);
or (n1861,n1862,n1865);
and (n1862,n1863,n1864);
xor (n1863,n1797,n1798);
and (n1864,n107,n163);
and (n1865,n1866,n1867);
xor (n1866,n1863,n1864);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
xor (n1869,n1803,n1804);
and (n1870,n106,n163);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
and (n1873,n1874,n1875);
xor (n1874,n1809,n1810);
and (n1875,n197,n163);
and (n1876,n135,n146);
or (n1877,n1878,n1881);
and (n1878,n1879,n1880);
xor (n1879,n1814,n1815);
and (n1880,n139,n146);
and (n1881,n1882,n1883);
xor (n1882,n1879,n1880);
or (n1883,n1884,n1887);
and (n1884,n1885,n1886);
xor (n1885,n1820,n1821);
and (n1886,n46,n146);
and (n1887,n1888,n1889);
xor (n1888,n1885,n1886);
or (n1889,n1890,n1893);
and (n1890,n1891,n1892);
xor (n1891,n1826,n1827);
and (n1892,n56,n146);
and (n1893,n1894,n1895);
xor (n1894,n1891,n1892);
or (n1895,n1896,n1899);
and (n1896,n1897,n1898);
xor (n1897,n1832,n1833);
and (n1898,n21,n146);
and (n1899,n1900,n1901);
xor (n1900,n1897,n1898);
or (n1901,n1902,n1905);
and (n1902,n1903,n1904);
xor (n1903,n1837,n1838);
and (n1904,n26,n146);
and (n1905,n1906,n1907);
xor (n1906,n1903,n1904);
or (n1907,n1908,n1911);
and (n1908,n1909,n1910);
xor (n1909,n1843,n1844);
and (n1910,n32,n146);
and (n1911,n1912,n1913);
xor (n1912,n1909,n1910);
or (n1913,n1914,n1917);
and (n1914,n1915,n1916);
xor (n1915,n1848,n1849);
and (n1916,n74,n146);
and (n1917,n1918,n1919);
xor (n1918,n1915,n1916);
or (n1919,n1920,n1922);
and (n1920,n1921,n573);
xor (n1921,n1854,n1855);
and (n1922,n1923,n1924);
xor (n1923,n1921,n573);
or (n1924,n1925,n1928);
and (n1925,n1926,n1927);
xor (n1926,n1860,n1861);
and (n1927,n107,n146);
and (n1928,n1929,n1930);
xor (n1929,n1926,n1927);
or (n1930,n1931,n1934);
and (n1931,n1932,n1933);
xor (n1932,n1866,n1867);
and (n1933,n106,n146);
and (n1934,n1935,n1936);
xor (n1935,n1932,n1933);
and (n1936,n1937,n1938);
xor (n1937,n1872,n1873);
and (n1938,n197,n146);
and (n1939,n139,n48);
or (n1940,n1941,n1944);
and (n1941,n1942,n1943);
xor (n1942,n1882,n1883);
and (n1943,n46,n48);
and (n1944,n1945,n1946);
xor (n1945,n1942,n1943);
or (n1946,n1947,n1950);
and (n1947,n1948,n1949);
xor (n1948,n1888,n1889);
and (n1949,n56,n48);
and (n1950,n1951,n1952);
xor (n1951,n1948,n1949);
or (n1952,n1953,n1955);
and (n1953,n1954,n282);
xor (n1954,n1894,n1895);
and (n1955,n1956,n1957);
xor (n1956,n1954,n282);
or (n1957,n1958,n1961);
and (n1958,n1959,n1960);
xor (n1959,n1900,n1901);
and (n1960,n26,n48);
and (n1961,n1962,n1963);
xor (n1962,n1959,n1960);
or (n1963,n1964,n1967);
and (n1964,n1965,n1966);
xor (n1965,n1906,n1907);
and (n1966,n32,n48);
and (n1967,n1968,n1969);
xor (n1968,n1965,n1966);
or (n1969,n1970,n1973);
and (n1970,n1971,n1972);
xor (n1971,n1912,n1913);
and (n1972,n74,n48);
and (n1973,n1974,n1975);
xor (n1974,n1971,n1972);
or (n1975,n1976,n1978);
and (n1976,n1977,n471);
xor (n1977,n1918,n1919);
and (n1978,n1979,n1980);
xor (n1979,n1977,n471);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
xor (n1982,n1923,n1924);
and (n1983,n107,n48);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1929,n1930);
and (n1989,n106,n48);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
and (n1992,n1993,n1994);
xor (n1993,n1935,n1936);
and (n1994,n197,n48);
and (n1995,n46,n65);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
xor (n1998,n1945,n1946);
and (n1999,n56,n65);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2005);
and (n2003,n2004,n220);
xor (n2004,n1951,n1952);
and (n2005,n2006,n2007);
xor (n2006,n2004,n220);
or (n2007,n2008,n2011);
and (n2008,n2009,n2010);
xor (n2009,n1956,n1957);
and (n2010,n26,n65);
and (n2011,n2012,n2013);
xor (n2012,n2009,n2010);
or (n2013,n2014,n2017);
and (n2014,n2015,n2016);
xor (n2015,n1962,n1963);
and (n2016,n32,n65);
and (n2017,n2018,n2019);
xor (n2018,n2015,n2016);
or (n2019,n2020,n2023);
and (n2020,n2021,n2022);
xor (n2021,n1968,n1969);
and (n2022,n74,n65);
and (n2023,n2024,n2025);
xor (n2024,n2021,n2022);
or (n2025,n2026,n2029);
and (n2026,n2027,n2028);
xor (n2027,n1974,n1975);
and (n2028,n73,n65);
and (n2029,n2030,n2031);
xor (n2030,n2027,n2028);
or (n2031,n2032,n2035);
and (n2032,n2033,n2034);
xor (n2033,n1979,n1980);
and (n2034,n107,n65);
and (n2035,n2036,n2037);
xor (n2036,n2033,n2034);
or (n2037,n2038,n2041);
and (n2038,n2039,n2040);
xor (n2039,n1985,n1986);
and (n2040,n106,n65);
and (n2041,n2042,n2043);
xor (n2042,n2039,n2040);
and (n2043,n2044,n2045);
xor (n2044,n1991,n1992);
and (n2045,n197,n65);
and (n2046,n56,n19);
or (n2047,n2048,n2050);
and (n2048,n2049,n22);
xor (n2049,n2001,n2002);
and (n2050,n2051,n2052);
xor (n2051,n2049,n22);
or (n2052,n2053,n2056);
and (n2053,n2054,n2055);
xor (n2054,n2006,n2007);
and (n2055,n26,n19);
and (n2056,n2057,n2058);
xor (n2057,n2054,n2055);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n2012,n2013);
and (n2061,n32,n19);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n2018,n2019);
and (n2067,n74,n19);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2073);
and (n2071,n2072,n410);
xor (n2072,n2024,n2025);
and (n2073,n2074,n2075);
xor (n2074,n2072,n410);
or (n2075,n2076,n2079);
and (n2076,n2077,n2078);
xor (n2077,n2030,n2031);
and (n2078,n107,n19);
and (n2079,n2080,n2081);
xor (n2080,n2077,n2078);
or (n2081,n2082,n2085);
and (n2082,n2083,n2084);
xor (n2083,n2036,n2037);
and (n2084,n106,n19);
and (n2085,n2086,n2087);
xor (n2086,n2083,n2084);
and (n2087,n2088,n2089);
xor (n2088,n2042,n2043);
and (n2089,n197,n19);
and (n2090,n21,n38);
or (n2091,n2092,n2095);
and (n2092,n2093,n2094);
xor (n2093,n2051,n2052);
and (n2094,n26,n38);
and (n2095,n2096,n2097);
xor (n2096,n2093,n2094);
or (n2097,n2098,n2101);
and (n2098,n2099,n2100);
xor (n2099,n2057,n2058);
and (n2100,n32,n38);
and (n2101,n2102,n2103);
xor (n2102,n2099,n2100);
or (n2103,n2104,n2107);
and (n2104,n2105,n2106);
xor (n2105,n2063,n2064);
and (n2106,n74,n38);
and (n2107,n2108,n2109);
xor (n2108,n2105,n2106);
or (n2109,n2110,n2113);
and (n2110,n2111,n2112);
xor (n2111,n2069,n2070);
and (n2112,n73,n38);
and (n2113,n2114,n2115);
xor (n2114,n2111,n2112);
or (n2115,n2116,n2119);
and (n2116,n2117,n2118);
xor (n2117,n2074,n2075);
and (n2118,n107,n38);
and (n2119,n2120,n2121);
xor (n2120,n2117,n2118);
or (n2121,n2122,n2125);
and (n2122,n2123,n2124);
xor (n2123,n2080,n2081);
and (n2124,n106,n38);
and (n2125,n2126,n2127);
xor (n2126,n2123,n2124);
and (n2127,n2128,n2129);
xor (n2128,n2086,n2087);
and (n2129,n197,n38);
and (n2130,n26,n82);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2096,n2097);
and (n2134,n32,n82);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2102,n2103);
and (n2140,n74,n82);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2108,n2109);
and (n2146,n73,n82);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2114,n2115);
and (n2152,n107,n82);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2158);
and (n2156,n2157,n404);
xor (n2157,n2120,n2121);
and (n2158,n2159,n2160);
xor (n2159,n2157,n404);
and (n2160,n2161,n2162);
xor (n2161,n2126,n2127);
and (n2162,n197,n82);
and (n2163,n32,n88);
or (n2164,n2165,n2168);
and (n2165,n2166,n2167);
xor (n2166,n2136,n2137);
and (n2167,n74,n88);
and (n2168,n2169,n2170);
xor (n2169,n2166,n2167);
or (n2170,n2171,n2174);
and (n2171,n2172,n2173);
xor (n2172,n2142,n2143);
and (n2173,n73,n88);
and (n2174,n2175,n2176);
xor (n2175,n2172,n2173);
or (n2176,n2177,n2180);
and (n2177,n2178,n2179);
xor (n2178,n2148,n2149);
and (n2179,n107,n88);
and (n2180,n2181,n2182);
xor (n2181,n2178,n2179);
or (n2182,n2183,n2186);
and (n2183,n2184,n2185);
xor (n2184,n2154,n2155);
and (n2185,n106,n88);
and (n2186,n2187,n2188);
xor (n2187,n2184,n2185);
and (n2188,n2189,n2190);
xor (n2189,n2159,n2160);
and (n2190,n197,n88);
and (n2191,n74,n99);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2169,n2170);
and (n2195,n73,n99);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2175,n2176);
and (n2201,n107,n99);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2181,n2182);
and (n2207,n106,n99);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
and (n2210,n2211,n2212);
xor (n2211,n2187,n2188);
and (n2212,n197,n99);
and (n2213,n73,n118);
or (n2214,n2215,n2218);
and (n2215,n2216,n2217);
xor (n2216,n2197,n2198);
and (n2217,n107,n118);
and (n2218,n2219,n2220);
xor (n2219,n2216,n2217);
or (n2220,n2221,n2224);
and (n2221,n2222,n2223);
xor (n2222,n2203,n2204);
and (n2223,n106,n118);
and (n2224,n2225,n2226);
xor (n2225,n2222,n2223);
and (n2226,n2227,n2228);
xor (n2227,n2209,n2210);
and (n2228,n197,n118);
endmodule
