module top (out,n19,n20,n24,n26,n28,n29,n30,n33,n34
        ,n38,n40,n42,n43,n46,n48,n50,n52,n53,n54
        ,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64
        ,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74
        ,n75,n76,n77,n78,n79,n80,n89,n90,n91,n99
        ,n100,n101,n108,n109,n110,n121,n122,n123,n127,n128
        ,n129,n138,n139,n140,n151,n152,n153,n162,n163,n164
        ,n168,n169,n170,n178,n179,n180,n183,n184,n185,n197
        ,n198,n199,n206,n207,n208,n212,n213,n214,n222,n223
        ,n224,n250,n251,n252,n263,n264,n265,n272,n273,n274
        ,n281,n282,n283,n325,n326,n327,n353,n354,n355,n390
        ,n391,n392,n399,n400,n401,n410,n411,n412,n828,n829
        ,n830,n891,n892,n893,n925,n926,n930,n932,n934,n937
        ,n938,n942,n944,n946,n947,n950,n952,n954,n956,n957
        ,n958,n959,n960,n961,n962,n963,n964,n965,n966,n967
        ,n968,n969,n970,n971,n972,n973,n974,n975,n976,n977
        ,n978,n979,n980,n981,n982,n983,n984,n987,n988,n991
        ,n992,n993,n998,n999,n1003,n1004,n1005);
output out;
input n19;
input n20;
input n24;
input n26;
input n28;
input n29;
input n30;
input n33;
input n34;
input n38;
input n40;
input n42;
input n43;
input n46;
input n48;
input n50;
input n52;
input n53;
input n54;
input n55;
input n56;
input n57;
input n58;
input n59;
input n60;
input n61;
input n62;
input n63;
input n64;
input n65;
input n66;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n89;
input n90;
input n91;
input n99;
input n100;
input n101;
input n108;
input n109;
input n110;
input n121;
input n122;
input n123;
input n127;
input n128;
input n129;
input n138;
input n139;
input n140;
input n151;
input n152;
input n153;
input n162;
input n163;
input n164;
input n168;
input n169;
input n170;
input n178;
input n179;
input n180;
input n183;
input n184;
input n185;
input n197;
input n198;
input n199;
input n206;
input n207;
input n208;
input n212;
input n213;
input n214;
input n222;
input n223;
input n224;
input n250;
input n251;
input n252;
input n263;
input n264;
input n265;
input n272;
input n273;
input n274;
input n281;
input n282;
input n283;
input n325;
input n326;
input n327;
input n353;
input n354;
input n355;
input n390;
input n391;
input n392;
input n399;
input n400;
input n401;
input n410;
input n411;
input n412;
input n828;
input n829;
input n830;
input n891;
input n892;
input n893;
input n925;
input n926;
input n930;
input n932;
input n934;
input n937;
input n938;
input n942;
input n944;
input n946;
input n947;
input n950;
input n952;
input n954;
input n956;
input n957;
input n958;
input n959;
input n960;
input n961;
input n962;
input n963;
input n964;
input n965;
input n966;
input n967;
input n968;
input n969;
input n970;
input n971;
input n972;
input n973;
input n974;
input n975;
input n976;
input n977;
input n978;
input n979;
input n980;
input n981;
input n982;
input n983;
input n984;
input n987;
input n988;
input n991;
input n992;
input n993;
input n998;
input n999;
input n1003;
input n1004;
input n1005;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n39;
wire n41;
wire n44;
wire n45;
wire n47;
wire n49;
wire n51;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n124;
wire n125;
wire n126;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n165;
wire n166;
wire n167;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n181;
wire n182;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n209;
wire n210;
wire n211;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n927;
wire n928;
wire n929;
wire n931;
wire n933;
wire n935;
wire n936;
wire n939;
wire n940;
wire n941;
wire n943;
wire n945;
wire n948;
wire n949;
wire n951;
wire n953;
wire n955;
wire n985;
wire n986;
wire n989;
wire n990;
wire n994;
wire n995;
wire n996;
wire n997;
wire n1000;
wire n1001;
wire n1002;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
xnor (out,n0,n1029);
nand (n0,n1,n917);
nor (n1,n2,n915);
and (n2,n3,n810);
nand (n3,n4,n809);
or (n4,n5,n495);
not (n5,n6);
or (n6,n7,n445);
xor (n7,n8,n364);
xor (n8,n9,n290);
xor (n9,n10,n186);
xor (n10,n11,n112);
nand (n11,n12,n103);
or (n12,n13,n82);
not (n13,n14);
nand (n14,n15,n81);
or (n15,n16,n31);
not (n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n30);
and (s0n17,notn17,n18);
and (s1n17,n30,n29);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,n19);
and (s1n18,n21,n20);
and (n21,n22,n27);
and (n22,n23,n25);
not (n23,n24);
not (n25,n26);
not (n27,n28);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n44);
and (s0n31,notn31,n32);
and (s1n31,n44,n43);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n35);
and (s0n32,notn32,n33);
and (s1n32,n35,n34);
and (n35,n36,n41);
and (n36,n37,n39);
not (n37,n38);
not (n39,n40);
not (n41,n42);
and (n44,n45,n47);
not (n45,n46);
or (n47,n48,n49);
and (n49,n50,n51);
or (n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80);
nand (n81,n31,n16);
nand (n82,n83,n94);
or (n83,n84,n92);
not (n84,n85);
nand (n85,n17,n86);
not (n86,n87);
wire s0n87,s1n87,notn87;
or (n87,s0n87,s1n87);
not(notn87,n30);
and (s0n87,notn87,n88);
and (s1n87,n30,n91);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n21);
and (s0n88,notn88,n89);
and (s1n88,n21,n90);
not (n92,n93);
nand (n93,n16,n87);
not (n94,n95);
nand (n95,n96,n102);
or (n96,n97,n86);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n30);
and (s0n97,notn97,n98);
and (s1n97,n30,n101);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n21);
and (s0n98,notn98,n99);
and (s1n98,n21,n100);
nand (n102,n86,n97);
nand (n103,n104,n95);
nand (n104,n105,n111);
or (n105,n16,n106);
wire s0n106,s1n106,notn106;
or (n106,s0n106,s1n106);
not(notn106,n44);
and (s0n106,notn106,n107);
and (s1n106,n44,n110);
wire s0n107,s1n107,notn107;
or (n107,s0n107,s1n107);
not(notn107,n35);
and (s0n107,notn107,n108);
and (s1n107,n35,n109);
nand (n111,n106,n16);
nor (n112,n113,n155);
not (n113,n114);
nand (n114,n115,n146);
or (n115,n116,n131);
not (n116,n117);
nand (n117,n118,n130);
or (n118,n119,n124);
wire s0n119,s1n119,notn119;
or (n119,s0n119,s1n119);
not(notn119,n30);
and (s0n119,notn119,n120);
and (s1n119,n30,n123);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n21);
and (s0n120,notn120,n121);
and (s1n120,n21,n122);
not (n124,n125);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n44);
and (s0n125,notn125,n126);
and (s1n125,n44,n129);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n35);
and (s0n126,notn126,n127);
and (s1n126,n35,n128);
nand (n130,n124,n119);
nand (n131,n132,n142);
not (n132,n133);
nand (n133,n134,n141);
or (n134,n135,n17);
not (n135,n136);
wire s0n136,s1n136,notn136;
or (n136,s0n136,s1n136);
not(notn136,n30);
and (s0n136,notn136,n137);
and (s1n136,n30,n140);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n21);
and (s0n137,notn137,n138);
and (s1n137,n21,n139);
nand (n141,n17,n135);
nand (n142,n143,n145);
or (n143,n144,n136);
not (n144,n119);
nand (n145,n144,n136);
nand (n146,n147,n133);
nand (n147,n148,n154);
or (n148,n144,n149);
wire s0n149,s1n149,notn149;
or (n149,s0n149,s1n149);
not(notn149,n44);
and (s0n149,notn149,n150);
and (s1n149,n44,n153);
wire s0n150,s1n150,notn150;
or (n150,s0n150,s1n150);
not(notn150,n35);
and (s0n150,notn150,n151);
and (s1n150,n35,n152);
nand (n154,n149,n144);
nand (n155,n156,n181);
or (n156,n157,n171);
not (n157,n158);
nand (n158,n159,n165);
not (n159,n160);
wire s0n160,s1n160,notn160;
or (n160,s0n160,s1n160);
not(notn160,n44);
and (s0n160,notn160,n161);
and (s1n160,n44,n164);
wire s0n161,s1n161,notn161;
or (n161,s0n161,s1n161);
not(notn161,n35);
and (s0n161,notn161,n162);
and (s1n161,n35,n163);
not (n165,n166);
wire s0n166,s1n166,notn166;
or (n166,s0n166,s1n166);
not(notn166,n30);
and (s0n166,notn166,n167);
and (s1n166,n30,n170);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n21);
and (s0n167,notn167,n168);
and (s1n167,n21,n169);
not (n171,n172);
nand (n172,n173,n175);
not (n173,n174);
and (n174,n160,n166);
not (n175,n176);
wire s0n176,s1n176,notn176;
or (n176,s0n176,s1n176);
not(notn176,n30);
and (s0n176,notn176,n177);
and (s1n176,n30,n180);
wire s0n177,s1n177,notn177;
or (n177,s0n177,s1n177);
not(notn177,n21);
and (s0n177,notn177,n178);
and (s1n177,n21,n179);
wire s0n181,s1n181,notn181;
or (n181,s0n181,s1n181);
not(notn181,n30);
and (s0n181,notn181,n182);
and (s1n181,n30,n185);
wire s0n182,s1n182,notn182;
or (n182,s0n182,s1n182);
not(notn182,n21);
and (s0n182,notn182,n183);
and (s1n182,n21,n184);
or (n186,n187,n289);
and (n187,n188,n255);
xor (n188,n189,n231);
nand (n189,n190,n216);
or (n190,n191,n201);
not (n191,n192);
nand (n192,n193,n200);
or (n193,n119,n194);
not (n194,n195);
wire s0n195,s1n195,notn195;
or (n195,s0n195,s1n195);
not(notn195,n30);
and (s0n195,notn195,n196);
and (s1n195,n30,n199);
wire s0n196,s1n196,notn196;
or (n196,s0n196,s1n196);
not(notn196,n21);
and (s0n196,notn196,n197);
and (s1n196,n21,n198);
nand (n200,n194,n119);
not (n201,n202);
nand (n202,n203,n215);
or (n203,n204,n209);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n30);
and (s0n204,notn204,n205);
and (s1n204,n30,n208);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n21);
and (s0n205,notn205,n206);
and (s1n205,n21,n207);
not (n209,n210);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n44);
and (s0n210,notn210,n211);
and (s1n210,n44,n214);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n35);
and (s0n211,notn211,n212);
and (s1n211,n35,n213);
nand (n215,n209,n204);
nand (n216,n217,n226);
nand (n217,n218,n225);
or (n218,n219,n220);
not (n219,n204);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n44);
and (s0n220,notn220,n221);
and (s1n220,n44,n224);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n35);
and (s0n221,notn221,n222);
and (s1n221,n35,n223);
nand (n225,n220,n219);
not (n226,n227);
nand (n227,n191,n228);
nand (n228,n229,n230);
or (n229,n194,n204);
nand (n230,n204,n194);
nand (n231,n232,n245);
or (n232,n233,n238);
not (n233,n234);
nor (n234,n235,n237);
and (n235,n236,n159);
not (n236,n181);
and (n237,n160,n181);
nand (n238,n239,n244);
or (n239,n240,n242);
not (n240,n241);
nand (n241,n181,n165);
not (n242,n243);
nand (n243,n236,n166);
xnor (n244,n176,n166);
nand (n245,n246,n254);
nand (n246,n247,n253);
or (n247,n236,n248);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n44);
and (s0n248,notn248,n249);
and (s1n248,n44,n252);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n35);
and (s0n249,notn249,n250);
and (s1n249,n35,n251);
nand (n253,n236,n248);
not (n254,n244);
nand (n255,n256,n276);
or (n256,n257,n267);
not (n257,n258);
nand (n258,n259,n266);
or (n259,n260,n204);
not (n260,n261);
wire s0n261,s1n261,notn261;
or (n261,s0n261,s1n261);
not(notn261,n30);
and (s0n261,notn261,n262);
and (s1n261,n30,n265);
wire s0n262,s1n262,notn262;
or (n262,s0n262,s1n262);
not(notn262,n21);
and (s0n262,notn262,n263);
and (s1n262,n21,n264);
nand (n266,n204,n260);
not (n267,n268);
nand (n268,n269,n275);
or (n269,n175,n270);
wire s0n270,s1n270,notn270;
or (n270,s0n270,s1n270);
not(notn270,n44);
and (s0n270,notn270,n271);
and (s1n270,n44,n274);
wire s0n271,s1n271,notn271;
or (n271,s0n271,s1n271);
not(notn271,n35);
and (s0n271,notn271,n272);
and (s1n271,n35,n273);
nand (n275,n270,n175);
nand (n276,n277,n285);
nand (n277,n278,n284);
or (n278,n175,n279);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n44);
and (s0n279,notn279,n280);
and (s1n279,n44,n283);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n35);
and (s0n280,notn280,n281);
and (s1n280,n35,n282);
nand (n284,n279,n175);
nor (n285,n286,n258);
nor (n286,n287,n288);
and (n287,n175,n261);
and (n288,n176,n260);
and (n289,n189,n231);
or (n290,n291,n363);
and (n291,n292,n362);
xor (n292,n293,n330);
or (n293,n294,n329);
and (n294,n295,n313);
xor (n295,n296,n305);
nand (n296,n297,n304);
or (n297,n298,n303);
not (n298,n299);
nand (n299,n300,n302);
or (n300,n176,n301);
not (n301,n248);
nand (n302,n301,n176);
not (n303,n285);
nand (n304,n277,n258);
nand (n305,n306,n308);
or (n306,n191,n307);
not (n307,n217);
nand (n308,n226,n309);
nand (n309,n310,n312);
or (n310,n204,n311);
not (n311,n270);
nand (n312,n311,n204);
nand (n313,n314,n320);
or (n314,n315,n82);
not (n315,n316);
nor (n316,n317,n318);
and (n317,n149,n17);
and (n318,n16,n319);
not (n319,n149);
nand (n320,n321,n95);
nand (n321,n322,n328);
or (n322,n16,n323);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n44);
and (s0n323,notn323,n324);
and (s1n323,n44,n327);
wire s0n324,s1n324,notn324;
or (n324,s0n324,s1n324);
not(notn324,n35);
and (s0n324,notn324,n325);
and (s1n324,n35,n326);
nand (n328,n323,n16);
and (n329,n296,n305);
or (n330,n331,n361);
and (n331,n332,n341);
xor (n332,n333,n334);
nor (n333,n159,n244);
nand (n334,n335,n340);
or (n335,n131,n336);
not (n336,n337);
nand (n337,n338,n339);
or (n338,n119,n209);
nand (n339,n209,n119);
nand (n340,n117,n133);
nand (n341,n342,n356);
or (n342,n343,n348);
not (n343,n344);
nand (n344,n345,n347);
or (n345,n97,n346);
not (n346,n31);
nand (n347,n346,n97);
not (n348,n349);
nor (n349,n350,n351);
not (n350,n97);
wire s0n351,s1n351,notn351;
or (n351,s0n351,s1n351);
not(notn351,n30);
and (s0n351,notn351,n352);
and (s1n351,n30,n355);
wire s0n352,s1n352,notn352;
or (n352,s0n352,s1n352);
not(notn352,n21);
and (s0n352,notn352,n353);
and (s1n352,n21,n354);
nand (n356,n357,n351);
nand (n357,n358,n360);
or (n358,n97,n359);
not (n359,n106);
nand (n360,n359,n97);
and (n361,n333,n334);
xor (n362,n188,n255);
and (n363,n293,n330);
xor (n364,n365,n429);
xor (n365,n366,n403);
xor (n366,n367,n382);
xor (n367,n368,n375);
nand (n368,n369,n371);
or (n369,n370,n238);
not (n370,n246);
nand (n371,n372,n254);
nand (n372,n373,n374);
or (n373,n236,n279);
nand (n374,n279,n236);
nand (n375,n376,n381);
or (n376,n257,n377);
not (n377,n378);
nand (n378,n379,n380);
or (n379,n175,n220);
nand (n380,n220,n175);
nand (n381,n268,n285);
nand (n382,n383,n394);
or (n383,n348,n384);
not (n384,n385);
nand (n385,n386,n393);
or (n386,n97,n387);
not (n387,n388);
wire s0n388,s1n388,notn388;
or (n388,s0n388,s1n388);
not(notn388,n44);
and (s0n388,notn388,n389);
and (s1n388,n44,n392);
wire s0n389,s1n389,notn389;
or (n389,s0n389,s1n389);
not(notn389,n35);
and (s0n389,notn389,n390);
and (s1n389,n35,n391);
nand (n393,n387,n97);
nand (n394,n395,n351);
nand (n395,n396,n402);
or (n396,n350,n397);
wire s0n397,s1n397,notn397;
or (n397,s0n397,s1n397);
not(notn397,n44);
and (s0n397,notn397,n398);
and (s1n397,n44,n401);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n35);
and (s0n398,notn398,n399);
and (s1n398,n35,n400);
nand (n402,n397,n350);
xor (n403,n404,n423);
xor (n404,n405,n415);
nor (n405,n159,n406);
nor (n406,n407,n413);
and (n407,n236,n408);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n30);
and (s0n408,notn408,n409);
and (s1n408,n30,n412);
wire s0n409,s1n409,notn409;
or (n409,s0n409,s1n409);
not(notn409,n21);
and (s0n409,notn409,n410);
and (s1n409,n21,n411);
and (n413,n181,n414);
not (n414,n408);
nand (n415,n416,n418);
or (n416,n417,n131);
not (n417,n147);
nand (n418,n419,n133);
nand (n419,n420,n422);
or (n420,n119,n421);
not (n421,n323);
nand (n422,n421,n119);
nand (n423,n424,n425);
or (n424,n201,n227);
nand (n425,n426,n192);
nand (n426,n427,n428);
or (n427,n219,n125);
nand (n428,n125,n219);
or (n429,n430,n444);
and (n430,n431,n440);
xor (n431,n432,n436);
nand (n432,n433,n435);
or (n433,n434,n82);
not (n434,n321);
nand (n435,n95,n14);
nand (n436,n437,n439);
or (n437,n438,n348);
not (n438,n357);
nand (n439,n385,n351);
nand (n440,n441,n443);
or (n441,n442,n113);
not (n442,n155);
or (n443,n155,n114);
and (n444,n432,n436);
or (n445,n446,n494);
and (n446,n447,n450);
xor (n447,n448,n449);
xor (n448,n431,n440);
xor (n449,n292,n362);
or (n450,n451,n493);
and (n451,n452,n492);
xor (n452,n453,n467);
and (n453,n454,n460);
nor (n454,n455,n175);
and (n455,n456,n459);
nand (n456,n457,n219);
not (n457,n458);
and (n458,n160,n261);
nand (n459,n159,n260);
nand (n460,n461,n466);
or (n461,n131,n462);
not (n462,n463);
nand (n463,n464,n465);
or (n464,n144,n220);
nand (n465,n220,n144);
nand (n466,n337,n133);
or (n467,n468,n491);
and (n468,n469,n484);
xor (n469,n470,n477);
nand (n470,n471,n476);
or (n471,n348,n472);
not (n472,n473);
nand (n473,n474,n475);
or (n474,n97,n421);
nand (n475,n421,n97);
nand (n476,n344,n351);
nand (n477,n478,n483);
or (n478,n479,n82);
not (n479,n480);
nand (n480,n481,n482);
or (n481,n16,n125);
nand (n482,n125,n16);
nand (n483,n316,n95);
nand (n484,n485,n490);
or (n485,n486,n227);
not (n486,n487);
nand (n487,n488,n489);
or (n488,n219,n279);
nand (n489,n279,n219);
nand (n490,n309,n192);
and (n491,n470,n477);
xor (n492,n332,n341);
and (n493,n453,n467);
and (n494,n448,n449);
not (n495,n496);
nand (n496,n497,n793,n799);
nand (n497,n498,n539,n646);
nand (n498,n499,n501);
not (n499,n500);
xor (n500,n447,n450);
not (n501,n502);
or (n502,n503,n538);
and (n503,n504,n537);
xor (n504,n505,n506);
xor (n505,n295,n313);
or (n506,n507,n536);
and (n507,n508,n517);
xor (n508,n509,n516);
nand (n509,n510,n515);
or (n510,n303,n511);
not (n511,n512);
nor (n512,n513,n514);
and (n513,n160,n176);
and (n514,n175,n159);
nand (n515,n258,n299);
xor (n516,n454,n460);
or (n517,n518,n535);
and (n518,n519,n528);
xor (n519,n520,n521);
and (n520,n258,n160);
nand (n521,n522,n527);
or (n522,n82,n523);
not (n523,n524);
nand (n524,n525,n526);
or (n525,n17,n209);
nand (n526,n209,n17);
nand (n527,n480,n95);
nand (n528,n529,n534);
or (n529,n348,n530);
not (n530,n531);
nor (n531,n532,n533);
and (n532,n149,n97);
and (n533,n350,n319);
nand (n534,n473,n351);
and (n535,n520,n521);
and (n536,n509,n516);
xor (n537,n452,n492);
and (n538,n505,n506);
not (n539,n540);
nand (n540,n541,n639);
nor (n541,n542,n609);
nor (n542,n543,n579);
xor (n543,n544,n578);
xor (n544,n545,n546);
xor (n545,n469,n484);
or (n546,n547,n577);
and (n547,n548,n563);
xor (n548,n549,n556);
nand (n549,n550,n555);
or (n550,n551,n227);
not (n551,n552);
nand (n552,n553,n554);
or (n553,n219,n248);
nand (n554,n248,n219);
nand (n555,n487,n192);
nand (n556,n557,n562);
or (n557,n558,n131);
not (n558,n559);
nand (n559,n560,n561);
or (n560,n144,n270);
nand (n561,n270,n144);
nand (n562,n463,n133);
and (n563,n564,n571);
nand (n564,n565,n570);
or (n565,n566,n82);
not (n566,n567);
nand (n567,n568,n569);
or (n568,n16,n220);
nand (n569,n220,n16);
nand (n570,n524,n95);
nor (n571,n572,n219);
and (n572,n573,n576);
nand (n573,n574,n144);
not (n574,n575);
and (n575,n160,n195);
nand (n576,n159,n194);
and (n577,n549,n556);
xor (n578,n508,n517);
or (n579,n580,n608);
and (n580,n581,n607);
xor (n581,n582,n606);
or (n582,n583,n605);
and (n583,n584,n598);
xor (n584,n585,n591);
nand (n585,n586,n590);
nand (n586,n587,n349);
nand (n587,n588,n589);
or (n588,n350,n125);
nand (n589,n125,n350);
nand (n590,n531,n351);
nand (n591,n592,n597);
or (n592,n593,n227);
not (n593,n594);
nand (n594,n595,n596);
or (n595,n204,n159);
or (n596,n160,n219);
nand (n597,n552,n192);
nand (n598,n599,n604);
or (n599,n600,n131);
not (n600,n601);
nand (n601,n602,n603);
or (n602,n144,n279);
nand (n603,n279,n144);
nand (n604,n559,n133);
and (n605,n585,n591);
xor (n606,n519,n528);
xor (n607,n548,n563);
and (n608,n582,n606);
nor (n609,n610,n611);
xor (n610,n581,n607);
or (n611,n612,n638);
and (n612,n613,n637);
xor (n613,n614,n618);
nand (n614,n615,n617);
or (n615,n571,n616);
not (n616,n564);
nand (n617,n616,n571);
or (n618,n619,n636);
and (n619,n620,n629);
xor (n620,n621,n622);
nor (n621,n159,n191);
nand (n622,n623,n628);
or (n623,n624,n82);
not (n624,n625);
nand (n625,n626,n627);
or (n626,n17,n311);
nand (n627,n311,n17);
nand (n628,n567,n95);
nand (n629,n630,n635);
or (n630,n631,n131);
not (n631,n632);
nand (n632,n633,n634);
or (n633,n144,n248);
nand (n634,n248,n144);
nand (n635,n601,n133);
and (n636,n621,n622);
xor (n637,n584,n598);
and (n638,n614,n618);
nand (n639,n640,n642);
not (n640,n641);
xor (n641,n504,n537);
not (n642,n643);
or (n643,n644,n645);
and (n644,n544,n578);
and (n645,n545,n546);
nand (n646,n647,n792);
or (n647,n648,n679);
not (n648,n649);
nand (n649,n650,n652);
not (n650,n651);
xor (n651,n613,n637);
not (n652,n653);
or (n653,n654,n678);
and (n654,n655,n677);
xor (n655,n656,n663);
nand (n656,n657,n662);
or (n657,n348,n658);
not (n658,n659);
nand (n659,n660,n661);
or (n660,n97,n209);
nand (n661,n97,n209);
nand (n662,n587,n351);
and (n663,n664,n671);
nand (n664,n665,n666);
or (n665,n94,n624);
nand (n666,n667,n668);
not (n667,n82);
nand (n668,n669,n670);
or (n669,n16,n279);
nand (n670,n279,n16);
nor (n671,n672,n144);
and (n672,n673,n676);
nand (n673,n674,n16);
not (n674,n675);
and (n675,n160,n136);
nand (n676,n159,n135);
xor (n677,n620,n629);
and (n678,n656,n663);
not (n679,n680);
nand (n680,n681,n791);
or (n681,n682,n710);
not (n682,n683);
nand (n683,n684,n686);
not (n684,n685);
xor (n685,n655,n677);
not (n686,n687);
or (n687,n688,n709);
and (n688,n689,n705);
xor (n689,n690,n697);
nand (n690,n691,n696);
or (n691,n692,n131);
not (n692,n693);
nor (n693,n694,n695);
and (n694,n144,n159);
and (n695,n160,n119);
nand (n696,n133,n632);
nand (n697,n698,n700);
or (n698,n699,n658);
not (n699,n351);
nand (n700,n701,n349);
nand (n701,n702,n704);
or (n702,n97,n703);
not (n703,n220);
nand (n704,n97,n703);
nand (n705,n706,n708);
or (n706,n671,n707);
not (n707,n664);
nand (n708,n707,n671);
and (n709,n690,n697);
not (n710,n711);
nand (n711,n712,n790);
or (n712,n713,n785);
nor (n713,n714,n784);
and (n714,n715,n751);
nand (n715,n716,n734);
not (n716,n717);
xor (n717,n718,n727);
xor (n718,n719,n720);
and (n719,n133,n160);
nand (n720,n721,n723);
or (n721,n699,n722);
not (n722,n701);
nand (n723,n724,n349);
nand (n724,n725,n726);
or (n725,n97,n311);
nand (n726,n311,n97);
nand (n727,n728,n733);
or (n728,n729,n82);
not (n729,n730);
nand (n730,n731,n732);
or (n731,n16,n248);
nand (n732,n248,n16);
nand (n733,n668,n95);
nand (n734,n735,n744);
not (n735,n736);
nand (n736,n737,n17);
or (n737,n738,n740);
not (n738,n739);
nand (n739,n86,n159);
not (n740,n741);
nand (n741,n742,n350);
not (n742,n743);
and (n743,n160,n87);
nand (n744,n745,n747);
or (n745,n699,n746);
not (n746,n724);
nand (n747,n748,n349);
nand (n748,n749,n750);
or (n749,n350,n279);
nand (n750,n279,n350);
nand (n751,n752,n783);
nand (n752,n753,n764);
or (n753,n754,n757);
nand (n754,n755,n756);
or (n755,n736,n744);
nand (n756,n744,n736);
nand (n757,n758,n763);
or (n758,n759,n82);
not (n759,n760);
nor (n760,n761,n762);
and (n761,n16,n159);
and (n762,n160,n17);
nand (n763,n95,n730);
or (n764,n765,n782);
and (n765,n766,n775);
xor (n766,n767,n768);
and (n767,n160,n95);
nand (n768,n769,n771);
or (n769,n699,n770);
not (n770,n748);
nand (n771,n772,n349);
nand (n772,n773,n774);
or (n773,n350,n248);
nand (n774,n248,n350);
nor (n775,n776,n779);
nor (n776,n777,n778);
and (n777,n349,n159);
and (n778,n772,n351);
nand (n779,n780,n97);
not (n780,n781);
and (n781,n160,n351);
and (n782,n767,n768);
nand (n783,n754,n757);
nor (n784,n716,n734);
nor (n785,n786,n787);
xor (n786,n689,n705);
or (n787,n788,n789);
and (n788,n718,n727);
and (n789,n719,n720);
nand (n790,n786,n787);
nand (n791,n685,n687);
nand (n792,n651,n653);
nand (n793,n794,n498);
or (n794,n795,n797);
not (n795,n796);
nand (n796,n641,n643);
not (n797,n798);
nand (n798,n500,n502);
nand (n799,n498,n800);
nor (n800,n801,n808);
nand (n801,n802,n807);
or (n802,n803,n805);
not (n803,n804);
nand (n804,n610,n611);
not (n805,n806);
nand (n806,n543,n579);
not (n807,n542);
not (n808,n639);
nand (n809,n7,n445);
not (n810,n811);
nand (n811,n812,n914);
not (n812,n813);
nor (n813,n814,n911);
xor (n814,n815,n847);
xor (n815,n816,n844);
xor (n816,n817,n841);
xor (n817,n818,n838);
xor (n818,n819,n831);
nor (n819,n820,n825);
and (n820,n821,n824);
nand (n821,n822,n236);
not (n822,n823);
and (n823,n160,n408);
nand (n824,n159,n414);
not (n825,n826);
wire s0n826,s1n826,notn826;
or (n826,s0n826,s1n826);
not(notn826,n30);
and (s0n826,notn826,n827);
and (s1n826,n30,n830);
wire s0n827,s1n827,notn827;
or (n827,s0n827,s1n827);
not(notn827,n21);
and (s0n827,notn827,n828);
and (s1n827,n21,n829);
nand (n831,n832,n834);
or (n832,n227,n833);
not (n833,n426);
nand (n834,n835,n192);
nand (n835,n836,n837);
or (n836,n204,n319);
nand (n837,n319,n204);
or (n838,n839,n840);
and (n839,n404,n423);
and (n840,n405,n415);
or (n841,n842,n843);
and (n842,n367,n382);
and (n843,n368,n375);
or (n844,n845,n846);
and (n845,n365,n429);
and (n846,n366,n403);
xor (n847,n848,n908);
xor (n848,n849,n881);
xor (n849,n850,n874);
xor (n850,n851,n858);
nand (n851,n852,n854);
or (n852,n853,n238);
not (n853,n372);
nand (n854,n254,n855);
nand (n855,n856,n857);
or (n856,n236,n270);
nand (n857,n270,n236);
nand (n858,n859,n869);
or (n859,n860,n863);
nor (n860,n861,n862);
and (n861,n826,n159);
and (n862,n825,n160);
nand (n863,n864,n406);
or (n864,n865,n867);
not (n865,n866);
nand (n866,n826,n414);
not (n867,n868);
nand (n868,n825,n408);
nand (n869,n870,n873);
nand (n870,n871,n872);
or (n871,n825,n248);
nand (n872,n248,n825);
not (n873,n406);
nand (n874,n875,n877);
or (n875,n876,n82);
not (n876,n104);
nand (n877,n878,n95);
nand (n878,n879,n880);
or (n879,n16,n388);
nand (n880,n388,n16);
xor (n881,n882,n902);
xor (n882,n883,n895);
nand (n883,n884,n886);
or (n884,n885,n348);
not (n885,n395);
nand (n886,n887,n351);
nand (n887,n888,n894);
or (n888,n350,n889);
wire s0n889,s1n889,notn889;
or (n889,s0n889,s1n889);
not(notn889,n44);
and (s0n889,notn889,n890);
and (s1n889,n44,n893);
wire s0n890,s1n890,notn890;
or (n890,s0n890,s1n890);
not(notn890,n35);
and (s0n890,notn890,n891);
and (s1n890,n35,n892);
nand (n894,n889,n350);
nand (n895,n896,n898);
nand (n896,n897,n419);
not (n897,n131);
nand (n898,n133,n899);
nand (n899,n900,n901);
or (n900,n119,n346);
nand (n901,n346,n119);
nand (n902,n903,n904);
or (n903,n303,n377);
nand (n904,n905,n258);
nand (n905,n906,n907);
or (n906,n175,n210);
nand (n907,n210,n175);
or (n908,n909,n910);
and (n909,n10,n186);
and (n910,n11,n112);
or (n911,n912,n913);
and (n912,n8,n364);
and (n913,n9,n290);
nand (n914,n814,n911);
and (n915,n916,n811);
not (n916,n3);
not (n917,n918);
or (n918,n919,n1016,n1028);
and (n919,n920,n1006);
xor (n920,n921,n1000);
xor (n921,n922,n994);
xor (n922,n923,n985);
and (n923,n924,n935);
wire s0n924,s1n924,notn924;
or (n924,s0n924,s1n924);
not(notn924,n927);
and (s0n924,notn924,n925);
and (s1n924,n927,n926);
and (n927,n928,n933);
and (n928,n929,n931);
not (n929,n930);
not (n931,n932);
not (n933,n934);
wire s0n935,s1n935,notn935;
or (n935,s0n935,s1n935);
not(notn935,n948);
and (s0n935,notn935,n936);
and (s1n935,n948,n947);
wire s0n936,s1n936,notn936;
or (n936,s0n936,s1n936);
not(notn936,n939);
and (s0n936,notn936,n937);
and (s1n936,n939,n938);
and (n939,n940,n945);
and (n940,n941,n943);
not (n941,n942);
not (n943,n944);
not (n945,n946);
and (n948,n949,n951);
not (n949,n950);
or (n951,n952,n953);
and (n953,n954,n955);
or (n955,n956,n957,n958,n959,n960,n961,n962,n963,n964,n965,n966,n967,n968,n969,n970,n971,n972,n973,n974,n975,n976,n977,n978,n979,n980,n981,n982,n983,n984);
and (n985,n986,n989);
wire s0n986,s1n986,notn986;
or (n986,s0n986,s1n986);
not(notn986,n927);
and (s0n986,notn986,n987);
and (s1n986,n927,n988);
wire s0n989,s1n989,notn989;
or (n989,s0n989,s1n989);
not(notn989,n948);
and (s0n989,notn989,n990);
and (s1n989,n948,n993);
wire s0n990,s1n990,notn990;
or (n990,s0n990,s1n990);
not(notn990,n939);
and (s0n990,notn990,n991);
and (s1n990,n939,n992);
and (n994,n995,n996);
and (n995,n986,n935);
and (n996,n997,n989);
wire s0n997,s1n997,notn997;
or (n997,s0n997,s1n997);
not(notn997,n927);
and (s0n997,notn997,n998);
and (s1n997,n927,n999);
and (n1000,n997,n1001);
wire s0n1001,s1n1001,notn1001;
or (n1001,s0n1001,s1n1001);
not(notn1001,n948);
and (s0n1001,notn1001,n1002);
and (s1n1001,n948,n1005);
wire s0n1002,s1n1002,notn1002;
or (n1002,s0n1002,s1n1002);
not(notn1002,n939);
and (s0n1002,notn1002,n1003);
and (s1n1002,n939,n1004);
not (n1006,n1007);
xor (n1007,n1008,n1015);
xor (n1008,n1009,n1012);
xor (n1009,n1010,n1011);
and (n1010,n88,n160);
and (n1011,n98,n248);
and (n1012,n1013,n1014);
and (n1013,n98,n160);
and (n1014,n352,n248);
and (n1015,n352,n279);
and (n1016,n1006,n1017);
or (n1017,n1018,n1022,n1027);
and (n1018,n1019,n1020);
xor (n1019,n995,n996);
not (n1020,n1021);
xor (n1021,n1013,n1014);
and (n1022,n1020,n1023);
or (n1023,n1024,n1025);
and (n1024,n997,n935);
not (n1025,n1026);
and (n1026,n352,n160);
and (n1027,n1019,n1023);
and (n1028,n920,n1017);
or (n1029,n1030,n1854);
and (n1030,n1031,n1780);
xor (n1031,n1032,n1760);
xor (n1032,n1033,n1693);
xor (n1033,n1034,n1668);
xor (n1034,n1035,n1607);
xor (n1035,n1036,n1577);
xor (n1036,n1037,n1523);
xor (n1037,n1038,n1488);
xor (n1038,n1039,n1439);
xor (n1039,n1040,n1399);
xor (n1040,n1041,n1356);
xor (n1041,n1042,n1311);
xor (n1042,n1043,n1272);
xor (n1043,n1044,n1161);
xor (n1044,n1045,n1129);
xor (n1045,n1046,n1128);
xor (n1046,n1047,n1103);
xor (n1047,n1048,n1102);
xor (n1048,n1049,n1083);
xor (n1049,n1050,n1082);
xor (n1050,n1051,n1069);
xor (n1051,n1052,n1068);
xor (n1052,n1053,n1061);
xor (n1053,n1054,n1060);
xor (n1054,n1055,n1056);
and (n1055,n917,n781);
and (n1056,n917,n1057);
xor (n1057,n1058,n1059);
and (n1058,n248,n351);
and (n1059,n160,n97);
and (n1060,n1055,n1056);
and (n1061,n917,n1062);
xor (n1062,n1063,n743);
xor (n1063,n1064,n1067);
xor (n1064,n1065,n1066);
and (n1065,n279,n351);
and (n1066,n248,n97);
and (n1067,n1058,n1059);
and (n1068,n1053,n1061);
and (n1069,n917,n1070);
xor (n1070,n1071,n762);
xor (n1071,n1072,n1081);
xor (n1072,n1073,n1080);
xor (n1073,n1074,n1077);
xor (n1074,n1075,n1076);
and (n1075,n270,n351);
and (n1076,n279,n97);
or (n1077,n1078,n1079);
and (n1078,n1065,n1066);
and (n1079,n1064,n1067);
and (n1080,n248,n87);
and (n1081,n1063,n743);
and (n1082,n1051,n1069);
and (n1083,n917,n1084);
xor (n1084,n1085,n675);
xor (n1085,n1086,n1101);
xor (n1086,n1087,n1100);
xor (n1087,n1088,n1097);
xor (n1088,n1089,n1096);
xor (n1089,n1090,n1093);
xor (n1090,n1091,n1092);
and (n1091,n220,n351);
and (n1092,n270,n97);
or (n1093,n1094,n1095);
and (n1094,n1075,n1076);
and (n1095,n1074,n1077);
and (n1096,n279,n87);
or (n1097,n1098,n1099);
and (n1098,n1073,n1080);
and (n1099,n1072,n1081);
and (n1100,n248,n17);
and (n1101,n1071,n762);
and (n1102,n1049,n1083);
and (n1103,n917,n1104);
xor (n1104,n1105,n695);
xor (n1105,n1106,n1127);
xor (n1106,n1107,n1126);
xor (n1107,n1108,n1123);
xor (n1108,n1109,n1122);
xor (n1109,n1110,n1119);
xor (n1110,n1111,n1118);
xor (n1111,n1112,n1115);
xor (n1112,n1113,n1114);
and (n1113,n210,n351);
and (n1114,n220,n97);
or (n1115,n1116,n1117);
and (n1116,n1091,n1092);
and (n1117,n1090,n1093);
and (n1118,n270,n87);
or (n1119,n1120,n1121);
and (n1120,n1089,n1096);
and (n1121,n1088,n1097);
and (n1122,n279,n17);
or (n1123,n1124,n1125);
and (n1124,n1087,n1100);
and (n1125,n1086,n1101);
and (n1126,n248,n136);
and (n1127,n1085,n675);
and (n1128,n1047,n1103);
not (n1129,n1130);
nand (n1130,n1131,n917);
xor (n1131,n1132,n575);
xor (n1132,n1133,n1160);
xor (n1133,n1134,n1159);
xor (n1134,n1135,n1156);
xor (n1135,n1136,n1155);
xor (n1136,n1137,n1152);
xor (n1137,n1138,n1151);
xor (n1138,n1139,n1148);
xor (n1139,n1140,n1147);
xor (n1140,n1141,n1144);
xor (n1141,n1142,n1143);
and (n1142,n125,n351);
and (n1143,n210,n97);
or (n1144,n1145,n1146);
and (n1145,n1113,n1114);
and (n1146,n1112,n1115);
and (n1147,n220,n87);
or (n1148,n1149,n1150);
and (n1149,n1111,n1118);
and (n1150,n1110,n1119);
and (n1151,n270,n17);
or (n1152,n1153,n1154);
and (n1153,n1109,n1122);
and (n1154,n1108,n1123);
and (n1155,n279,n136);
or (n1156,n1157,n1158);
and (n1157,n1107,n1126);
and (n1158,n1106,n1127);
and (n1159,n248,n119);
and (n1160,n1105,n695);
or (n1161,n1162,n1163);
and (n1162,n1045,n1129);
and (n1163,n1044,n1164);
or (n1164,n1162,n1165);
and (n1165,n1044,n1166);
or (n1166,n1162,n1167);
and (n1167,n1044,n1168);
or (n1168,n1162,n1169);
and (n1169,n1044,n1170);
or (n1170,n1162,n1171);
and (n1171,n1044,n1172);
or (n1172,n1162,n1173);
and (n1173,n1044,n1174);
or (n1174,n1162,n1175);
and (n1175,n1044,n1176);
or (n1176,n1177,n1261);
and (n1177,n1178,n1260);
xor (n1178,n1046,n1179);
or (n1179,n1180,n1249);
and (n1180,n1181,n1248);
xor (n1181,n1048,n1182);
or (n1182,n1183,n1237);
and (n1183,n1184,n1236);
xor (n1184,n1050,n1185);
or (n1185,n1186,n1224);
and (n1186,n1187,n1223);
xor (n1187,n1052,n1188);
or (n1188,n1189,n1211);
and (n1189,n1190,n1210);
xor (n1190,n1054,n1191);
or (n1191,n1192,n1196);
and (n1192,n1055,n1193);
and (n1193,n1194,n1057);
xor (n1194,n1195,n1017);
xor (n1195,n920,n1006);
and (n1196,n1197,n1198);
xor (n1197,n1055,n1193);
or (n1198,n1199,n1204);
and (n1199,n1200,n1201);
and (n1200,n1194,n781);
and (n1201,n1202,n1057);
xor (n1202,n1203,n1023);
xor (n1203,n1019,n1020);
and (n1204,n1205,n1206);
xor (n1205,n1200,n1201);
and (n1206,n1207,n1208);
and (n1207,n1202,n781);
and (n1208,n1209,n1057);
xor (n1209,n1024,n1026);
and (n1210,n1194,n1062);
and (n1211,n1212,n1213);
xor (n1212,n1190,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1197,n1198);
and (n1216,n1202,n1062);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
and (n1219,n1220,n1221);
xor (n1220,n1205,n1206);
not (n1221,n1222);
nand (n1222,n1062,n1209);
and (n1223,n1194,n1070);
and (n1224,n1225,n1226);
xor (n1225,n1187,n1223);
or (n1226,n1227,n1230);
and (n1227,n1228,n1229);
xor (n1228,n1212,n1213);
and (n1229,n1202,n1070);
and (n1230,n1231,n1232);
xor (n1231,n1228,n1229);
and (n1232,n1233,n1234);
xor (n1233,n1218,n1219);
not (n1234,n1235);
nand (n1235,n1070,n1209);
and (n1236,n1194,n1084);
and (n1237,n1238,n1239);
xor (n1238,n1184,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1225,n1226);
and (n1242,n1202,n1084);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
and (n1245,n1246,n1247);
xor (n1246,n1231,n1232);
and (n1247,n1084,n1209);
and (n1248,n1194,n1104);
and (n1249,n1250,n1251);
xor (n1250,n1181,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1238,n1239);
and (n1254,n1104,n1202);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
and (n1257,n1258,n1259);
xor (n1258,n1244,n1245);
and (n1259,n1104,n1209);
and (n1260,n1131,n1194);
and (n1261,n1262,n1263);
xor (n1262,n1178,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1250,n1251);
and (n1266,n1202,n1131);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
and (n1269,n1270,n1271);
xor (n1270,n1256,n1257);
and (n1271,n1131,n1209);
not (n1272,n1273);
nand (n1273,n1274,n917);
xor (n1274,n1275,n1310);
xor (n1275,n1276,n1309);
xor (n1276,n1277,n1308);
xor (n1277,n1278,n1305);
xor (n1278,n1279,n1304);
xor (n1279,n1280,n1301);
xor (n1280,n1281,n1300);
xor (n1281,n1282,n1297);
xor (n1282,n1283,n1296);
xor (n1283,n1284,n1293);
xor (n1284,n1285,n1292);
xor (n1285,n1286,n1289);
xor (n1286,n1287,n1288);
and (n1287,n149,n351);
and (n1288,n125,n97);
or (n1289,n1290,n1291);
and (n1290,n1142,n1143);
and (n1291,n1141,n1144);
and (n1292,n210,n87);
or (n1293,n1294,n1295);
and (n1294,n1140,n1147);
and (n1295,n1139,n1148);
and (n1296,n220,n17);
or (n1297,n1298,n1299);
and (n1298,n1138,n1151);
and (n1299,n1137,n1152);
and (n1300,n270,n136);
or (n1301,n1302,n1303);
and (n1302,n1136,n1155);
and (n1303,n1135,n1156);
and (n1304,n279,n119);
or (n1305,n1306,n1307);
and (n1306,n1134,n1159);
and (n1307,n1133,n1160);
and (n1308,n248,n195);
and (n1309,n1132,n575);
and (n1310,n160,n204);
or (n1311,n1312,n1314);
and (n1312,n1313,n1272);
xor (n1313,n1044,n1164);
and (n1314,n1315,n1316);
xor (n1315,n1313,n1272);
or (n1316,n1317,n1319);
and (n1317,n1318,n1272);
xor (n1318,n1044,n1166);
and (n1319,n1320,n1321);
xor (n1320,n1318,n1272);
or (n1321,n1322,n1324);
and (n1322,n1323,n1272);
xor (n1323,n1044,n1168);
and (n1324,n1325,n1326);
xor (n1325,n1323,n1272);
or (n1326,n1327,n1329);
and (n1327,n1328,n1272);
xor (n1328,n1044,n1170);
and (n1329,n1330,n1331);
xor (n1330,n1328,n1272);
or (n1331,n1332,n1334);
and (n1332,n1333,n1272);
xor (n1333,n1044,n1172);
and (n1334,n1335,n1336);
xor (n1335,n1333,n1272);
or (n1336,n1337,n1339);
and (n1337,n1338,n1272);
xor (n1338,n1044,n1174);
and (n1339,n1340,n1341);
xor (n1340,n1338,n1272);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1044,n1176);
and (n1344,n1274,n1194);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1351);
and (n1348,n1349,n1350);
xor (n1349,n1262,n1263);
and (n1350,n1202,n1274);
and (n1351,n1352,n1353);
xor (n1352,n1349,n1350);
and (n1353,n1354,n1355);
xor (n1354,n1268,n1269);
and (n1355,n1209,n1274);
not (n1356,n1357);
nand (n1357,n1358,n917);
xor (n1358,n1359,n458);
xor (n1359,n1360,n1398);
xor (n1360,n1361,n1397);
xor (n1361,n1362,n1394);
xor (n1362,n1363,n1393);
xor (n1363,n1364,n1390);
xor (n1364,n1365,n1389);
xor (n1365,n1366,n1386);
xor (n1366,n1367,n1385);
xor (n1367,n1368,n1382);
xor (n1368,n1369,n1381);
xor (n1369,n1370,n1378);
xor (n1370,n1371,n1377);
xor (n1371,n1372,n1374);
xor (n1372,n1373,n532);
and (n1373,n323,n351);
or (n1374,n1375,n1376);
and (n1375,n1287,n1288);
and (n1376,n1286,n1289);
and (n1377,n125,n87);
or (n1378,n1379,n1380);
and (n1379,n1285,n1292);
and (n1380,n1284,n1293);
and (n1381,n210,n17);
or (n1382,n1383,n1384);
and (n1383,n1283,n1296);
and (n1384,n1282,n1297);
and (n1385,n220,n136);
or (n1386,n1387,n1388);
and (n1387,n1281,n1300);
and (n1388,n1280,n1301);
and (n1389,n270,n119);
or (n1390,n1391,n1392);
and (n1391,n1279,n1304);
and (n1392,n1278,n1305);
and (n1393,n279,n195);
or (n1394,n1395,n1396);
and (n1395,n1277,n1308);
and (n1396,n1276,n1309);
and (n1397,n248,n204);
and (n1398,n1275,n1310);
or (n1399,n1400,n1402);
and (n1400,n1401,n1356);
xor (n1401,n1315,n1316);
and (n1402,n1403,n1404);
xor (n1403,n1401,n1356);
or (n1404,n1405,n1407);
and (n1405,n1406,n1356);
xor (n1406,n1320,n1321);
and (n1407,n1408,n1409);
xor (n1408,n1406,n1356);
or (n1409,n1410,n1412);
and (n1410,n1411,n1356);
xor (n1411,n1325,n1326);
and (n1412,n1413,n1414);
xor (n1413,n1411,n1356);
or (n1414,n1415,n1417);
and (n1415,n1416,n1356);
xor (n1416,n1330,n1331);
and (n1417,n1418,n1419);
xor (n1418,n1416,n1356);
or (n1419,n1420,n1422);
and (n1420,n1421,n1356);
xor (n1421,n1335,n1336);
and (n1422,n1423,n1424);
xor (n1423,n1421,n1356);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1340,n1341);
and (n1427,n1358,n1194);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1346,n1347);
and (n1433,n1358,n1202);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
and (n1436,n1437,n1438);
xor (n1437,n1352,n1353);
and (n1438,n1358,n1209);
and (n1439,n917,n1440);
xor (n1440,n1441,n513);
xor (n1441,n1442,n1487);
xor (n1442,n1443,n1486);
xor (n1443,n1444,n1483);
xor (n1444,n1445,n1482);
xor (n1445,n1446,n1479);
xor (n1446,n1447,n1478);
xor (n1447,n1448,n1475);
xor (n1448,n1449,n1474);
xor (n1449,n1450,n1471);
xor (n1450,n1451,n1470);
xor (n1451,n1452,n1467);
xor (n1452,n1453,n1466);
xor (n1453,n1454,n1463);
xor (n1454,n1455,n1462);
xor (n1455,n1456,n1459);
xor (n1456,n1457,n1458);
and (n1457,n31,n351);
and (n1458,n323,n97);
or (n1459,n1460,n1461);
and (n1460,n1373,n532);
and (n1461,n1372,n1374);
and (n1462,n149,n87);
or (n1463,n1464,n1465);
and (n1464,n1371,n1377);
and (n1465,n1370,n1378);
and (n1466,n125,n17);
or (n1467,n1468,n1469);
and (n1468,n1369,n1381);
and (n1469,n1368,n1382);
and (n1470,n210,n136);
or (n1471,n1472,n1473);
and (n1472,n1367,n1385);
and (n1473,n1366,n1386);
and (n1474,n220,n119);
or (n1475,n1476,n1477);
and (n1476,n1365,n1389);
and (n1477,n1364,n1390);
and (n1478,n270,n195);
or (n1479,n1480,n1481);
and (n1480,n1363,n1393);
and (n1481,n1362,n1394);
and (n1482,n279,n204);
or (n1483,n1484,n1485);
and (n1484,n1361,n1397);
and (n1485,n1360,n1398);
and (n1486,n248,n261);
and (n1487,n1359,n458);
or (n1488,n1489,n1491);
and (n1489,n1490,n1439);
xor (n1490,n1403,n1404);
and (n1491,n1492,n1493);
xor (n1492,n1490,n1439);
or (n1493,n1494,n1496);
and (n1494,n1495,n1439);
xor (n1495,n1408,n1409);
and (n1496,n1497,n1498);
xor (n1497,n1495,n1439);
or (n1498,n1499,n1501);
and (n1499,n1500,n1439);
xor (n1500,n1413,n1414);
and (n1501,n1502,n1503);
xor (n1502,n1500,n1439);
or (n1503,n1504,n1506);
and (n1504,n1505,n1439);
xor (n1505,n1418,n1419);
and (n1506,n1507,n1508);
xor (n1507,n1505,n1439);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1423,n1424);
and (n1511,n1194,n1440);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1429,n1430);
and (n1517,n1202,n1440);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
and (n1520,n1521,n1522);
xor (n1521,n1435,n1436);
and (n1522,n1209,n1440);
and (n1523,n917,n1524);
xor (n1524,n1525,n174);
xor (n1525,n1526,n1576);
xor (n1526,n1527,n1575);
xor (n1527,n1528,n1572);
xor (n1528,n1529,n1571);
xor (n1529,n1530,n1568);
xor (n1530,n1531,n1567);
xor (n1531,n1532,n1564);
xor (n1532,n1533,n1563);
xor (n1533,n1534,n1560);
xor (n1534,n1535,n1559);
xor (n1535,n1536,n1556);
xor (n1536,n1537,n1555);
xor (n1537,n1538,n1552);
xor (n1538,n1539,n317);
xor (n1539,n1540,n1549);
xor (n1540,n1541,n1548);
xor (n1541,n1542,n1545);
xor (n1542,n1543,n1544);
and (n1543,n106,n351);
and (n1544,n31,n97);
or (n1545,n1546,n1547);
and (n1546,n1457,n1458);
and (n1547,n1456,n1459);
and (n1548,n323,n87);
or (n1549,n1550,n1551);
and (n1550,n1455,n1462);
and (n1551,n1454,n1463);
or (n1552,n1553,n1554);
and (n1553,n1453,n1466);
and (n1554,n1452,n1467);
and (n1555,n125,n136);
or (n1556,n1557,n1558);
and (n1557,n1451,n1470);
and (n1558,n1450,n1471);
and (n1559,n210,n119);
or (n1560,n1561,n1562);
and (n1561,n1449,n1474);
and (n1562,n1448,n1475);
and (n1563,n220,n195);
or (n1564,n1565,n1566);
and (n1565,n1447,n1478);
and (n1566,n1446,n1479);
and (n1567,n270,n204);
or (n1568,n1569,n1570);
and (n1569,n1445,n1482);
and (n1570,n1444,n1483);
and (n1571,n279,n261);
or (n1572,n1573,n1574);
and (n1573,n1443,n1486);
and (n1574,n1442,n1487);
and (n1575,n248,n176);
and (n1576,n1441,n513);
or (n1577,n1578,n1580);
and (n1578,n1579,n1523);
xor (n1579,n1492,n1493);
and (n1580,n1581,n1582);
xor (n1581,n1579,n1523);
or (n1582,n1583,n1585);
and (n1583,n1584,n1523);
xor (n1584,n1497,n1498);
and (n1585,n1586,n1587);
xor (n1586,n1584,n1523);
or (n1587,n1588,n1590);
and (n1588,n1589,n1523);
xor (n1589,n1502,n1503);
and (n1590,n1591,n1592);
xor (n1591,n1589,n1523);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1507,n1508);
and (n1595,n1194,n1524);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1513,n1514);
and (n1601,n1202,n1524);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
and (n1604,n1605,n1606);
xor (n1605,n1519,n1520);
and (n1606,n1209,n1524);
and (n1607,n917,n1608);
xor (n1608,n1609,n237);
xor (n1609,n1610,n1667);
xor (n1610,n1611,n1666);
xor (n1611,n1612,n1663);
xor (n1612,n1613,n1662);
xor (n1613,n1614,n1659);
xor (n1614,n1615,n1658);
xor (n1615,n1616,n1655);
xor (n1616,n1617,n1654);
xor (n1617,n1618,n1651);
xor (n1618,n1619,n1650);
xor (n1619,n1620,n1647);
xor (n1620,n1621,n1646);
xor (n1621,n1622,n1643);
xor (n1622,n1623,n1642);
xor (n1623,n1624,n1639);
xor (n1624,n1625,n1638);
xor (n1625,n1626,n1635);
xor (n1626,n1627,n1634);
xor (n1627,n1628,n1631);
xor (n1628,n1629,n1630);
and (n1629,n388,n351);
and (n1630,n106,n97);
or (n1631,n1632,n1633);
and (n1632,n1543,n1544);
and (n1633,n1542,n1545);
and (n1634,n31,n87);
or (n1635,n1636,n1637);
and (n1636,n1541,n1548);
and (n1637,n1540,n1549);
and (n1638,n323,n17);
or (n1639,n1640,n1641);
and (n1640,n1539,n317);
and (n1641,n1538,n1552);
and (n1642,n149,n136);
or (n1643,n1644,n1645);
and (n1644,n1537,n1555);
and (n1645,n1536,n1556);
and (n1646,n125,n119);
or (n1647,n1648,n1649);
and (n1648,n1535,n1559);
and (n1649,n1534,n1560);
and (n1650,n210,n195);
or (n1651,n1652,n1653);
and (n1652,n1533,n1563);
and (n1653,n1532,n1564);
and (n1654,n220,n204);
or (n1655,n1656,n1657);
and (n1656,n1531,n1567);
and (n1657,n1530,n1568);
and (n1658,n270,n261);
or (n1659,n1660,n1661);
and (n1660,n1529,n1571);
and (n1661,n1528,n1572);
and (n1662,n279,n176);
or (n1663,n1664,n1665);
and (n1664,n1527,n1575);
and (n1665,n1526,n1576);
and (n1666,n248,n166);
and (n1667,n1525,n174);
or (n1668,n1669,n1671);
and (n1669,n1670,n1607);
xor (n1670,n1581,n1582);
and (n1671,n1672,n1673);
xor (n1672,n1670,n1607);
or (n1673,n1674,n1676);
and (n1674,n1675,n1607);
xor (n1675,n1586,n1587);
and (n1676,n1677,n1678);
xor (n1677,n1675,n1607);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1591,n1592);
and (n1681,n1194,n1608);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1597,n1598);
and (n1687,n1202,n1608);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
and (n1690,n1691,n1692);
xor (n1691,n1603,n1604);
and (n1692,n1209,n1608);
and (n1693,n917,n1694);
xor (n1694,n1695,n823);
xor (n1695,n1696,n1759);
xor (n1696,n1697,n1758);
xor (n1697,n1698,n1755);
xor (n1698,n1699,n1754);
xor (n1699,n1700,n1751);
xor (n1700,n1701,n1750);
xor (n1701,n1702,n1747);
xor (n1702,n1703,n1746);
xor (n1703,n1704,n1743);
xor (n1704,n1705,n1742);
xor (n1705,n1706,n1739);
xor (n1706,n1707,n1738);
xor (n1707,n1708,n1735);
xor (n1708,n1709,n1734);
xor (n1709,n1710,n1731);
xor (n1710,n1711,n1730);
xor (n1711,n1712,n1727);
xor (n1712,n1713,n1726);
xor (n1713,n1714,n1723);
xor (n1714,n1715,n1722);
xor (n1715,n1716,n1719);
xor (n1716,n1717,n1718);
and (n1717,n397,n351);
and (n1718,n388,n97);
or (n1719,n1720,n1721);
and (n1720,n1629,n1630);
and (n1721,n1628,n1631);
and (n1722,n106,n87);
or (n1723,n1724,n1725);
and (n1724,n1627,n1634);
and (n1725,n1626,n1635);
and (n1726,n31,n17);
or (n1727,n1728,n1729);
and (n1728,n1625,n1638);
and (n1729,n1624,n1639);
and (n1730,n323,n136);
or (n1731,n1732,n1733);
and (n1732,n1623,n1642);
and (n1733,n1622,n1643);
and (n1734,n149,n119);
or (n1735,n1736,n1737);
and (n1736,n1621,n1646);
and (n1737,n1620,n1647);
and (n1738,n125,n195);
or (n1739,n1740,n1741);
and (n1740,n1619,n1650);
and (n1741,n1618,n1651);
and (n1742,n210,n204);
or (n1743,n1744,n1745);
and (n1744,n1617,n1654);
and (n1745,n1616,n1655);
and (n1746,n220,n261);
or (n1747,n1748,n1749);
and (n1748,n1615,n1658);
and (n1749,n1614,n1659);
and (n1750,n270,n176);
or (n1751,n1752,n1753);
and (n1752,n1613,n1662);
and (n1753,n1612,n1663);
and (n1754,n279,n166);
or (n1755,n1756,n1757);
and (n1756,n1611,n1666);
and (n1757,n1610,n1667);
and (n1758,n248,n181);
and (n1759,n1609,n237);
or (n1760,n1761,n1763);
and (n1761,n1762,n1693);
xor (n1762,n1672,n1673);
and (n1763,n1764,n1765);
xor (n1764,n1762,n1693);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1677,n1678);
and (n1768,n1194,n1694);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1683,n1684);
and (n1774,n1202,n1694);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
and (n1777,n1778,n1779);
xor (n1778,n1689,n1690);
and (n1779,n1209,n1694);
and (n1780,n917,n1781);
xor (n1781,n1782,n1853);
xor (n1782,n1783,n1852);
xor (n1783,n1784,n1851);
xor (n1784,n1785,n1848);
xor (n1785,n1786,n1847);
xor (n1786,n1787,n1844);
xor (n1787,n1788,n1843);
xor (n1788,n1789,n1840);
xor (n1789,n1790,n1839);
xor (n1790,n1791,n1836);
xor (n1791,n1792,n1835);
xor (n1792,n1793,n1832);
xor (n1793,n1794,n1831);
xor (n1794,n1795,n1828);
xor (n1795,n1796,n1827);
xor (n1796,n1797,n1824);
xor (n1797,n1798,n1823);
xor (n1798,n1799,n1820);
xor (n1799,n1800,n1819);
xor (n1800,n1801,n1816);
xor (n1801,n1802,n1815);
xor (n1802,n1803,n1812);
xor (n1803,n1804,n1811);
xor (n1804,n1805,n1808);
xor (n1805,n1806,n1807);
and (n1806,n889,n351);
and (n1807,n397,n97);
or (n1808,n1809,n1810);
and (n1809,n1717,n1718);
and (n1810,n1716,n1719);
and (n1811,n388,n87);
or (n1812,n1813,n1814);
and (n1813,n1715,n1722);
and (n1814,n1714,n1723);
and (n1815,n106,n17);
or (n1816,n1817,n1818);
and (n1817,n1713,n1726);
and (n1818,n1712,n1727);
and (n1819,n31,n136);
or (n1820,n1821,n1822);
and (n1821,n1711,n1730);
and (n1822,n1710,n1731);
and (n1823,n323,n119);
or (n1824,n1825,n1826);
and (n1825,n1709,n1734);
and (n1826,n1708,n1735);
and (n1827,n149,n195);
or (n1828,n1829,n1830);
and (n1829,n1707,n1738);
and (n1830,n1706,n1739);
and (n1831,n125,n204);
or (n1832,n1833,n1834);
and (n1833,n1705,n1742);
and (n1834,n1704,n1743);
and (n1835,n210,n261);
or (n1836,n1837,n1838);
and (n1837,n1703,n1746);
and (n1838,n1702,n1747);
and (n1839,n220,n176);
or (n1840,n1841,n1842);
and (n1841,n1701,n1750);
and (n1842,n1700,n1751);
and (n1843,n270,n166);
or (n1844,n1845,n1846);
and (n1845,n1699,n1754);
and (n1846,n1698,n1755);
and (n1847,n279,n181);
or (n1848,n1849,n1850);
and (n1849,n1697,n1758);
and (n1850,n1696,n1759);
and (n1851,n248,n408);
and (n1852,n1695,n823);
and (n1853,n160,n826);
and (n1854,n1855,n1856);
xor (n1855,n1031,n1780);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n1764,n1765);
and (n1859,n1194,n1781);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1770,n1771);
and (n1865,n1202,n1781);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
and (n1868,n1869,n1870);
xor (n1869,n1776,n1777);
and (n1870,n1209,n1781);
endmodule
