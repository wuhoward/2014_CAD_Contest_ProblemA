module top (out,n3,n7,n9,n10,n12,n14,n15,n35,n36
        ,n44,n45,n47,n48,n65,n66,n68,n77,n78,n87
        ,n98,n99,n106,n112,n125,n134,n139,n157,n201);
output out;
input n3;
input n7;
input n9;
input n10;
input n12;
input n14;
input n15;
input n35;
input n36;
input n44;
input n45;
input n47;
input n48;
input n65;
input n66;
input n68;
input n77;
input n78;
input n87;
input n98;
input n99;
input n106;
input n112;
input n125;
input n134;
input n139;
input n157;
input n201;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n8;
wire n11;
wire n13;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n46;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
xor (out,n0,n395);
nand (n0,n1,n16);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
xor (n5,n6,n11);
and (n6,n7,n8);
wire s0n8,s1n8,notn8;
or (n8,s0n8,s1n8);
not(notn8,n3);
and (s0n8,notn8,n9);
and (s1n8,n3,n10);
and (n11,n12,n13);
wire s0n13,s1n13,notn13;
or (n13,s0n13,s1n13);
not(notn13,n3);
and (s0n13,notn13,n14);
and (s1n13,n3,n15);
nand (n16,n17,n2);
nand (n17,n18,n394);
or (n18,n19,n225);
not (n19,n20);
or (n20,n21,n224);
and (n21,n22,n181);
or (n22,n23,n180);
and (n23,n24,n149);
xor (n24,n25,n116);
or (n25,n26,n115);
and (n26,n27,n90);
xor (n27,n28,n59);
nand (n28,n29,n54);
or (n29,n30,n39);
not (n30,n31);
nand (n31,n32,n37);
or (n32,n33,n12);
not (n33,n34);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n3);
and (s0n34,notn34,n35);
and (s1n34,n3,n36);
or (n37,n34,n38);
not (n38,n12);
nand (n39,n40,n51);
nor (n40,n41,n49);
and (n41,n42,n46);
not (n42,n43);
wire s0n43,s1n43,notn43;
or (n43,s0n43,s1n43);
not(notn43,n3);
and (s0n43,notn43,n44);
and (s1n43,n3,n45);
wire s0n46,s1n46,notn46;
or (n46,s0n46,s1n46);
not(notn46,n3);
and (s0n46,notn46,n47);
and (s1n46,n3,n48);
and (n49,n43,n50);
not (n50,n46);
nand (n51,n52,n53);
or (n52,n42,n34);
nand (n53,n34,n42);
or (n54,n40,n55);
nor (n55,n56,n57);
and (n56,n7,n33);
and (n57,n58,n34);
not (n58,n7);
nand (n59,n60,n84);
or (n60,n61,n71);
not (n61,n62);
nand (n62,n63,n69);
or (n63,n64,n67);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n3);
and (s0n64,notn64,n65);
and (s1n64,n3,n66);
not (n67,n68);
or (n69,n70,n68);
not (n70,n64);
not (n71,n72);
and (n72,n73,n80);
nand (n73,n74,n79);
or (n74,n75,n64);
not (n75,n76);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n3);
and (s0n76,notn76,n77);
and (s1n76,n3,n78);
nand (n79,n64,n75);
not (n80,n81);
nand (n81,n82,n83);
or (n82,n75,n13);
nand (n83,n13,n75);
nand (n84,n81,n85);
nor (n85,n86,n88);
and (n86,n87,n64);
and (n88,n89,n70);
not (n89,n87);
nand (n90,n91,n109);
or (n91,n92,n104);
nand (n92,n93,n101);
not (n93,n94);
nand (n94,n95,n100);
or (n95,n96,n64);
not (n96,n97);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n3);
and (s0n97,notn97,n98);
and (s1n97,n3,n99);
nand (n100,n64,n96);
nand (n101,n102,n103);
or (n102,n96,n46);
nand (n103,n46,n96);
nor (n104,n105,n107);
and (n105,n50,n106);
and (n107,n46,n108);
not (n108,n106);
or (n109,n93,n110);
nor (n110,n111,n113);
and (n111,n50,n112);
and (n113,n46,n114);
not (n114,n112);
and (n115,n28,n59);
xor (n116,n117,n143);
xor (n117,n118,n126);
and (n118,n119,n12);
not (n119,n120);
nand (n120,n34,n121);
not (n121,n122);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n3);
and (s0n122,notn122,1'b0);
and (s1n122,n3,n124);
and (n124,n125,n36);
nand (n126,n127,n136);
or (n127,n128,n131);
not (n128,n129);
nor (n129,n130,n8);
not (n130,n13);
nor (n131,n132,n135);
and (n132,n133,n13);
not (n133,n134);
and (n135,n134,n130);
or (n136,n137,n142);
nor (n137,n138,n140);
and (n138,n130,n139);
and (n140,n13,n141);
not (n141,n139);
not (n142,n8);
nand (n143,n144,n145);
or (n144,n39,n55);
or (n145,n40,n146);
nor (n146,n147,n148);
and (n147,n106,n33);
and (n148,n108,n34);
xor (n149,n150,n166);
xor (n150,n151,n160);
nand (n151,n152,n154);
or (n152,n71,n153);
not (n153,n85);
or (n154,n80,n155);
nor (n155,n156,n158);
and (n156,n70,n157);
and (n158,n64,n159);
not (n159,n157);
nand (n160,n161,n162);
or (n161,n92,n110);
or (n162,n93,n163);
nor (n163,n164,n165);
and (n164,n50,n68);
and (n165,n46,n67);
and (n166,n167,n172);
nor (n167,n168,n33);
nor (n168,n169,n171);
and (n169,n50,n170);
nand (n170,n43,n12);
and (n171,n42,n38);
nand (n172,n173,n178);
or (n173,n174,n128);
not (n174,n175);
nor (n175,n176,n177);
and (n176,n157,n13);
and (n177,n159,n130);
nand (n178,n179,n8);
not (n179,n131);
and (n180,n25,n116);
xor (n181,n182,n207);
xor (n182,n183,n204);
xor (n183,n184,n196);
xor (n184,n185,n192);
nand (n185,n186,n187);
or (n186,n146,n39);
nand (n187,n188,n191);
nor (n188,n189,n190);
and (n189,n112,n34);
and (n190,n114,n33);
not (n191,n40);
nor (n192,n120,n193);
nor (n193,n194,n195);
and (n194,n122,n58);
and (n195,n121,n7);
nand (n196,n197,n198);
or (n197,n128,n137);
or (n198,n199,n142);
nor (n199,n200,n202);
and (n200,n130,n201);
and (n202,n13,n203);
not (n203,n201);
or (n204,n205,n206);
and (n205,n150,n166);
and (n206,n151,n160);
xor (n207,n208,n221);
xor (n208,n209,n215);
nand (n209,n210,n211);
or (n210,n92,n163);
or (n211,n93,n212);
nor (n212,n213,n214);
and (n213,n50,n87);
and (n214,n46,n89);
nand (n215,n216,n217);
or (n216,n71,n155);
or (n217,n218,n80);
nor (n218,n219,n220);
and (n219,n70,n134);
and (n220,n64,n133);
or (n221,n222,n223);
and (n222,n117,n143);
and (n223,n118,n126);
nor (n224,n22,n181);
not (n225,n226);
nand (n226,n227,n393);
or (n227,n228,n388);
nor (n228,n229,n386);
and (n229,n230,n375);
or (n230,n231,n374);
and (n231,n232,n290);
xor (n232,n233,n273);
or (n233,n234,n272);
and (n234,n235,n257);
xor (n235,n236,n246);
nand (n236,n237,n242);
or (n237,n238,n71);
not (n238,n239);
nor (n239,n240,n241);
and (n240,n108,n70);
and (n241,n106,n64);
nand (n242,n81,n243);
nor (n243,n244,n245);
and (n244,n112,n64);
and (n245,n70,n114);
nand (n246,n247,n252);
or (n247,n248,n93);
not (n248,n249);
nor (n249,n250,n251);
and (n250,n7,n46);
and (n251,n58,n50);
nand (n252,n253,n254);
not (n253,n92);
nand (n254,n255,n256);
or (n255,n50,n12);
or (n256,n46,n38);
xor (n257,n258,n263);
and (n258,n259,n46);
nand (n259,n260,n262);
or (n260,n64,n261);
and (n261,n12,n97);
or (n262,n97,n12);
nand (n263,n264,n268);
or (n264,n128,n265);
nor (n265,n266,n267);
and (n266,n130,n68);
and (n267,n13,n67);
or (n268,n269,n142);
nor (n269,n270,n271);
and (n270,n87,n130);
and (n271,n89,n13);
and (n272,n236,n246);
xor (n273,n274,n279);
xor (n274,n275,n278);
nand (n275,n276,n277);
or (n276,n248,n92);
or (n277,n93,n104);
and (n278,n258,n263);
xor (n279,n280,n286);
xor (n280,n281,n282);
and (n281,n191,n12);
nand (n282,n283,n284);
or (n283,n142,n174);
nand (n284,n285,n129);
not (n285,n269);
nand (n286,n287,n289);
or (n287,n288,n71);
not (n288,n243);
nand (n289,n81,n62);
or (n290,n291,n373);
and (n291,n292,n313);
xor (n292,n293,n312);
or (n293,n294,n311);
and (n294,n295,n304);
xor (n295,n296,n297);
and (n296,n94,n12);
nand (n297,n298,n303);
or (n298,n299,n71);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n7,n64);
and (n302,n58,n70);
nand (n303,n239,n81);
nand (n304,n305,n310);
or (n305,n128,n306);
not (n306,n307);
nor (n307,n308,n309);
and (n308,n114,n130);
and (n309,n112,n13);
or (n310,n265,n142);
and (n311,n296,n297);
xor (n312,n235,n257);
or (n313,n314,n372);
and (n314,n315,n371);
xor (n315,n316,n330);
nor (n316,n317,n325);
not (n317,n318);
nand (n318,n319,n324);
or (n319,n320,n128);
not (n320,n321);
nand (n321,n322,n323);
or (n322,n108,n13);
nand (n323,n13,n108);
nand (n324,n307,n8);
nand (n325,n326,n64);
nand (n326,n327,n329);
or (n327,n13,n328);
and (n328,n12,n76);
or (n329,n76,n12);
nand (n330,n331,n369);
or (n331,n332,n355);
not (n332,n333);
nand (n333,n334,n354);
or (n334,n335,n344);
nor (n335,n336,n343);
nand (n336,n337,n342);
or (n337,n338,n128);
not (n338,n339);
nand (n339,n340,n341);
or (n340,n58,n13);
nand (n341,n13,n58);
nand (n342,n321,n8);
nor (n343,n80,n38);
nand (n344,n345,n352);
nand (n345,n346,n351);
or (n346,n347,n128);
not (n347,n348);
nand (n348,n349,n350);
or (n349,n130,n12);
or (n350,n13,n38);
nand (n351,n339,n8);
nor (n352,n353,n130);
and (n353,n12,n8);
nand (n354,n336,n343);
not (n355,n356);
nand (n356,n357,n365);
not (n357,n358);
nand (n358,n359,n364);
or (n359,n360,n71);
not (n360,n361);
nand (n361,n362,n363);
or (n362,n70,n12);
or (n363,n64,n38);
nand (n364,n81,n300);
nor (n365,n366,n368);
and (n366,n317,n367);
not (n367,n325);
and (n368,n318,n325);
nand (n369,n370,n358);
not (n370,n365);
xor (n371,n295,n304);
and (n372,n316,n330);
and (n373,n293,n312);
and (n374,n233,n273);
or (n375,n376,n383);
xor (n376,n377,n382);
xor (n377,n378,n379);
xor (n378,n167,n172);
or (n379,n380,n381);
and (n380,n280,n286);
and (n381,n281,n282);
xor (n382,n27,n90);
or (n383,n384,n385);
and (n384,n274,n279);
and (n385,n275,n278);
not (n386,n387);
nand (n387,n376,n383);
nor (n388,n389,n390);
xor (n389,n24,n149);
or (n390,n391,n392);
and (n391,n377,n382);
and (n392,n378,n379);
nand (n393,n389,n390);
or (n394,n226,n20);
wire s0n395,s1n395,notn395;
or (n395,s0n395,s1n395);
not(notn395,n3);
and (s0n395,notn395,n396);
and (s1n395,n3,n5);
xor (n396,n397,n602);
xor (n397,n398,n600);
xor (n398,n399,n599);
xor (n399,n400,n590);
xor (n400,n401,n589);
xor (n401,n402,n574);
xor (n402,n403,n573);
xor (n403,n404,n553);
xor (n404,n405,n552);
xor (n405,n406,n526);
xor (n406,n407,n525);
xor (n407,n408,n496);
xor (n408,n409,n495);
xor (n409,n410,n457);
xor (n410,n411,n456);
xor (n411,n412,n415);
xor (n412,n413,n414);
and (n413,n201,n8);
and (n414,n139,n13);
or (n415,n416,n419);
and (n416,n417,n418);
and (n417,n139,n8);
and (n418,n134,n13);
and (n419,n420,n421);
xor (n420,n417,n418);
or (n421,n422,n424);
and (n422,n423,n176);
and (n423,n134,n8);
and (n424,n425,n426);
xor (n425,n423,n176);
or (n426,n427,n430);
and (n427,n428,n429);
and (n428,n157,n8);
and (n429,n87,n13);
and (n430,n431,n432);
xor (n431,n428,n429);
or (n432,n433,n436);
and (n433,n434,n435);
and (n434,n87,n8);
and (n435,n68,n13);
and (n436,n437,n438);
xor (n437,n434,n435);
or (n438,n439,n441);
and (n439,n440,n309);
and (n440,n68,n8);
and (n441,n442,n443);
xor (n442,n440,n309);
or (n443,n444,n447);
and (n444,n445,n446);
and (n445,n112,n8);
and (n446,n106,n13);
and (n447,n448,n449);
xor (n448,n445,n446);
or (n449,n450,n453);
and (n450,n451,n452);
and (n451,n106,n8);
and (n452,n7,n13);
and (n453,n454,n455);
xor (n454,n451,n452);
and (n455,n6,n11);
and (n456,n134,n76);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n420,n421);
and (n460,n157,n76);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n425,n426);
and (n466,n87,n76);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n431,n432);
and (n472,n68,n76);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n437,n438);
and (n478,n112,n76);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n442,n443);
and (n484,n106,n76);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n448,n449);
and (n490,n7,n76);
and (n491,n492,n493);
xor (n492,n489,n490);
and (n493,n494,n328);
xor (n494,n454,n455);
and (n495,n157,n64);
or (n496,n497,n499);
and (n497,n498,n86);
xor (n498,n462,n463);
and (n499,n500,n501);
xor (n500,n498,n86);
or (n501,n502,n505);
and (n502,n503,n504);
xor (n503,n468,n469);
and (n504,n68,n64);
and (n505,n506,n507);
xor (n506,n503,n504);
or (n507,n508,n510);
and (n508,n509,n244);
xor (n509,n474,n475);
and (n510,n511,n512);
xor (n511,n509,n244);
or (n512,n513,n515);
and (n513,n514,n241);
xor (n514,n480,n481);
and (n515,n516,n517);
xor (n516,n514,n241);
or (n517,n518,n520);
and (n518,n519,n301);
xor (n519,n486,n487);
and (n520,n521,n522);
xor (n521,n519,n301);
and (n522,n523,n524);
xor (n523,n492,n493);
and (n524,n12,n64);
and (n525,n87,n97);
or (n526,n527,n530);
and (n527,n528,n529);
xor (n528,n500,n501);
and (n529,n68,n97);
and (n530,n531,n532);
xor (n531,n528,n529);
or (n532,n533,n536);
and (n533,n534,n535);
xor (n534,n506,n507);
and (n535,n112,n97);
and (n536,n537,n538);
xor (n537,n534,n535);
or (n538,n539,n542);
and (n539,n540,n541);
xor (n540,n511,n512);
and (n541,n106,n97);
and (n542,n543,n544);
xor (n543,n540,n541);
or (n544,n545,n548);
and (n545,n546,n547);
xor (n546,n516,n517);
and (n547,n7,n97);
and (n548,n549,n550);
xor (n549,n546,n547);
and (n550,n551,n261);
xor (n551,n521,n522);
and (n552,n68,n46);
or (n553,n554,n557);
and (n554,n555,n556);
xor (n555,n531,n532);
and (n556,n112,n46);
and (n557,n558,n559);
xor (n558,n555,n556);
or (n559,n560,n563);
and (n560,n561,n562);
xor (n561,n537,n538);
and (n562,n106,n46);
and (n563,n564,n565);
xor (n564,n561,n562);
or (n565,n566,n568);
and (n566,n567,n250);
xor (n567,n543,n544);
and (n568,n569,n570);
xor (n569,n567,n250);
and (n570,n571,n572);
xor (n571,n549,n550);
and (n572,n12,n46);
and (n573,n112,n43);
or (n574,n575,n578);
and (n575,n576,n577);
xor (n576,n558,n559);
and (n577,n106,n43);
and (n578,n579,n580);
xor (n579,n576,n577);
or (n580,n581,n584);
and (n581,n582,n583);
xor (n582,n564,n565);
and (n583,n7,n43);
and (n584,n585,n586);
xor (n585,n582,n583);
and (n586,n587,n588);
xor (n587,n569,n570);
not (n588,n170);
and (n589,n106,n34);
or (n590,n591,n594);
and (n591,n592,n593);
xor (n592,n579,n580);
and (n593,n7,n34);
and (n594,n595,n596);
xor (n595,n592,n593);
and (n596,n597,n598);
xor (n597,n585,n586);
and (n598,n12,n34);
and (n599,n7,n122);
and (n600,n601,n602);
xor (n601,n595,n596);
and (n602,n12,n122);
endmodule
