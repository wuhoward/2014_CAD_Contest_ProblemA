module top (out,n3,n4,n5,n22,n24,n32,n34,n43,n51
        ,n52,n57,n61,n70,n71,n77,n81,n87,n97,n109
        ,n120,n131,n143,n154,n181,n200);
output out;
input n3;
input n4;
input n5;
input n22;
input n24;
input n32;
input n34;
input n43;
input n51;
input n52;
input n57;
input n61;
input n70;
input n71;
input n77;
input n81;
input n87;
input n97;
input n109;
input n120;
input n131;
input n143;
input n154;
input n181;
input n200;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
xnor (out,n0,n466);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n463);
nand (n7,n8,n462);
or (n8,n9,n254);
not (n9,n10);
nor (n10,n11,n253);
not (n11,n12);
nand (n12,n13,n216);
xor (n13,n14,n169);
xor (n14,n15,n90);
xor (n15,n16,n64);
xor (n16,n17,n46);
nand (n17,n18,n39);
or (n18,n19,n27);
not (n19,n20);
nand (n20,n21,n25);
or (n21,n22,n23);
not (n23,n24);
or (n25,n26,n24);
not (n26,n22);
not (n27,n28);
and (n28,n29,n36);
not (n29,n30);
nand (n30,n31,n35);
or (n31,n32,n33);
not (n33,n34);
nand (n35,n32,n33);
nand (n36,n37,n38);
or (n37,n32,n26);
nand (n38,n26,n32);
nand (n39,n40,n30);
not (n40,n41);
nor (n41,n42,n44);
and (n42,n26,n43);
and (n44,n22,n45);
not (n45,n43);
nand (n46,n47,n58);
or (n47,n48,n55);
nor (n48,n49,n53);
and (n49,n50,n52);
not (n50,n51);
and (n53,n51,n54);
not (n54,n52);
nand (n55,n51,n56);
not (n56,n57);
or (n58,n59,n56);
nor (n59,n60,n62);
and (n60,n50,n61);
and (n62,n51,n63);
not (n63,n61);
nand (n64,n65,n84);
or (n65,n66,n79);
nand (n66,n67,n74);
nor (n67,n68,n72);
and (n68,n69,n71);
not (n69,n70);
and (n72,n70,n73);
not (n73,n71);
nand (n74,n75,n78);
or (n75,n71,n76);
not (n76,n77);
nand (n78,n76,n71);
nor (n79,n80,n82);
and (n80,n76,n81);
and (n82,n77,n83);
not (n83,n81);
or (n84,n67,n85);
nor (n85,n86,n88);
and (n86,n76,n87);
and (n88,n77,n89);
not (n89,n87);
or (n90,n91,n168);
and (n91,n92,n133);
xor (n92,n93,n101);
nand (n93,n94,n100);
or (n94,n66,n95);
nor (n95,n96,n98);
and (n96,n76,n97);
and (n98,n77,n99);
not (n99,n97);
or (n100,n79,n67);
xor (n101,n102,n110);
and (n102,n103,n22);
nand (n103,n104,n105);
or (n104,n34,n32);
nand (n105,n106,n108);
or (n106,n107,n33);
not (n107,n32);
not (n108,n109);
nand (n110,n111,n126);
or (n111,n112,n116);
not (n112,n113);
nand (n113,n114,n115);
or (n114,n70,n89);
or (n115,n69,n87);
not (n116,n117);
nor (n117,n118,n122);
nand (n118,n119,n121);
or (n119,n50,n120);
nand (n121,n50,n120);
nor (n122,n123,n124);
and (n123,n69,n120);
and (n124,n70,n125);
not (n125,n120);
or (n126,n127,n128);
not (n127,n118);
nor (n128,n129,n132);
and (n129,n130,n70);
not (n130,n131);
and (n132,n131,n69);
or (n133,n134,n167);
and (n134,n135,n149);
xor (n135,n136,n137);
and (n136,n30,n109);
nand (n137,n138,n145);
or (n138,n56,n139);
not (n139,n140);
nor (n140,n141,n144);
and (n141,n142,n50);
not (n142,n143);
and (n144,n51,n143);
or (n145,n146,n55);
nor (n146,n147,n148);
and (n147,n50,n131);
and (n148,n51,n130);
nand (n149,n150,n163);
or (n150,n151,n160);
nand (n151,n152,n156);
nand (n152,n153,n155);
or (n153,n154,n33);
nand (n155,n33,n154);
not (n156,n157);
nand (n157,n158,n159);
or (n158,n76,n154);
nand (n159,n76,n154);
nor (n160,n161,n162);
and (n161,n33,n24);
and (n162,n34,n23);
or (n163,n156,n164);
nor (n164,n165,n166);
and (n165,n45,n34);
and (n166,n43,n33);
and (n167,n136,n137);
and (n168,n93,n101);
xor (n169,n170,n195);
xor (n170,n171,n172);
and (n171,n102,n110);
or (n172,n173,n194);
and (n173,n174,n191);
xor (n174,n175,n184);
nand (n175,n176,n183);
or (n176,n156,n177);
not (n177,n178);
nand (n178,n179,n182);
or (n179,n34,n180);
not (n180,n181);
or (n182,n33,n181);
or (n183,n164,n151);
nand (n184,n185,n190);
or (n185,n186,n27);
not (n186,n187);
nand (n187,n188,n189);
or (n188,n22,n108);
or (n189,n26,n109);
nand (n190,n20,n30);
nand (n191,n192,n193);
or (n192,n139,n55);
or (n193,n48,n56);
and (n194,n175,n184);
xor (n195,n196,n209);
xor (n196,n197,n203);
nor (n197,n198,n108);
nor (n198,n199,n201);
and (n199,n26,n200);
and (n201,n22,n202);
not (n202,n200);
nand (n203,n204,n205);
or (n204,n128,n116);
nand (n205,n206,n118);
nand (n206,n207,n208);
or (n207,n70,n142);
or (n208,n69,n143);
nand (n209,n210,n211);
or (n210,n177,n151);
nand (n211,n212,n157);
not (n212,n213);
nor (n213,n214,n215);
and (n214,n33,n97);
and (n215,n34,n99);
or (n216,n217,n252);
and (n217,n218,n251);
xor (n218,n219,n220);
xor (n219,n174,n191);
or (n220,n221,n250);
and (n221,n222,n236);
xor (n222,n223,n230);
nand (n223,n224,n229);
or (n224,n225,n116);
not (n225,n226);
nand (n226,n227,n228);
or (n227,n70,n83);
or (n228,n69,n81);
nand (n229,n118,n113);
nand (n230,n231,n235);
or (n231,n66,n232);
nor (n232,n233,n234);
and (n233,n181,n76);
and (n234,n77,n180);
or (n235,n67,n95);
and (n236,n237,n243);
nor (n237,n238,n33);
nor (n238,n239,n241);
and (n239,n240,n108);
nand (n240,n77,n154);
and (n241,n76,n242);
not (n242,n154);
nand (n243,n244,n249);
or (n244,n55,n245);
not (n245,n246);
nor (n246,n247,n248);
and (n247,n51,n87);
and (n248,n89,n50);
or (n249,n146,n56);
and (n250,n223,n230);
xor (n251,n92,n133);
and (n252,n219,n220);
nor (n253,n13,n216);
not (n254,n255);
nor (n255,n256,n454);
and (n256,n257,n437);
or (n257,n258,n436);
and (n258,n259,n327);
xor (n259,n260,n307);
or (n260,n261,n306);
and (n261,n262,n289);
xor (n262,n263,n272);
nand (n263,n264,n268);
or (n264,n66,n265);
nor (n265,n266,n267);
and (n266,n76,n24);
and (n267,n77,n23);
or (n268,n67,n269);
nor (n269,n270,n271);
and (n270,n76,n43);
and (n271,n77,n45);
and (n272,n273,n283);
nand (n273,n274,n279);
or (n274,n55,n275);
not (n275,n276);
nor (n276,n277,n278);
and (n277,n51,n97);
and (n278,n99,n50);
nand (n279,n280,n57);
nand (n280,n281,n282);
or (n281,n81,n50);
nand (n282,n50,n81);
not (n283,n284);
nand (n284,n285,n77);
nand (n285,n286,n287);
or (n286,n70,n71);
nand (n287,n288,n108);
or (n288,n73,n69);
xor (n289,n290,n296);
xor (n290,n291,n292);
and (n291,n157,n109);
nand (n292,n293,n294);
or (n293,n56,n245);
or (n294,n295,n55);
not (n295,n280);
nand (n296,n297,n302);
or (n297,n298,n116);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n70,n181);
and (n301,n180,n69);
nand (n302,n118,n303);
nand (n303,n304,n305);
or (n304,n70,n99);
or (n305,n69,n97);
and (n306,n263,n272);
xor (n307,n308,n313);
xor (n308,n309,n310);
xor (n309,n237,n243);
or (n310,n311,n312);
and (n311,n290,n296);
and (n312,n291,n292);
xor (n313,n314,n324);
xor (n314,n315,n321);
nand (n315,n316,n320);
or (n316,n151,n317);
nor (n317,n318,n319);
and (n318,n33,n109);
and (n319,n34,n108);
or (n320,n160,n156);
nand (n321,n322,n323);
or (n322,n225,n127);
nand (n323,n117,n303);
nand (n324,n325,n326);
or (n325,n66,n269);
or (n326,n67,n232);
or (n327,n328,n435);
and (n328,n329,n353);
xor (n329,n330,n352);
or (n330,n331,n351);
and (n331,n332,n347);
xor (n332,n333,n340);
nand (n333,n334,n339);
or (n334,n335,n116);
not (n335,n336);
nand (n336,n337,n338);
or (n337,n70,n45);
or (n338,n69,n43);
nand (n339,n118,n299);
nand (n340,n341,n346);
or (n341,n342,n66);
not (n342,n343);
nand (n343,n344,n345);
or (n344,n108,n77);
or (n345,n76,n109);
or (n346,n67,n265);
nand (n347,n348,n350);
or (n348,n283,n349);
not (n349,n273);
or (n350,n273,n284);
and (n351,n333,n340);
xor (n352,n262,n289);
or (n353,n354,n434);
and (n354,n355,n376);
xor (n355,n356,n375);
or (n356,n357,n374);
and (n357,n358,n367);
xor (n358,n359,n360);
nor (n359,n67,n108);
nand (n360,n361,n366);
or (n361,n362,n116);
not (n362,n363);
nor (n363,n364,n365);
and (n364,n23,n69);
and (n365,n70,n24);
nand (n366,n118,n336);
nand (n367,n368,n373);
or (n368,n55,n369);
not (n369,n370);
nor (n370,n371,n372);
and (n371,n180,n50);
and (n372,n51,n181);
or (n373,n275,n56);
and (n374,n359,n360);
xor (n375,n332,n347);
or (n376,n377,n433);
and (n377,n378,n432);
xor (n378,n379,n393);
nor (n379,n380,n388);
not (n380,n381);
nand (n381,n382,n383);
or (n382,n56,n369);
nand (n383,n384,n387);
nor (n384,n385,n386);
and (n385,n45,n50);
and (n386,n51,n43);
not (n387,n55);
nand (n388,n389,n70);
nand (n389,n390,n391);
or (n390,n120,n51);
or (n391,n392,n109);
and (n392,n51,n120);
nand (n393,n394,n431);
or (n394,n395,n419);
not (n395,n396);
nand (n396,n397,n418);
or (n397,n398,n407);
nor (n398,n399,n400);
and (n399,n118,n109);
nand (n400,n401,n403);
or (n401,n56,n402);
not (n402,n384);
nand (n403,n404,n387);
nand (n404,n405,n406);
or (n405,n23,n51);
or (n406,n50,n24);
nand (n407,n408,n411);
not (n408,n409);
nand (n409,n410,n51);
nand (n410,n109,n57);
nand (n411,n412,n414);
or (n412,n56,n413);
not (n413,n404);
nand (n414,n415,n387);
nor (n415,n416,n417);
and (n416,n108,n50);
and (n417,n51,n109);
nand (n418,n399,n400);
not (n419,n420);
nand (n420,n421,n425);
nor (n421,n422,n423);
and (n422,n388,n381);
and (n423,n424,n380);
not (n424,n388);
nor (n425,n426,n430);
and (n426,n117,n427);
nand (n427,n428,n429);
or (n428,n70,n108);
or (n429,n69,n109);
and (n430,n118,n363);
or (n431,n421,n425);
xor (n432,n358,n367);
and (n433,n379,n393);
and (n434,n356,n375);
and (n435,n330,n352);
and (n436,n260,n307);
nor (n437,n438,n449);
nor (n438,n439,n440);
xor (n439,n218,n251);
or (n440,n441,n448);
and (n441,n442,n447);
xor (n442,n443,n446);
or (n443,n444,n445);
and (n444,n314,n324);
and (n445,n315,n321);
xor (n446,n135,n149);
xor (n447,n222,n236);
and (n448,n443,n446);
nor (n449,n450,n451);
xor (n450,n442,n447);
or (n451,n452,n453);
and (n452,n308,n313);
and (n453,n309,n310);
not (n454,n455);
nand (n455,n456,n461);
or (n456,n457,n459);
not (n457,n458);
nand (n458,n450,n451);
not (n459,n460);
nand (n460,n439,n440);
not (n461,n438);
or (n462,n255,n10);
not (n463,n464);
nand (n464,n465,n3);
not (n465,n4);
wire s0n466,s1n466,notn466;
or (n466,s0n466,s1n466);
not(notn466,n4);
and (s0n466,notn466,n467);
and (s1n466,n4,1'b0);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n3);
and (s0n467,notn467,n5);
and (s1n467,n3,n468);
xor (n468,n469,n732);
xor (n469,n470,n729);
xor (n470,n471,n728);
xor (n471,n472,n720);
xor (n472,n473,n719);
xor (n473,n474,n704);
xor (n474,n475,n703);
xor (n475,n476,n683);
xor (n476,n477,n682);
xor (n477,n478,n655);
xor (n478,n479,n654);
xor (n479,n480,n622);
xor (n480,n481,n621);
xor (n481,n482,n584);
xor (n482,n483,n583);
xor (n483,n484,n539);
xor (n484,n485,n538);
xor (n485,n486,n489);
xor (n486,n487,n488);
and (n487,n200,n109);
and (n488,n22,n24);
or (n489,n490,n493);
and (n490,n491,n492);
and (n491,n22,n109);
and (n492,n32,n24);
and (n493,n494,n495);
xor (n494,n491,n492);
or (n495,n496,n499);
and (n496,n497,n498);
and (n497,n32,n109);
and (n498,n34,n24);
and (n499,n500,n501);
xor (n500,n497,n498);
or (n501,n502,n505);
and (n502,n503,n504);
and (n503,n34,n109);
and (n504,n154,n24);
and (n505,n506,n507);
xor (n506,n503,n504);
or (n507,n508,n511);
and (n508,n509,n510);
and (n509,n154,n109);
and (n510,n77,n24);
and (n511,n512,n513);
xor (n512,n509,n510);
or (n513,n514,n517);
and (n514,n515,n516);
and (n515,n77,n109);
and (n516,n71,n24);
and (n517,n518,n519);
xor (n518,n515,n516);
or (n519,n520,n522);
and (n520,n521,n365);
and (n521,n71,n109);
and (n522,n523,n524);
xor (n523,n521,n365);
or (n524,n525,n528);
and (n525,n526,n527);
and (n526,n70,n109);
and (n527,n120,n24);
and (n528,n529,n530);
xor (n529,n526,n527);
or (n530,n531,n534);
and (n531,n532,n533);
and (n532,n120,n109);
and (n533,n51,n24);
and (n534,n535,n536);
xor (n535,n532,n533);
and (n536,n417,n537);
and (n537,n57,n24);
and (n538,n32,n43);
or (n539,n540,n543);
and (n540,n541,n542);
xor (n541,n494,n495);
and (n542,n34,n43);
and (n543,n544,n545);
xor (n544,n541,n542);
or (n545,n546,n549);
and (n546,n547,n548);
xor (n547,n500,n501);
and (n548,n154,n43);
and (n549,n550,n551);
xor (n550,n547,n548);
or (n551,n552,n555);
and (n552,n553,n554);
xor (n553,n506,n507);
and (n554,n77,n43);
and (n555,n556,n557);
xor (n556,n553,n554);
or (n557,n558,n561);
and (n558,n559,n560);
xor (n559,n512,n513);
and (n560,n71,n43);
and (n561,n562,n563);
xor (n562,n559,n560);
or (n563,n564,n567);
and (n564,n565,n566);
xor (n565,n518,n519);
and (n566,n70,n43);
and (n567,n568,n569);
xor (n568,n565,n566);
or (n569,n570,n573);
and (n570,n571,n572);
xor (n571,n523,n524);
and (n572,n120,n43);
and (n573,n574,n575);
xor (n574,n571,n572);
or (n575,n576,n578);
and (n576,n577,n386);
xor (n577,n529,n530);
and (n578,n579,n580);
xor (n579,n577,n386);
and (n580,n581,n582);
xor (n581,n535,n536);
and (n582,n57,n43);
and (n583,n34,n181);
or (n584,n585,n588);
and (n585,n586,n587);
xor (n586,n544,n545);
and (n587,n154,n181);
and (n588,n589,n590);
xor (n589,n586,n587);
or (n590,n591,n594);
and (n591,n592,n593);
xor (n592,n550,n551);
and (n593,n77,n181);
and (n594,n595,n596);
xor (n595,n592,n593);
or (n596,n597,n600);
and (n597,n598,n599);
xor (n598,n556,n557);
and (n599,n71,n181);
and (n600,n601,n602);
xor (n601,n598,n599);
or (n602,n603,n605);
and (n603,n604,n300);
xor (n604,n562,n563);
and (n605,n606,n607);
xor (n606,n604,n300);
or (n607,n608,n611);
and (n608,n609,n610);
xor (n609,n568,n569);
and (n610,n120,n181);
and (n611,n612,n613);
xor (n612,n609,n610);
or (n613,n614,n616);
and (n614,n615,n372);
xor (n615,n574,n575);
and (n616,n617,n618);
xor (n617,n615,n372);
and (n618,n619,n620);
xor (n619,n579,n580);
and (n620,n57,n181);
and (n621,n154,n97);
or (n622,n623,n626);
and (n623,n624,n625);
xor (n624,n589,n590);
and (n625,n77,n97);
and (n626,n627,n628);
xor (n627,n624,n625);
or (n628,n629,n632);
and (n629,n630,n631);
xor (n630,n595,n596);
and (n631,n71,n97);
and (n632,n633,n634);
xor (n633,n630,n631);
or (n634,n635,n638);
and (n635,n636,n637);
xor (n636,n601,n602);
and (n637,n70,n97);
and (n638,n639,n640);
xor (n639,n636,n637);
or (n640,n641,n644);
and (n641,n642,n643);
xor (n642,n606,n607);
and (n643,n120,n97);
and (n644,n645,n646);
xor (n645,n642,n643);
or (n646,n647,n649);
and (n647,n648,n277);
xor (n648,n612,n613);
and (n649,n650,n651);
xor (n650,n648,n277);
and (n651,n652,n653);
xor (n652,n617,n618);
and (n653,n57,n97);
and (n654,n77,n81);
or (n655,n656,n659);
and (n656,n657,n658);
xor (n657,n627,n628);
and (n658,n71,n81);
and (n659,n660,n661);
xor (n660,n657,n658);
or (n661,n662,n665);
and (n662,n663,n664);
xor (n663,n633,n634);
and (n664,n70,n81);
and (n665,n666,n667);
xor (n666,n663,n664);
or (n667,n668,n671);
and (n668,n669,n670);
xor (n669,n639,n640);
and (n670,n120,n81);
and (n671,n672,n673);
xor (n672,n669,n670);
or (n673,n674,n677);
and (n674,n675,n676);
xor (n675,n645,n646);
and (n676,n51,n81);
and (n677,n678,n679);
xor (n678,n675,n676);
and (n679,n680,n681);
xor (n680,n650,n651);
and (n681,n57,n81);
and (n682,n71,n87);
or (n683,n684,n687);
and (n684,n685,n686);
xor (n685,n660,n661);
and (n686,n70,n87);
and (n687,n688,n689);
xor (n688,n685,n686);
or (n689,n690,n693);
and (n690,n691,n692);
xor (n691,n666,n667);
and (n692,n120,n87);
and (n693,n694,n695);
xor (n694,n691,n692);
or (n695,n696,n698);
and (n696,n697,n247);
xor (n697,n672,n673);
and (n698,n699,n700);
xor (n699,n697,n247);
and (n700,n701,n702);
xor (n701,n678,n679);
and (n702,n57,n87);
and (n703,n70,n131);
or (n704,n705,n708);
and (n705,n706,n707);
xor (n706,n688,n689);
and (n707,n120,n131);
and (n708,n709,n710);
xor (n709,n706,n707);
or (n710,n711,n714);
and (n711,n712,n713);
xor (n712,n694,n695);
and (n713,n51,n131);
and (n714,n715,n716);
xor (n715,n712,n713);
and (n716,n717,n718);
xor (n717,n699,n700);
and (n718,n57,n131);
and (n719,n120,n143);
or (n720,n721,n723);
and (n721,n722,n144);
xor (n722,n709,n710);
and (n723,n724,n725);
xor (n724,n722,n144);
and (n725,n726,n727);
xor (n726,n715,n716);
and (n727,n57,n143);
and (n728,n51,n52);
and (n729,n730,n731);
xor (n730,n724,n725);
and (n731,n57,n52);
and (n732,n57,n61);
endmodule
