module top (out,n9,n12,n13,n17,n20,n21,n25,n33,n36
        ,n37,n41,n47,n61,n62,n128,n131,n168,n176,n177
        ,n223,n281,n282,n334,n339,n385,n386,n423,n492,n556
        ,n650,n723,n808);
output out;
input n9;
input n12;
input n13;
input n17;
input n20;
input n21;
input n25;
input n33;
input n36;
input n37;
input n41;
input n47;
input n61;
input n62;
input n128;
input n131;
input n168;
input n176;
input n177;
input n223;
input n281;
input n282;
input n334;
input n339;
input n385;
input n386;
input n423;
input n492;
input n556;
input n650;
input n723;
input n808;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n10;
wire n11;
wire n14;
wire n15;
wire n16;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n335;
wire n336;
wire n337;
wire n338;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
xor (out,n0,n1465);
xor (n0,n1,n148);
xor (n1,n2,n107);
xor (n2,n3,n95);
xor (n3,n4,n51);
or (n4,n5,n48,n50);
and (n5,n6,n46);
or (n6,n7,n29,n45);
and (n7,n8,n14);
and (n8,n9,n10);
not (n10,n11);
and (n11,n12,n13);
xnor (n14,n15,n26);
nor (n15,n16,n24);
and (n16,n17,n18);
and (n18,n19,n22);
xor (n19,n20,n21);
not (n22,n23);
xor (n23,n21,n9);
and (n24,n25,n23);
and (n26,n20,n27);
not (n27,n28);
and (n28,n21,n9);
and (n29,n14,n30);
xnor (n30,n31,n42);
nor (n31,n32,n40);
and (n32,n33,n34);
and (n34,n35,n38);
xor (n35,n36,n37);
not (n38,n39);
xor (n39,n37,n20);
and (n40,n41,n39);
and (n42,n36,n43);
not (n43,n44);
and (n44,n37,n20);
and (n45,n8,n30);
and (n46,n47,n36);
and (n48,n46,n49);
and (n49,n33,n36);
and (n50,n6,n49);
or (n51,n52,n91,n94);
and (n52,n53,n81);
or (n53,n54,n78,n80);
and (n54,n55,n76);
or (n55,n56,n70,n75);
and (n56,n57,n63);
not (n57,n58);
and (n58,n13,n59);
not (n59,n60);
and (n60,n61,n62);
xnor (n63,n64,n8);
not (n64,n65);
and (n65,n25,n66);
and (n66,n67,n68);
xor (n67,n9,n12);
not (n68,n69);
xor (n69,n12,n13);
and (n70,n63,n71);
xnor (n71,n72,n26);
nor (n72,n73,n74);
and (n73,n41,n18);
and (n74,n17,n23);
and (n75,n57,n71);
xor (n76,n77,n30);
xor (n77,n8,n14);
and (n78,n76,n79);
not (n79,n46);
and (n80,n55,n79);
xor (n81,n82,n87);
xor (n82,n83,n84);
not (n83,n8);
xnor (n84,n85,n26);
not (n85,n86);
and (n86,n25,n18);
xnor (n87,n88,n42);
nor (n88,n89,n90);
and (n89,n41,n34);
and (n90,n17,n39);
and (n91,n81,n92);
xor (n92,n93,n49);
xor (n93,n6,n46);
and (n94,n53,n92);
xnor (n95,n96,n100);
or (n96,n97,n98,n99);
and (n97,n83,n84);
and (n98,n84,n87);
and (n99,n83,n87);
xor (n100,n101,n106);
xor (n101,n26,n102);
xnor (n102,n103,n42);
nor (n103,n104,n105);
and (n104,n17,n34);
and (n105,n25,n39);
and (n106,n41,n36);
and (n107,n108,n146);
or (n108,n109,n142,n145);
and (n109,n110,n138);
or (n110,n111,n132,n137);
and (n111,n112,n124);
or (n112,n113,n118,n123);
and (n113,n58,n114);
xnor (n114,n115,n8);
nor (n115,n116,n117);
and (n116,n17,n66);
and (n117,n25,n69);
and (n118,n114,n119);
xnor (n119,n120,n26);
nor (n120,n121,n122);
and (n121,n33,n18);
and (n122,n41,n23);
and (n123,n58,n119);
or (n124,n125,n130);
xnor (n125,n126,n42);
nor (n126,n127,n129);
and (n127,n128,n34);
and (n129,n47,n39);
and (n130,n131,n36);
and (n132,n124,n133);
xnor (n133,n134,n42);
nor (n134,n135,n136);
and (n135,n47,n34);
and (n136,n33,n39);
and (n137,n112,n133);
and (n138,n139,n140);
and (n139,n128,n36);
xor (n140,n141,n71);
xor (n141,n57,n63);
and (n142,n138,n143);
xor (n143,n144,n79);
xor (n144,n55,n76);
and (n145,n110,n143);
xor (n146,n147,n92);
xor (n147,n53,n81);
or (n148,n149,n201);
and (n149,n150,n151);
xor (n150,n108,n146);
and (n151,n152,n199);
or (n152,n153,n196,n198);
and (n153,n154,n194);
or (n154,n155,n191,n193);
and (n155,n156,n170);
or (n156,n157,n166,n169);
and (n157,n158,n162);
xnor (n158,n159,n26);
nor (n159,n160,n161);
and (n160,n47,n18);
and (n161,n33,n23);
xnor (n162,n163,n42);
nor (n163,n164,n165);
and (n164,n131,n34);
and (n165,n128,n39);
and (n166,n162,n167);
and (n167,n168,n36);
and (n169,n158,n167);
or (n170,n171,n185,n190);
and (n171,n172,n178);
not (n172,n173);
and (n173,n62,n174);
not (n174,n175);
and (n175,n176,n177);
xnor (n178,n179,n58);
not (n179,n180);
and (n180,n25,n181);
and (n181,n182,n183);
xor (n182,n13,n61);
not (n183,n184);
xor (n184,n61,n62);
and (n185,n178,n186);
xnor (n186,n187,n8);
nor (n187,n188,n189);
and (n188,n41,n66);
and (n189,n17,n69);
and (n190,n172,n186);
and (n191,n170,n192);
xnor (n192,n125,n130);
and (n193,n156,n192);
xor (n194,n195,n133);
xor (n195,n112,n124);
and (n196,n194,n197);
xor (n197,n139,n140);
and (n198,n154,n197);
xor (n199,n200,n143);
xor (n200,n110,n138);
and (n201,n202,n203);
xor (n202,n150,n151);
or (n203,n204,n249);
and (n204,n205,n206);
xor (n205,n152,n199);
and (n206,n207,n247);
or (n207,n208,n243,n246);
and (n208,n209,n241);
or (n209,n210,n237,n240);
and (n210,n211,n225);
or (n211,n212,n221,n224);
and (n212,n213,n217);
xnor (n213,n214,n26);
nor (n214,n215,n216);
and (n215,n128,n18);
and (n216,n47,n23);
xnor (n217,n218,n42);
nor (n218,n219,n220);
and (n219,n168,n34);
and (n220,n131,n39);
and (n221,n217,n222);
and (n222,n223,n36);
and (n224,n213,n222);
or (n225,n226,n231,n236);
and (n226,n173,n227);
xnor (n227,n228,n58);
nor (n228,n229,n230);
and (n229,n17,n181);
and (n230,n25,n184);
and (n231,n227,n232);
xnor (n232,n233,n8);
nor (n233,n234,n235);
and (n234,n33,n66);
and (n235,n41,n69);
and (n236,n173,n232);
and (n237,n225,n238);
xor (n238,n239,n167);
xor (n239,n158,n162);
and (n240,n211,n238);
xor (n241,n242,n119);
xor (n242,n58,n114);
and (n243,n241,n244);
xor (n244,n245,n192);
xor (n245,n156,n170);
and (n246,n209,n244);
xor (n247,n248,n197);
xor (n248,n154,n194);
and (n249,n250,n251);
xor (n250,n205,n206);
or (n251,n252,n366);
and (n252,n253,n254);
xor (n253,n207,n247);
or (n254,n255,n362,n365);
and (n255,n256,n302);
or (n256,n257,n298,n301);
and (n257,n258,n296);
or (n258,n259,n275);
or (n259,n260,n269,n274);
and (n260,n261,n265);
xnor (n261,n262,n8);
nor (n262,n263,n264);
and (n263,n47,n66);
and (n264,n33,n69);
xnor (n265,n266,n26);
nor (n266,n267,n268);
and (n267,n131,n18);
and (n268,n128,n23);
and (n269,n265,n270);
xnor (n270,n271,n42);
nor (n271,n272,n273);
and (n272,n223,n34);
and (n273,n168,n39);
and (n274,n261,n270);
or (n275,n276,n290,n295);
and (n276,n277,n283);
not (n277,n278);
and (n278,n177,n279);
not (n279,n280);
and (n280,n281,n282);
xnor (n283,n284,n173);
not (n284,n285);
and (n285,n25,n286);
and (n286,n287,n288);
xor (n287,n62,n176);
not (n288,n289);
xor (n289,n176,n177);
and (n290,n283,n291);
xnor (n291,n292,n58);
nor (n292,n293,n294);
and (n293,n41,n181);
and (n294,n17,n184);
and (n295,n277,n291);
xor (n296,n297,n186);
xor (n297,n172,n178);
and (n298,n296,n299);
xor (n299,n300,n238);
xor (n300,n211,n225);
and (n301,n258,n299);
or (n302,n303,n358,n361);
and (n303,n304,n354);
or (n304,n305,n350,n353);
and (n305,n306,n341);
or (n306,n307,n337,n340);
and (n307,n308,n320);
or (n308,n309,n314,n319);
and (n309,n278,n310);
xnor (n310,n311,n173);
nor (n311,n312,n313);
and (n312,n17,n286);
and (n313,n25,n289);
and (n314,n310,n315);
xnor (n315,n316,n58);
nor (n316,n317,n318);
and (n317,n33,n181);
and (n318,n41,n184);
and (n319,n278,n315);
or (n320,n321,n330,n336);
and (n321,n322,n326);
xnor (n322,n323,n8);
nor (n323,n324,n325);
and (n324,n128,n66);
and (n325,n47,n69);
xnor (n326,n327,n26);
nor (n327,n328,n329);
and (n328,n168,n18);
and (n329,n131,n23);
and (n330,n326,n331);
xnor (n331,n332,n42);
nor (n332,n333,n335);
and (n333,n334,n34);
and (n335,n223,n39);
and (n336,n322,n331);
and (n337,n320,n338);
and (n338,n339,n36);
and (n340,n308,n338);
or (n341,n342,n346,n349);
and (n342,n343,n344);
and (n343,n334,n36);
xor (n344,n345,n270);
xor (n345,n261,n265);
and (n346,n344,n347);
xor (n347,n348,n291);
xor (n348,n277,n283);
and (n349,n343,n347);
and (n350,n341,n351);
xor (n351,n352,n222);
xor (n352,n213,n217);
and (n353,n306,n351);
and (n354,n355,n357);
xor (n355,n356,n232);
xor (n356,n173,n227);
xnor (n357,n259,n275);
and (n358,n354,n359);
xor (n359,n360,n299);
xor (n360,n258,n296);
and (n361,n304,n359);
and (n362,n302,n363);
xor (n363,n364,n244);
xor (n364,n209,n241);
and (n365,n256,n363);
and (n366,n367,n368);
xor (n367,n253,n254);
or (n368,n369,n445);
and (n369,n370,n372);
xor (n370,n371,n363);
xor (n371,n256,n302);
and (n372,n373,n443);
or (n373,n374,n440,n442);
and (n374,n375,n438);
or (n375,n376,n434,n437);
and (n376,n377,n425);
or (n377,n378,n416,n424);
and (n378,n379,n400);
or (n379,n380,n394,n399);
and (n380,n381,n387);
not (n381,n382);
and (n382,n282,n383);
not (n383,n384);
and (n384,n385,n386);
xnor (n387,n388,n278);
not (n388,n389);
and (n389,n25,n390);
and (n390,n391,n392);
xor (n391,n177,n281);
not (n392,n393);
xor (n393,n281,n282);
and (n394,n387,n395);
xnor (n395,n396,n173);
nor (n396,n397,n398);
and (n397,n41,n286);
and (n398,n17,n289);
and (n399,n381,n395);
or (n400,n401,n410,n415);
and (n401,n402,n406);
xnor (n402,n403,n58);
nor (n403,n404,n405);
and (n404,n47,n181);
and (n405,n33,n184);
xnor (n406,n407,n8);
nor (n407,n408,n409);
and (n408,n131,n66);
and (n409,n128,n69);
and (n410,n406,n411);
xnor (n411,n412,n26);
nor (n412,n413,n414);
and (n413,n223,n18);
and (n414,n168,n23);
and (n415,n402,n411);
and (n416,n400,n417);
and (n417,n418,n422);
xnor (n418,n419,n42);
nor (n419,n420,n421);
and (n420,n339,n34);
and (n421,n334,n39);
and (n422,n423,n36);
and (n424,n379,n417);
or (n425,n426,n431,n433);
and (n426,n427,n429);
xor (n427,n428,n315);
xor (n428,n278,n310);
xor (n429,n430,n331);
xor (n430,n322,n326);
and (n431,n429,n432);
not (n432,n338);
and (n433,n427,n432);
and (n434,n425,n435);
xor (n435,n436,n347);
xor (n436,n343,n344);
and (n437,n377,n435);
xor (n438,n439,n351);
xor (n439,n306,n341);
and (n440,n438,n441);
xor (n441,n355,n357);
and (n442,n375,n441);
xor (n443,n444,n359);
xor (n444,n304,n354);
and (n445,n446,n447);
xor (n446,n370,n372);
or (n447,n448,n516);
and (n448,n449,n450);
xor (n449,n373,n443);
and (n450,n451,n514);
or (n451,n452,n510,n513);
and (n452,n453,n508);
or (n453,n454,n503,n507);
and (n454,n455,n494);
or (n455,n456,n485,n493);
and (n456,n457,n469);
or (n457,n458,n463,n468);
and (n458,n382,n459);
xnor (n459,n460,n278);
nor (n460,n461,n462);
and (n461,n17,n390);
and (n462,n25,n393);
and (n463,n459,n464);
xnor (n464,n465,n173);
nor (n465,n466,n467);
and (n466,n33,n286);
and (n467,n41,n289);
and (n468,n382,n464);
or (n469,n470,n479,n484);
and (n470,n471,n475);
xnor (n471,n472,n58);
nor (n472,n473,n474);
and (n473,n128,n181);
and (n474,n47,n184);
xnor (n475,n476,n8);
nor (n476,n477,n478);
and (n477,n168,n66);
and (n478,n131,n69);
and (n479,n475,n480);
xnor (n480,n481,n26);
nor (n481,n482,n483);
and (n482,n334,n18);
and (n483,n223,n23);
and (n484,n471,n480);
and (n485,n469,n486);
or (n486,n487,n491);
xnor (n487,n488,n42);
nor (n488,n489,n490);
and (n489,n423,n34);
and (n490,n339,n39);
and (n491,n492,n36);
and (n493,n457,n486);
or (n494,n495,n500,n502);
and (n495,n496,n498);
xor (n496,n497,n395);
xor (n497,n381,n387);
xor (n498,n499,n411);
xor (n499,n402,n406);
and (n500,n498,n501);
xor (n501,n418,n422);
and (n502,n496,n501);
and (n503,n494,n504);
xor (n504,n505,n429);
xor (n505,n338,n506);
not (n506,n427);
and (n507,n455,n504);
xor (n508,n509,n338);
xor (n509,n308,n320);
and (n510,n508,n511);
xor (n511,n512,n435);
xor (n512,n377,n425);
and (n513,n453,n511);
xor (n514,n515,n441);
xor (n515,n375,n438);
and (n516,n517,n518);
xor (n517,n449,n450);
or (n518,n519,n597);
and (n519,n520,n521);
xor (n520,n451,n514);
and (n521,n522,n595);
or (n522,n523,n591,n594);
and (n523,n524,n589);
or (n524,n525,n585,n588);
and (n525,n526,n576);
or (n526,n527,n558,n575);
and (n527,n528,n544);
or (n528,n529,n538,n543);
and (n529,n530,n531);
not (n530,n386);
xnor (n531,n532,n382);
not (n532,n533);
and (n533,n25,n534);
and (n534,n535,n536);
xor (n535,n282,n385);
not (n536,n537);
xor (n537,n385,n386);
and (n538,n531,n539);
xnor (n539,n540,n278);
nor (n540,n541,n542);
and (n541,n41,n390);
and (n542,n17,n393);
and (n543,n530,n539);
or (n544,n545,n554,n557);
and (n545,n546,n550);
xnor (n546,n547,n26);
nor (n547,n548,n549);
and (n548,n339,n18);
and (n549,n334,n23);
xnor (n550,n551,n42);
nor (n551,n552,n553);
and (n552,n492,n34);
and (n553,n423,n39);
and (n554,n550,n555);
and (n555,n556,n36);
and (n557,n546,n555);
and (n558,n544,n559);
or (n559,n560,n569,n574);
and (n560,n561,n565);
xnor (n561,n562,n173);
nor (n562,n563,n564);
and (n563,n47,n286);
and (n564,n33,n289);
xnor (n565,n566,n58);
nor (n566,n567,n568);
and (n567,n131,n181);
and (n568,n128,n184);
and (n569,n565,n570);
xnor (n570,n571,n8);
nor (n571,n572,n573);
and (n572,n223,n66);
and (n573,n168,n69);
and (n574,n561,n570);
and (n575,n528,n559);
or (n576,n577,n582,n584);
and (n577,n578,n580);
xor (n578,n579,n464);
xor (n579,n382,n459);
xor (n580,n581,n480);
xor (n581,n471,n475);
and (n582,n580,n583);
xnor (n583,n487,n491);
and (n584,n578,n583);
and (n585,n576,n586);
xor (n586,n587,n501);
xor (n587,n496,n498);
and (n588,n526,n586);
xor (n589,n590,n417);
xor (n590,n379,n400);
and (n591,n589,n592);
xor (n592,n593,n504);
xor (n593,n455,n494);
and (n594,n524,n592);
xor (n595,n596,n511);
xor (n596,n453,n508);
and (n597,n598,n599);
xor (n598,n520,n521);
or (n599,n600,n672);
and (n600,n601,n602);
xor (n601,n522,n595);
and (n602,n603,n670);
or (n603,n604,n666,n669);
and (n604,n605,n664);
or (n605,n606,n658,n663);
and (n606,n607,n653);
or (n607,n608,n637,n652);
and (n608,n609,n625);
or (n609,n610,n619,n624);
and (n610,n611,n615);
xnor (n611,n612,n173);
nor (n612,n613,n614);
and (n613,n128,n286);
and (n614,n47,n289);
xnor (n615,n616,n58);
nor (n616,n617,n618);
and (n617,n168,n181);
and (n618,n131,n184);
and (n619,n615,n620);
xnor (n620,n621,n8);
nor (n621,n622,n623);
and (n622,n334,n66);
and (n623,n223,n69);
and (n624,n611,n620);
or (n625,n626,n631,n636);
and (n626,n386,n627);
xnor (n627,n628,n382);
nor (n628,n629,n630);
and (n629,n17,n534);
and (n630,n25,n537);
and (n631,n627,n632);
xnor (n632,n633,n278);
nor (n633,n634,n635);
and (n634,n33,n390);
and (n635,n41,n393);
and (n636,n386,n632);
and (n637,n625,n638);
or (n638,n639,n648,n651);
and (n639,n640,n644);
xnor (n640,n641,n26);
nor (n641,n642,n643);
and (n642,n423,n18);
and (n643,n339,n23);
xnor (n644,n645,n42);
nor (n645,n646,n647);
and (n646,n556,n34);
and (n647,n492,n39);
and (n648,n644,n649);
and (n649,n650,n36);
and (n651,n640,n649);
and (n652,n609,n638);
or (n653,n654,n656);
xor (n654,n655,n555);
xor (n655,n546,n550);
xor (n656,n657,n570);
xor (n657,n561,n565);
and (n658,n653,n659);
xor (n659,n660,n662);
xor (n660,n661,n580);
not (n661,n578);
not (n662,n583);
and (n663,n607,n659);
xor (n664,n665,n486);
xor (n665,n457,n469);
and (n666,n664,n667);
xor (n667,n668,n586);
xor (n668,n526,n576);
and (n669,n605,n667);
xor (n670,n671,n592);
xor (n671,n524,n589);
and (n672,n673,n674);
xor (n673,n601,n602);
or (n674,n675,n754);
and (n675,n676,n677);
xor (n676,n603,n670);
and (n677,n678,n752);
or (n678,n679,n748,n751);
and (n679,n680,n744);
or (n680,n681,n740,n743);
and (n681,n682,n730);
or (n682,n683,n716,n729);
and (n683,n684,n700);
or (n684,n685,n694,n699);
and (n685,n686,n690);
xnor (n686,n687,n278);
nor (n687,n688,n689);
and (n688,n47,n390);
and (n689,n33,n393);
xnor (n690,n691,n173);
nor (n691,n692,n693);
and (n692,n131,n286);
and (n693,n128,n289);
and (n694,n690,n695);
xnor (n695,n696,n58);
nor (n696,n697,n698);
and (n697,n223,n181);
and (n698,n168,n184);
and (n699,n686,n695);
or (n700,n701,n710,n715);
and (n701,n702,n706);
xnor (n702,n703,n8);
nor (n703,n704,n705);
and (n704,n339,n66);
and (n705,n334,n69);
xnor (n706,n707,n26);
nor (n707,n708,n709);
and (n708,n492,n18);
and (n709,n423,n23);
and (n710,n706,n711);
xnor (n711,n712,n42);
nor (n712,n713,n714);
and (n713,n650,n34);
and (n714,n556,n39);
and (n715,n702,n711);
and (n716,n700,n717);
and (n717,n718,n725);
xnor (n718,n719,n386);
not (n719,n720);
and (n720,n25,n721);
and (n721,n722,n724);
xor (n722,n386,n723);
not (n724,n723);
xnor (n725,n726,n382);
nor (n726,n727,n728);
and (n727,n41,n534);
and (n728,n17,n537);
and (n729,n684,n717);
or (n730,n731,n736,n739);
and (n731,n732,n734);
xor (n732,n733,n620);
xor (n733,n611,n615);
xor (n734,n735,n632);
xor (n735,n386,n627);
and (n736,n734,n737);
xor (n737,n738,n649);
xor (n738,n640,n644);
and (n739,n732,n737);
and (n740,n730,n741);
xor (n741,n742,n539);
xor (n742,n530,n531);
and (n743,n682,n741);
and (n744,n745,n747);
xor (n745,n746,n638);
xor (n746,n609,n625);
xnor (n747,n654,n656);
and (n748,n744,n749);
xor (n749,n750,n559);
xor (n750,n528,n544);
and (n751,n680,n749);
xor (n752,n753,n667);
xor (n753,n605,n664);
and (n754,n755,n756);
xor (n755,n676,n677);
or (n756,n757,n836);
and (n757,n758,n759);
xor (n758,n678,n752);
or (n759,n760,n832,n835);
and (n760,n761,n830);
or (n761,n762,n827,n829);
and (n762,n763,n825);
or (n763,n764,n821,n824);
and (n764,n765,n811);
or (n765,n766,n799,n810);
and (n766,n767,n783);
or (n767,n768,n777,n782);
and (n768,n769,n773);
xnor (n769,n770,n386);
nor (n770,n771,n772);
and (n771,n17,n721);
and (n772,n25,n723);
xnor (n773,n774,n382);
nor (n774,n775,n776);
and (n775,n33,n534);
and (n776,n41,n537);
and (n777,n773,n778);
xnor (n778,n779,n278);
nor (n779,n780,n781);
and (n780,n128,n390);
and (n781,n47,n393);
and (n782,n769,n778);
or (n783,n784,n793,n798);
and (n784,n785,n789);
xnor (n785,n786,n173);
nor (n786,n787,n788);
and (n787,n168,n286);
and (n788,n131,n289);
xnor (n789,n790,n58);
nor (n790,n791,n792);
and (n791,n334,n181);
and (n792,n223,n184);
and (n793,n789,n794);
xnor (n794,n795,n8);
nor (n795,n796,n797);
and (n796,n423,n66);
and (n797,n339,n69);
and (n798,n785,n794);
and (n799,n783,n800);
and (n800,n801,n805);
xnor (n801,n802,n26);
nor (n802,n803,n804);
and (n803,n556,n18);
and (n804,n492,n23);
xnor (n805,n806,n42);
nor (n806,n807,n809);
and (n807,n808,n34);
and (n809,n650,n39);
and (n810,n767,n800);
or (n811,n812,n817,n820);
and (n812,n813,n815);
not (n813,n814);
nand (n814,n808,n36);
xor (n815,n816,n695);
xor (n816,n686,n690);
and (n817,n815,n818);
xor (n818,n819,n711);
xor (n819,n702,n706);
and (n820,n813,n818);
and (n821,n811,n822);
xor (n822,n823,n737);
xor (n823,n732,n734);
and (n824,n765,n822);
xor (n825,n826,n741);
xor (n826,n682,n730);
and (n827,n825,n828);
xor (n828,n745,n747);
and (n829,n763,n828);
xor (n830,n831,n749);
xor (n831,n680,n744);
and (n832,n830,n833);
xor (n833,n834,n659);
xor (n834,n607,n653);
and (n835,n761,n833);
and (n836,n837,n838);
xor (n837,n758,n759);
or (n838,n839,n916);
and (n839,n840,n842);
xor (n840,n841,n833);
xor (n841,n761,n830);
and (n842,n843,n914);
or (n843,n844,n910,n913);
and (n844,n845,n905);
or (n845,n846,n902,n904);
and (n846,n847,n893);
or (n847,n848,n875,n892);
and (n848,n849,n863);
or (n849,n850,n859,n862);
and (n850,n851,n855);
xnor (n851,n852,n8);
nor (n852,n853,n854);
and (n853,n492,n66);
and (n854,n423,n69);
xnor (n855,n856,n26);
nor (n856,n857,n858);
and (n857,n650,n18);
and (n858,n556,n23);
and (n859,n855,n860);
xnor (n860,n861,n42);
nand (n861,n808,n39);
and (n862,n851,n860);
or (n863,n864,n873,n874);
and (n864,n865,n869);
xnor (n865,n866,n386);
nor (n866,n867,n868);
and (n867,n41,n721);
and (n868,n17,n723);
xnor (n869,n870,n382);
nor (n870,n871,n872);
and (n871,n47,n534);
and (n872,n33,n537);
and (n873,n869,n42);
and (n874,n865,n42);
and (n875,n863,n876);
or (n876,n877,n886,n891);
and (n877,n878,n882);
xnor (n878,n879,n278);
nor (n879,n880,n881);
and (n880,n131,n390);
and (n881,n128,n393);
xnor (n882,n883,n173);
nor (n883,n884,n885);
and (n884,n223,n286);
and (n885,n168,n289);
and (n886,n882,n887);
xnor (n887,n888,n58);
nor (n888,n889,n890);
and (n889,n339,n181);
and (n890,n334,n184);
and (n891,n878,n887);
and (n892,n849,n876);
or (n893,n894,n899,n901);
and (n894,n895,n897);
xor (n895,n896,n778);
xor (n896,n769,n773);
xor (n897,n898,n794);
xor (n898,n785,n789);
and (n899,n897,n900);
xor (n900,n801,n805);
and (n901,n895,n900);
and (n902,n893,n903);
xor (n903,n718,n725);
and (n904,n847,n903);
and (n905,n906,n908);
xor (n906,n907,n800);
xor (n907,n767,n783);
xor (n908,n909,n818);
xor (n909,n813,n815);
and (n910,n905,n911);
xor (n911,n912,n717);
xor (n912,n684,n700);
and (n913,n845,n911);
xor (n914,n915,n828);
xor (n915,n763,n825);
and (n916,n917,n918);
xor (n917,n840,n842);
or (n918,n919,n926);
and (n919,n920,n921);
xor (n920,n843,n914);
and (n921,n922,n924);
xor (n922,n923,n911);
xor (n923,n845,n905);
xor (n924,n925,n822);
xor (n925,n765,n811);
and (n926,n927,n928);
xor (n927,n920,n921);
or (n928,n929,n992);
and (n929,n930,n936);
xor (n930,n931,n934);
xor (n931,n911,n932);
xor (n932,n925,n933);
not (n933,n734);
xor (n934,n923,n935);
xnor (n935,n732,n737);
or (n936,n937,n989,n991);
and (n937,n938,n987);
or (n938,n939,n983,n986);
and (n939,n940,n978);
or (n940,n941,n974,n977);
and (n941,n942,n958);
or (n942,n943,n952,n957);
and (n943,n944,n948);
xnor (n944,n945,n386);
nor (n945,n946,n947);
and (n946,n33,n721);
and (n947,n41,n723);
xnor (n948,n949,n382);
nor (n949,n950,n951);
and (n950,n128,n534);
and (n951,n47,n537);
and (n952,n948,n953);
xnor (n953,n954,n278);
nor (n954,n955,n956);
and (n955,n168,n390);
and (n956,n131,n393);
and (n957,n944,n953);
or (n958,n959,n968,n973);
and (n959,n960,n964);
xnor (n960,n961,n173);
nor (n961,n962,n963);
and (n962,n334,n286);
and (n963,n223,n289);
xnor (n964,n965,n58);
nor (n965,n966,n967);
and (n966,n423,n181);
and (n967,n339,n184);
and (n968,n964,n969);
xnor (n969,n970,n8);
nor (n970,n971,n972);
and (n971,n556,n66);
and (n972,n492,n69);
and (n973,n960,n969);
and (n974,n958,n975);
xor (n975,n976,n860);
xor (n976,n851,n855);
and (n977,n942,n975);
and (n978,n979,n981);
xor (n979,n980,n42);
xor (n980,n865,n869);
xor (n981,n982,n887);
xor (n982,n878,n882);
and (n983,n978,n984);
xor (n984,n985,n900);
xor (n985,n895,n897);
and (n986,n940,n984);
xor (n987,n988,n903);
xor (n988,n847,n893);
and (n989,n987,n990);
xor (n990,n906,n908);
and (n991,n938,n990);
and (n992,n993,n994);
xor (n993,n930,n936);
or (n994,n995,n1049);
and (n995,n996,n998);
xor (n996,n997,n990);
xor (n997,n938,n987);
or (n998,n999,n1045,n1048);
and (n999,n1000,n1043);
or (n1000,n1001,n1040,n1042);
and (n1001,n1002,n1038);
or (n1002,n1003,n1032,n1037);
and (n1003,n1004,n1016);
or (n1004,n1005,n1014,n1015);
and (n1005,n1006,n1010);
xnor (n1006,n1007,n386);
nor (n1007,n1008,n1009);
and (n1008,n47,n721);
and (n1009,n33,n723);
xnor (n1010,n1011,n382);
nor (n1011,n1012,n1013);
and (n1012,n131,n534);
and (n1013,n128,n537);
and (n1014,n1010,n26);
and (n1015,n1006,n26);
or (n1016,n1017,n1026,n1031);
and (n1017,n1018,n1022);
xnor (n1018,n1019,n278);
nor (n1019,n1020,n1021);
and (n1020,n223,n390);
and (n1021,n168,n393);
xnor (n1022,n1023,n173);
nor (n1023,n1024,n1025);
and (n1024,n339,n286);
and (n1025,n334,n289);
and (n1026,n1022,n1027);
xnor (n1027,n1028,n58);
nor (n1028,n1029,n1030);
and (n1029,n492,n181);
and (n1030,n423,n184);
and (n1031,n1018,n1027);
and (n1032,n1016,n1033);
xnor (n1033,n1034,n26);
nor (n1034,n1035,n1036);
and (n1035,n808,n18);
and (n1036,n650,n23);
and (n1037,n1004,n1033);
xor (n1038,n1039,n975);
xor (n1039,n942,n958);
and (n1040,n1038,n1041);
xor (n1041,n979,n981);
and (n1042,n1002,n1041);
xor (n1043,n1044,n876);
xor (n1044,n849,n863);
and (n1045,n1043,n1046);
xor (n1046,n1047,n984);
xor (n1047,n940,n978);
and (n1048,n1000,n1046);
and (n1049,n1050,n1051);
xor (n1050,n996,n998);
or (n1051,n1052,n1122);
and (n1052,n1053,n1055);
xor (n1053,n1054,n1046);
xor (n1054,n1000,n1043);
or (n1055,n1056,n1118,n1121);
and (n1056,n1057,n1113);
or (n1057,n1058,n1109,n1112);
and (n1058,n1059,n1099);
or (n1059,n1060,n1093,n1098);
and (n1060,n1061,n1077);
or (n1061,n1062,n1071,n1076);
and (n1062,n1063,n1067);
xnor (n1063,n1064,n173);
nor (n1064,n1065,n1066);
and (n1065,n423,n286);
and (n1066,n339,n289);
xnor (n1067,n1068,n58);
nor (n1068,n1069,n1070);
and (n1069,n556,n181);
and (n1070,n492,n184);
and (n1071,n1067,n1072);
xnor (n1072,n1073,n8);
nor (n1073,n1074,n1075);
and (n1074,n808,n66);
and (n1075,n650,n69);
and (n1076,n1063,n1072);
or (n1077,n1078,n1087,n1092);
and (n1078,n1079,n1083);
xnor (n1079,n1080,n386);
nor (n1080,n1081,n1082);
and (n1081,n128,n721);
and (n1082,n47,n723);
xnor (n1083,n1084,n382);
nor (n1084,n1085,n1086);
and (n1085,n168,n534);
and (n1086,n131,n537);
and (n1087,n1083,n1088);
xnor (n1088,n1089,n278);
nor (n1089,n1090,n1091);
and (n1090,n334,n390);
and (n1091,n223,n393);
and (n1092,n1079,n1088);
and (n1093,n1077,n1094);
xnor (n1094,n1095,n8);
nor (n1095,n1096,n1097);
and (n1096,n650,n66);
and (n1097,n556,n69);
and (n1098,n1061,n1094);
or (n1099,n1100,n1105,n1108);
and (n1100,n1101,n1103);
xnor (n1101,n1102,n26);
nand (n1102,n808,n23);
xor (n1103,n1104,n26);
xor (n1104,n1006,n1010);
and (n1105,n1103,n1106);
xor (n1106,n1107,n1027);
xor (n1107,n1018,n1022);
and (n1108,n1101,n1106);
and (n1109,n1099,n1110);
xor (n1110,n1111,n969);
xor (n1111,n960,n964);
and (n1112,n1059,n1110);
and (n1113,n1114,n1116);
xor (n1114,n1115,n953);
xor (n1115,n944,n948);
xor (n1116,n1117,n1033);
xor (n1117,n1004,n1016);
and (n1118,n1113,n1119);
xor (n1119,n1120,n1041);
xor (n1120,n1002,n1038);
and (n1121,n1057,n1119);
and (n1122,n1123,n1124);
xor (n1123,n1053,n1055);
or (n1124,n1125,n1177);
and (n1125,n1126,n1128);
xor (n1126,n1127,n1119);
xor (n1127,n1057,n1113);
or (n1128,n1129,n1174,n1176);
and (n1129,n1130,n1172);
or (n1130,n1131,n1168,n1171);
and (n1131,n1132,n1166);
or (n1132,n1133,n1162,n1165);
and (n1133,n1134,n1150);
or (n1134,n1135,n1144,n1149);
and (n1135,n1136,n1140);
xnor (n1136,n1137,n278);
nor (n1137,n1138,n1139);
and (n1138,n339,n390);
and (n1139,n334,n393);
xnor (n1140,n1141,n173);
nor (n1141,n1142,n1143);
and (n1142,n492,n286);
and (n1143,n423,n289);
and (n1144,n1140,n1145);
xnor (n1145,n1146,n58);
nor (n1146,n1147,n1148);
and (n1147,n650,n181);
and (n1148,n556,n184);
and (n1149,n1136,n1145);
or (n1150,n1151,n1160,n1161);
and (n1151,n1152,n1156);
xnor (n1152,n1153,n386);
nor (n1153,n1154,n1155);
and (n1154,n131,n721);
and (n1155,n128,n723);
xnor (n1156,n1157,n382);
nor (n1157,n1158,n1159);
and (n1158,n223,n534);
and (n1159,n168,n537);
and (n1160,n1156,n8);
and (n1161,n1152,n8);
and (n1162,n1150,n1163);
xor (n1163,n1164,n1072);
xor (n1164,n1063,n1067);
and (n1165,n1134,n1163);
xor (n1166,n1167,n1094);
xor (n1167,n1061,n1077);
and (n1168,n1166,n1169);
xor (n1169,n1170,n1106);
xor (n1170,n1101,n1103);
and (n1171,n1132,n1169);
xor (n1172,n1173,n1110);
xor (n1173,n1059,n1099);
and (n1174,n1172,n1175);
xor (n1175,n1114,n1116);
and (n1176,n1130,n1175);
and (n1177,n1178,n1179);
xor (n1178,n1126,n1128);
or (n1179,n1180,n1218);
and (n1180,n1181,n1183);
xor (n1181,n1182,n1175);
xor (n1182,n1130,n1172);
and (n1183,n1184,n1216);
or (n1184,n1185,n1212,n1215);
and (n1185,n1186,n1210);
or (n1186,n1187,n1206,n1209);
and (n1187,n1188,n1204);
or (n1188,n1189,n1198,n1203);
and (n1189,n1190,n1194);
xnor (n1190,n1191,n386);
nor (n1191,n1192,n1193);
and (n1192,n168,n721);
and (n1193,n131,n723);
xnor (n1194,n1195,n382);
nor (n1195,n1196,n1197);
and (n1196,n334,n534);
and (n1197,n223,n537);
and (n1198,n1194,n1199);
xnor (n1199,n1200,n278);
nor (n1200,n1201,n1202);
and (n1201,n423,n390);
and (n1202,n339,n393);
and (n1203,n1190,n1199);
xnor (n1204,n1205,n8);
nand (n1205,n808,n69);
and (n1206,n1204,n1207);
xor (n1207,n1208,n1145);
xor (n1208,n1136,n1140);
and (n1209,n1188,n1207);
xor (n1210,n1211,n1088);
xor (n1211,n1079,n1083);
and (n1212,n1210,n1213);
xor (n1213,n1214,n1163);
xor (n1214,n1134,n1150);
and (n1215,n1186,n1213);
xor (n1216,n1217,n1169);
xor (n1217,n1132,n1166);
and (n1218,n1219,n1220);
xor (n1219,n1181,n1183);
or (n1220,n1221,n1273);
and (n1221,n1222,n1223);
xor (n1222,n1184,n1216);
and (n1223,n1224,n1271);
or (n1224,n1225,n1267,n1270);
and (n1225,n1226,n1260);
or (n1226,n1227,n1254,n1259);
and (n1227,n1228,n1242);
or (n1228,n1229,n1238,n1241);
and (n1229,n1230,n1234);
xnor (n1230,n1231,n278);
nor (n1231,n1232,n1233);
and (n1232,n492,n390);
and (n1233,n423,n393);
xnor (n1234,n1235,n173);
nor (n1235,n1236,n1237);
and (n1236,n650,n286);
and (n1237,n556,n289);
and (n1238,n1234,n1239);
xnor (n1239,n1240,n58);
nand (n1240,n808,n184);
and (n1241,n1230,n1239);
or (n1242,n1243,n1252,n1253);
and (n1243,n1244,n1248);
xnor (n1244,n1245,n386);
nor (n1245,n1246,n1247);
and (n1246,n223,n721);
and (n1247,n168,n723);
xnor (n1248,n1249,n382);
nor (n1249,n1250,n1251);
and (n1250,n339,n534);
and (n1251,n334,n537);
and (n1252,n1248,n58);
and (n1253,n1244,n58);
and (n1254,n1242,n1255);
xnor (n1255,n1256,n173);
nor (n1256,n1257,n1258);
and (n1257,n556,n286);
and (n1258,n492,n289);
and (n1259,n1228,n1255);
and (n1260,n1261,n1265);
xnor (n1261,n1262,n58);
nor (n1262,n1263,n1264);
and (n1263,n808,n181);
and (n1264,n650,n184);
xor (n1265,n1266,n1199);
xor (n1266,n1190,n1194);
and (n1267,n1260,n1268);
xor (n1268,n1269,n8);
xor (n1269,n1152,n1156);
and (n1270,n1226,n1268);
xor (n1271,n1272,n1213);
xor (n1272,n1186,n1210);
and (n1273,n1274,n1275);
xor (n1274,n1222,n1223);
or (n1275,n1276,n1283);
and (n1276,n1277,n1278);
xor (n1277,n1224,n1271);
and (n1278,n1279,n1281);
xor (n1279,n1280,n1207);
xor (n1280,n1188,n1204);
xor (n1281,n1282,n1268);
xor (n1282,n1226,n1260);
and (n1283,n1284,n1285);
xor (n1284,n1277,n1278);
or (n1285,n1286,n1319);
and (n1286,n1287,n1288);
xor (n1287,n1279,n1281);
or (n1288,n1289,n1316,n1318);
and (n1289,n1290,n1314);
or (n1290,n1291,n1310,n1313);
and (n1291,n1292,n1308);
or (n1292,n1293,n1302,n1307);
and (n1293,n1294,n1298);
xnor (n1294,n1295,n386);
nor (n1295,n1296,n1297);
and (n1296,n334,n721);
and (n1297,n223,n723);
xnor (n1298,n1299,n382);
nor (n1299,n1300,n1301);
and (n1300,n423,n534);
and (n1301,n339,n537);
and (n1302,n1298,n1303);
xnor (n1303,n1304,n278);
nor (n1304,n1305,n1306);
and (n1305,n556,n390);
and (n1306,n492,n393);
and (n1307,n1294,n1303);
xor (n1308,n1309,n1239);
xor (n1309,n1230,n1234);
and (n1310,n1308,n1311);
xor (n1311,n1312,n58);
xor (n1312,n1244,n1248);
and (n1313,n1292,n1311);
xor (n1314,n1315,n1255);
xor (n1315,n1228,n1242);
and (n1316,n1314,n1317);
xor (n1317,n1261,n1265);
and (n1318,n1290,n1317);
and (n1319,n1320,n1321);
xor (n1320,n1287,n1288);
or (n1321,n1322,n1355);
and (n1322,n1323,n1325);
xor (n1323,n1324,n1317);
xor (n1324,n1290,n1314);
and (n1325,n1326,n1353);
or (n1326,n1327,n1347,n1352);
and (n1327,n1328,n1340);
or (n1328,n1329,n1338,n1339);
and (n1329,n1330,n1334);
xnor (n1330,n1331,n386);
nor (n1331,n1332,n1333);
and (n1332,n339,n721);
and (n1333,n334,n723);
xnor (n1334,n1335,n382);
nor (n1335,n1336,n1337);
and (n1336,n492,n534);
and (n1337,n423,n537);
and (n1338,n1334,n173);
and (n1339,n1330,n173);
and (n1340,n1341,n1345);
xnor (n1341,n1342,n278);
nor (n1342,n1343,n1344);
and (n1343,n650,n390);
and (n1344,n556,n393);
xnor (n1345,n1346,n173);
nand (n1346,n808,n289);
and (n1347,n1340,n1348);
xnor (n1348,n1349,n173);
nor (n1349,n1350,n1351);
and (n1350,n808,n286);
and (n1351,n650,n289);
and (n1352,n1328,n1348);
xor (n1353,n1354,n1311);
xor (n1354,n1292,n1308);
and (n1355,n1356,n1357);
xor (n1356,n1323,n1325);
or (n1357,n1358,n1365);
and (n1358,n1359,n1360);
xor (n1359,n1326,n1353);
and (n1360,n1361,n1363);
xor (n1361,n1362,n1303);
xor (n1362,n1294,n1298);
xor (n1363,n1364,n1348);
xor (n1364,n1328,n1340);
and (n1365,n1366,n1367);
xor (n1366,n1359,n1360);
or (n1367,n1368,n1393);
and (n1368,n1369,n1370);
xor (n1369,n1361,n1363);
or (n1370,n1371,n1390,n1392);
and (n1371,n1372,n1388);
or (n1372,n1373,n1382,n1387);
and (n1373,n1374,n1378);
xnor (n1374,n1375,n386);
nor (n1375,n1376,n1377);
and (n1376,n423,n721);
and (n1377,n339,n723);
xnor (n1378,n1379,n382);
nor (n1379,n1380,n1381);
and (n1380,n556,n534);
and (n1381,n492,n537);
and (n1382,n1378,n1383);
xnor (n1383,n1384,n278);
nor (n1384,n1385,n1386);
and (n1385,n808,n390);
and (n1386,n650,n393);
and (n1387,n1374,n1383);
xor (n1388,n1389,n173);
xor (n1389,n1330,n1334);
and (n1390,n1388,n1391);
xor (n1391,n1341,n1345);
and (n1392,n1372,n1391);
and (n1393,n1394,n1395);
xor (n1394,n1369,n1370);
or (n1395,n1396,n1414);
and (n1396,n1397,n1399);
xor (n1397,n1398,n1391);
xor (n1398,n1372,n1388);
and (n1399,n1400,n1412);
or (n1400,n1401,n1410,n1411);
and (n1401,n1402,n1406);
xnor (n1402,n1403,n386);
nor (n1403,n1404,n1405);
and (n1404,n492,n721);
and (n1405,n423,n723);
xnor (n1406,n1407,n382);
nor (n1407,n1408,n1409);
and (n1408,n650,n534);
and (n1409,n556,n537);
and (n1410,n1406,n278);
and (n1411,n1402,n278);
xor (n1412,n1413,n1383);
xor (n1413,n1374,n1378);
and (n1414,n1415,n1416);
xor (n1415,n1397,n1399);
or (n1416,n1417,n1424);
and (n1417,n1418,n1419);
xor (n1418,n1400,n1412);
and (n1419,n1420,n1422);
xnor (n1420,n1421,n278);
nand (n1421,n808,n393);
xor (n1422,n1423,n278);
xor (n1423,n1402,n1406);
and (n1424,n1425,n1426);
xor (n1425,n1418,n1419);
or (n1426,n1427,n1438);
and (n1427,n1428,n1429);
xor (n1428,n1420,n1422);
and (n1429,n1430,n1434);
xnor (n1430,n1431,n386);
nor (n1431,n1432,n1433);
and (n1432,n556,n721);
and (n1433,n492,n723);
xnor (n1434,n1435,n382);
nor (n1435,n1436,n1437);
and (n1436,n808,n534);
and (n1437,n650,n537);
and (n1438,n1439,n1440);
xor (n1439,n1428,n1429);
or (n1440,n1441,n1448);
and (n1441,n1442,n1443);
xor (n1442,n1430,n1434);
and (n1443,n1444,n382);
xnor (n1444,n1445,n386);
nor (n1445,n1446,n1447);
and (n1446,n650,n721);
and (n1447,n556,n723);
and (n1448,n1449,n1450);
xor (n1449,n1442,n1443);
or (n1450,n1451,n1455);
and (n1451,n1452,n1454);
xnor (n1452,n1453,n382);
nand (n1453,n808,n537);
xor (n1454,n1444,n382);
and (n1455,n1456,n1457);
xor (n1456,n1452,n1454);
and (n1457,n1458,n1462);
xnor (n1458,n1459,n386);
nor (n1459,n1460,n1461);
and (n1460,n808,n721);
and (n1461,n650,n723);
and (n1462,n1463,n386);
xnor (n1463,n1464,n386);
nand (n1464,n808,n723);
xor (n1465,n1466,n1508);
xor (n1466,n1467,n1479);
xor (n1467,n1468,n1478);
xor (n1468,n1469,n1472);
or (n1469,n98,n1470,n1471);
and (n1470,n87,n49);
and (n1471,n84,n49);
or (n1472,n1473,n1476);
or (n1473,n1474,n29,n1475);
and (n1474,n83,n14);
and (n1475,n83,n30);
xor (n1476,n1477,n49);
xor (n1477,n84,n87);
not (n1478,n100);
or (n1479,n1480,n1505,n1507);
and (n1480,n1481,n1488);
or (n1481,n1482,n1486,n1487);
and (n1482,n1483,n139);
or (n1483,n70,n1484,n1485);
and (n1484,n71,n133);
and (n1485,n63,n133);
and (n1486,n139,n46);
and (n1487,n1483,n46);
or (n1488,n1489,n1501,n1504);
and (n1489,n1490,n1500);
or (n1490,n1491,n1497,n1499);
and (n1491,n1492,n1495);
or (n1492,n1493,n118,n1494);
and (n1493,n57,n114);
and (n1494,n57,n119);
xor (n1495,n1496,n133);
xor (n1496,n63,n71);
and (n1497,n1495,n1498);
not (n1498,n139);
and (n1499,n1492,n1498);
not (n1500,n76);
and (n1501,n1500,n1502);
xor (n1502,n1503,n46);
xor (n1503,n1483,n139);
and (n1504,n1490,n1502);
and (n1505,n1488,n1506);
xnor (n1506,n1473,n1476);
and (n1507,n1481,n1506);
or (n1508,n1509,n1531);
and (n1509,n1510,n1512);
xor (n1510,n1511,n1506);
xor (n1511,n1481,n1488);
and (n1512,n1513,n1529);
or (n1513,n1514,n1525,n1528);
and (n1514,n1515,n1523);
or (n1515,n1516,n1521,n1522);
and (n1516,n1517,n1520);
or (n1517,n185,n1518,n1519);
and (n1518,n186,n158);
and (n1519,n178,n158);
or (n1520,n162,n167);
and (n1521,n1520,n125);
and (n1522,n1517,n125);
and (n1523,n130,n1524);
not (n1524,n241);
and (n1525,n1523,n1526);
xor (n1526,n1527,n1498);
xor (n1527,n1492,n1495);
and (n1528,n1515,n1526);
xor (n1529,n1530,n1502);
xor (n1530,n1490,n1500);
and (n1531,n1532,n1533);
xor (n1532,n1510,n1512);
or (n1533,n1534,n1554);
and (n1534,n1535,n1536);
xor (n1535,n1513,n1529);
and (n1536,n1537,n1552);
or (n1537,n1538,n1549,n1551);
and (n1538,n1539,n1547);
or (n1539,n1540,n1544,n1546);
and (n1540,n211,n1541);
or (n1541,n1542,n231,n1543);
and (n1542,n172,n227);
and (n1543,n172,n232);
and (n1544,n1541,n1545);
xnor (n1545,n162,n167);
and (n1546,n211,n1545);
xor (n1547,n1548,n125);
xor (n1548,n1517,n1520);
and (n1549,n1547,n1550);
xor (n1550,n130,n1524);
and (n1551,n1539,n1550);
xor (n1552,n1553,n1526);
xor (n1553,n1515,n1523);
and (n1554,n1555,n1556);
xor (n1555,n1535,n1536);
or (n1556,n1557,n1580);
and (n1557,n1558,n1559);
xor (n1558,n1537,n1552);
and (n1559,n1560,n1578);
or (n1560,n1561,n1574,n1577);
and (n1561,n1562,n1572);
or (n1562,n1563,n1570,n1571);
and (n1563,n1564,n1567);
or (n1564,n269,n1565,n1566);
and (n1565,n270,n343);
and (n1566,n265,n343);
or (n1567,n290,n1568,n1569);
and (n1568,n291,n261);
and (n1569,n283,n261);
and (n1570,n1567,n351);
and (n1571,n1564,n351);
xor (n1572,n1573,n158);
xor (n1573,n178,n186);
and (n1574,n1572,n1575);
xor (n1575,n1576,n1545);
xor (n1576,n211,n1541);
and (n1577,n1562,n1575);
xor (n1578,n1579,n1550);
xor (n1579,n1539,n1547);
and (n1580,n1581,n1582);
xor (n1581,n1558,n1559);
or (n1582,n1583,n1632);
and (n1583,n1584,n1585);
xor (n1584,n1560,n1578);
or (n1585,n1586,n1628,n1631);
and (n1586,n1587,n1598);
or (n1587,n1588,n1594,n1597);
and (n1588,n1589,n1593);
or (n1589,n1590,n320);
or (n1590,n1591,n314,n1592);
and (n1591,n277,n310);
and (n1592,n277,n315);
not (n1593,n355);
and (n1594,n1593,n1595);
xor (n1595,n1596,n351);
xor (n1596,n1564,n1567);
and (n1597,n1589,n1595);
or (n1598,n1599,n1624,n1627);
and (n1599,n1600,n1620);
or (n1600,n1601,n1616,n1619);
and (n1601,n1602,n1612);
or (n1602,n1603,n1610,n1611);
and (n1603,n1604,n1607);
or (n1604,n394,n1605,n1606);
and (n1605,n395,n402);
and (n1606,n387,n402);
or (n1607,n410,n1608,n1609);
and (n1608,n411,n418);
and (n1609,n406,n418);
and (n1610,n1607,n422);
and (n1611,n1604,n422);
or (n1612,n1613,n1614,n1615);
and (n1613,n338,n506);
and (n1614,n506,n429);
and (n1615,n338,n429);
and (n1616,n1612,n1617);
xor (n1617,n1618,n343);
xor (n1618,n265,n270);
and (n1619,n1602,n1617);
and (n1620,n1621,n1623);
xor (n1621,n1622,n261);
xor (n1622,n283,n291);
xnor (n1623,n1590,n320);
and (n1624,n1620,n1625);
xor (n1625,n1626,n1595);
xor (n1626,n1589,n1593);
and (n1627,n1600,n1625);
and (n1628,n1598,n1629);
xor (n1629,n1630,n1575);
xor (n1630,n1562,n1572);
and (n1631,n1587,n1629);
and (n1632,n1633,n1634);
xor (n1633,n1584,n1585);
or (n1634,n1635,n1669);
and (n1635,n1636,n1638);
xor (n1636,n1637,n1629);
xor (n1637,n1587,n1598);
and (n1638,n1639,n1667);
or (n1639,n1640,n1664,n1666);
and (n1640,n1641,n1662);
or (n1641,n1642,n1660,n1661);
and (n1642,n1643,n1651);
or (n1643,n1644,n1648,n1650);
and (n1644,n1645,n469);
or (n1645,n1646,n463,n1647);
and (n1646,n381,n459);
and (n1647,n381,n464);
and (n1648,n469,n1649);
and (n1649,n487,n491);
and (n1650,n1645,n1649);
or (n1651,n1652,n1657,n1659);
and (n1652,n1653,n1655);
xor (n1653,n1654,n402);
xor (n1654,n387,n395);
xor (n1655,n1656,n418);
xor (n1656,n406,n411);
and (n1657,n1655,n1658);
not (n1658,n422);
and (n1659,n1653,n1658);
and (n1660,n1651,n504);
and (n1661,n1643,n504);
xor (n1662,n1663,n1617);
xor (n1663,n1602,n1612);
and (n1664,n1662,n1665);
xor (n1665,n1621,n1623);
and (n1666,n1641,n1665);
xor (n1667,n1668,n1625);
xor (n1668,n1600,n1620);
and (n1669,n1670,n1671);
xor (n1670,n1636,n1638);
or (n1671,n1672,n1706);
and (n1672,n1673,n1674);
xor (n1673,n1639,n1667);
and (n1674,n1675,n1704);
or (n1675,n1676,n1700,n1703);
and (n1676,n1677,n1698);
or (n1677,n1678,n1694,n1697);
and (n1678,n1679,n1690);
or (n1679,n1680,n1687,n1689);
and (n1680,n1681,n1684);
or (n1681,n538,n1682,n1683);
and (n1682,n539,n561);
and (n1683,n531,n561);
or (n1684,n569,n1685,n1686);
and (n1685,n570,n546);
and (n1686,n565,n546);
and (n1687,n1684,n1688);
or (n1688,n550,n555);
and (n1689,n1681,n1688);
or (n1690,n1691,n1692,n1693);
and (n1691,n661,n580);
and (n1692,n580,n662);
and (n1693,n661,n662);
and (n1694,n1690,n1695);
xor (n1695,n1696,n1658);
xor (n1696,n1653,n1655);
and (n1697,n1679,n1695);
xor (n1698,n1699,n422);
xor (n1699,n1604,n1607);
and (n1700,n1698,n1701);
xor (n1701,n1702,n504);
xor (n1702,n1643,n1651);
and (n1703,n1677,n1701);
xor (n1704,n1705,n1665);
xor (n1705,n1641,n1662);
and (n1706,n1707,n1708);
xor (n1707,n1673,n1674);
or (n1708,n1709,n1741);
and (n1709,n1710,n1711);
xor (n1710,n1675,n1704);
and (n1711,n1712,n1739);
or (n1712,n1713,n1735,n1738);
and (n1713,n1714,n1733);
or (n1714,n1715,n1731,n1732);
and (n1715,n1716,n1722);
or (n1716,n1717,n1721,n652);
and (n1717,n609,n1718);
or (n1718,n1719,n631,n1720);
and (n1719,n530,n627);
and (n1720,n530,n632);
and (n1721,n1718,n638);
or (n1722,n1723,n1728,n1730);
and (n1723,n1724,n1726);
xor (n1724,n1725,n561);
xor (n1725,n531,n539);
xor (n1726,n1727,n546);
xor (n1727,n565,n570);
and (n1728,n1726,n1729);
xnor (n1729,n550,n555);
and (n1730,n1724,n1729);
and (n1731,n1722,n659);
and (n1732,n1716,n659);
xor (n1733,n1734,n1649);
xor (n1734,n1645,n469);
and (n1735,n1733,n1736);
xor (n1736,n1737,n1695);
xor (n1737,n1679,n1690);
and (n1738,n1714,n1736);
xor (n1739,n1740,n1701);
xor (n1740,n1677,n1698);
and (n1741,n1742,n1743);
xor (n1742,n1710,n1711);
or (n1743,n1744,n1764);
and (n1744,n1745,n1746);
xor (n1745,n1712,n1739);
and (n1746,n1747,n1762);
or (n1747,n1748,n1758,n1761);
and (n1748,n1749,n1756);
or (n1749,n1750,n1752,n1755);
and (n1750,n682,n1751);
or (n1751,n732,n737);
and (n1752,n1751,n1753);
xor (n1753,n1754,n1729);
xor (n1754,n1724,n1726);
and (n1755,n682,n1753);
xor (n1756,n1757,n1688);
xor (n1757,n1681,n1684);
and (n1758,n1756,n1759);
xor (n1759,n1760,n659);
xor (n1760,n1716,n1722);
and (n1761,n1749,n1759);
xor (n1762,n1763,n1736);
xor (n1763,n1714,n1733);
and (n1764,n1765,n1766);
xor (n1765,n1745,n1746);
or (n1766,n1767,n1783);
and (n1767,n1768,n1769);
xor (n1768,n1747,n1762);
and (n1769,n1770,n1781);
or (n1770,n1771,n1777,n1780);
and (n1771,n1772,n1775);
or (n1772,n764,n1773,n1774);
and (n1773,n811,n933);
and (n1774,n765,n933);
xor (n1775,n1776,n638);
xor (n1776,n609,n1718);
and (n1777,n1775,n1778);
xor (n1778,n1779,n1753);
xor (n1779,n682,n1751);
and (n1780,n1772,n1778);
xor (n1781,n1782,n1759);
xor (n1782,n1749,n1756);
and (n1783,n1784,n1785);
xor (n1784,n1768,n1769);
or (n1785,n1786,n1794);
and (n1786,n1787,n1788);
xor (n1787,n1770,n1781);
and (n1788,n1789,n1792);
or (n1789,n844,n1790,n1791);
and (n1790,n905,n935);
and (n1791,n845,n935);
xor (n1792,n1793,n1778);
xor (n1793,n1772,n1775);
and (n1794,n1795,n1796);
xor (n1795,n1787,n1788);
or (n1796,n1797,n926);
and (n1797,n1798,n1799);
xor (n1798,n1789,n1792);
or (n1799,n1800,n1801,n1802);
and (n1800,n911,n932);
and (n1801,n932,n934);
and (n1802,n911,n934);
endmodule
