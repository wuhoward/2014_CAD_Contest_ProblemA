module top (out,n12,n15,n16,n20,n23,n24,n28,n36,n39
        ,n40,n44,n54,n57,n58,n62,n69,n72,n73,n77
        ,n85,n88,n89,n93,n103,n106,n107,n111,n116,n323
        ,n415,n488,n573);
output out;
input n12;
input n15;
input n16;
input n20;
input n23;
input n24;
input n28;
input n36;
input n39;
input n40;
input n44;
input n54;
input n57;
input n58;
input n62;
input n69;
input n72;
input n73;
input n77;
input n85;
input n88;
input n89;
input n93;
input n103;
input n106;
input n107;
input n111;
input n116;
input n323;
input n415;
input n488;
input n573;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n17;
wire n18;
wire n19;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
xor (out,n0,n1230);
xor (n0,n1,n364);
xor (n1,n2,n288);
xor (n2,n3,n241);
or (n3,n4,n192,n240);
and (n4,n5,n182);
or (n5,n6,n152,n181);
and (n6,n7,n118);
or (n7,n8,n98,n117);
and (n8,n9,n49);
or (n9,n10,n32,n48);
and (n10,n11,n17);
and (n11,n12,n13);
not (n13,n14);
and (n14,n15,n16);
xnor (n17,n18,n29);
nor (n18,n19,n27);
and (n19,n20,n21);
and (n21,n22,n25);
xor (n22,n23,n24);
not (n25,n26);
xor (n26,n24,n12);
and (n27,n28,n26);
and (n29,n23,n30);
not (n30,n31);
and (n31,n24,n12);
and (n32,n17,n33);
xnor (n33,n34,n45);
nor (n34,n35,n43);
and (n35,n36,n37);
and (n37,n38,n41);
xor (n38,n39,n40);
not (n41,n42);
xor (n42,n40,n23);
and (n43,n44,n42);
and (n45,n39,n46);
not (n46,n47);
and (n47,n40,n23);
and (n48,n11,n33);
or (n49,n50,n81,n97);
and (n50,n51,n66);
xnor (n51,n52,n63);
nor (n52,n53,n61);
and (n53,n54,n55);
and (n55,n56,n59);
xor (n56,n57,n58);
not (n59,n60);
xor (n60,n58,n39);
and (n61,n62,n60);
and (n63,n57,n64);
not (n64,n65);
and (n65,n58,n39);
xnor (n66,n67,n78);
nor (n67,n68,n76);
and (n68,n69,n70);
and (n70,n71,n74);
xor (n71,n72,n73);
not (n74,n75);
xor (n75,n73,n57);
and (n76,n77,n75);
and (n78,n72,n79);
not (n79,n80);
and (n80,n73,n57);
and (n81,n66,n82);
xnor (n82,n83,n94);
nor (n83,n84,n92);
and (n84,n85,n86);
and (n86,n87,n90);
xor (n87,n88,n89);
not (n90,n91);
xor (n91,n89,n72);
and (n92,n93,n91);
and (n94,n88,n95);
not (n95,n96);
and (n96,n89,n72);
and (n97,n51,n82);
and (n98,n49,n99);
or (n99,n100,n115);
xnor (n100,n101,n112);
nor (n101,n102,n110);
and (n102,n103,n104);
and (n104,n105,n108);
xor (n105,n106,n107);
not (n108,n109);
xor (n109,n107,n88);
and (n110,n111,n109);
and (n112,n106,n113);
not (n113,n114);
and (n114,n107,n88);
and (n115,n116,n106);
and (n117,n9,n99);
or (n118,n119,n144,n151);
and (n119,n120,n130);
xor (n120,n121,n126);
xor (n121,n122,n123);
not (n122,n11);
xnor (n123,n124,n29);
not (n124,n125);
and (n125,n28,n21);
xnor (n126,n127,n45);
nor (n127,n128,n129);
and (n128,n44,n37);
and (n129,n20,n42);
xor (n130,n131,n140);
xor (n131,n132,n136);
xnor (n132,n133,n63);
nor (n133,n134,n135);
and (n134,n62,n55);
and (n135,n36,n60);
xnor (n136,n137,n78);
nor (n137,n138,n139);
and (n138,n77,n70);
and (n139,n54,n75);
xnor (n140,n141,n94);
nor (n141,n142,n143);
and (n142,n93,n86);
and (n143,n69,n91);
and (n144,n130,n145);
xor (n145,n146,n150);
xnor (n146,n147,n112);
nor (n147,n148,n149);
and (n148,n111,n104);
and (n149,n85,n109);
and (n150,n103,n106);
and (n151,n120,n145);
and (n152,n118,n153);
xor (n153,n154,n167);
xor (n154,n155,n156);
and (n155,n111,n106);
not (n156,n157);
xor (n157,n158,n163);
xor (n158,n29,n159);
xnor (n159,n160,n45);
nor (n160,n161,n162);
and (n161,n20,n37);
and (n162,n28,n42);
xnor (n163,n164,n63);
nor (n164,n165,n166);
and (n165,n36,n55);
and (n166,n44,n60);
xor (n167,n168,n177);
xor (n168,n169,n173);
xnor (n169,n170,n78);
nor (n170,n171,n172);
and (n171,n54,n70);
and (n172,n62,n75);
xnor (n173,n174,n94);
nor (n174,n175,n176);
and (n175,n69,n86);
and (n176,n77,n91);
xnor (n177,n178,n112);
nor (n178,n179,n180);
and (n179,n85,n104);
and (n180,n93,n109);
and (n181,n7,n153);
xor (n182,n183,n155);
xor (n183,n184,n188);
or (n184,n185,n186,n187);
and (n185,n29,n159);
and (n186,n159,n163);
and (n187,n29,n163);
or (n188,n189,n190,n191);
and (n189,n169,n173);
and (n190,n173,n177);
and (n191,n169,n177);
and (n192,n182,n193);
xor (n193,n194,n213);
xor (n194,n195,n208);
or (n195,n196,n205,n207);
and (n196,n197,n201);
or (n197,n198,n199,n200);
and (n198,n122,n123);
and (n199,n123,n126);
and (n200,n122,n126);
or (n201,n202,n203,n204);
and (n202,n132,n136);
and (n203,n136,n140);
and (n204,n132,n140);
and (n205,n201,n206);
and (n206,n146,n150);
and (n207,n197,n206);
or (n208,n209,n210,n212);
and (n209,n157,n167);
and (n210,n167,n211);
not (n211,n155);
and (n212,n157,n211);
xor (n213,n214,n230);
xor (n214,n215,n216);
and (n215,n85,n106);
xor (n216,n217,n226);
xor (n217,n218,n222);
xnor (n218,n219,n78);
nor (n219,n220,n221);
and (n220,n62,n70);
and (n221,n36,n75);
xnor (n222,n223,n94);
nor (n223,n224,n225);
and (n224,n77,n86);
and (n225,n54,n91);
xnor (n226,n227,n112);
nor (n227,n228,n229);
and (n228,n93,n104);
and (n229,n69,n109);
xor (n230,n231,n236);
xor (n231,n232,n233);
not (n232,n29);
xnor (n233,n234,n45);
not (n234,n235);
and (n235,n28,n37);
xnor (n236,n237,n63);
nor (n237,n238,n239);
and (n238,n44,n55);
and (n239,n20,n60);
and (n240,n5,n193);
xor (n241,n242,n268);
xor (n242,n243,n247);
or (n243,n244,n245,n246);
and (n244,n195,n208);
and (n245,n208,n213);
and (n246,n195,n213);
xor (n247,n248,n257);
xor (n248,n249,n253);
or (n249,n250,n251,n252);
and (n250,n184,n188);
and (n251,n188,n155);
and (n252,n184,n155);
or (n253,n254,n255,n256);
and (n254,n215,n216);
and (n255,n216,n230);
and (n256,n215,n230);
xor (n257,n258,n267);
xor (n258,n259,n263);
xnor (n259,n260,n94);
nor (n260,n261,n262);
and (n261,n54,n86);
and (n262,n62,n91);
xnor (n263,n264,n112);
nor (n264,n265,n266);
and (n265,n69,n104);
and (n266,n77,n109);
and (n267,n93,n106);
xor (n268,n269,n279);
xor (n269,n270,n275);
xor (n270,n45,n271);
xnor (n271,n272,n63);
nor (n272,n273,n274);
and (n273,n20,n55);
and (n274,n28,n60);
xnor (n275,n276,n78);
nor (n276,n277,n278);
and (n277,n36,n70);
and (n278,n44,n75);
xnor (n279,n280,n284);
or (n280,n281,n282,n283);
and (n281,n218,n222);
and (n282,n222,n226);
and (n283,n218,n226);
or (n284,n285,n286,n287);
and (n285,n232,n233);
and (n286,n233,n236);
and (n287,n232,n236);
and (n288,n289,n362);
or (n289,n290,n358,n361);
and (n290,n291,n356);
or (n291,n292,n352,n355);
and (n292,n293,n343);
or (n293,n294,n325,n342);
and (n294,n295,n311);
or (n295,n296,n305,n310);
and (n296,n297,n298);
not (n297,n16);
xnor (n298,n299,n11);
not (n299,n300);
and (n300,n28,n301);
and (n301,n302,n303);
xor (n302,n12,n15);
not (n303,n304);
xor (n304,n15,n16);
and (n305,n298,n306);
xnor (n306,n307,n29);
nor (n307,n308,n309);
and (n308,n44,n21);
and (n309,n20,n26);
and (n310,n297,n306);
or (n311,n312,n321,n324);
and (n312,n313,n317);
xnor (n313,n314,n94);
nor (n314,n315,n316);
and (n315,n111,n86);
and (n316,n85,n91);
xnor (n317,n318,n112);
nor (n318,n319,n320);
and (n319,n116,n104);
and (n320,n103,n109);
and (n321,n317,n322);
and (n322,n323,n106);
and (n324,n313,n322);
and (n325,n311,n326);
or (n326,n327,n336,n341);
and (n327,n328,n332);
xnor (n328,n329,n45);
nor (n329,n330,n331);
and (n330,n62,n37);
and (n331,n36,n42);
xnor (n332,n333,n63);
nor (n333,n334,n335);
and (n334,n77,n55);
and (n335,n54,n60);
and (n336,n332,n337);
xnor (n337,n338,n78);
nor (n338,n339,n340);
and (n339,n93,n70);
and (n340,n69,n75);
and (n341,n328,n337);
and (n342,n295,n326);
or (n343,n344,n349,n351);
and (n344,n345,n347);
xor (n345,n346,n33);
xor (n346,n11,n17);
xor (n347,n348,n82);
xor (n348,n51,n66);
and (n349,n347,n350);
xnor (n350,n100,n115);
and (n351,n345,n350);
and (n352,n343,n353);
xor (n353,n354,n145);
xor (n354,n120,n130);
and (n355,n293,n353);
xor (n356,n357,n206);
xor (n357,n197,n201);
and (n358,n356,n359);
xor (n359,n360,n153);
xor (n360,n7,n118);
and (n361,n291,n359);
xor (n362,n363,n193);
xor (n363,n5,n182);
or (n364,n365,n437);
and (n365,n366,n367);
xor (n366,n289,n362);
and (n367,n368,n435);
or (n368,n369,n431,n434);
and (n369,n370,n429);
or (n370,n371,n423,n428);
and (n371,n372,n418);
or (n372,n373,n402,n417);
and (n373,n374,n390);
or (n374,n375,n384,n389);
and (n375,n376,n380);
xnor (n376,n377,n45);
nor (n377,n378,n379);
and (n378,n54,n37);
and (n379,n62,n42);
xnor (n380,n381,n63);
nor (n381,n382,n383);
and (n382,n69,n55);
and (n383,n77,n60);
and (n384,n380,n385);
xnor (n385,n386,n78);
nor (n386,n387,n388);
and (n387,n85,n70);
and (n388,n93,n75);
and (n389,n376,n385);
or (n390,n391,n396,n401);
and (n391,n16,n392);
xnor (n392,n393,n11);
nor (n393,n394,n395);
and (n394,n20,n301);
and (n395,n28,n304);
and (n396,n392,n397);
xnor (n397,n398,n29);
nor (n398,n399,n400);
and (n399,n36,n21);
and (n400,n44,n26);
and (n401,n16,n397);
and (n402,n390,n403);
or (n403,n404,n413,n416);
and (n404,n405,n409);
xnor (n405,n406,n94);
nor (n406,n407,n408);
and (n407,n103,n86);
and (n408,n111,n91);
xnor (n409,n410,n112);
nor (n410,n411,n412);
and (n411,n323,n104);
and (n412,n116,n109);
and (n413,n409,n414);
and (n414,n415,n106);
and (n416,n405,n414);
and (n417,n374,n403);
or (n418,n419,n421);
xor (n419,n420,n322);
xor (n420,n313,n317);
xor (n421,n422,n337);
xor (n422,n328,n332);
and (n423,n418,n424);
xor (n424,n425,n427);
xor (n425,n426,n347);
not (n426,n345);
not (n427,n350);
and (n428,n372,n424);
xor (n429,n430,n99);
xor (n430,n9,n49);
and (n431,n429,n432);
xor (n432,n433,n353);
xor (n433,n293,n343);
and (n434,n370,n432);
xor (n435,n436,n359);
xor (n436,n291,n356);
and (n437,n438,n439);
xor (n438,n366,n367);
or (n439,n440,n519);
and (n440,n441,n442);
xor (n441,n368,n435);
and (n442,n443,n517);
or (n443,n444,n513,n516);
and (n444,n445,n509);
or (n445,n446,n505,n508);
and (n446,n447,n495);
or (n447,n448,n481,n494);
and (n448,n449,n465);
or (n449,n450,n459,n464);
and (n450,n451,n455);
xnor (n451,n452,n29);
nor (n452,n453,n454);
and (n453,n62,n21);
and (n454,n36,n26);
xnor (n455,n456,n45);
nor (n456,n457,n458);
and (n457,n77,n37);
and (n458,n54,n42);
and (n459,n455,n460);
xnor (n460,n461,n63);
nor (n461,n462,n463);
and (n462,n93,n55);
and (n463,n69,n60);
and (n464,n451,n460);
or (n465,n466,n475,n480);
and (n466,n467,n471);
xnor (n467,n468,n78);
nor (n468,n469,n470);
and (n469,n111,n70);
and (n470,n85,n75);
xnor (n471,n472,n94);
nor (n472,n473,n474);
and (n473,n116,n86);
and (n474,n103,n91);
and (n475,n471,n476);
xnor (n476,n477,n112);
nor (n477,n478,n479);
and (n478,n415,n104);
and (n479,n323,n109);
and (n480,n467,n476);
and (n481,n465,n482);
and (n482,n483,n490);
xnor (n483,n484,n16);
not (n484,n485);
and (n485,n28,n486);
and (n486,n487,n489);
xor (n487,n16,n488);
not (n489,n488);
xnor (n490,n491,n11);
nor (n491,n492,n493);
and (n492,n44,n301);
and (n493,n20,n304);
and (n494,n449,n482);
or (n495,n496,n501,n504);
and (n496,n497,n499);
xor (n497,n498,n385);
xor (n498,n376,n380);
xor (n499,n500,n397);
xor (n500,n16,n392);
and (n501,n499,n502);
xor (n502,n503,n414);
xor (n503,n405,n409);
and (n504,n497,n502);
and (n505,n495,n506);
xor (n506,n507,n306);
xor (n507,n297,n298);
and (n508,n447,n506);
and (n509,n510,n512);
xor (n510,n511,n403);
xor (n511,n374,n390);
xnor (n512,n419,n421);
and (n513,n509,n514);
xor (n514,n515,n326);
xor (n515,n295,n311);
and (n516,n445,n514);
xor (n517,n518,n432);
xor (n518,n370,n429);
and (n519,n520,n521);
xor (n520,n441,n442);
or (n521,n522,n601);
and (n522,n523,n524);
xor (n523,n443,n517);
or (n524,n525,n597,n600);
and (n525,n526,n595);
or (n526,n527,n592,n594);
and (n527,n528,n590);
or (n528,n529,n586,n589);
and (n529,n530,n576);
or (n530,n531,n564,n575);
and (n531,n532,n548);
or (n532,n533,n542,n547);
and (n533,n534,n538);
xnor (n534,n535,n16);
nor (n535,n536,n537);
and (n536,n20,n486);
and (n537,n28,n488);
xnor (n538,n539,n11);
nor (n539,n540,n541);
and (n540,n36,n301);
and (n541,n44,n304);
and (n542,n538,n543);
xnor (n543,n544,n29);
nor (n544,n545,n546);
and (n545,n54,n21);
and (n546,n62,n26);
and (n547,n534,n543);
or (n548,n549,n558,n563);
and (n549,n550,n554);
xnor (n550,n551,n45);
nor (n551,n552,n553);
and (n552,n69,n37);
and (n553,n77,n42);
xnor (n554,n555,n63);
nor (n555,n556,n557);
and (n556,n85,n55);
and (n557,n93,n60);
and (n558,n554,n559);
xnor (n559,n560,n78);
nor (n560,n561,n562);
and (n561,n103,n70);
and (n562,n111,n75);
and (n563,n550,n559);
and (n564,n548,n565);
and (n565,n566,n570);
xnor (n566,n567,n94);
nor (n567,n568,n569);
and (n568,n323,n86);
and (n569,n116,n91);
xnor (n570,n571,n112);
nor (n571,n572,n574);
and (n572,n573,n104);
and (n574,n415,n109);
and (n575,n532,n565);
or (n576,n577,n582,n585);
and (n577,n578,n580);
not (n578,n579);
nand (n579,n573,n106);
xor (n580,n581,n460);
xor (n581,n451,n455);
and (n582,n580,n583);
xor (n583,n584,n476);
xor (n584,n467,n471);
and (n585,n578,n583);
and (n586,n576,n587);
xor (n587,n588,n502);
xor (n588,n497,n499);
and (n589,n530,n587);
xor (n590,n591,n506);
xor (n591,n447,n495);
and (n592,n590,n593);
xor (n593,n510,n512);
and (n594,n528,n593);
xor (n595,n596,n514);
xor (n596,n445,n509);
and (n597,n595,n598);
xor (n598,n599,n424);
xor (n599,n372,n418);
and (n600,n526,n598);
and (n601,n602,n603);
xor (n602,n523,n524);
or (n603,n604,n681);
and (n604,n605,n607);
xor (n605,n606,n598);
xor (n606,n526,n595);
and (n607,n608,n679);
or (n608,n609,n675,n678);
and (n609,n610,n670);
or (n610,n611,n667,n669);
and (n611,n612,n658);
or (n612,n613,n640,n657);
and (n613,n614,n628);
or (n614,n615,n624,n627);
and (n615,n616,n620);
xnor (n616,n617,n78);
nor (n617,n618,n619);
and (n618,n116,n70);
and (n619,n103,n75);
xnor (n620,n621,n94);
nor (n621,n622,n623);
and (n622,n415,n86);
and (n623,n323,n91);
and (n624,n620,n625);
xnor (n625,n626,n112);
nand (n626,n573,n109);
and (n627,n616,n625);
or (n628,n629,n638,n639);
and (n629,n630,n634);
xnor (n630,n631,n16);
nor (n631,n632,n633);
and (n632,n44,n486);
and (n633,n20,n488);
xnor (n634,n635,n11);
nor (n635,n636,n637);
and (n636,n62,n301);
and (n637,n36,n304);
and (n638,n634,n112);
and (n639,n630,n112);
and (n640,n628,n641);
or (n641,n642,n651,n656);
and (n642,n643,n647);
xnor (n643,n644,n29);
nor (n644,n645,n646);
and (n645,n77,n21);
and (n646,n54,n26);
xnor (n647,n648,n45);
nor (n648,n649,n650);
and (n649,n93,n37);
and (n650,n69,n42);
and (n651,n647,n652);
xnor (n652,n653,n63);
nor (n653,n654,n655);
and (n654,n111,n55);
and (n655,n85,n60);
and (n656,n643,n652);
and (n657,n614,n641);
or (n658,n659,n664,n666);
and (n659,n660,n662);
xor (n660,n661,n543);
xor (n661,n534,n538);
xor (n662,n663,n559);
xor (n663,n550,n554);
and (n664,n662,n665);
xor (n665,n566,n570);
and (n666,n660,n665);
and (n667,n658,n668);
xor (n668,n483,n490);
and (n669,n612,n668);
and (n670,n671,n673);
xor (n671,n672,n565);
xor (n672,n532,n548);
xor (n673,n674,n583);
xor (n674,n578,n580);
and (n675,n670,n676);
xor (n676,n677,n482);
xor (n677,n449,n465);
and (n678,n610,n676);
xor (n679,n680,n593);
xor (n680,n528,n590);
and (n681,n682,n683);
xor (n682,n605,n607);
or (n683,n684,n691);
and (n684,n685,n686);
xor (n685,n608,n679);
and (n686,n687,n689);
xor (n687,n688,n676);
xor (n688,n610,n670);
xor (n689,n690,n587);
xor (n690,n530,n576);
and (n691,n692,n693);
xor (n692,n685,n686);
or (n693,n694,n757);
and (n694,n695,n701);
xor (n695,n696,n699);
xor (n696,n676,n697);
xor (n697,n690,n698);
not (n698,n499);
xor (n699,n688,n700);
xnor (n700,n497,n502);
or (n701,n702,n754,n756);
and (n702,n703,n752);
or (n703,n704,n748,n751);
and (n704,n705,n743);
or (n705,n706,n739,n742);
and (n706,n707,n723);
or (n707,n708,n717,n722);
and (n708,n709,n713);
xnor (n709,n710,n16);
nor (n710,n711,n712);
and (n711,n36,n486);
and (n712,n44,n488);
xnor (n713,n714,n11);
nor (n714,n715,n716);
and (n715,n54,n301);
and (n716,n62,n304);
and (n717,n713,n718);
xnor (n718,n719,n29);
nor (n719,n720,n721);
and (n720,n69,n21);
and (n721,n77,n26);
and (n722,n709,n718);
or (n723,n724,n733,n738);
and (n724,n725,n729);
xnor (n725,n726,n45);
nor (n726,n727,n728);
and (n727,n85,n37);
and (n728,n93,n42);
xnor (n729,n730,n63);
nor (n730,n731,n732);
and (n731,n103,n55);
and (n732,n111,n60);
and (n733,n729,n734);
xnor (n734,n735,n78);
nor (n735,n736,n737);
and (n736,n323,n70);
and (n737,n116,n75);
and (n738,n725,n734);
and (n739,n723,n740);
xor (n740,n741,n625);
xor (n741,n616,n620);
and (n742,n707,n740);
and (n743,n744,n746);
xor (n744,n745,n112);
xor (n745,n630,n634);
xor (n746,n747,n652);
xor (n747,n643,n647);
and (n748,n743,n749);
xor (n749,n750,n665);
xor (n750,n660,n662);
and (n751,n705,n749);
xor (n752,n753,n668);
xor (n753,n612,n658);
and (n754,n752,n755);
xor (n755,n671,n673);
and (n756,n703,n755);
and (n757,n758,n759);
xor (n758,n695,n701);
or (n759,n760,n814);
and (n760,n761,n763);
xor (n761,n762,n755);
xor (n762,n703,n752);
or (n763,n764,n810,n813);
and (n764,n765,n808);
or (n765,n766,n805,n807);
and (n766,n767,n803);
or (n767,n768,n797,n802);
and (n768,n769,n781);
or (n769,n770,n779,n780);
and (n770,n771,n775);
xnor (n771,n772,n16);
nor (n772,n773,n774);
and (n773,n62,n486);
and (n774,n36,n488);
xnor (n775,n776,n11);
nor (n776,n777,n778);
and (n777,n77,n301);
and (n778,n54,n304);
and (n779,n775,n94);
and (n780,n771,n94);
or (n781,n782,n791,n796);
and (n782,n783,n787);
xnor (n783,n784,n29);
nor (n784,n785,n786);
and (n785,n93,n21);
and (n786,n69,n26);
xnor (n787,n788,n45);
nor (n788,n789,n790);
and (n789,n111,n37);
and (n790,n85,n42);
and (n791,n787,n792);
xnor (n792,n793,n63);
nor (n793,n794,n795);
and (n794,n116,n55);
and (n795,n103,n60);
and (n796,n783,n792);
and (n797,n781,n798);
xnor (n798,n799,n94);
nor (n799,n800,n801);
and (n800,n573,n86);
and (n801,n415,n91);
and (n802,n769,n798);
xor (n803,n804,n740);
xor (n804,n707,n723);
and (n805,n803,n806);
xor (n806,n744,n746);
and (n807,n767,n806);
xor (n808,n809,n641);
xor (n809,n614,n628);
and (n810,n808,n811);
xor (n811,n812,n749);
xor (n812,n705,n743);
and (n813,n765,n811);
and (n814,n815,n816);
xor (n815,n761,n763);
or (n816,n817,n887);
and (n817,n818,n820);
xor (n818,n819,n811);
xor (n819,n765,n808);
or (n820,n821,n883,n886);
and (n821,n822,n878);
or (n822,n823,n874,n877);
and (n823,n824,n864);
or (n824,n825,n858,n863);
and (n825,n826,n842);
or (n826,n827,n836,n841);
and (n827,n828,n832);
xnor (n828,n829,n45);
nor (n829,n830,n831);
and (n830,n103,n37);
and (n831,n111,n42);
xnor (n832,n833,n63);
nor (n833,n834,n835);
and (n834,n323,n55);
and (n835,n116,n60);
and (n836,n832,n837);
xnor (n837,n838,n78);
nor (n838,n839,n840);
and (n839,n573,n70);
and (n840,n415,n75);
and (n841,n828,n837);
or (n842,n843,n852,n857);
and (n843,n844,n848);
xnor (n844,n845,n16);
nor (n845,n846,n847);
and (n846,n54,n486);
and (n847,n62,n488);
xnor (n848,n849,n11);
nor (n849,n850,n851);
and (n850,n69,n301);
and (n851,n77,n304);
and (n852,n848,n853);
xnor (n853,n854,n29);
nor (n854,n855,n856);
and (n855,n85,n21);
and (n856,n93,n26);
and (n857,n844,n853);
and (n858,n842,n859);
xnor (n859,n860,n78);
nor (n860,n861,n862);
and (n861,n415,n70);
and (n862,n323,n75);
and (n863,n826,n859);
or (n864,n865,n870,n873);
and (n865,n866,n868);
xnor (n866,n867,n94);
nand (n867,n573,n91);
xor (n868,n869,n94);
xor (n869,n771,n775);
and (n870,n868,n871);
xor (n871,n872,n792);
xor (n872,n783,n787);
and (n873,n866,n871);
and (n874,n864,n875);
xor (n875,n876,n734);
xor (n876,n725,n729);
and (n877,n824,n875);
and (n878,n879,n881);
xor (n879,n880,n718);
xor (n880,n709,n713);
xor (n881,n882,n798);
xor (n882,n769,n781);
and (n883,n878,n884);
xor (n884,n885,n806);
xor (n885,n767,n803);
and (n886,n822,n884);
and (n887,n888,n889);
xor (n888,n818,n820);
or (n889,n890,n942);
and (n890,n891,n893);
xor (n891,n892,n884);
xor (n892,n822,n878);
or (n893,n894,n939,n941);
and (n894,n895,n937);
or (n895,n896,n933,n936);
and (n896,n897,n931);
or (n897,n898,n927,n930);
and (n898,n899,n915);
or (n899,n900,n909,n914);
and (n900,n901,n905);
xnor (n901,n902,n29);
nor (n902,n903,n904);
and (n903,n111,n21);
and (n904,n85,n26);
xnor (n905,n906,n45);
nor (n906,n907,n908);
and (n907,n116,n37);
and (n908,n103,n42);
and (n909,n905,n910);
xnor (n910,n911,n63);
nor (n911,n912,n913);
and (n912,n415,n55);
and (n913,n323,n60);
and (n914,n901,n910);
or (n915,n916,n925,n926);
and (n916,n917,n921);
xnor (n917,n918,n16);
nor (n918,n919,n920);
and (n919,n77,n486);
and (n920,n54,n488);
xnor (n921,n922,n11);
nor (n922,n923,n924);
and (n923,n93,n301);
and (n924,n69,n304);
and (n925,n921,n78);
and (n926,n917,n78);
and (n927,n915,n928);
xor (n928,n929,n837);
xor (n929,n828,n832);
and (n930,n899,n928);
xor (n931,n932,n859);
xor (n932,n826,n842);
and (n933,n931,n934);
xor (n934,n935,n871);
xor (n935,n866,n868);
and (n936,n897,n934);
xor (n937,n938,n875);
xor (n938,n824,n864);
and (n939,n937,n940);
xor (n940,n879,n881);
and (n941,n895,n940);
and (n942,n943,n944);
xor (n943,n891,n893);
or (n944,n945,n983);
and (n945,n946,n948);
xor (n946,n947,n940);
xor (n947,n895,n937);
and (n948,n949,n981);
or (n949,n950,n977,n980);
and (n950,n951,n975);
or (n951,n952,n971,n974);
and (n952,n953,n969);
or (n953,n954,n963,n968);
and (n954,n955,n959);
xnor (n955,n956,n16);
nor (n956,n957,n958);
and (n957,n69,n486);
and (n958,n77,n488);
xnor (n959,n960,n11);
nor (n960,n961,n962);
and (n961,n85,n301);
and (n962,n93,n304);
and (n963,n959,n964);
xnor (n964,n965,n29);
nor (n965,n966,n967);
and (n966,n103,n21);
and (n967,n111,n26);
and (n968,n955,n964);
xnor (n969,n970,n78);
nand (n970,n573,n75);
and (n971,n969,n972);
xor (n972,n973,n910);
xor (n973,n901,n905);
and (n974,n953,n972);
xor (n975,n976,n853);
xor (n976,n844,n848);
and (n977,n975,n978);
xor (n978,n979,n928);
xor (n979,n899,n915);
and (n980,n951,n978);
xor (n981,n982,n934);
xor (n982,n897,n931);
and (n983,n984,n985);
xor (n984,n946,n948);
or (n985,n986,n1038);
and (n986,n987,n988);
xor (n987,n949,n981);
and (n988,n989,n1036);
or (n989,n990,n1032,n1035);
and (n990,n991,n1025);
or (n991,n992,n1019,n1024);
and (n992,n993,n1007);
or (n993,n994,n1003,n1006);
and (n994,n995,n999);
xnor (n995,n996,n29);
nor (n996,n997,n998);
and (n997,n116,n21);
and (n998,n103,n26);
xnor (n999,n1000,n45);
nor (n1000,n1001,n1002);
and (n1001,n415,n37);
and (n1002,n323,n42);
and (n1003,n999,n1004);
xnor (n1004,n1005,n63);
nand (n1005,n573,n60);
and (n1006,n995,n1004);
or (n1007,n1008,n1017,n1018);
and (n1008,n1009,n1013);
xnor (n1009,n1010,n16);
nor (n1010,n1011,n1012);
and (n1011,n93,n486);
and (n1012,n69,n488);
xnor (n1013,n1014,n11);
nor (n1014,n1015,n1016);
and (n1015,n111,n301);
and (n1016,n85,n304);
and (n1017,n1013,n63);
and (n1018,n1009,n63);
and (n1019,n1007,n1020);
xnor (n1020,n1021,n45);
nor (n1021,n1022,n1023);
and (n1022,n323,n37);
and (n1023,n116,n42);
and (n1024,n993,n1020);
and (n1025,n1026,n1030);
xnor (n1026,n1027,n63);
nor (n1027,n1028,n1029);
and (n1028,n573,n55);
and (n1029,n415,n60);
xor (n1030,n1031,n964);
xor (n1031,n955,n959);
and (n1032,n1025,n1033);
xor (n1033,n1034,n78);
xor (n1034,n917,n921);
and (n1035,n991,n1033);
xor (n1036,n1037,n978);
xor (n1037,n951,n975);
and (n1038,n1039,n1040);
xor (n1039,n987,n988);
or (n1040,n1041,n1048);
and (n1041,n1042,n1043);
xor (n1042,n989,n1036);
and (n1043,n1044,n1046);
xor (n1044,n1045,n972);
xor (n1045,n953,n969);
xor (n1046,n1047,n1033);
xor (n1047,n991,n1025);
and (n1048,n1049,n1050);
xor (n1049,n1042,n1043);
or (n1050,n1051,n1084);
and (n1051,n1052,n1053);
xor (n1052,n1044,n1046);
or (n1053,n1054,n1081,n1083);
and (n1054,n1055,n1079);
or (n1055,n1056,n1075,n1078);
and (n1056,n1057,n1073);
or (n1057,n1058,n1067,n1072);
and (n1058,n1059,n1063);
xnor (n1059,n1060,n16);
nor (n1060,n1061,n1062);
and (n1061,n85,n486);
and (n1062,n93,n488);
xnor (n1063,n1064,n11);
nor (n1064,n1065,n1066);
and (n1065,n103,n301);
and (n1066,n111,n304);
and (n1067,n1063,n1068);
xnor (n1068,n1069,n29);
nor (n1069,n1070,n1071);
and (n1070,n323,n21);
and (n1071,n116,n26);
and (n1072,n1059,n1068);
xor (n1073,n1074,n1004);
xor (n1074,n995,n999);
and (n1075,n1073,n1076);
xor (n1076,n1077,n63);
xor (n1077,n1009,n1013);
and (n1078,n1057,n1076);
xor (n1079,n1080,n1020);
xor (n1080,n993,n1007);
and (n1081,n1079,n1082);
xor (n1082,n1026,n1030);
and (n1083,n1055,n1082);
and (n1084,n1085,n1086);
xor (n1085,n1052,n1053);
or (n1086,n1087,n1120);
and (n1087,n1088,n1090);
xor (n1088,n1089,n1082);
xor (n1089,n1055,n1079);
and (n1090,n1091,n1118);
or (n1091,n1092,n1112,n1117);
and (n1092,n1093,n1105);
or (n1093,n1094,n1103,n1104);
and (n1094,n1095,n1099);
xnor (n1095,n1096,n16);
nor (n1096,n1097,n1098);
and (n1097,n111,n486);
and (n1098,n85,n488);
xnor (n1099,n1100,n11);
nor (n1100,n1101,n1102);
and (n1101,n116,n301);
and (n1102,n103,n304);
and (n1103,n1099,n45);
and (n1104,n1095,n45);
and (n1105,n1106,n1110);
xnor (n1106,n1107,n29);
nor (n1107,n1108,n1109);
and (n1108,n415,n21);
and (n1109,n323,n26);
xnor (n1110,n1111,n45);
nand (n1111,n573,n42);
and (n1112,n1105,n1113);
xnor (n1113,n1114,n45);
nor (n1114,n1115,n1116);
and (n1115,n573,n37);
and (n1116,n415,n42);
and (n1117,n1093,n1113);
xor (n1118,n1119,n1076);
xor (n1119,n1057,n1073);
and (n1120,n1121,n1122);
xor (n1121,n1088,n1090);
or (n1122,n1123,n1130);
and (n1123,n1124,n1125);
xor (n1124,n1091,n1118);
and (n1125,n1126,n1128);
xor (n1126,n1127,n1068);
xor (n1127,n1059,n1063);
xor (n1128,n1129,n1113);
xor (n1129,n1093,n1105);
and (n1130,n1131,n1132);
xor (n1131,n1124,n1125);
or (n1132,n1133,n1158);
and (n1133,n1134,n1135);
xor (n1134,n1126,n1128);
or (n1135,n1136,n1155,n1157);
and (n1136,n1137,n1153);
or (n1137,n1138,n1147,n1152);
and (n1138,n1139,n1143);
xnor (n1139,n1140,n16);
nor (n1140,n1141,n1142);
and (n1141,n103,n486);
and (n1142,n111,n488);
xnor (n1143,n1144,n11);
nor (n1144,n1145,n1146);
and (n1145,n323,n301);
and (n1146,n116,n304);
and (n1147,n1143,n1148);
xnor (n1148,n1149,n29);
nor (n1149,n1150,n1151);
and (n1150,n573,n21);
and (n1151,n415,n26);
and (n1152,n1139,n1148);
xor (n1153,n1154,n45);
xor (n1154,n1095,n1099);
and (n1155,n1153,n1156);
xor (n1156,n1106,n1110);
and (n1157,n1137,n1156);
and (n1158,n1159,n1160);
xor (n1159,n1134,n1135);
or (n1160,n1161,n1179);
and (n1161,n1162,n1164);
xor (n1162,n1163,n1156);
xor (n1163,n1137,n1153);
and (n1164,n1165,n1177);
or (n1165,n1166,n1175,n1176);
and (n1166,n1167,n1171);
xnor (n1167,n1168,n16);
nor (n1168,n1169,n1170);
and (n1169,n116,n486);
and (n1170,n103,n488);
xnor (n1171,n1172,n11);
nor (n1172,n1173,n1174);
and (n1173,n415,n301);
and (n1174,n323,n304);
and (n1175,n1171,n29);
and (n1176,n1167,n29);
xor (n1177,n1178,n1148);
xor (n1178,n1139,n1143);
and (n1179,n1180,n1181);
xor (n1180,n1162,n1164);
or (n1181,n1182,n1189);
and (n1182,n1183,n1184);
xor (n1183,n1165,n1177);
and (n1184,n1185,n1187);
xnor (n1185,n1186,n29);
nand (n1186,n573,n26);
xor (n1187,n1188,n29);
xor (n1188,n1167,n1171);
and (n1189,n1190,n1191);
xor (n1190,n1183,n1184);
or (n1191,n1192,n1203);
and (n1192,n1193,n1194);
xor (n1193,n1185,n1187);
and (n1194,n1195,n1199);
xnor (n1195,n1196,n16);
nor (n1196,n1197,n1198);
and (n1197,n323,n486);
and (n1198,n116,n488);
xnor (n1199,n1200,n11);
nor (n1200,n1201,n1202);
and (n1201,n573,n301);
and (n1202,n415,n304);
and (n1203,n1204,n1205);
xor (n1204,n1193,n1194);
or (n1205,n1206,n1213);
and (n1206,n1207,n1208);
xor (n1207,n1195,n1199);
and (n1208,n1209,n11);
xnor (n1209,n1210,n16);
nor (n1210,n1211,n1212);
and (n1211,n415,n486);
and (n1212,n323,n488);
and (n1213,n1214,n1215);
xor (n1214,n1207,n1208);
or (n1215,n1216,n1220);
and (n1216,n1217,n1219);
xnor (n1217,n1218,n11);
nand (n1218,n573,n304);
xor (n1219,n1209,n11);
and (n1220,n1221,n1222);
xor (n1221,n1217,n1219);
and (n1222,n1223,n1227);
xnor (n1223,n1224,n16);
nor (n1224,n1225,n1226);
and (n1225,n573,n486);
and (n1226,n415,n488);
and (n1227,n1228,n16);
xnor (n1228,n1229,n16);
nand (n1229,n573,n488);
xor (n1230,n1231,n1334);
xor (n1231,n1232,n1302);
xor (n1232,n1233,n1283);
or (n1233,n1234,n1274,n1282);
and (n1234,n1235,n1256);
or (n1235,n1236,n1254,n1255);
and (n1236,n1237,n1245);
or (n1237,n1238,n1242,n1244);
and (n1238,n1239,n49);
or (n1239,n1240,n32,n1241);
and (n1240,n122,n17);
and (n1241,n122,n33);
and (n1242,n49,n1243);
and (n1243,n100,n115);
and (n1244,n1239,n1243);
or (n1245,n1246,n1251,n1253);
and (n1246,n1247,n1249);
xor (n1247,n1248,n132);
xor (n1248,n123,n126);
xor (n1249,n1250,n146);
xor (n1250,n136,n140);
and (n1251,n1249,n1252);
not (n1252,n150);
and (n1253,n1247,n1252);
and (n1254,n1245,n153);
and (n1255,n1237,n153);
xor (n1256,n1257,n1272);
xor (n1257,n1258,n1268);
or (n1258,n1259,n1266,n1267);
and (n1259,n1260,n1263);
or (n1260,n199,n1261,n1262);
and (n1261,n126,n132);
and (n1262,n123,n132);
or (n1263,n203,n1264,n1265);
and (n1264,n140,n146);
and (n1265,n136,n146);
and (n1266,n1263,n150);
and (n1267,n1260,n150);
or (n1268,n1269,n1270,n1271);
and (n1269,n155,n156);
and (n1270,n156,n167);
and (n1271,n155,n167);
xor (n1272,n1273,n215);
xor (n1273,n222,n226);
and (n1274,n1256,n1275);
xor (n1275,n1276,n1278);
xor (n1276,n1277,n218);
xor (n1277,n233,n236);
xnor (n1278,n1279,n188);
or (n1279,n1280,n186,n1281);
and (n1280,n232,n159);
and (n1281,n232,n163);
and (n1282,n1235,n1275);
xor (n1283,n1284,n1290);
xor (n1284,n1285,n1289);
or (n1285,n1286,n1287,n1288);
and (n1286,n1258,n1268);
and (n1287,n1268,n1272);
and (n1288,n1258,n1272);
and (n1289,n1276,n1278);
xor (n1290,n1291,n1294);
xor (n1291,n1292,n1293);
or (n1292,n1279,n188);
not (n1293,n269);
xor (n1294,n1295,n257);
xor (n1295,n1296,n1299);
or (n1296,n282,n1297,n1298);
and (n1297,n226,n215);
and (n1298,n222,n215);
or (n1299,n286,n1300,n1301);
and (n1300,n236,n218);
and (n1301,n233,n218);
and (n1302,n1303,n1332);
or (n1303,n1304,n1328,n1331);
and (n1304,n1305,n1326);
or (n1305,n1306,n1322,n1325);
and (n1306,n1307,n1318);
or (n1307,n1308,n1315,n1317);
and (n1308,n1309,n1312);
or (n1309,n305,n1310,n1311);
and (n1310,n306,n328);
and (n1311,n298,n328);
or (n1312,n336,n1313,n1314);
and (n1313,n337,n313);
and (n1314,n332,n313);
and (n1315,n1312,n1316);
or (n1316,n317,n322);
and (n1317,n1309,n1316);
or (n1318,n1319,n1320,n1321);
and (n1319,n426,n347);
and (n1320,n347,n427);
and (n1321,n426,n427);
and (n1322,n1318,n1323);
xor (n1323,n1324,n1252);
xor (n1324,n1247,n1249);
and (n1325,n1307,n1323);
xor (n1326,n1327,n150);
xor (n1327,n1260,n1263);
and (n1328,n1326,n1329);
xor (n1329,n1330,n153);
xor (n1330,n1237,n1245);
and (n1331,n1305,n1329);
xor (n1332,n1333,n1275);
xor (n1333,n1235,n1256);
or (n1334,n1335,n1367);
and (n1335,n1336,n1337);
xor (n1336,n1303,n1332);
and (n1337,n1338,n1365);
or (n1338,n1339,n1361,n1364);
and (n1339,n1340,n1359);
or (n1340,n1341,n1357,n1358);
and (n1341,n1342,n1348);
or (n1342,n1343,n1347,n417);
and (n1343,n374,n1344);
or (n1344,n1345,n396,n1346);
and (n1345,n297,n392);
and (n1346,n297,n397);
and (n1347,n1344,n403);
or (n1348,n1349,n1354,n1356);
and (n1349,n1350,n1352);
xor (n1350,n1351,n328);
xor (n1351,n298,n306);
xor (n1352,n1353,n313);
xor (n1353,n332,n337);
and (n1354,n1352,n1355);
xnor (n1355,n317,n322);
and (n1356,n1350,n1355);
and (n1357,n1348,n424);
and (n1358,n1342,n424);
xor (n1359,n1360,n1243);
xor (n1360,n1239,n49);
and (n1361,n1359,n1362);
xor (n1362,n1363,n1323);
xor (n1363,n1307,n1318);
and (n1364,n1340,n1362);
xor (n1365,n1366,n1329);
xor (n1366,n1305,n1326);
and (n1367,n1368,n1369);
xor (n1368,n1336,n1337);
or (n1369,n1370,n1390);
and (n1370,n1371,n1372);
xor (n1371,n1338,n1365);
and (n1372,n1373,n1388);
or (n1373,n1374,n1384,n1387);
and (n1374,n1375,n1382);
or (n1375,n1376,n1378,n1381);
and (n1376,n447,n1377);
or (n1377,n497,n502);
and (n1378,n1377,n1379);
xor (n1379,n1380,n1355);
xor (n1380,n1350,n1352);
and (n1381,n447,n1379);
xor (n1382,n1383,n1316);
xor (n1383,n1309,n1312);
and (n1384,n1382,n1385);
xor (n1385,n1386,n424);
xor (n1386,n1342,n1348);
and (n1387,n1375,n1385);
xor (n1388,n1389,n1362);
xor (n1389,n1340,n1359);
and (n1390,n1391,n1392);
xor (n1391,n1371,n1372);
or (n1392,n1393,n1409);
and (n1393,n1394,n1395);
xor (n1394,n1373,n1388);
and (n1395,n1396,n1407);
or (n1396,n1397,n1403,n1406);
and (n1397,n1398,n1401);
or (n1398,n529,n1399,n1400);
and (n1399,n576,n698);
and (n1400,n530,n698);
xor (n1401,n1402,n403);
xor (n1402,n374,n1344);
and (n1403,n1401,n1404);
xor (n1404,n1405,n1379);
xor (n1405,n447,n1377);
and (n1406,n1398,n1404);
xor (n1407,n1408,n1385);
xor (n1408,n1375,n1382);
and (n1409,n1410,n1411);
xor (n1410,n1394,n1395);
or (n1411,n1412,n1420);
and (n1412,n1413,n1414);
xor (n1413,n1396,n1407);
and (n1414,n1415,n1418);
or (n1415,n609,n1416,n1417);
and (n1416,n670,n700);
and (n1417,n610,n700);
xor (n1418,n1419,n1404);
xor (n1419,n1398,n1401);
and (n1420,n1421,n1422);
xor (n1421,n1413,n1414);
or (n1422,n1423,n691);
and (n1423,n1424,n1425);
xor (n1424,n1415,n1418);
or (n1425,n1426,n1427,n1428);
and (n1426,n676,n697);
and (n1427,n697,n699);
and (n1428,n676,n699);
endmodule
