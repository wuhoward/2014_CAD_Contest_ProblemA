module top (out,n14,n16,n17,n21,n25,n27,n28,n30,n33
        ,n38,n40,n42,n45,n56,n58,n59,n61,n68,n70
        ,n73,n80,n82,n89,n98,n100,n101,n103,n106,n110
        ,n112,n114,n117,n122,n124,n126,n129,n146,n164,n165
        ,n195,n197,n199,n205,n324,n388,n464,n646,n765);
output out;
input n14;
input n16;
input n17;
input n21;
input n25;
input n27;
input n28;
input n30;
input n33;
input n38;
input n40;
input n42;
input n45;
input n56;
input n58;
input n59;
input n61;
input n68;
input n70;
input n73;
input n80;
input n82;
input n89;
input n98;
input n100;
input n101;
input n103;
input n106;
input n110;
input n112;
input n114;
input n117;
input n122;
input n124;
input n126;
input n129;
input n146;
input n164;
input n165;
input n195;
input n197;
input n199;
input n205;
input n324;
input n388;
input n464;
input n646;
input n765;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n24;
wire n26;
wire n29;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n41;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n102;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n111;
wire n113;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n125;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n198;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
xor (out,n0,n2338);
xnor (n0,n1,n2248);
nand (n1,n2,n598);
nand (n2,n3,n508);
nand (n3,n4,n369,n507);
nand (n4,n5,n223);
xor (n5,n6,n184);
xor (n6,n7,n91);
xor (n7,n8,n74);
xor (n8,n9,n47);
nand (n9,n10,n34,n46);
nand (n10,n11,n22);
xor (n11,n12,n21);
or (n12,n13,n18);
and (n13,n14,n15);
xor (n15,n16,n17);
and (n18,n14,n19);
nor (n19,n15,n20);
xnor (n20,n21,n16);
xor (n22,n23,n33);
or (n23,n24,n29);
and (n24,n25,n26);
xor (n26,n27,n28);
and (n29,n30,n31);
nor (n31,n26,n32);
xnor (n32,n33,n27);
nand (n34,n35,n22);
xor (n35,n36,n45);
or (n36,n37,n41);
and (n37,n38,n39);
xor (n39,n40,n33);
and (n41,n42,n43);
nor (n43,n39,n44);
xnor (n44,n45,n40);
nand (n46,n11,n35);
xor (n47,n48,n64);
xor (n48,n49,n53);
xor (n49,n50,n45);
or (n50,n51,n52);
and (n51,n30,n39);
and (n52,n38,n43);
xor (n53,n54,n28);
or (n54,n55,n60);
and (n55,n56,n57);
xor (n57,n58,n59);
and (n60,n61,n62);
nor (n62,n57,n63);
xnor (n63,n28,n58);
xor (n64,n65,n73);
or (n65,n66,n69);
and (n66,n42,n67);
xor (n67,n68,n45);
and (n69,n70,n71);
nor (n71,n67,n72);
xnor (n72,n73,n68);
xor (n74,n75,n86);
xor (n75,n76,n85);
xor (n76,n77,n59);
or (n77,n78,n81);
and (n78,n14,n79);
xor (n79,n80,n21);
and (n81,n82,n83);
nor (n83,n79,n84);
xnor (n84,n59,n80);
not (n85,n11);
xor (n86,n87,n33);
or (n87,n88,n90);
and (n88,n89,n26);
and (n90,n25,n31);
nand (n91,n92,n147,n183);
nand (n92,n93,n131);
nand (n93,n94,n118,n130);
nand (n94,n95,n107);
xor (n95,n96,n106);
or (n96,n97,n102);
and (n97,n98,n99);
xor (n99,n100,n101);
and (n102,n103,n104);
nor (n104,n99,n105);
xnor (n105,n106,n100);
xor (n107,n108,n117);
or (n108,n109,n113);
and (n109,n110,n111);
xor (n111,n112,n106);
and (n113,n114,n115);
nor (n115,n111,n116);
xnor (n116,n117,n112);
nand (n118,n119,n107);
xor (n119,n120,n129);
or (n120,n121,n125);
and (n121,n122,n123);
xor (n123,n124,n117);
and (n125,n126,n127);
nor (n127,n123,n128);
xnor (n128,n129,n124);
nand (n130,n95,n119);
xor (n131,n132,n142);
xor (n132,n133,n137);
xor (n133,n134,n28);
or (n134,n135,n136);
and (n135,n61,n57);
and (n136,n89,n62);
not (n137,n138);
xor (n138,n139,n59);
or (n139,n140,n141);
and (n140,n82,n79);
and (n141,n56,n83);
xor (n142,n143,n73);
or (n143,n144,n145);
and (n144,n70,n67);
and (n145,n146,n71);
nand (n147,n148,n131);
nand (n148,n149,n169,n182);
nand (n149,n150,n129);
xor (n150,n151,n159);
xor (n151,n152,n155);
xor (n152,n153,n21);
or (n153,n13,n154);
and (n154,n82,n19);
xor (n155,n156,n59);
or (n156,n157,n158);
and (n157,n56,n79);
and (n158,n61,n83);
not (n159,n160);
xor (n160,n161,n17);
or (n161,n162,n166);
and (n162,n14,n163);
xor (n163,n164,n165);
and (n166,n14,n167);
nor (n167,n163,n168);
xnor (n168,n17,n164);
nand (n169,n170,n129);
nand (n170,n171,n176,n181);
nand (n171,n172,n160);
xor (n172,n173,n59);
or (n173,n174,n175);
and (n174,n61,n79);
and (n175,n89,n83);
nand (n176,n177,n160);
xor (n177,n178,n28);
or (n178,n179,n180);
and (n179,n25,n57);
and (n180,n30,n62);
nand (n181,n172,n177);
nand (n182,n150,n170);
nand (n183,n93,n148);
xor (n184,n185,n213);
xor (n185,n186,n190);
nand (n186,n187,n188,n189);
nand (n187,n133,n137);
nand (n188,n142,n137);
nand (n189,n133,n142);
nand (n190,n191,n207,n212);
nand (n191,n192,n202);
xor (n192,n193,n101);
or (n193,n194,n198);
and (n194,n195,n196);
xor (n196,n197,n73);
and (n198,n199,n200);
nor (n200,n196,n201);
xnor (n201,n101,n197);
xor (n202,n203,n106);
or (n203,n204,n206);
and (n204,n205,n99);
and (n206,n98,n104);
nand (n207,n208,n202);
xor (n208,n209,n117);
or (n209,n210,n211);
and (n210,n103,n111);
and (n211,n110,n115);
nand (n212,n192,n208);
xor (n213,n214,n219);
xor (n214,n138,n215);
xor (n215,n216,n101);
or (n216,n217,n218);
and (n217,n146,n196);
and (n218,n195,n200);
xor (n219,n220,n106);
or (n220,n221,n222);
and (n221,n199,n99);
and (n222,n205,n104);
xor (n223,n224,n340);
xor (n224,n225,n287);
xor (n225,n226,n249);
xor (n226,n227,n239);
nand (n227,n228,n233,n238);
nand (n228,n229,n129);
xor (n229,n230,n129);
or (n230,n231,n232);
and (n231,n114,n123);
and (n232,n122,n127);
nand (n233,n234,n129);
nand (n234,n235,n236,n237);
nand (n235,n152,n155);
nand (n236,n159,n155);
nand (n237,n152,n159);
nand (n238,n229,n234);
xor (n239,n240,n129);
xor (n240,n241,n245);
xor (n241,n242,n117);
or (n242,n243,n244);
and (n243,n98,n111);
and (n244,n103,n115);
xor (n245,n246,n129);
or (n246,n247,n248);
and (n247,n110,n123);
and (n248,n114,n127);
nand (n249,n250,n269,n286);
nand (n250,n251,n267);
nand (n251,n252,n261,n266);
nand (n252,n253,n257);
xor (n253,n254,n28);
or (n254,n255,n256);
and (n255,n89,n57);
and (n256,n25,n62);
xor (n257,n258,n33);
or (n258,n259,n260);
and (n259,n30,n26);
and (n260,n38,n31);
nand (n261,n262,n257);
xor (n262,n263,n45);
or (n263,n264,n265);
and (n264,n42,n39);
and (n265,n70,n43);
nand (n266,n253,n262);
xor (n267,n268,n35);
xor (n268,n11,n22);
nand (n269,n270,n267);
nand (n270,n271,n280,n285);
nand (n271,n272,n276);
xor (n272,n273,n101);
or (n273,n274,n275);
and (n274,n199,n196);
and (n275,n205,n200);
xor (n276,n277,n21);
or (n277,n278,n279);
and (n278,n82,n15);
and (n279,n56,n19);
nand (n280,n281,n276);
xor (n281,n282,n73);
or (n282,n283,n284);
and (n283,n146,n67);
and (n284,n195,n71);
nand (n285,n272,n281);
nand (n286,n251,n270);
nand (n287,n288,n292,n339);
nand (n288,n289,n291);
xor (n289,n290,n208);
xor (n290,n192,n202);
xor (n291,n230,n234);
nand (n292,n293,n291);
nand (n293,n294,n313,n338);
nand (n294,n295,n297);
xor (n295,n296,n262);
xor (n296,n253,n257);
nand (n297,n298,n307,n312);
nand (n298,n299,n303);
xor (n299,n300,n33);
or (n300,n301,n302);
and (n301,n38,n26);
and (n302,n42,n31);
xor (n303,n304,n45);
or (n304,n305,n306);
and (n305,n70,n39);
and (n306,n146,n43);
nand (n307,n308,n303);
xor (n308,n309,n101);
or (n309,n310,n311);
and (n310,n205,n196);
and (n311,n98,n200);
nand (n312,n299,n308);
nand (n313,n314,n297);
nand (n314,n315,n325,n337);
nand (n315,n316,n320);
xor (n316,n317,n117);
or (n317,n318,n319);
and (n318,n114,n111);
and (n319,n122,n115);
xor (n320,n321,n129);
or (n321,n322,n323);
and (n322,n126,n123);
and (n323,n324,n127);
nand (n325,n326,n320);
nand (n326,n327,n332,n336);
not (n327,n328);
xor (n328,n329,n59);
or (n329,n330,n331);
and (n330,n89,n79);
and (n331,n25,n83);
nand (n332,n333,n328);
xor (n333,n334,n17);
or (n334,n162,n335);
and (n335,n82,n167);
not (n336,n333);
nand (n337,n316,n326);
nand (n338,n295,n314);
nand (n339,n289,n293);
nand (n340,n341,n365,n368);
nand (n341,n342,n344);
xor (n342,n343,n270);
xor (n343,n251,n267);
nand (n344,n345,n361,n364);
nand (n345,n346,n359);
nand (n346,n347,n353,n358);
nand (n347,n348,n349);
not (n348,n276);
xor (n349,n350,n73);
or (n350,n351,n352);
and (n351,n195,n67);
and (n352,n199,n71);
nand (n353,n354,n349);
xor (n354,n355,n106);
or (n355,n356,n357);
and (n356,n103,n99);
and (n357,n110,n104);
nand (n358,n348,n354);
xor (n359,n360,n281);
xor (n360,n272,n276);
nand (n361,n362,n359);
xor (n362,n363,n119);
xor (n363,n95,n107);
nand (n364,n346,n362);
nand (n365,n366,n344);
xor (n366,n367,n148);
xor (n367,n93,n131);
nand (n368,n342,n366);
nand (n369,n370,n223);
nand (n370,n371,n422,n506);
nand (n371,n372,n420);
nand (n372,n373,n416,n419);
nand (n373,n374,n414);
nand (n374,n375,n396,n413);
nand (n375,n129,n376);
nand (n376,n377,n390,n395);
nand (n377,n378,n382);
xor (n378,n379,n21);
or (n379,n380,n381);
and (n380,n56,n15);
and (n381,n61,n19);
not (n382,n383);
xnor (n383,n384,n165);
nor (n384,n385,n389);
and (n385,n14,n386);
and (n386,n387,n165);
not (n387,n388);
and (n389,n14,n388);
nand (n390,n391,n382);
xor (n391,n392,n28);
or (n392,n393,n394);
and (n393,n30,n57);
and (n394,n38,n62);
nand (n395,n378,n391);
nand (n396,n397,n376);
nand (n397,n398,n407,n412);
nand (n398,n399,n403);
xor (n399,n400,n33);
or (n400,n401,n402);
and (n401,n42,n26);
and (n402,n70,n31);
xor (n403,n404,n45);
or (n404,n405,n406);
and (n405,n146,n39);
and (n406,n195,n43);
nand (n407,n408,n403);
xor (n408,n409,n73);
or (n409,n410,n411);
and (n410,n199,n67);
and (n411,n205,n71);
nand (n412,n399,n408);
nand (n413,n129,n397);
xor (n414,n415,n170);
xor (n415,n150,n129);
nand (n416,n417,n414);
xor (n417,n418,n314);
xor (n418,n295,n297);
nand (n419,n374,n417);
xor (n420,n421,n293);
xor (n421,n289,n291);
nand (n422,n423,n420);
nand (n423,n424,n502,n505);
nand (n424,n425,n450);
nand (n425,n426,n431,n449);
nand (n426,n427,n429);
xor (n427,n428,n308);
xor (n428,n299,n303);
xor (n429,n430,n177);
xor (n430,n172,n160);
nand (n431,n432,n429);
nand (n432,n433,n443,n448);
nand (n433,n434,n438);
xor (n434,n435,n101);
or (n435,n436,n437);
and (n436,n98,n196);
and (n437,n103,n200);
and (n438,n129,n439);
xor (n439,n440,n59);
or (n440,n441,n442);
and (n441,n25,n79);
and (n442,n30,n83);
nand (n443,n444,n438);
xor (n444,n445,n106);
or (n445,n446,n447);
and (n446,n110,n99);
and (n447,n114,n104);
nand (n448,n434,n444);
nand (n449,n427,n432);
nand (n450,n451,n479,n501);
nand (n451,n452,n454);
xor (n452,n453,n354);
xor (n453,n348,n349);
nand (n454,n455,n465,n478);
nand (n455,n456,n460);
xor (n456,n457,n117);
or (n457,n458,n459);
and (n458,n122,n111);
and (n459,n126,n115);
xor (n460,n461,n129);
or (n461,n462,n463);
and (n462,n324,n123);
and (n463,n464,n127);
nand (n465,n466,n460);
nand (n466,n467,n476,n477);
nand (n467,n468,n472);
xor (n468,n469,n17);
or (n469,n470,n471);
and (n470,n82,n163);
and (n471,n56,n167);
xor (n472,n473,n21);
or (n473,n474,n475);
and (n474,n61,n15);
and (n475,n89,n19);
nand (n476,n383,n472);
nand (n477,n468,n383);
nand (n478,n456,n466);
nand (n479,n480,n454);
nand (n480,n481,n499,n500);
nand (n481,n482,n498);
nand (n482,n483,n492,n497);
nand (n483,n484,n488);
xor (n484,n485,n28);
or (n485,n486,n487);
and (n486,n38,n57);
and (n487,n42,n62);
xor (n488,n489,n33);
or (n489,n490,n491);
and (n490,n70,n26);
and (n491,n146,n31);
nand (n492,n493,n488);
xor (n493,n494,n45);
or (n494,n495,n496);
and (n495,n195,n39);
and (n496,n199,n43);
nand (n497,n484,n493);
xor (n498,n327,n333);
nand (n499,n129,n498);
nand (n500,n482,n129);
nand (n501,n452,n480);
nand (n502,n503,n450);
xor (n503,n504,n362);
xor (n504,n346,n359);
nand (n505,n425,n503);
nand (n506,n372,n423);
nand (n507,n5,n370);
xor (n508,n509,n594);
xor (n509,n510,n514);
nand (n510,n511,n512,n513);
nand (n511,n7,n91);
nand (n512,n184,n91);
nand (n513,n7,n184);
xor (n514,n515,n560);
xor (n515,n516,n556);
xor (n516,n517,n536);
xor (n517,n518,n522);
nand (n518,n519,n520,n521);
nand (n519,n241,n245);
nand (n520,n129,n245);
nand (n521,n241,n129);
xor (n522,n523,n532);
xor (n523,n524,n528);
xor (n524,n525,n129);
or (n525,n526,n527);
and (n526,n103,n123);
and (n527,n110,n127);
not (n528,n529);
xor (n529,n530,n59);
or (n530,n78,n531);
and (n531,n14,n83);
xor (n532,n533,n106);
or (n533,n534,n535);
and (n534,n195,n99);
and (n535,n199,n104);
xor (n536,n537,n542);
xor (n537,n129,n538);
nand (n538,n539,n540,n541);
nand (n539,n76,n85);
nand (n540,n86,n85);
nand (n541,n76,n86);
xor (n542,n543,n552);
xor (n543,n544,n548);
xor (n544,n545,n45);
or (n545,n546,n547);
and (n546,n25,n39);
and (n547,n30,n43);
xor (n548,n549,n28);
or (n549,n550,n551);
and (n550,n82,n57);
and (n551,n56,n62);
xor (n552,n553,n33);
or (n553,n554,n555);
and (n554,n61,n26);
and (n555,n89,n31);
nand (n556,n557,n558,n559);
nand (n557,n227,n239);
nand (n558,n249,n239);
nand (n559,n227,n249);
xor (n560,n561,n570);
xor (n561,n562,n566);
nand (n562,n563,n564,n565);
nand (n563,n9,n47);
nand (n564,n74,n47);
nand (n565,n9,n74);
nand (n566,n567,n568,n569);
nand (n567,n186,n190);
nand (n568,n213,n190);
nand (n569,n186,n213);
xor (n570,n571,n590);
xor (n571,n572,n576);
nand (n572,n573,n574,n575);
nand (n573,n49,n53);
nand (n574,n64,n53);
nand (n575,n49,n64);
xor (n576,n577,n586);
xor (n577,n578,n582);
xor (n578,n579,n73);
or (n579,n580,n581);
and (n580,n38,n67);
and (n581,n42,n71);
xor (n582,n583,n101);
or (n583,n584,n585);
and (n584,n70,n196);
and (n585,n146,n200);
xor (n586,n587,n117);
or (n587,n588,n589);
and (n588,n205,n111);
and (n589,n98,n115);
nand (n590,n591,n592,n593);
nand (n591,n138,n215);
nand (n592,n219,n215);
nand (n593,n138,n219);
nand (n594,n595,n596,n597);
nand (n595,n225,n287);
nand (n596,n340,n287);
nand (n597,n225,n340);
nand (n598,n599,n2246);
nand (n599,n600,n845);
nor (n600,n601,n843);
nor (n601,n602,n836);
nand (n602,n603,n826);
nand (n603,n604,n814,n825);
nand (n604,n605,n706);
nand (n605,n606,n633,n705);
nand (n606,n607,n609);
xor (n607,n608,n432);
xor (n608,n427,n429);
nand (n609,n610,n629,n632);
nand (n610,n611,n627);
nand (n611,n612,n621,n626);
nand (n612,n129,n613);
and (n613,n614,n617);
xnor (n614,n615,n165);
nor (n615,n616,n389);
and (n616,n82,n386);
xor (n617,n618,n17);
or (n618,n619,n620);
and (n619,n56,n163);
and (n620,n61,n167);
nand (n621,n622,n613);
xor (n622,n623,n106);
or (n623,n624,n625);
and (n624,n114,n99);
and (n625,n122,n104);
nand (n626,n129,n622);
xor (n627,n628,n444);
xor (n628,n434,n438);
nand (n629,n630,n627);
xor (n630,n631,n466);
xor (n631,n456,n460);
nand (n632,n611,n630);
nand (n633,n634,n609);
nand (n634,n635,n701,n704);
nand (n635,n636,n665);
nand (n636,n637,n647,n664);
nand (n637,n638,n642);
xor (n638,n639,n117);
or (n639,n640,n641);
and (n640,n126,n111);
and (n641,n324,n115);
xor (n642,n643,n129);
or (n643,n644,n645);
and (n644,n464,n123);
and (n645,n646,n127);
nand (n647,n648,n642);
nand (n648,n649,n658,n663);
nand (n649,n650,n654);
xor (n650,n651,n59);
or (n651,n652,n653);
and (n652,n30,n79);
and (n653,n38,n83);
xor (n654,n655,n21);
or (n655,n656,n657);
and (n656,n89,n15);
and (n657,n25,n19);
nand (n658,n659,n654);
xor (n659,n660,n28);
or (n660,n661,n662);
and (n661,n42,n57);
and (n662,n70,n62);
nand (n663,n650,n659);
nand (n664,n638,n648);
nand (n665,n666,n685,n700);
nand (n666,n667,n669);
xor (n667,n668,n383);
xor (n668,n468,n472);
nand (n669,n670,n679,n684);
nand (n670,n671,n675);
xor (n671,n672,n33);
or (n672,n673,n674);
and (n673,n146,n26);
and (n674,n195,n31);
xor (n675,n676,n45);
or (n676,n677,n678);
and (n677,n199,n39);
and (n678,n205,n43);
nand (n679,n680,n675);
xor (n680,n681,n73);
or (n681,n682,n683);
and (n682,n98,n67);
and (n683,n103,n71);
nand (n684,n671,n680);
nand (n685,n686,n669);
nand (n686,n687,n693,n699);
nand (n687,n688,n692);
xor (n688,n689,n101);
or (n689,n690,n691);
and (n690,n110,n196);
and (n691,n114,n200);
xor (n692,n614,n617);
nand (n693,n694,n692);
and (n694,n129,n695);
xor (n695,n696,n17);
or (n696,n697,n698);
and (n697,n61,n163);
and (n698,n89,n167);
nand (n699,n688,n694);
nand (n700,n667,n686);
nand (n701,n702,n665);
xor (n702,n703,n129);
xor (n703,n482,n498);
nand (n704,n636,n702);
nand (n705,n607,n634);
nand (n706,n707,n737,n813);
nand (n707,n708,n710);
xor (n708,n709,n480);
xor (n709,n452,n454);
xor (n710,n711,n716);
xor (n711,n712,n714);
xor (n712,n713,n326);
xor (n713,n316,n320);
xor (n714,n715,n397);
xor (n715,n129,n376);
nand (n716,n717,n733,n736);
nand (n717,n718,n731);
nand (n718,n719,n728,n730);
nand (n719,n720,n724);
xor (n720,n721,n73);
or (n721,n722,n723);
and (n722,n205,n67);
and (n723,n98,n71);
xor (n724,n725,n101);
or (n725,n726,n727);
and (n726,n103,n196);
and (n727,n110,n200);
nand (n728,n729,n724);
xor (n729,n129,n439);
nand (n730,n720,n729);
xor (n731,n732,n408);
xor (n732,n399,n403);
nand (n733,n734,n731);
xor (n734,n735,n391);
xor (n735,n378,n382);
nand (n736,n718,n734);
nand (n737,n738,n710);
nand (n738,n739,n752,n812);
nand (n739,n740,n750);
nand (n740,n741,n746,n749);
nand (n741,n742,n744);
xor (n742,n743,n493);
xor (n743,n484,n488);
xor (n744,n745,n622);
xor (n745,n129,n613);
nand (n746,n747,n744);
xor (n747,n748,n729);
xor (n748,n720,n724);
nand (n749,n742,n747);
xor (n750,n751,n734);
xor (n751,n718,n731);
nand (n752,n753,n750);
nand (n753,n754,n808,n811);
nand (n754,n755,n772);
nand (n755,n756,n766,n771);
nand (n756,n757,n761);
xor (n757,n758,n106);
or (n758,n759,n760);
and (n759,n122,n99);
and (n760,n126,n104);
xor (n761,n762,n129);
or (n762,n763,n764);
and (n763,n646,n123);
and (n764,n765,n127);
nand (n766,n767,n761);
xor (n767,n768,n117);
or (n768,n769,n770);
and (n769,n324,n111);
and (n770,n464,n115);
nand (n771,n757,n767);
nand (n772,n773,n792,n807);
nand (n773,n774,n790);
nand (n774,n775,n784,n789);
nand (n775,n776,n780);
xor (n776,n777,n59);
or (n777,n778,n779);
and (n778,n38,n79);
and (n779,n42,n83);
xnor (n780,n781,n165);
nor (n781,n782,n783);
and (n782,n56,n386);
and (n783,n82,n388);
nand (n784,n785,n780);
xor (n785,n786,n21);
or (n786,n787,n788);
and (n787,n25,n15);
and (n788,n30,n19);
nand (n789,n776,n785);
xor (n790,n791,n659);
xor (n791,n650,n654);
nand (n792,n793,n790);
nand (n793,n794,n801,n806);
nand (n794,n795,n799);
xor (n795,n796,n28);
or (n796,n797,n798);
and (n797,n70,n57);
and (n798,n146,n62);
xnor (n799,n800,n129);
nand (n800,n765,n123);
nand (n801,n802,n799);
xor (n802,n803,n33);
or (n803,n804,n805);
and (n804,n195,n26);
and (n805,n199,n31);
nand (n806,n795,n802);
nand (n807,n774,n793);
nand (n808,n809,n772);
xor (n809,n810,n648);
xor (n810,n638,n642);
nand (n811,n755,n809);
nand (n812,n740,n753);
nand (n813,n708,n738);
nand (n814,n815,n706);
xor (n815,n816,n823);
xor (n816,n817,n821);
nand (n817,n818,n819,n820);
nand (n818,n712,n714);
nand (n819,n716,n714);
nand (n820,n712,n716);
xor (n821,n822,n417);
xor (n822,n374,n414);
xor (n823,n824,n503);
xor (n824,n425,n450);
nand (n825,n605,n815);
xor (n826,n827,n832);
xor (n827,n828,n830);
xor (n828,n829,n366);
xor (n829,n342,n344);
xor (n830,n831,n423);
xor (n831,n372,n420);
nand (n832,n833,n834,n835);
nand (n833,n817,n821);
nand (n834,n823,n821);
nand (n835,n817,n823);
nor (n836,n837,n841);
nand (n837,n838,n839,n840);
nand (n838,n828,n830);
nand (n839,n832,n830);
nand (n840,n828,n832);
xor (n841,n842,n370);
xor (n842,n5,n223);
not (n843,n844);
nand (n844,n837,n841);
nand (n845,n846,n848);
nor (n846,n847,n836);
nor (n847,n603,n826);
nand (n848,n849,n1231);
nor (n849,n850,n1225);
nor (n850,n851,n1201);
nor (n851,n852,n1199);
nor (n852,n853,n1176);
nand (n853,n854,n1148);
nand (n854,n855,n1110,n1147);
nand (n855,n856,n976);
nand (n856,n857,n914,n975);
nand (n857,n858,n902);
nand (n858,n859,n889,n901);
nand (n859,n860,n874);
xor (n860,n861,n870);
xor (n861,n862,n866);
xor (n862,n863,n59);
or (n863,n864,n865);
and (n864,n42,n79);
and (n865,n70,n83);
xor (n866,n867,n21);
or (n867,n868,n869);
and (n868,n30,n15);
and (n869,n38,n19);
xor (n870,n871,n28);
or (n871,n872,n873);
and (n872,n146,n57);
and (n873,n195,n62);
nand (n874,n875,n885,n888);
nand (n875,n876,n880);
xor (n876,n877,n28);
or (n877,n878,n879);
and (n878,n195,n57);
and (n879,n199,n62);
xor (n880,n117,n881);
xor (n881,n882,n17);
or (n882,n883,n884);
and (n883,n25,n163);
and (n884,n30,n167);
nand (n885,n886,n880);
xnor (n886,n887,n117);
nand (n887,n765,n111);
nand (n888,n876,n886);
nand (n889,n890,n874);
xor (n890,n891,n897);
xor (n891,n892,n896);
xor (n892,n893,n33);
or (n893,n894,n895);
and (n894,n199,n26);
and (n895,n205,n31);
and (n896,n117,n881);
xor (n897,n898,n45);
or (n898,n899,n900);
and (n899,n98,n39);
and (n900,n103,n43);
nand (n901,n860,n890);
xor (n902,n903,n912);
xor (n903,n904,n908);
xor (n904,n905,n117);
or (n905,n906,n907);
and (n906,n464,n111);
and (n907,n646,n115);
nand (n908,n909,n910,n911);
nand (n909,n892,n896);
nand (n910,n897,n896);
nand (n911,n892,n897);
xor (n912,n913,n785);
xor (n913,n776,n780);
nand (n914,n915,n902);
nand (n915,n916,n952,n974);
nand (n916,n917,n933);
nand (n917,n918,n927,n932);
nand (n918,n919,n923);
xor (n919,n920,n33);
or (n920,n921,n922);
and (n921,n205,n26);
and (n922,n98,n31);
xor (n923,n924,n45);
or (n924,n925,n926);
and (n925,n103,n39);
and (n926,n110,n43);
nand (n927,n928,n923);
xor (n928,n929,n73);
or (n929,n930,n931);
and (n930,n114,n67);
and (n931,n122,n71);
nand (n932,n919,n928);
xor (n933,n934,n943);
xor (n934,n935,n939);
xor (n935,n936,n73);
or (n936,n937,n938);
and (n937,n110,n67);
and (n938,n114,n71);
xor (n939,n940,n101);
or (n940,n941,n942);
and (n941,n122,n196);
and (n942,n126,n200);
xor (n943,n944,n948);
xnor (n944,n945,n165);
nor (n945,n946,n947);
and (n946,n61,n386);
and (n947,n56,n388);
xor (n948,n949,n17);
or (n949,n950,n951);
and (n950,n89,n163);
and (n951,n25,n167);
nand (n952,n953,n933);
nand (n953,n954,n968,n973);
nand (n954,n955,n959);
xor (n955,n956,n101);
or (n956,n957,n958);
and (n957,n126,n196);
and (n958,n324,n200);
and (n959,n960,n964);
xor (n960,n961,n17);
or (n961,n962,n963);
and (n962,n30,n163);
and (n963,n38,n167);
xnor (n964,n965,n165);
nor (n965,n966,n967);
and (n966,n25,n386);
and (n967,n89,n388);
nand (n968,n969,n959);
xor (n969,n970,n106);
or (n970,n971,n972);
and (n971,n464,n99);
and (n972,n646,n104);
nand (n973,n955,n969);
nand (n974,n917,n953);
nand (n975,n858,n915);
nand (n976,n977,n1042,n1109);
nand (n977,n978,n990);
xor (n978,n979,n988);
xor (n979,n980,n984);
nand (n980,n981,n982,n983);
nand (n981,n862,n866);
nand (n982,n870,n866);
nand (n983,n862,n870);
nand (n984,n985,n986,n987);
nand (n985,n935,n939);
nand (n986,n943,n939);
nand (n987,n935,n943);
xor (n988,n989,n802);
xor (n989,n795,n799);
xor (n990,n991,n1034);
xor (n991,n992,n1020);
nand (n992,n993,n1002,n1019);
nand (n993,n994,n998);
xor (n994,n995,n106);
or (n995,n996,n997);
and (n996,n324,n99);
and (n997,n464,n104);
xor (n998,n999,n117);
or (n999,n1000,n1001);
and (n1000,n646,n111);
and (n1001,n765,n115);
nand (n1002,n1003,n998);
nand (n1003,n1004,n1013,n1018);
nand (n1004,n1005,n1009);
xnor (n1005,n1006,n165);
nor (n1006,n1007,n1008);
and (n1007,n89,n386);
and (n1008,n61,n388);
xor (n1009,n1010,n59);
or (n1010,n1011,n1012);
and (n1011,n70,n79);
and (n1012,n146,n83);
nand (n1013,n1014,n1009);
xor (n1014,n1015,n21);
or (n1015,n1016,n1017);
and (n1016,n38,n15);
and (n1017,n42,n19);
nand (n1018,n1005,n1014);
nand (n1019,n994,n1003);
xor (n1020,n1021,n1030);
xor (n1021,n1022,n1026);
xor (n1022,n1023,n45);
or (n1023,n1024,n1025);
and (n1024,n205,n39);
and (n1025,n98,n43);
xor (n1026,n1027,n73);
or (n1027,n1028,n1029);
and (n1028,n103,n67);
and (n1029,n110,n71);
xor (n1030,n1031,n101);
or (n1031,n1032,n1033);
and (n1032,n114,n196);
and (n1033,n122,n200);
xor (n1034,n1035,n1038);
xor (n1035,n1036,n1037);
xor (n1036,n129,n695);
and (n1037,n944,n948);
xor (n1038,n1039,n106);
or (n1039,n1040,n1041);
and (n1040,n126,n99);
and (n1041,n324,n104);
nand (n1042,n1043,n990);
nand (n1043,n1044,n1086,n1108);
nand (n1044,n1045,n1047);
xor (n1045,n1046,n1003);
xor (n1046,n994,n998);
nand (n1047,n1048,n1068,n1085);
nand (n1048,n1049,n1066);
nand (n1049,n1050,n1060,n1065);
nand (n1050,n1051,n1056);
and (n1051,n1052,n106);
xnor (n1052,n1053,n165);
nor (n1053,n1054,n1055);
and (n1054,n30,n386);
and (n1055,n25,n388);
xor (n1056,n1057,n33);
or (n1057,n1058,n1059);
and (n1058,n98,n26);
and (n1059,n103,n31);
nand (n1060,n1061,n1056);
xor (n1061,n1062,n45);
or (n1062,n1063,n1064);
and (n1063,n110,n39);
and (n1064,n114,n43);
nand (n1065,n1051,n1061);
xor (n1066,n1067,n1014);
xor (n1067,n1005,n1009);
nand (n1068,n1069,n1066);
nand (n1069,n1070,n1079,n1084);
nand (n1070,n1071,n1075);
xor (n1071,n1072,n59);
or (n1072,n1073,n1074);
and (n1073,n146,n79);
and (n1074,n195,n83);
xor (n1075,n1076,n21);
or (n1076,n1077,n1078);
and (n1077,n42,n15);
and (n1078,n70,n19);
nand (n1079,n1080,n1075);
xor (n1080,n1081,n28);
or (n1081,n1082,n1083);
and (n1082,n199,n57);
and (n1083,n205,n62);
nand (n1084,n1071,n1080);
nand (n1085,n1049,n1069);
nand (n1086,n1087,n1047);
nand (n1087,n1088,n1104,n1107);
nand (n1088,n1089,n1102);
nand (n1089,n1090,n1099,n1101);
nand (n1090,n1091,n1095);
xor (n1091,n1092,n73);
or (n1092,n1093,n1094);
and (n1093,n122,n67);
and (n1094,n126,n71);
xor (n1095,n1096,n101);
or (n1096,n1097,n1098);
and (n1097,n324,n196);
and (n1098,n464,n200);
nand (n1099,n1100,n1095);
xor (n1100,n960,n964);
nand (n1101,n1091,n1100);
xor (n1102,n1103,n886);
xor (n1103,n876,n880);
nand (n1104,n1105,n1102);
xor (n1105,n1106,n928);
xor (n1106,n919,n923);
nand (n1107,n1089,n1105);
nand (n1108,n1045,n1087);
nand (n1109,n978,n1043);
nand (n1110,n1111,n976);
xor (n1111,n1112,n1135);
xor (n1112,n1113,n1125);
xor (n1113,n1114,n1121);
xor (n1114,n1115,n1119);
nand (n1115,n1116,n1117,n1118);
nand (n1116,n1022,n1026);
nand (n1117,n1030,n1026);
nand (n1118,n1022,n1030);
xor (n1119,n1120,n680);
xor (n1120,n671,n675);
nand (n1121,n1122,n1123,n1124);
nand (n1122,n1036,n1037);
nand (n1123,n1038,n1037);
nand (n1124,n1036,n1038);
xor (n1125,n1126,n1133);
xor (n1126,n1127,n1129);
xor (n1127,n1128,n694);
xor (n1128,n688,n692);
nand (n1129,n1130,n1131,n1132);
nand (n1130,n904,n908);
nand (n1131,n912,n908);
nand (n1132,n904,n912);
xor (n1133,n1134,n767);
xor (n1134,n757,n761);
xor (n1135,n1136,n1143);
xor (n1136,n1137,n1139);
xor (n1137,n1138,n793);
xor (n1138,n774,n790);
nand (n1139,n1140,n1141,n1142);
nand (n1140,n980,n984);
nand (n1141,n988,n984);
nand (n1142,n980,n988);
nand (n1143,n1144,n1145,n1146);
nand (n1144,n992,n1020);
nand (n1145,n1034,n1020);
nand (n1146,n992,n1034);
nand (n1147,n856,n1111);
xor (n1148,n1149,n1172);
xor (n1149,n1150,n1162);
xor (n1150,n1151,n1158);
xor (n1151,n1152,n1154);
xor (n1152,n1153,n686);
xor (n1153,n667,n669);
nand (n1154,n1155,n1156,n1157);
nand (n1155,n1115,n1119);
nand (n1156,n1121,n1119);
nand (n1157,n1115,n1121);
nand (n1158,n1159,n1160,n1161);
nand (n1159,n1127,n1129);
nand (n1160,n1133,n1129);
nand (n1161,n1127,n1133);
xor (n1162,n1163,n1168);
xor (n1163,n1164,n1166);
xor (n1164,n1165,n747);
xor (n1165,n742,n744);
xor (n1166,n1167,n809);
xor (n1167,n755,n772);
nand (n1168,n1169,n1170,n1171);
nand (n1169,n1137,n1139);
nand (n1170,n1143,n1139);
nand (n1171,n1137,n1143);
nand (n1172,n1173,n1174,n1175);
nand (n1173,n1113,n1125);
nand (n1174,n1135,n1125);
nand (n1175,n1113,n1135);
nor (n1176,n1177,n1181);
nand (n1177,n1178,n1179,n1180);
nand (n1178,n1150,n1162);
nand (n1179,n1172,n1162);
nand (n1180,n1150,n1172);
xor (n1181,n1182,n1191);
xor (n1182,n1183,n1187);
nand (n1183,n1184,n1185,n1186);
nand (n1184,n1152,n1154);
nand (n1185,n1158,n1154);
nand (n1186,n1152,n1158);
nand (n1187,n1188,n1189,n1190);
nand (n1188,n1164,n1166);
nand (n1189,n1168,n1166);
nand (n1190,n1164,n1168);
xor (n1191,n1192,n1197);
xor (n1192,n1193,n1195);
xor (n1193,n1194,n630);
xor (n1194,n611,n627);
xor (n1195,n1196,n702);
xor (n1196,n636,n665);
xor (n1197,n1198,n753);
xor (n1198,n740,n750);
not (n1199,n1200);
nand (n1200,n1177,n1181);
not (n1201,n1202);
nor (n1202,n1203,n1218);
nor (n1203,n1204,n1208);
nand (n1204,n1205,n1206,n1207);
nand (n1205,n1183,n1187);
nand (n1206,n1191,n1187);
nand (n1207,n1183,n1191);
xor (n1208,n1209,n1214);
xor (n1209,n1210,n1212);
xor (n1210,n1211,n634);
xor (n1211,n607,n609);
xor (n1212,n1213,n738);
xor (n1213,n708,n710);
nand (n1214,n1215,n1216,n1217);
nand (n1215,n1193,n1195);
nand (n1216,n1197,n1195);
nand (n1217,n1193,n1197);
nor (n1218,n1219,n1223);
nand (n1219,n1220,n1221,n1222);
nand (n1220,n1210,n1212);
nand (n1221,n1214,n1212);
nand (n1222,n1210,n1214);
xor (n1223,n1224,n815);
xor (n1224,n605,n706);
not (n1225,n1226);
nor (n1226,n1227,n1229);
nor (n1227,n1228,n1218);
nand (n1228,n1204,n1208);
not (n1229,n1230);
nand (n1230,n1219,n1223);
nand (n1231,n1232,n2242);
nand (n1232,n1233,n1818);
nor (n1233,n1234,n1803);
nor (n1234,n1235,n1524);
nand (n1235,n1236,n1501);
nor (n1236,n1237,n1478);
nor (n1237,n1238,n1450);
nand (n1238,n1239,n1378,n1449);
nand (n1239,n1240,n1280);
xor (n1240,n1241,n1268);
xor (n1241,n1242,n1244);
xor (n1242,n1243,n1100);
xor (n1243,n1091,n1095);
nand (n1244,n1245,n1254,n1267);
nand (n1245,n1246,n1250);
xor (n1246,n1247,n73);
or (n1247,n1248,n1249);
and (n1248,n126,n67);
and (n1249,n324,n71);
xor (n1250,n1251,n101);
or (n1251,n1252,n1253);
and (n1252,n464,n196);
and (n1253,n646,n200);
nand (n1254,n1255,n1250);
xor (n1255,n1256,n1265);
xor (n1256,n1257,n1261);
xor (n1257,n1258,n17);
or (n1258,n1259,n1260);
and (n1259,n38,n163);
and (n1260,n42,n167);
xor (n1261,n1262,n59);
or (n1262,n1263,n1264);
and (n1263,n195,n79);
and (n1264,n199,n83);
xnor (n1265,n1266,n106);
nand (n1266,n765,n99);
nand (n1267,n1246,n1255);
xor (n1268,n1269,n1278);
xor (n1269,n1270,n1274);
xor (n1270,n1271,n106);
or (n1271,n1272,n1273);
and (n1272,n646,n99);
and (n1273,n765,n104);
nand (n1274,n1275,n1276,n1277);
nand (n1275,n1257,n1261);
nand (n1276,n1265,n1261);
nand (n1277,n1257,n1265);
xor (n1278,n1279,n1080);
xor (n1279,n1071,n1075);
nand (n1280,n1281,n1335,n1377);
nand (n1281,n1282,n1284);
xor (n1282,n1283,n1255);
xor (n1283,n1246,n1250);
xor (n1284,n1285,n1324);
xor (n1285,n1286,n1302);
nand (n1286,n1287,n1296,n1301);
nand (n1287,n1288,n1292);
xor (n1288,n1289,n59);
or (n1289,n1290,n1291);
and (n1290,n199,n79);
and (n1291,n205,n83);
xor (n1292,n1293,n21);
or (n1293,n1294,n1295);
and (n1294,n146,n15);
and (n1295,n195,n19);
nand (n1296,n1297,n1292);
xor (n1297,n1298,n28);
or (n1298,n1299,n1300);
and (n1299,n98,n57);
and (n1300,n103,n62);
nand (n1301,n1288,n1297);
nand (n1302,n1303,n1318,n1323);
nand (n1303,n1304,n1313);
xor (n1304,n1305,n1309);
xnor (n1305,n1306,n165);
nor (n1306,n1307,n1308);
and (n1307,n38,n386);
and (n1308,n30,n388);
xor (n1309,n1310,n17);
or (n1310,n1311,n1312);
and (n1311,n42,n163);
and (n1312,n70,n167);
and (n1313,n1314,n101);
xnor (n1314,n1315,n165);
nor (n1315,n1316,n1317);
and (n1316,n42,n386);
and (n1317,n38,n388);
nand (n1318,n1319,n1313);
xor (n1319,n1320,n33);
or (n1320,n1321,n1322);
and (n1321,n110,n26);
and (n1322,n114,n31);
nand (n1323,n1304,n1319);
xor (n1324,n1325,n1331);
xor (n1325,n1326,n1330);
xor (n1326,n1327,n33);
or (n1327,n1328,n1329);
and (n1328,n103,n26);
and (n1329,n110,n31);
and (n1330,n1305,n1309);
xor (n1331,n1332,n45);
or (n1332,n1333,n1334);
and (n1333,n114,n39);
and (n1334,n122,n43);
nand (n1335,n1336,n1284);
nand (n1336,n1337,n1361,n1376);
nand (n1337,n1338,n1359);
nand (n1338,n1339,n1353,n1358);
nand (n1339,n1340,n1349);
and (n1340,n1341,n1345);
xnor (n1341,n1342,n165);
nor (n1342,n1343,n1344);
and (n1343,n70,n386);
and (n1344,n42,n388);
xor (n1345,n1346,n17);
or (n1346,n1347,n1348);
and (n1347,n146,n163);
and (n1348,n195,n167);
xor (n1349,n1350,n33);
or (n1350,n1351,n1352);
and (n1351,n114,n26);
and (n1352,n122,n31);
nand (n1353,n1354,n1349);
xor (n1354,n1355,n45);
or (n1355,n1356,n1357);
and (n1356,n126,n39);
and (n1357,n324,n43);
nand (n1358,n1340,n1354);
xor (n1359,n1360,n1319);
xor (n1360,n1304,n1313);
nand (n1361,n1362,n1359);
xor (n1362,n1363,n1372);
xor (n1363,n1364,n1368);
xor (n1364,n1365,n45);
or (n1365,n1366,n1367);
and (n1366,n122,n39);
and (n1367,n126,n43);
xor (n1368,n1369,n73);
or (n1369,n1370,n1371);
and (n1370,n324,n67);
and (n1371,n464,n71);
xor (n1372,n1373,n101);
or (n1373,n1374,n1375);
and (n1374,n646,n196);
and (n1375,n765,n200);
nand (n1376,n1338,n1362);
nand (n1377,n1282,n1336);
nand (n1378,n1379,n1280);
xor (n1379,n1380,n1406);
xor (n1380,n1381,n1385);
nand (n1381,n1382,n1383,n1384);
nand (n1382,n1286,n1302);
nand (n1383,n1324,n1302);
nand (n1384,n1286,n1324);
xor (n1385,n1386,n1404);
xor (n1386,n1387,n1400);
nand (n1387,n1388,n1394,n1399);
nand (n1388,n1389,n1393);
xor (n1389,n1390,n21);
or (n1390,n1391,n1392);
and (n1391,n70,n15);
and (n1392,n146,n19);
xor (n1393,n1052,n106);
nand (n1394,n1395,n1393);
xor (n1395,n1396,n28);
or (n1396,n1397,n1398);
and (n1397,n205,n57);
and (n1398,n98,n62);
nand (n1399,n1389,n1395);
nand (n1400,n1401,n1402,n1403);
nand (n1401,n1326,n1330);
nand (n1402,n1331,n1330);
nand (n1403,n1326,n1331);
xor (n1404,n1405,n1061);
xor (n1405,n1051,n1056);
nand (n1406,n1407,n1414,n1448);
nand (n1407,n1408,n1412);
nand (n1408,n1409,n1410,n1411);
nand (n1409,n1364,n1368);
nand (n1410,n1372,n1368);
nand (n1411,n1364,n1372);
xor (n1412,n1413,n1395);
xor (n1413,n1389,n1393);
nand (n1414,n1415,n1412);
nand (n1415,n1416,n1433,n1447);
nand (n1416,n1417,n1431);
nand (n1417,n1418,n1427,n1430);
nand (n1418,n1419,n1423);
xor (n1419,n1420,n17);
or (n1420,n1421,n1422);
and (n1421,n70,n163);
and (n1422,n146,n167);
xor (n1423,n1424,n59);
or (n1424,n1425,n1426);
and (n1425,n205,n79);
and (n1426,n98,n83);
nand (n1427,n1428,n1423);
xnor (n1428,n1429,n101);
nand (n1429,n765,n196);
nand (n1430,n1419,n1428);
xor (n1431,n1432,n1297);
xor (n1432,n1288,n1292);
nand (n1433,n1434,n1431);
nand (n1434,n1435,n1441,n1446);
nand (n1435,n1436,n1440);
xor (n1436,n1437,n21);
or (n1437,n1438,n1439);
and (n1438,n195,n15);
and (n1439,n199,n19);
xor (n1440,n1314,n101);
nand (n1441,n1442,n1440);
xor (n1442,n1443,n28);
or (n1443,n1444,n1445);
and (n1444,n103,n57);
and (n1445,n110,n62);
nand (n1446,n1436,n1442);
nand (n1447,n1417,n1434);
nand (n1448,n1408,n1415);
nand (n1449,n1240,n1379);
xor (n1450,n1451,n1474);
xor (n1451,n1452,n1464);
xor (n1452,n1453,n1460);
xor (n1453,n1454,n1456);
xor (n1454,n1455,n969);
xor (n1455,n955,n959);
nand (n1456,n1457,n1458,n1459);
nand (n1457,n1270,n1274);
nand (n1458,n1278,n1274);
nand (n1459,n1270,n1278);
nand (n1460,n1461,n1462,n1463);
nand (n1461,n1387,n1400);
nand (n1462,n1404,n1400);
nand (n1463,n1387,n1404);
xor (n1464,n1465,n1470);
xor (n1465,n1466,n1468);
xor (n1466,n1467,n1069);
xor (n1467,n1049,n1066);
xor (n1468,n1469,n1105);
xor (n1469,n1089,n1102);
nand (n1470,n1471,n1472,n1473);
nand (n1471,n1242,n1244);
nand (n1472,n1268,n1244);
nand (n1473,n1242,n1268);
nand (n1474,n1475,n1476,n1477);
nand (n1475,n1381,n1385);
nand (n1476,n1406,n1385);
nand (n1477,n1381,n1406);
nor (n1478,n1479,n1483);
nand (n1479,n1480,n1481,n1482);
nand (n1480,n1452,n1464);
nand (n1481,n1474,n1464);
nand (n1482,n1452,n1474);
xor (n1483,n1484,n1493);
xor (n1484,n1485,n1489);
nand (n1485,n1486,n1487,n1488);
nand (n1486,n1454,n1456);
nand (n1487,n1460,n1456);
nand (n1488,n1454,n1460);
nand (n1489,n1490,n1491,n1492);
nand (n1490,n1466,n1468);
nand (n1491,n1470,n1468);
nand (n1492,n1466,n1470);
xor (n1493,n1494,n1499);
xor (n1494,n1495,n1497);
xor (n1495,n1496,n890);
xor (n1496,n860,n874);
xor (n1497,n1498,n953);
xor (n1498,n917,n933);
xor (n1499,n1500,n1087);
xor (n1500,n1045,n1047);
nor (n1501,n1502,n1517);
nor (n1502,n1503,n1507);
nand (n1503,n1504,n1505,n1506);
nand (n1504,n1485,n1489);
nand (n1505,n1493,n1489);
nand (n1506,n1485,n1493);
xor (n1507,n1508,n1513);
xor (n1508,n1509,n1511);
xor (n1509,n1510,n915);
xor (n1510,n858,n902);
xor (n1511,n1512,n1043);
xor (n1512,n978,n990);
nand (n1513,n1514,n1515,n1516);
nand (n1514,n1495,n1497);
nand (n1515,n1499,n1497);
nand (n1516,n1495,n1499);
nor (n1517,n1518,n1522);
nand (n1518,n1519,n1520,n1521);
nand (n1519,n1509,n1511);
nand (n1520,n1513,n1511);
nand (n1521,n1509,n1513);
xor (n1522,n1523,n1111);
xor (n1523,n856,n976);
nor (n1524,n1525,n1797);
nor (n1525,n1526,n1773);
nor (n1526,n1527,n1771);
nor (n1527,n1528,n1746);
nand (n1528,n1529,n1708);
nand (n1529,n1530,n1655,n1707);
nand (n1530,n1531,n1582);
xor (n1531,n1532,n1569);
xor (n1532,n1533,n1554);
nand (n1533,n1534,n1548,n1553);
nand (n1534,n1535,n1544);
and (n1535,n1536,n1540);
xnor (n1536,n1537,n165);
nor (n1537,n1538,n1539);
and (n1538,n195,n386);
and (n1539,n146,n388);
xor (n1540,n1541,n17);
or (n1541,n1542,n1543);
and (n1542,n199,n163);
and (n1543,n205,n167);
xor (n1544,n1545,n33);
or (n1545,n1546,n1547);
and (n1546,n126,n26);
and (n1547,n324,n31);
nand (n1548,n1549,n1544);
xor (n1549,n1550,n45);
or (n1550,n1551,n1552);
and (n1551,n464,n39);
and (n1552,n646,n43);
nand (n1553,n1535,n1549);
xor (n1554,n1555,n1564);
xor (n1555,n1556,n1560);
xor (n1556,n1557,n59);
or (n1557,n1558,n1559);
and (n1558,n98,n79);
and (n1559,n103,n83);
xor (n1560,n1561,n21);
or (n1561,n1562,n1563);
and (n1562,n199,n15);
and (n1563,n205,n19);
and (n1564,n1565,n73);
xnor (n1565,n1566,n165);
nor (n1566,n1567,n1568);
and (n1567,n146,n386);
and (n1568,n70,n388);
nand (n1569,n1570,n1576,n1581);
nand (n1570,n1571,n1575);
xor (n1571,n1572,n21);
or (n1572,n1573,n1574);
and (n1573,n205,n15);
and (n1574,n98,n19);
xor (n1575,n1565,n73);
nand (n1576,n1577,n1575);
xor (n1577,n1578,n28);
or (n1578,n1579,n1580);
and (n1579,n114,n57);
and (n1580,n122,n62);
nand (n1581,n1571,n1577);
xor (n1582,n1583,n1619);
xor (n1583,n1584,n1595);
xor (n1584,n1585,n1591);
xor (n1585,n1586,n1590);
xor (n1586,n1587,n28);
or (n1587,n1588,n1589);
and (n1588,n110,n57);
and (n1589,n114,n62);
xor (n1590,n1341,n1345);
xor (n1591,n1592,n33);
or (n1592,n1593,n1594);
and (n1593,n122,n26);
and (n1594,n126,n31);
xor (n1595,n1596,n1605);
xor (n1596,n1597,n1601);
xor (n1597,n1598,n45);
or (n1598,n1599,n1600);
and (n1599,n324,n39);
and (n1600,n464,n43);
xor (n1601,n1602,n73);
or (n1602,n1603,n1604);
and (n1603,n646,n67);
and (n1604,n765,n71);
nand (n1605,n1606,n1613,n1618);
nand (n1606,n1607,n1611);
xor (n1607,n1608,n17);
or (n1608,n1609,n1610);
and (n1609,n195,n163);
and (n1610,n199,n167);
xnor (n1611,n1612,n73);
nand (n1612,n765,n67);
nand (n1613,n1614,n1611);
xor (n1614,n1615,n59);
or (n1615,n1616,n1617);
and (n1616,n103,n79);
and (n1617,n110,n83);
nand (n1618,n1607,n1614);
nand (n1619,n1620,n1640,n1654);
nand (n1620,n1621,n1623);
xor (n1621,n1622,n1614);
xor (n1622,n1607,n1611);
nand (n1623,n1624,n1633,n1639);
nand (n1624,n1625,n1629);
xor (n1625,n1626,n59);
or (n1626,n1627,n1628);
and (n1627,n110,n79);
and (n1628,n114,n83);
xor (n1629,n1630,n21);
or (n1630,n1631,n1632);
and (n1631,n98,n15);
and (n1632,n103,n19);
nand (n1633,n1634,n1629);
and (n1634,n1635,n45);
xnor (n1635,n1636,n165);
nor (n1636,n1637,n1638);
and (n1637,n199,n386);
and (n1638,n195,n388);
nand (n1639,n1625,n1634);
nand (n1640,n1641,n1623);
nand (n1641,n1642,n1648,n1653);
nand (n1642,n1643,n1647);
xor (n1643,n1644,n28);
or (n1644,n1645,n1646);
and (n1645,n122,n57);
and (n1646,n126,n62);
xor (n1647,n1536,n1540);
nand (n1648,n1649,n1647);
xor (n1649,n1650,n33);
or (n1650,n1651,n1652);
and (n1651,n324,n26);
and (n1652,n464,n31);
nand (n1653,n1643,n1649);
nand (n1654,n1621,n1641);
nand (n1655,n1656,n1582);
nand (n1656,n1657,n1662,n1706);
nand (n1657,n1658,n1660);
xor (n1658,n1659,n1549);
xor (n1659,n1535,n1544);
xor (n1660,n1661,n1577);
xor (n1661,n1571,n1575);
nand (n1662,n1663,n1660);
nand (n1663,n1664,n1683,n1705);
nand (n1664,n1665,n1669);
xor (n1665,n1666,n45);
or (n1666,n1667,n1668);
and (n1667,n646,n39);
and (n1668,n765,n43);
nand (n1669,n1670,n1677,n1682);
nand (n1670,n1671,n1675);
xor (n1671,n1672,n17);
or (n1672,n1673,n1674);
and (n1673,n205,n163);
and (n1674,n98,n167);
xnor (n1675,n1676,n45);
nand (n1676,n765,n39);
nand (n1677,n1678,n1675);
xor (n1678,n1679,n59);
or (n1679,n1680,n1681);
and (n1680,n114,n79);
and (n1681,n122,n83);
nand (n1682,n1671,n1678);
nand (n1683,n1684,n1669);
nand (n1684,n1685,n1699,n1704);
nand (n1685,n1686,n1690);
xor (n1686,n1687,n21);
or (n1687,n1688,n1689);
and (n1688,n103,n15);
and (n1689,n110,n19);
and (n1690,n1691,n1695);
xnor (n1691,n1692,n165);
nor (n1692,n1693,n1694);
and (n1693,n205,n386);
and (n1694,n199,n388);
xor (n1695,n1696,n17);
or (n1696,n1697,n1698);
and (n1697,n98,n163);
and (n1698,n103,n167);
nand (n1699,n1700,n1690);
xor (n1700,n1701,n28);
or (n1701,n1702,n1703);
and (n1702,n126,n57);
and (n1703,n324,n62);
nand (n1704,n1686,n1700);
nand (n1705,n1665,n1684);
nand (n1706,n1658,n1663);
nand (n1707,n1531,n1656);
xor (n1708,n1709,n1724);
xor (n1709,n1710,n1720);
xor (n1710,n1711,n1718);
xor (n1711,n1712,n1716);
nand (n1712,n1713,n1714,n1715);
nand (n1713,n1556,n1560);
nand (n1714,n1564,n1560);
nand (n1715,n1556,n1564);
xor (n1716,n1717,n1354);
xor (n1717,n1340,n1349);
xor (n1718,n1719,n1442);
xor (n1719,n1436,n1440);
nand (n1720,n1721,n1722,n1723);
nand (n1721,n1584,n1595);
nand (n1722,n1619,n1595);
nand (n1723,n1584,n1619);
xor (n1724,n1725,n1734);
xor (n1725,n1726,n1730);
nand (n1726,n1727,n1728,n1729);
nand (n1727,n1597,n1601);
nand (n1728,n1605,n1601);
nand (n1729,n1597,n1605);
nand (n1730,n1731,n1732,n1733);
nand (n1731,n1533,n1554);
nand (n1732,n1569,n1554);
nand (n1733,n1533,n1569);
xor (n1734,n1735,n1744);
xor (n1735,n1736,n1740);
xor (n1736,n1737,n73);
or (n1737,n1738,n1739);
and (n1738,n464,n67);
and (n1739,n646,n71);
nand (n1740,n1741,n1742,n1743);
nand (n1741,n1586,n1590);
nand (n1742,n1591,n1590);
nand (n1743,n1586,n1591);
xor (n1744,n1745,n1428);
xor (n1745,n1419,n1423);
nor (n1746,n1747,n1751);
nand (n1747,n1748,n1749,n1750);
nand (n1748,n1710,n1720);
nand (n1749,n1724,n1720);
nand (n1750,n1710,n1724);
xor (n1751,n1752,n1759);
xor (n1752,n1753,n1755);
xor (n1753,n1754,n1362);
xor (n1754,n1338,n1359);
nand (n1755,n1756,n1757,n1758);
nand (n1756,n1726,n1730);
nand (n1757,n1734,n1730);
nand (n1758,n1726,n1734);
xor (n1759,n1760,n1769);
xor (n1760,n1761,n1765);
nand (n1761,n1762,n1763,n1764);
nand (n1762,n1736,n1740);
nand (n1763,n1744,n1740);
nand (n1764,n1736,n1744);
nand (n1765,n1766,n1767,n1768);
nand (n1766,n1712,n1716);
nand (n1767,n1718,n1716);
nand (n1768,n1712,n1718);
xor (n1769,n1770,n1434);
xor (n1770,n1417,n1431);
not (n1771,n1772);
nand (n1772,n1747,n1751);
not (n1773,n1774);
nor (n1774,n1775,n1790);
nor (n1775,n1776,n1780);
nand (n1776,n1777,n1778,n1779);
nand (n1777,n1753,n1755);
nand (n1778,n1759,n1755);
nand (n1779,n1753,n1759);
xor (n1780,n1781,n1788);
xor (n1781,n1782,n1784);
xor (n1782,n1783,n1415);
xor (n1783,n1408,n1412);
nand (n1784,n1785,n1786,n1787);
nand (n1785,n1761,n1765);
nand (n1786,n1769,n1765);
nand (n1787,n1761,n1769);
xor (n1788,n1789,n1336);
xor (n1789,n1282,n1284);
nor (n1790,n1791,n1795);
nand (n1791,n1792,n1793,n1794);
nand (n1792,n1782,n1784);
nand (n1793,n1788,n1784);
nand (n1794,n1782,n1788);
xor (n1795,n1796,n1379);
xor (n1796,n1240,n1280);
not (n1797,n1798);
nor (n1798,n1799,n1801);
nor (n1799,n1800,n1790);
nand (n1800,n1776,n1780);
not (n1801,n1802);
nand (n1802,n1791,n1795);
not (n1803,n1804);
nor (n1804,n1805,n1812);
nor (n1805,n1806,n1811);
nor (n1806,n1807,n1809);
nor (n1807,n1808,n1478);
nand (n1808,n1238,n1450);
not (n1809,n1810);
nand (n1810,n1479,n1483);
not (n1811,n1501);
not (n1812,n1813);
nor (n1813,n1814,n1816);
nor (n1814,n1815,n1517);
nand (n1815,n1503,n1507);
not (n1816,n1817);
nand (n1817,n1518,n1522);
nand (n1818,n1819,n1823);
nor (n1819,n1820,n1235);
nand (n1820,n1821,n1774);
nor (n1821,n1822,n1746);
nor (n1822,n1529,n1708);
nand (n1823,n1824,n2135);
nor (n1824,n1825,n2120);
nor (n1825,n1826,n1991);
nand (n1826,n1827,n1968);
nor (n1827,n1828,n1945);
nor (n1828,n1829,n1918);
nand (n1829,n1830,n1875,n1917);
nand (n1830,n1831,n1843);
xor (n1831,n1832,n1838);
xor (n1832,n1833,n1834);
xor (n1833,n1691,n1695);
xor (n1834,n1835,n33);
or (n1835,n1836,n1837);
and (n1836,n646,n26);
and (n1837,n765,n31);
and (n1838,n33,n1839);
xor (n1839,n1840,n17);
or (n1840,n1841,n1842);
and (n1841,n103,n163);
and (n1842,n110,n167);
nand (n1843,n1844,n1861,n1874);
nand (n1844,n1845,n1846);
xor (n1845,n33,n1839);
nand (n1846,n1847,n1856,n1860);
nand (n1847,n1848,n1852);
xor (n1848,n1849,n59);
or (n1849,n1850,n1851);
and (n1850,n324,n79);
and (n1851,n464,n83);
xor (n1852,n1853,n21);
or (n1853,n1854,n1855);
and (n1854,n122,n15);
and (n1855,n126,n19);
nand (n1856,n1857,n1852);
and (n1857,n28,n1858);
xnor (n1858,n1859,n28);
nand (n1859,n765,n57);
nand (n1860,n1848,n1857);
nand (n1861,n1862,n1846);
xor (n1862,n1863,n1870);
xor (n1863,n1864,n1868);
xnor (n1864,n1865,n165);
nor (n1865,n1866,n1867);
and (n1866,n98,n386);
and (n1867,n205,n388);
xnor (n1868,n1869,n33);
nand (n1869,n765,n26);
xor (n1870,n1871,n59);
or (n1871,n1872,n1873);
and (n1872,n126,n79);
and (n1873,n324,n83);
nand (n1874,n1845,n1862);
nand (n1875,n1876,n1843);
xor (n1876,n1877,n1896);
xor (n1877,n1878,n1882);
nand (n1878,n1879,n1880,n1881);
nand (n1879,n1864,n1868);
nand (n1880,n1870,n1868);
nand (n1881,n1864,n1870);
xor (n1882,n1883,n1892);
xor (n1883,n1884,n1888);
xor (n1884,n1885,n59);
or (n1885,n1886,n1887);
and (n1886,n122,n79);
and (n1887,n126,n83);
xor (n1888,n1889,n21);
or (n1889,n1890,n1891);
and (n1890,n110,n15);
and (n1891,n114,n19);
xor (n1892,n1893,n28);
or (n1893,n1894,n1895);
and (n1894,n324,n57);
and (n1895,n464,n62);
nand (n1896,n1897,n1911,n1916);
nand (n1897,n1898,n1902);
xor (n1898,n1899,n21);
or (n1899,n1900,n1901);
and (n1900,n114,n15);
and (n1901,n122,n19);
and (n1902,n1903,n1907);
xnor (n1903,n1904,n165);
nor (n1904,n1905,n1906);
and (n1905,n103,n386);
and (n1906,n98,n388);
xor (n1907,n1908,n17);
or (n1908,n1909,n1910);
and (n1909,n110,n163);
and (n1910,n114,n167);
nand (n1911,n1912,n1902);
xor (n1912,n1913,n28);
or (n1913,n1914,n1915);
and (n1914,n464,n57);
and (n1915,n646,n62);
nand (n1916,n1898,n1912);
nand (n1917,n1831,n1876);
xor (n1918,n1919,n1933);
xor (n1919,n1920,n1929);
xor (n1920,n1921,n1927);
xor (n1921,n1922,n1926);
xor (n1922,n1923,n33);
or (n1923,n1924,n1925);
and (n1924,n464,n26);
and (n1925,n646,n31);
xor (n1926,n1635,n45);
xor (n1927,n1928,n1678);
xor (n1928,n1671,n1675);
nand (n1929,n1930,n1931,n1932);
nand (n1930,n1878,n1882);
nand (n1931,n1896,n1882);
nand (n1932,n1878,n1896);
xor (n1933,n1934,n1943);
xor (n1934,n1935,n1939);
nand (n1935,n1936,n1937,n1938);
nand (n1936,n1833,n1834);
nand (n1937,n1838,n1834);
nand (n1938,n1833,n1838);
nand (n1939,n1940,n1941,n1942);
nand (n1940,n1884,n1888);
nand (n1941,n1892,n1888);
nand (n1942,n1884,n1892);
xor (n1943,n1944,n1700);
xor (n1944,n1686,n1690);
nor (n1945,n1946,n1950);
nand (n1946,n1947,n1948,n1949);
nand (n1947,n1920,n1929);
nand (n1948,n1933,n1929);
nand (n1949,n1920,n1933);
xor (n1950,n1951,n1958);
xor (n1951,n1952,n1954);
xor (n1952,n1953,n1684);
xor (n1953,n1665,n1669);
nand (n1954,n1955,n1956,n1957);
nand (n1955,n1935,n1939);
nand (n1956,n1943,n1939);
nand (n1957,n1935,n1943);
xor (n1958,n1959,n1964);
xor (n1959,n1960,n1962);
xor (n1960,n1961,n1634);
xor (n1961,n1625,n1629);
xor (n1962,n1963,n1649);
xor (n1963,n1643,n1647);
nand (n1964,n1965,n1966,n1967);
nand (n1965,n1922,n1926);
nand (n1966,n1927,n1926);
nand (n1967,n1922,n1927);
nor (n1968,n1969,n1984);
nor (n1969,n1970,n1974);
nand (n1970,n1971,n1972,n1973);
nand (n1971,n1952,n1954);
nand (n1972,n1958,n1954);
nand (n1973,n1952,n1958);
xor (n1974,n1975,n1982);
xor (n1975,n1976,n1978);
xor (n1976,n1977,n1641);
xor (n1977,n1621,n1623);
nand (n1978,n1979,n1980,n1981);
nand (n1979,n1960,n1962);
nand (n1980,n1964,n1962);
nand (n1981,n1960,n1964);
xor (n1982,n1983,n1663);
xor (n1983,n1658,n1660);
nor (n1984,n1985,n1989);
nand (n1985,n1986,n1987,n1988);
nand (n1986,n1976,n1978);
nand (n1987,n1982,n1978);
nand (n1988,n1976,n1982);
xor (n1989,n1990,n1656);
xor (n1990,n1531,n1582);
nor (n1991,n1992,n2114);
nor (n1992,n1993,n2090);
nor (n1993,n1994,n2087);
nor (n1994,n1995,n2063);
nand (n1995,n1996,n2035);
or (n1996,n1997,n2021,n2034);
and (n1997,n1998,n2007);
xor (n1998,n1999,n2003);
xnor (n1999,n2000,n165);
nor (n2000,n2001,n2002);
and (n2001,n114,n386);
and (n2002,n110,n388);
xnor (n2003,n2004,n17);
nor (n2004,n2005,n2006);
and (n2005,n126,n167);
and (n2006,n122,n163);
or (n2007,n2008,n2015,n2020);
and (n2008,n2009,n2011);
not (n2009,n2010);
nand (n2010,n765,n79);
xnor (n2011,n2012,n165);
nor (n2012,n2013,n2014);
and (n2013,n122,n386);
and (n2014,n114,n388);
and (n2015,n2011,n2016);
xnor (n2016,n2017,n17);
nor (n2017,n2018,n2019);
and (n2018,n324,n167);
and (n2019,n126,n163);
and (n2020,n2009,n2016);
and (n2021,n2007,n2022);
xor (n2022,n2023,n2030);
xor (n2023,n2024,n2026);
and (n2024,n59,n2025);
xnor (n2025,n2010,n59);
xnor (n2026,n2027,n21);
nor (n2027,n2028,n2029);
and (n2028,n464,n19);
and (n2029,n324,n15);
xnor (n2030,n2031,n59);
nor (n2031,n2032,n2033);
and (n2032,n765,n83);
and (n2033,n646,n79);
and (n2034,n1998,n2022);
xor (n2035,n2036,n2052);
xor (n2036,n2037,n2041);
or (n2037,n2038,n2039,n2040);
and (n2038,n2024,n2026);
and (n2039,n2026,n2030);
and (n2040,n2024,n2030);
xor (n2041,n2042,n2048);
xor (n2042,n2043,n2044);
and (n2043,n1999,n2003);
xnor (n2044,n2045,n21);
nor (n2045,n2046,n2047);
and (n2046,n324,n19);
and (n2047,n126,n15);
xnor (n2048,n2049,n59);
nor (n2049,n2050,n2051);
and (n2050,n646,n83);
and (n2051,n464,n79);
xor (n2052,n2053,n2059);
xor (n2053,n2054,n2055);
not (n2054,n1859);
xnor (n2055,n2056,n165);
nor (n2056,n2057,n2058);
and (n2057,n110,n386);
and (n2058,n103,n388);
xnor (n2059,n2060,n17);
nor (n2060,n2061,n2062);
and (n2061,n122,n167);
and (n2062,n114,n163);
nor (n2063,n2064,n2068);
or (n2064,n2065,n2066,n2067);
and (n2065,n2037,n2041);
and (n2066,n2041,n2052);
and (n2067,n2037,n2052);
xor (n2068,n2069,n2076);
xor (n2069,n2070,n2074);
or (n2070,n2071,n2072,n2073);
and (n2071,n2043,n2044);
and (n2072,n2044,n2048);
and (n2073,n2043,n2048);
xor (n2074,n2075,n1857);
xor (n2075,n1848,n1852);
xor (n2076,n2077,n2083);
xor (n2077,n2078,n2082);
xor (n2078,n2079,n28);
or (n2079,n2080,n2081);
and (n2080,n646,n57);
and (n2081,n765,n62);
xor (n2082,n1903,n1907);
or (n2083,n2084,n2085,n2086);
and (n2084,n2054,n2055);
and (n2085,n2055,n2059);
and (n2086,n2054,n2059);
not (n2087,n2088);
not (n2088,n2089);
and (n2089,n2064,n2068);
not (n2090,n2091);
nor (n2091,n2092,n2107);
nor (n2092,n2093,n2097);
nand (n2093,n2094,n2095,n2096);
nand (n2094,n2070,n2074);
nand (n2095,n2076,n2074);
nand (n2096,n2070,n2076);
xor (n2097,n2098,n2105);
xor (n2098,n2099,n2101);
xor (n2099,n2100,n1912);
xor (n2100,n1898,n1902);
nand (n2101,n2102,n2103,n2104);
nand (n2102,n2078,n2082);
nand (n2103,n2083,n2082);
nand (n2104,n2078,n2083);
xor (n2105,n2106,n1862);
xor (n2106,n1845,n1846);
nor (n2107,n2108,n2112);
nand (n2108,n2109,n2110,n2111);
nand (n2109,n2099,n2101);
nand (n2110,n2105,n2101);
nand (n2111,n2099,n2105);
xor (n2112,n2113,n1876);
xor (n2113,n1831,n1843);
not (n2114,n2115);
nor (n2115,n2116,n2118);
nor (n2116,n2117,n2107);
nand (n2117,n2093,n2097);
not (n2118,n2119);
nand (n2119,n2108,n2112);
not (n2120,n2121);
nor (n2121,n2122,n2129);
nor (n2122,n2123,n2128);
nor (n2123,n2124,n2126);
nor (n2124,n2125,n1945);
nand (n2125,n1829,n1918);
not (n2126,n2127);
nand (n2127,n1946,n1950);
not (n2128,n1968);
not (n2129,n2130);
nor (n2130,n2131,n2133);
nor (n2131,n2132,n1984);
nand (n2132,n1970,n1974);
not (n2133,n2134);
nand (n2134,n1985,n1989);
nand (n2135,n2136,n2140);
nor (n2136,n2137,n1826);
nand (n2137,n2138,n2091);
nor (n2138,n2139,n2063);
nor (n2139,n1996,n2035);
or (n2140,n2141,n2163);
and (n2141,n2142,n2144);
xor (n2142,n2143,n2022);
xor (n2143,n1998,n2007);
or (n2144,n2145,n2159,n2162);
and (n2145,n2146,n2155);
and (n2146,n2147,n2151);
xnor (n2147,n2148,n165);
nor (n2148,n2149,n2150);
and (n2149,n126,n386);
and (n2150,n122,n388);
xnor (n2151,n2152,n17);
nor (n2152,n2153,n2154);
and (n2153,n464,n167);
and (n2154,n324,n163);
xnor (n2155,n2156,n21);
nor (n2156,n2157,n2158);
and (n2157,n646,n19);
and (n2158,n464,n15);
and (n2159,n2155,n2160);
xor (n2160,n2161,n2016);
xor (n2161,n2009,n2011);
and (n2162,n2146,n2160);
and (n2163,n2164,n2165);
xor (n2164,n2142,n2144);
or (n2165,n2166,n2181);
and (n2166,n2167,n2179);
or (n2167,n2168,n2173,n2178);
and (n2168,n2169,n2170);
xor (n2169,n2147,n2151);
and (n2170,n21,n2171);
xnor (n2171,n2172,n21);
nand (n2172,n765,n15);
and (n2173,n2170,n2174);
xnor (n2174,n2175,n21);
nor (n2175,n2176,n2177);
and (n2176,n765,n19);
and (n2177,n646,n15);
and (n2178,n2169,n2174);
xor (n2179,n2180,n2160);
xor (n2180,n2146,n2155);
and (n2181,n2182,n2183);
xor (n2182,n2167,n2179);
or (n2183,n2184,n2200);
and (n2184,n2185,n2187);
xor (n2185,n2186,n2174);
xor (n2186,n2169,n2170);
or (n2187,n2188,n2194,n2199);
and (n2188,n2189,n2190);
not (n2189,n2172);
xnor (n2190,n2191,n165);
nor (n2191,n2192,n2193);
and (n2192,n324,n386);
and (n2193,n126,n388);
and (n2194,n2190,n2195);
xnor (n2195,n2196,n17);
nor (n2196,n2197,n2198);
and (n2197,n646,n167);
and (n2198,n464,n163);
and (n2199,n2189,n2195);
and (n2200,n2201,n2202);
xor (n2201,n2185,n2187);
or (n2202,n2203,n2214);
and (n2203,n2204,n2206);
xor (n2204,n2205,n2195);
xor (n2205,n2189,n2190);
and (n2206,n2207,n2210);
and (n2207,n17,n2208);
xnor (n2208,n2209,n17);
nand (n2209,n765,n163);
xnor (n2210,n2211,n165);
nor (n2211,n2212,n2213);
and (n2212,n464,n386);
and (n2213,n324,n388);
and (n2214,n2215,n2216);
xor (n2215,n2204,n2206);
or (n2216,n2217,n2223);
and (n2217,n2218,n2222);
xnor (n2218,n2219,n17);
nor (n2219,n2220,n2221);
and (n2220,n765,n167);
and (n2221,n646,n163);
xor (n2222,n2207,n2210);
and (n2223,n2224,n2225);
xor (n2224,n2218,n2222);
or (n2225,n2226,n2232);
and (n2226,n2227,n2231);
xnor (n2227,n2228,n165);
nor (n2228,n2229,n2230);
and (n2229,n646,n386);
and (n2230,n464,n388);
not (n2231,n2209);
and (n2232,n2233,n2234);
xor (n2233,n2227,n2231);
and (n2234,n2235,n2239);
xnor (n2235,n2236,n165);
nor (n2236,n2237,n2238);
and (n2237,n765,n386);
and (n2238,n646,n388);
and (n2239,n2240,n165);
xnor (n2240,n2241,n165);
nand (n2241,n765,n388);
not (n2242,n2243);
nand (n2243,n2244,n1202);
nor (n2244,n2245,n1176);
nor (n2245,n854,n1148);
not (n2246,n2247);
nor (n2247,n3,n508);
nand (n2248,n2249,n2337);
not (n2249,n2250);
nor (n2250,n2251,n2255);
nand (n2251,n2252,n2253,n2254);
nand (n2252,n510,n514);
nand (n2253,n594,n514);
nand (n2254,n510,n594);
xor (n2255,n2256,n2333);
xor (n2256,n2257,n2303);
xor (n2257,n2258,n2273);
xor (n2258,n2259,n2269);
xor (n2259,n2260,n2265);
xor (n2260,n2261,n129);
xor (n2261,n2262,n106);
or (n2262,n2263,n2264);
and (n2263,n146,n99);
and (n2264,n195,n104);
nand (n2265,n2266,n2267,n2268);
nand (n2266,n544,n548);
nand (n2267,n552,n548);
nand (n2268,n544,n552);
nand (n2269,n2270,n2271,n2272);
nand (n2270,n572,n576);
nand (n2271,n590,n576);
nand (n2272,n572,n590);
xor (n2273,n2274,n2299);
xor (n2274,n2275,n2285);
xor (n2275,n2276,n2281);
xor (n2276,n528,n2277);
xor (n2277,n2278,n28);
or (n2278,n2279,n2280);
and (n2279,n14,n57);
and (n2280,n82,n62);
xor (n2281,n2282,n45);
or (n2282,n2283,n2284);
and (n2283,n89,n39);
and (n2284,n25,n43);
xor (n2285,n2286,n2295);
xor (n2286,n2287,n2291);
xor (n2287,n2288,n33);
or (n2288,n2289,n2290);
and (n2289,n56,n26);
and (n2290,n61,n31);
xor (n2291,n2292,n73);
or (n2292,n2293,n2294);
and (n2293,n30,n67);
and (n2294,n38,n71);
xor (n2295,n2296,n101);
or (n2296,n2297,n2298);
and (n2297,n42,n196);
and (n2298,n70,n200);
nand (n2299,n2300,n2301,n2302);
nand (n2300,n578,n582);
nand (n2301,n586,n582);
nand (n2302,n578,n586);
xor (n2303,n2304,n2329);
xor (n2304,n2305,n2309);
nand (n2305,n2306,n2307,n2308);
nand (n2306,n518,n522);
nand (n2307,n536,n522);
nand (n2308,n518,n536);
xor (n2309,n2310,n2325);
xor (n2310,n2311,n2315);
nand (n2311,n2312,n2313,n2314);
nand (n2312,n524,n528);
nand (n2313,n532,n528);
nand (n2314,n524,n532);
xor (n2315,n2316,n529);
xor (n2316,n2317,n2321);
xor (n2317,n2318,n117);
or (n2318,n2319,n2320);
and (n2319,n199,n111);
and (n2320,n205,n115);
xor (n2321,n2322,n129);
or (n2322,n2323,n2324);
and (n2323,n98,n123);
and (n2324,n103,n127);
nand (n2325,n2326,n2327,n2328);
nand (n2326,n129,n538);
nand (n2327,n542,n538);
nand (n2328,n129,n542);
nand (n2329,n2330,n2331,n2332);
nand (n2330,n562,n566);
nand (n2331,n570,n566);
nand (n2332,n562,n570);
nand (n2333,n2334,n2335,n2336);
nand (n2334,n516,n556);
nand (n2335,n560,n556);
nand (n2336,n516,n560);
nand (n2337,n2251,n2255);
xor (n2338,n2339,n2664);
xor (n2339,n2340,n2463);
xor (n2340,n2341,n2409);
xor (n2341,n2342,n2383);
or (n2342,n2343,n2366,n2382);
and (n2343,n2344,n2355);
xor (n2344,n2345,n570);
xor (n2345,n2346,n566);
or (n2346,n2347,n2352,n2354);
and (n2347,n2348,n47);
or (n2348,n2349,n2350,n2351);
and (n2349,n85,n22);
not (n2350,n34);
and (n2351,n85,n35);
and (n2352,n47,n2353);
not (n2353,n74);
and (n2354,n2348,n2353);
or (n2355,n2356,n2359,n2365);
and (n2356,n2357,n184);
xor (n2357,n2358,n2353);
xor (n2358,n2348,n47);
and (n2359,n184,n2360);
or (n2360,n2361,n2362,n2364);
not (n2361,n286);
and (n2362,n270,n2363);
not (n2363,n267);
and (n2364,n251,n2363);
and (n2365,n2357,n2360);
and (n2366,n2355,n2367);
xor (n2367,n2368,n2377);
xor (n2368,n2369,n2373);
or (n2369,n2370,n2371,n2372);
and (n2370,n11,n76);
not (n2371,n541);
and (n2372,n11,n86);
xor (n2373,n2374,n2376);
xor (n2374,n542,n2375);
not (n2375,n522);
not (n2376,n519);
or (n2377,n2378,n2379,n2381);
and (n2378,n85,n240);
and (n2379,n240,n2380);
not (n2380,n92);
and (n2381,n85,n2380);
and (n2382,n2344,n2367);
xor (n2383,n2384,n2393);
xor (n2384,n2385,n2389);
or (n2385,n2386,n2387,n2388);
and (n2386,n2346,n566);
not (n2387,n2331);
and (n2388,n2346,n570);
or (n2389,n2390,n2391,n2392);
and (n2390,n2369,n2373);
and (n2391,n2373,n2377);
and (n2392,n2369,n2377);
xor (n2393,n2394,n2401);
xor (n2394,n2395,n2269);
xor (n2395,n2396,n2397);
xor (n2396,n2265,n2299);
or (n2397,n2398,n2399,n2400);
and (n2398,n529,n532);
not (n2399,n2314);
and (n2400,n529,n524);
xor (n2401,n2402,n2407);
xor (n2402,n2275,n2403);
or (n2403,n2404,n2405,n2406);
and (n2404,n542,n2375);
and (n2405,n2375,n2376);
and (n2406,n542,n2376);
xor (n2407,n2408,n2316);
xor (n2408,n2261,n2285);
or (n2409,n2410,n2425,n2462);
and (n2410,n2411,n2423);
or (n2411,n2412,n2419,n2422);
and (n2412,n2413,n2417);
or (n2413,n2414,n2415,n2416);
and (n2414,n229,n289);
and (n2415,n289,n367);
and (n2416,n229,n367);
xor (n2417,n2418,n2380);
xor (n2418,n85,n240);
and (n2419,n2417,n2420);
and (n2420,n344,n2421);
not (n2421,n342);
and (n2422,n2413,n2420);
xor (n2423,n2424,n2367);
xor (n2424,n2344,n2355);
and (n2425,n2423,n2426);
or (n2426,n2427,n2447,n2461);
and (n2427,n2428,n2445);
or (n2428,n2429,n2434,n2444);
and (n2429,n2430,n293);
or (n2430,n2431,n2432,n2433);
and (n2431,n160,n152);
not (n2432,n235);
and (n2433,n160,n155);
and (n2434,n293,n2435);
or (n2435,n2436,n2441,n2443);
and (n2436,n159,n2437);
or (n2437,n2438,n2439,n2440);
and (n2438,n159,n172);
not (n2439,n181);
and (n2440,n159,n177);
and (n2441,n2437,n2442);
not (n2442,n150);
and (n2443,n159,n2442);
and (n2444,n2430,n2435);
xor (n2445,n2446,n2360);
xor (n2446,n2357,n184);
and (n2447,n2445,n2448);
or (n2448,n2449,n2453,n2460);
and (n2449,n2450,n2452);
xor (n2450,n2451,n367);
xor (n2451,n229,n289);
not (n2452,n829);
and (n2453,n2452,n2454);
or (n2454,n2455,n2458,n2459);
and (n2455,n2456,n417);
and (n2456,n427,n2457);
not (n2457,n429);
and (n2458,n417,n503);
and (n2459,n2456,n503);
and (n2460,n2450,n2454);
and (n2461,n2428,n2448);
and (n2462,n2411,n2426);
or (n2463,n2464,n2539,n2663);
and (n2464,n2465,n2537);
or (n2465,n2466,n2533,n2536);
and (n2466,n2467,n2469);
xor (n2467,n2468,n2420);
xor (n2468,n2413,n2417);
or (n2469,n2470,n2504,n2532);
and (n2470,n2471,n2502);
or (n2471,n2472,n2490,n2501);
and (n2472,n2473,n2482);
and (n2473,n2474,n452);
or (n2474,n2475,n2480,n2481);
and (n2475,n2476,n456);
or (n2476,n2477,n2478,n2479);
and (n2477,n382,n468);
not (n2478,n467);
and (n2479,n382,n472);
not (n2480,n455);
and (n2481,n2476,n460);
or (n2482,n2483,n2488,n2489);
and (n2483,n397,n2484);
or (n2484,n2485,n2486,n2487);
and (n2485,n382,n434);
not (n2486,n448);
and (n2487,n382,n444);
and (n2488,n2484,n712);
and (n2489,n397,n712);
and (n2490,n2482,n2491);
or (n2491,n2492,n2498,n2500);
and (n2492,n2493,n2494);
not (n2493,n608);
or (n2494,n2495,n2496,n2497);
and (n2495,n383,n378);
not (n2496,n395);
and (n2497,n383,n391);
and (n2498,n2494,n2499);
not (n2499,n481);
and (n2500,n2493,n2499);
and (n2501,n2473,n2491);
xor (n2502,n2503,n2435);
xor (n2503,n2430,n293);
and (n2504,n2502,n2505);
or (n2505,n2506,n2528,n2531);
and (n2506,n2507,n2509);
xor (n2507,n2508,n2442);
xor (n2508,n159,n2437);
or (n2509,n2510,n2519,n2527);
and (n2510,n2511,n2518);
or (n2511,n2512,n2514,n2517);
and (n2512,n731,n2513);
not (n2513,n719);
and (n2514,n2513,n2515);
xor (n2515,n2516,n444);
xor (n2516,n382,n434);
and (n2517,n731,n2515);
xor (n2518,n2474,n452);
and (n2519,n2518,n2520);
or (n2520,n2521,n2525,n2526);
and (n2521,n2522,n2523);
not (n2522,n734);
xor (n2523,n2524,n460);
xor (n2524,n2476,n456);
and (n2525,n2523,n703);
and (n2526,n2522,n703);
and (n2527,n2511,n2520);
and (n2528,n2509,n2529);
xor (n2529,n2530,n503);
xor (n2530,n2456,n417);
and (n2531,n2507,n2529);
and (n2532,n2471,n2505);
and (n2533,n2469,n2534);
xor (n2534,n2535,n2448);
xor (n2535,n2428,n2445);
and (n2536,n2467,n2534);
xor (n2537,n2538,n2426);
xor (n2538,n2411,n2423);
and (n2539,n2537,n2540);
or (n2540,n2541,n2574,n2662);
and (n2541,n2542,n2572);
or (n2542,n2543,n2568,n2571);
and (n2543,n2544,n2546);
xor (n2544,n2545,n2454);
xor (n2545,n2450,n2452);
or (n2546,n2547,n2564,n2567);
and (n2547,n2548,n2550);
xor (n2548,n2549,n2491);
xor (n2549,n2473,n2482);
or (n2550,n2551,n2556,n2563);
and (n2551,n2552,n2554);
xor (n2552,n2553,n712);
xor (n2553,n397,n2484);
xor (n2554,n2555,n2499);
xor (n2555,n2493,n2494);
and (n2556,n2554,n2557);
and (n2557,n636,n2558);
or (n2558,n2559,n2560,n2562);
not (n2559,n685);
and (n2560,n686,n2561);
not (n2561,n667);
and (n2562,n669,n2561);
and (n2563,n2552,n2557);
and (n2564,n2550,n2565);
xor (n2565,n2566,n2529);
xor (n2566,n2507,n2509);
and (n2567,n2548,n2565);
and (n2568,n2546,n2569);
xor (n2569,n2570,n2505);
xor (n2570,n2471,n2502);
and (n2571,n2544,n2569);
xor (n2572,n2573,n2534);
xor (n2573,n2467,n2469);
and (n2574,n2572,n2575);
or (n2575,n2576,n2633,n2661);
and (n2576,n2577,n2579);
xor (n2577,n2578,n2569);
xor (n2578,n2544,n2546);
or (n2579,n2580,n2612,n2632);
and (n2580,n2581,n2610);
or (n2581,n2582,n2595,n2609);
and (n2582,n2583,n2593);
or (n2583,n2584,n2591,n2592);
and (n2584,n2585,n2589);
or (n2585,n2586,n2587,n2588);
and (n2586,n439,n622);
and (n2587,n622,n742);
and (n2588,n439,n742);
xor (n2589,n2590,n2515);
xor (n2590,n731,n2513);
and (n2591,n2589,n753);
and (n2592,n2585,n753);
xor (n2593,n2594,n2520);
xor (n2594,n2511,n2518);
and (n2595,n2593,n2596);
or (n2596,n2597,n2606,n2608);
and (n2597,n2598,n2604);
or (n2598,n2599,n2600,n2603);
and (n2599,n748,n613);
and (n2600,n613,n2601);
xor (n2601,n2602,n742);
xor (n2602,n439,n622);
and (n2603,n748,n2601);
xor (n2604,n2605,n703);
xor (n2605,n2522,n2523);
and (n2606,n2604,n2607);
xor (n2607,n636,n2558);
and (n2608,n2598,n2607);
and (n2609,n2583,n2596);
xor (n2610,n2611,n2565);
xor (n2611,n2548,n2550);
and (n2612,n2610,n2613);
or (n2613,n2614,n2628,n2631);
and (n2614,n2615,n2617);
xor (n2615,n2616,n2557);
xor (n2616,n2552,n2554);
or (n2617,n2618,n2626,n2627);
and (n2618,n2619,n2621);
xor (n2619,n2620,n753);
xor (n2620,n2585,n2589);
or (n2621,n2622,n2623,n2625);
not (n2622,n1185);
and (n2623,n1158,n2624);
not (n2624,n1152);
and (n2625,n1154,n2624);
and (n2626,n2621,n1187);
and (n2627,n2619,n1187);
and (n2628,n2617,n2629);
xor (n2629,n2630,n2596);
xor (n2630,n2583,n2593);
and (n2631,n2615,n2629);
and (n2632,n2581,n2613);
and (n2633,n2579,n2634);
or (n2634,n2635,n2637);
xor (n2635,n2636,n2613);
xor (n2636,n2581,n2610);
or (n2637,n2638,n2654,n2660);
and (n2638,n2639,n2652);
or (n2639,n2640,n2648,n2651);
and (n2640,n2641,n2643);
xor (n2641,n2642,n2607);
xor (n2642,n2598,n2604);
or (n2643,n2644,n2646,n2647);
and (n2644,n2645,n1172);
not (n2645,n1150);
not (n2646,n1179);
and (n2647,n2645,n1162);
and (n2648,n2643,n2649);
xor (n2649,n2650,n1187);
xor (n2650,n2619,n2621);
and (n2651,n2641,n2649);
xor (n2652,n2653,n2629);
xor (n2653,n2615,n2617);
and (n2654,n2652,n2655);
or (n2655,n2656,n2658);
or (n2656,n854,n2657);
not (n2657,n1148);
xor (n2658,n2659,n2649);
xor (n2659,n2641,n2643);
and (n2660,n2639,n2655);
and (n2661,n2577,n2634);
and (n2662,n2542,n2575);
and (n2663,n2465,n2540);
and (n2664,n2665,n2667);
xor (n2665,n2666,n2540);
xor (n2666,n2465,n2537);
or (n2667,n2668,n2670);
xor (n2668,n2669,n2575);
xor (n2669,n2542,n2572);
and (n2670,n2671,n2672);
not (n2671,n2668);
and (n2672,n2673,n2675);
xor (n2673,n2674,n2634);
xor (n2674,n2577,n2579);
and (n2675,n2676,n2677);
xnor (n2676,n2635,n2637);
and (n2677,n2678,n2680);
xor (n2678,n2679,n2655);
xor (n2679,n2639,n2652);
and (n2680,n2681,n2682);
xnor (n2681,n2656,n2658);
and (n2682,n2683,n1232);
not (n2683,n2684);
nand (n2684,n2685,n853);
not (n2685,n2245);
endmodule
