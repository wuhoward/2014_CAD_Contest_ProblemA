module top (out,n23,n28,n29,n30,n32,n33,n44,n47,n50
        ,n53,n56,n59,n62,n65,n68,n70,n73,n84,n94
        ,n99,n102,n105,n108,n111,n114,n117,n120,n123,n126
        ,n129,n131,n133,n141,n155,n160,n193,n198,n201,n204
        ,n207,n220,n265,n276,n288,n293,n296,n299,n302,n305
        ,n308,n324,n397,n407,n440,n445,n448,n635);
output out;
input n23;
input n28;
input n29;
input n30;
input n32;
input n33;
input n44;
input n47;
input n50;
input n53;
input n56;
input n59;
input n62;
input n65;
input n68;
input n70;
input n73;
input n84;
input n94;
input n99;
input n102;
input n105;
input n108;
input n111;
input n114;
input n117;
input n120;
input n123;
input n126;
input n129;
input n131;
input n133;
input n141;
input n155;
input n160;
input n193;
input n198;
input n201;
input n204;
input n207;
input n220;
input n265;
input n276;
input n288;
input n293;
input n296;
input n299;
input n302;
input n305;
input n308;
input n324;
input n397;
input n407;
input n440;
input n445;
input n448;
input n635;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n31;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n63;
wire n64;
wire n66;
wire n67;
wire n69;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n103;
wire n104;
wire n106;
wire n107;
wire n109;
wire n110;
wire n112;
wire n113;
wire n115;
wire n116;
wire n118;
wire n119;
wire n121;
wire n122;
wire n124;
wire n125;
wire n127;
wire n128;
wire n130;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n194;
wire n195;
wire n196;
wire n197;
wire n199;
wire n200;
wire n202;
wire n203;
wire n205;
wire n206;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n289;
wire n290;
wire n291;
wire n292;
wire n294;
wire n295;
wire n297;
wire n298;
wire n300;
wire n301;
wire n303;
wire n304;
wire n306;
wire n307;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n441;
wire n442;
wire n443;
wire n444;
wire n446;
wire n447;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
xor (out,n0,n2220);
nand (n0,n1,n2219);
or (n1,n2,n1076);
not (n2,n3);
nor (n3,n4,n1075);
not (n4,n5);
nand (n5,n6,n1008);
xor (n6,n7,n880);
xor (n7,n8,n657);
xor (n8,n9,n599);
xor (n9,n10,n430);
or (n10,n11,n429);
and (n11,n12,n367);
xor (n12,n13,n241);
xor (n13,n14,n186);
xor (n14,n15,n147);
nand (n15,n16,n136);
or (n16,n17,n90);
nand (n17,n18,n80);
or (n18,n19,n77);
and (n19,n20,n74);
wire s0n20,s1n20,notn20;
or (n20,s0n20,s1n20);
not(notn20,n71);
and (s0n20,notn20,n21);
and (s1n20,n71,n40);
wire s0n21,s1n21,notn21;
or (n21,s0n21,s1n21);
not(notn21,n24);
and (s0n21,notn21,1'b0);
and (s1n21,n24,n23);
or (n24,n25,n36);
or (n25,n26,n34);
nor (n26,n27,n29,n30,n31,n33);
not (n27,n28);
not (n31,n32);
nor (n34,n28,n35,n30,n31,n33);
not (n35,n29);
or (n36,n37,n39);
and (n37,n27,n29,n30,n31,n38);
not (n38,n33);
nor (n39,n27,n35,n30,n31,n33);
xor (n40,n41,n42);
not (n41,n23);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n57);
not (n55,n56);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n66);
not (n64,n65);
and (n66,n67,n69);
not (n67,n68);
not (n69,n70);
and (n71,n72,n73);
or (n72,n26,n37);
wire s0n74,s1n74,notn74;
or (n74,s0n74,s1n74);
not(notn74,n71);
and (s0n74,notn74,n75);
and (s1n74,n71,n76);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n24);
and (s0n75,notn75,1'b0);
and (s1n75,n24,n44);
xor (n76,n43,n45);
and (n77,n78,n79);
not (n78,n20);
not (n79,n74);
nand (n80,n81,n88);
or (n81,n78,n82);
wire s0n82,s1n82,notn82;
or (n82,s0n82,s1n82);
not(notn82,n71);
and (s0n82,notn82,n83);
and (s1n82,n71,n85);
wire s0n83,s1n83,notn83;
or (n83,s0n83,s1n83);
not(notn83,n24);
and (s0n83,notn83,1'b0);
and (s1n83,n24,n84);
xor (n85,n86,n87);
not (n86,n84);
and (n87,n41,n42);
or (n88,n89,n20);
not (n89,n82);
nor (n90,n91,n134);
and (n91,n89,n92);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n132);
and (s0n92,notn92,n93);
and (s1n92,n132,n95);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n24);
and (s0n93,notn93,1'b0);
and (s1n93,n24,n94);
xor (n95,n96,n97);
not (n96,n94);
and (n97,n98,n100);
not (n98,n99);
and (n100,n101,n103);
not (n101,n102);
and (n103,n104,n106);
not (n104,n105);
and (n106,n107,n109);
not (n107,n108);
and (n109,n110,n112);
not (n110,n111);
and (n112,n113,n115);
not (n113,n114);
and (n115,n116,n118);
not (n116,n117);
and (n118,n119,n121);
not (n119,n120);
and (n121,n122,n124);
not (n122,n123);
and (n124,n125,n127);
not (n125,n126);
and (n127,n128,n130);
not (n128,n129);
not (n130,n131);
and (n132,n72,n133);
and (n134,n82,n135);
not (n135,n92);
or (n136,n18,n137);
nor (n137,n138,n145);
and (n138,n89,n139);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n132);
and (s0n139,notn139,n140);
and (s1n139,n132,n142);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n24);
and (s0n140,notn140,1'b0);
and (s1n140,n24,n141);
xor (n142,n143,n144);
not (n143,n141);
and (n144,n96,n97);
and (n145,n82,n146);
not (n146,n139);
nand (n147,n148,n177);
or (n148,n149,n170);
or (n149,n150,n167);
nor (n150,n151,n165);
and (n151,n152,n162);
not (n152,n153);
wire s0n153,s1n153,notn153;
or (n153,s0n153,s1n153);
not(notn153,n71);
and (s0n153,notn153,n154);
and (s1n153,n71,n156);
wire s0n154,s1n154,notn154;
or (n154,s0n154,s1n154);
not(notn154,n24);
and (s0n154,notn154,1'b0);
and (s1n154,n24,n155);
xor (n156,n157,n158);
not (n157,n155);
and (n158,n159,n161);
not (n159,n160);
and (n161,n86,n87);
wire s0n162,s1n162,notn162;
or (n162,s0n162,s1n162);
not(notn162,n71);
and (s0n162,notn162,n163);
and (s1n162,n71,n164);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n24);
and (s0n163,notn163,1'b0);
and (s1n163,n24,n160);
xor (n164,n159,n161);
and (n165,n166,n153);
not (n166,n162);
nor (n167,n168,n169);
and (n168,n162,n82);
and (n169,n166,n89);
nor (n170,n171,n175);
and (n171,n152,n172);
wire s0n172,s1n172,notn172;
or (n172,s0n172,s1n172);
not(notn172,n132);
and (s0n172,notn172,n173);
and (s1n172,n132,n174);
wire s0n173,s1n173,notn173;
or (n173,s0n173,s1n173);
not(notn173,n24);
and (s0n173,notn173,1'b0);
and (s1n173,n24,n102);
xor (n174,n101,n103);
and (n175,n153,n176);
not (n176,n172);
or (n177,n178,n179);
not (n178,n167);
nor (n179,n180,n184);
and (n180,n152,n181);
wire s0n181,s1n181,notn181;
or (n181,s0n181,s1n181);
not(notn181,n132);
and (s0n181,notn181,n182);
and (s1n181,n132,n183);
wire s0n182,s1n182,notn182;
or (n182,s0n182,s1n182);
not(notn182,n24);
and (s0n182,notn182,1'b0);
and (s1n182,n24,n99);
xor (n183,n98,n100);
and (n184,n153,n185);
not (n185,n181);
nand (n186,n187,n232);
or (n187,n188,n225);
or (n188,n189,n215);
nor (n189,n190,n212);
and (n190,n191,n209);
wire s0n191,s1n191,notn191;
or (n191,s0n191,s1n191);
not(notn191,n71);
and (s0n191,notn191,n192);
and (s1n191,n71,n194);
wire s0n192,s1n192,notn192;
or (n192,s0n192,s1n192);
not(notn192,n24);
and (s0n192,notn192,1'b0);
and (s1n192,n24,n193);
xor (n194,n195,n196);
not (n195,n193);
and (n196,n197,n199);
not (n197,n198);
and (n199,n200,n202);
not (n200,n201);
and (n202,n203,n205);
not (n203,n204);
and (n205,n206,n208);
not (n206,n207);
and (n208,n157,n158);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n71);
and (s0n209,notn209,n210);
and (s1n209,n71,n211);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n24);
and (s0n210,notn210,1'b0);
and (s1n210,n24,n198);
xor (n211,n197,n199);
and (n212,n213,n214);
not (n213,n191);
not (n214,n209);
nor (n215,n216,n224);
and (n216,n191,n217);
not (n217,n218);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n71);
and (s0n218,notn218,n219);
and (s1n218,n71,n221);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n24);
and (s0n219,notn219,1'b0);
and (s1n219,n24,n220);
xor (n221,n222,n223);
not (n222,n220);
and (n223,n195,n196);
and (n224,n213,n218);
nor (n225,n226,n230);
and (n226,n217,n227);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n132);
and (s0n227,notn227,n228);
and (s1n227,n132,n229);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n24);
and (s0n228,notn228,1'b0);
and (s1n228,n24,n120);
xor (n229,n119,n121);
and (n230,n218,n231);
not (n231,n227);
or (n232,n233,n234);
not (n233,n189);
nor (n234,n235,n239);
and (n235,n236,n217);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n132);
and (s0n236,notn236,n237);
and (s1n236,n132,n238);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n24);
and (s0n237,notn237,1'b0);
and (s1n237,n24,n117);
xor (n238,n116,n118);
and (n239,n240,n218);
not (n240,n236);
xor (n241,n242,n330);
xor (n242,n243,n282);
nand (n243,n244,n271);
or (n244,n245,n261);
nand (n245,n246,n253);
nor (n246,n247,n251);
and (n247,n248,n74);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n71);
and (s0n248,notn248,n249);
and (s1n248,n71,n250);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n24);
and (s0n249,notn249,1'b0);
and (s1n249,n24,n47);
xor (n250,n46,n48);
and (n251,n252,n79);
not (n252,n248);
not (n253,n254);
nor (n254,n255,n259);
and (n255,n256,n248);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n71);
and (s0n256,notn256,n257);
and (s1n256,n71,n258);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n24);
and (s0n257,notn257,1'b0);
and (s1n257,n24,n50);
xor (n258,n49,n51);
and (n259,n260,n252);
not (n260,n256);
nor (n261,n262,n269);
and (n262,n79,n263);
wire s0n263,s1n263,notn263;
or (n263,s0n263,s1n263);
not(notn263,n132);
and (s0n263,notn263,n264);
and (s1n263,n132,n266);
wire s0n264,s1n264,notn264;
or (n264,s0n264,s1n264);
not(notn264,n24);
and (s0n264,notn264,1'b0);
and (s1n264,n24,n265);
xor (n266,n267,n268);
not (n267,n265);
and (n268,n143,n144);
and (n269,n74,n270);
not (n270,n263);
or (n271,n272,n253);
nor (n272,n273,n280);
and (n273,n79,n274);
wire s0n274,s1n274,notn274;
or (n274,s0n274,s1n274);
not(notn274,n132);
and (s0n274,notn274,n275);
and (s1n274,n132,n277);
wire s0n275,s1n275,notn275;
or (n275,s0n275,s1n275);
not(notn275,n24);
and (s0n275,notn275,1'b0);
and (s1n275,n24,n276);
xor (n277,n278,n279);
not (n278,n276);
and (n279,n267,n268);
and (n280,n74,n281);
not (n281,n274);
nand (n282,n283,n319);
or (n283,n284,n316);
nor (n284,n285,n314);
and (n285,n286,n310);
wire s0n286,s1n286,notn286;
or (n286,s0n286,s1n286);
not(notn286,n132);
and (s0n286,notn286,n287);
and (s1n286,n132,n289);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n24);
and (s0n287,notn287,1'b0);
and (s1n287,n24,n288);
xor (n289,n290,n291);
not (n290,n288);
and (n291,n292,n294);
not (n292,n293);
and (n294,n295,n297);
not (n295,n296);
and (n297,n298,n300);
not (n298,n299);
and (n300,n301,n303);
not (n301,n302);
and (n303,n304,n306);
not (n304,n305);
and (n306,n307,n309);
not (n307,n308);
and (n309,n278,n279);
not (n310,n311);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n71);
and (s0n311,notn311,n312);
and (s1n311,n71,n313);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n24);
and (s0n312,notn312,1'b0);
and (s1n312,n24,n68);
xor (n313,n67,n69);
and (n314,n315,n311);
not (n315,n286);
nand (n316,n311,n317);
not (n317,n318);
wire s0n318,s1n318,notn318;
or (n318,s0n318,s1n318);
not(notn318,n24);
and (s0n318,notn318,1'b0);
and (s1n318,n24,n70);
or (n319,n320,n317);
nor (n320,n321,n328);
and (n321,n322,n310);
wire s0n322,s1n322,notn322;
or (n322,s0n322,s1n322);
not(notn322,n132);
and (s0n322,notn322,n323);
and (s1n322,n132,n325);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n24);
and (s0n323,notn323,1'b0);
and (s1n323,n24,n324);
xor (n325,n326,n327);
not (n326,n324);
and (n327,n290,n291);
and (n328,n329,n311);
not (n329,n322);
nand (n330,n331,n359);
or (n331,n332,n352);
nand (n332,n333,n344);
not (n333,n334);
nand (n334,n335,n343);
or (n335,n336,n340);
not (n336,n337);
wire s0n337,s1n337,notn337;
or (n337,s0n337,s1n337);
not(notn337,n71);
and (s0n337,notn337,n338);
and (s1n337,n71,n339);
wire s0n338,s1n338,notn338;
or (n338,s0n338,s1n338);
not(notn338,n24);
and (s0n338,notn338,1'b0);
and (s1n338,n24,n62);
xor (n339,n61,n63);
wire s0n340,s1n340,notn340;
or (n340,s0n340,s1n340);
not(notn340,n71);
and (s0n340,notn340,n341);
and (s1n340,n71,n342);
wire s0n341,s1n341,notn341;
or (n341,s0n341,s1n341);
not(notn341,n24);
and (s0n341,notn341,1'b0);
and (s1n341,n24,n59);
xor (n342,n58,n60);
nand (n343,n340,n336);
nor (n344,n345,n351);
and (n345,n346,n350);
not (n346,n347);
wire s0n347,s1n347,notn347;
or (n347,s0n347,s1n347);
not(notn347,n71);
and (s0n347,notn347,n348);
and (s1n347,n71,n349);
wire s0n348,s1n348,notn348;
or (n348,s0n348,s1n348);
not(notn348,n24);
and (s0n348,notn348,1'b0);
and (s1n348,n24,n56);
xor (n349,n55,n57);
not (n350,n340);
and (n351,n347,n340);
nor (n352,n353,n357);
and (n353,n354,n346);
wire s0n354,s1n354,notn354;
or (n354,s0n354,s1n354);
not(notn354,n132);
and (s0n354,notn354,n355);
and (s1n354,n132,n356);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n24);
and (s0n355,notn355,1'b0);
and (s1n355,n24,n302);
xor (n356,n301,n303);
and (n357,n358,n347);
not (n358,n354);
or (n359,n360,n333);
nor (n360,n361,n365);
and (n361,n362,n346);
wire s0n362,s1n362,notn362;
or (n362,s0n362,s1n362);
not(notn362,n132);
and (s0n362,notn362,n363);
and (s1n362,n132,n364);
wire s0n363,s1n363,notn363;
or (n363,s0n363,s1n363);
not(notn363,n24);
and (s0n363,notn363,1'b0);
and (s1n363,n24,n299);
xor (n364,n298,n300);
and (n365,n366,n347);
not (n366,n362);
or (n367,n368,n428);
and (n368,n369,n390);
xor (n369,n370,n380);
nand (n370,n371,n379);
or (n371,n149,n372);
nor (n372,n373,n377);
and (n373,n152,n374);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n132);
and (s0n374,notn374,n375);
and (s1n374,n132,n376);
wire s0n375,s1n375,notn375;
or (n375,s0n375,s1n375);
not(notn375,n24);
and (s0n375,notn375,1'b0);
and (s1n375,n24,n105);
xor (n376,n104,n106);
and (n377,n153,n378);
not (n378,n374);
or (n379,n178,n170);
nand (n380,n381,n389);
or (n381,n188,n382);
nor (n382,n383,n387);
and (n383,n384,n217);
wire s0n384,s1n384,notn384;
or (n384,s0n384,s1n384);
not(notn384,n132);
and (s0n384,notn384,n385);
and (s1n384,n132,n386);
wire s0n385,s1n385,notn385;
or (n385,s0n385,s1n385);
not(notn385,n24);
and (s0n385,notn385,1'b0);
and (s1n385,n24,n123);
xor (n386,n122,n124);
and (n387,n388,n218);
not (n388,n384);
or (n389,n233,n225);
nand (n390,n391,n420);
or (n391,n392,n413);
nand (n392,n393,n403);
nor (n393,n394,n401);
and (n394,n217,n395);
wire s0n395,s1n395,notn395;
or (n395,s0n395,s1n395);
not(notn395,n71);
and (s0n395,notn395,n396);
and (s1n395,n71,n398);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n24);
and (s0n396,notn396,1'b0);
and (s1n396,n24,n397);
xor (n398,n399,n400);
not (n399,n397);
and (n400,n222,n223);
and (n401,n218,n402);
not (n402,n395);
nand (n403,n404,n411);
or (n404,n402,n405);
wire s0n405,s1n405,notn405;
or (n405,s0n405,s1n405);
not(notn405,n71);
and (s0n405,notn405,n406);
and (s1n405,n71,n408);
wire s0n406,s1n406,notn406;
or (n406,s0n406,s1n406);
not(notn406,n24);
and (s0n406,notn406,1'b0);
and (s1n406,n24,n407);
xor (n408,n409,n410);
not (n409,n407);
and (n410,n399,n400);
or (n411,n395,n412);
not (n412,n405);
nor (n413,n414,n418);
and (n414,n415,n412);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n132);
and (s0n415,notn415,n416);
and (s1n415,n132,n417);
wire s0n416,s1n416,notn416;
or (n416,s0n416,s1n416);
not(notn416,n24);
and (s0n416,notn416,1'b0);
and (s1n416,n24,n129);
xor (n417,n128,n130);
and (n418,n419,n405);
not (n419,n415);
or (n420,n393,n421);
nor (n421,n422,n426);
and (n422,n423,n412);
wire s0n423,s1n423,notn423;
or (n423,s0n423,s1n423);
not(notn423,n132);
and (s0n423,notn423,n424);
and (s1n423,n132,n425);
wire s0n424,s1n424,notn424;
or (n424,s0n424,s1n424);
not(notn424,n24);
and (s0n424,notn424,1'b0);
and (s1n424,n24,n126);
xor (n425,n125,n127);
and (n426,n427,n405);
not (n427,n423);
and (n428,n370,n380);
and (n429,n13,n241);
xor (n430,n431,n572);
xor (n431,n432,n505);
xor (n432,n433,n481);
xor (n433,n434,n457);
nor (n434,n435,n455);
and (n435,n436,n453);
nand (n436,n437,n450);
not (n437,n438);
wire s0n438,s1n438,notn438;
or (n438,s0n438,s1n438);
not(notn438,n71);
and (s0n438,notn438,n439);
and (s1n438,n71,n441);
wire s0n439,s1n439,notn439;
or (n439,s0n439,s1n439);
not(notn439,n24);
and (s0n439,notn439,1'b0);
and (s1n439,n24,n440);
xor (n441,n442,n443);
not (n442,n440);
and (n443,n444,n446);
not (n444,n445);
and (n446,n447,n449);
not (n447,n448);
and (n449,n409,n410);
wire s0n450,s1n450,notn450;
or (n450,s0n450,s1n450);
not(notn450,n71);
and (s0n450,notn450,n451);
and (s1n450,n71,n452);
wire s0n451,s1n451,notn451;
or (n451,s0n451,s1n451);
not(notn451,n24);
and (s0n451,notn451,1'b0);
and (s1n451,n24,n445);
xor (n452,n444,n446);
nand (n453,n438,n454);
not (n454,n450);
not (n455,n456);
wire s0n456,s1n456,notn456;
or (n456,s0n456,s1n456);
not(notn456,n24);
and (s0n456,notn456,1'b0);
and (s1n456,n24,n131);
nand (n457,n458,n477);
or (n458,n459,n470);
nand (n459,n460,n467);
nor (n460,n461,n465);
and (n461,n310,n462);
wire s0n462,s1n462,notn462;
or (n462,s0n462,s1n462);
not(notn462,n71);
and (s0n462,notn462,n463);
and (s1n462,n71,n464);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n24);
and (s0n463,notn463,1'b0);
and (s1n463,n24,n65);
xor (n464,n64,n66);
and (n465,n311,n466);
not (n466,n462);
nand (n467,n468,n469);
or (n468,n336,n462);
nand (n469,n336,n462);
nor (n470,n471,n475);
and (n471,n472,n336);
wire s0n472,s1n472,notn472;
or (n472,s0n472,s1n472);
not(notn472,n132);
and (s0n472,notn472,n473);
and (s1n472,n132,n474);
wire s0n473,s1n473,notn473;
or (n473,s0n473,s1n473);
not(notn473,n24);
and (s0n473,notn473,1'b0);
and (s1n473,n24,n293);
xor (n474,n292,n294);
and (n475,n476,n337);
not (n476,n472);
or (n477,n460,n478);
nor (n478,n479,n480);
and (n479,n286,n336);
and (n480,n315,n337);
nand (n481,n482,n501);
or (n482,n483,n494);
nand (n483,n484,n491);
or (n484,n485,n489);
and (n485,n347,n486);
wire s0n486,s1n486,notn486;
or (n486,s0n486,s1n486);
not(notn486,n71);
and (s0n486,notn486,n487);
and (s1n486,n71,n488);
wire s0n487,s1n487,notn487;
or (n487,s0n487,s1n487);
not(notn487,n24);
and (s0n487,notn487,1'b0);
and (s1n487,n24,n53);
xor (n488,n52,n54);
and (n489,n346,n490);
not (n490,n486);
nor (n491,n492,n493);
and (n492,n256,n486);
and (n493,n260,n490);
nor (n494,n495,n499);
and (n495,n496,n260);
wire s0n496,s1n496,notn496;
or (n496,s0n496,s1n496);
not(notn496,n132);
and (s0n496,notn496,n497);
and (s1n496,n132,n498);
wire s0n497,s1n497,notn497;
or (n497,s0n497,s1n497);
not(notn497,n24);
and (s0n497,notn497,1'b0);
and (s1n497,n24,n305);
xor (n498,n304,n306);
and (n499,n500,n256);
not (n500,n496);
or (n501,n502,n484);
nor (n502,n503,n504);
and (n503,n354,n260);
and (n504,n358,n256);
xor (n505,n506,n562);
xor (n506,n507,n533);
nand (n507,n508,n528);
or (n508,n509,n525);
not (n509,n510);
nor (n510,n511,n517);
nand (n511,n512,n516);
or (n512,n152,n513);
wire s0n513,s1n513,notn513;
or (n513,s0n513,s1n513);
not(notn513,n71);
and (s0n513,notn513,n514);
and (s1n513,n71,n515);
wire s0n514,s1n514,notn514;
or (n514,s0n514,s1n514);
not(notn514,n24);
and (s0n514,notn514,1'b0);
and (s1n514,n24,n207);
xor (n515,n206,n208);
nand (n516,n152,n513);
nor (n517,n518,n523);
and (n518,n519,n513);
not (n519,n520);
wire s0n520,s1n520,notn520;
or (n520,s0n520,s1n520);
not(notn520,n71);
and (s0n520,notn520,n521);
and (s1n520,n71,n522);
wire s0n521,s1n521,notn521;
or (n521,s0n521,s1n521);
not(notn521,n24);
and (s0n521,notn521,1'b0);
and (s1n521,n24,n204);
xor (n522,n203,n205);
and (n523,n524,n520);
not (n524,n513);
nor (n525,n526,n527);
and (n526,n519,n374);
and (n527,n520,n378);
or (n528,n529,n530);
not (n529,n511);
nor (n530,n531,n532);
and (n531,n519,n172);
and (n532,n520,n176);
nand (n533,n534,n554);
or (n534,n535,n547);
not (n535,n536);
and (n536,n537,n544);
nor (n537,n538,n543);
and (n538,n520,n539);
not (n539,n540);
wire s0n540,s1n540,notn540;
or (n540,s0n540,s1n540);
not(notn540,n71);
and (s0n540,notn540,n541);
and (s1n540,n71,n542);
wire s0n541,s1n541,notn541;
or (n541,s0n541,s1n541);
not(notn541,n24);
and (s0n541,notn541,1'b0);
and (s1n541,n24,n201);
xor (n542,n200,n202);
and (n543,n519,n540);
nand (n544,n545,n546);
or (n545,n539,n209);
or (n546,n214,n540);
nor (n547,n548,n552);
and (n548,n214,n549);
wire s0n549,s1n549,notn549;
or (n549,s0n549,s1n549);
not(notn549,n132);
and (s0n549,notn549,n550);
and (s1n549,n132,n551);
wire s0n550,s1n550,notn550;
or (n550,s0n550,s1n550);
not(notn550,n24);
and (s0n550,notn550,1'b0);
and (s1n550,n24,n111);
xor (n551,n110,n112);
and (n552,n209,n553);
not (n553,n549);
or (n554,n555,n537);
nor (n555,n556,n560);
and (n556,n214,n557);
wire s0n557,s1n557,notn557;
or (n557,s0n557,s1n557);
not(notn557,n132);
and (s0n557,notn557,n558);
and (s1n557,n132,n559);
wire s0n558,s1n558,notn558;
or (n558,s0n558,s1n558);
not(notn558,n24);
and (s0n558,notn558,1'b0);
and (s1n558,n24,n108);
xor (n559,n107,n109);
and (n560,n209,n561);
not (n561,n557);
nand (n562,n563,n564);
or (n563,n245,n272);
or (n564,n565,n253);
nor (n565,n566,n570);
and (n566,n79,n567);
wire s0n567,s1n567,notn567;
or (n567,s0n567,s1n567);
not(notn567,n132);
and (s0n567,notn567,n568);
and (s1n567,n132,n569);
wire s0n568,s1n568,notn568;
or (n568,s0n568,s1n568);
not(notn568,n24);
and (s0n568,notn568,1'b0);
and (s1n568,n24,n308);
xor (n569,n307,n309);
and (n570,n74,n571);
not (n571,n567);
xor (n572,n573,n590);
xor (n573,n574,n580);
nand (n574,n575,n576);
or (n575,n149,n179);
or (n576,n178,n577);
nor (n577,n578,n579);
and (n578,n152,n92);
and (n579,n153,n135);
nand (n580,n581,n582);
or (n581,n188,n234);
or (n582,n233,n583);
nor (n583,n584,n588);
and (n584,n217,n585);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n132);
and (s0n585,notn585,n586);
and (s1n585,n132,n587);
wire s0n586,s1n586,notn586;
or (n586,s0n586,s1n586);
not(notn586,n24);
and (s0n586,notn586,1'b0);
and (s1n586,n24,n114);
xor (n587,n113,n115);
and (n588,n218,n589);
not (n589,n585);
nand (n590,n591,n595);
or (n591,n392,n592);
nor (n592,n593,n594);
and (n593,n384,n412);
and (n594,n388,n405);
or (n595,n393,n596);
nor (n596,n597,n598);
and (n597,n412,n227);
and (n598,n405,n231);
xor (n599,n600,n626);
xor (n600,n601,n623);
or (n601,n602,n622);
and (n602,n603,n616);
xor (n603,n604,n610);
nand (n604,n605,n609);
or (n605,n483,n606);
nor (n606,n607,n608);
and (n607,n567,n260);
and (n608,n571,n256);
or (n609,n494,n484);
nand (n610,n611,n615);
or (n611,n509,n612);
nor (n612,n613,n614);
and (n613,n519,n557);
and (n614,n520,n561);
or (n615,n529,n525);
nand (n616,n617,n621);
or (n617,n535,n618);
nor (n618,n619,n620);
and (n619,n214,n585);
and (n620,n209,n589);
or (n621,n547,n537);
and (n622,n604,n610);
or (n623,n624,n625);
and (n624,n14,n186);
and (n625,n15,n147);
xor (n626,n627,n651);
xor (n627,n628,n641);
nand (n628,n629,n630);
or (n629,n320,n316);
or (n630,n631,n317);
nor (n631,n632,n639);
and (n632,n633,n310);
wire s0n633,s1n633,notn633;
or (n633,s0n633,s1n633);
not(notn633,n132);
and (s0n633,notn633,n634);
and (s1n633,n132,n636);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n24);
and (s0n634,notn634,1'b0);
and (s1n634,n24,n635);
xor (n636,n637,n638);
not (n637,n635);
and (n638,n326,n327);
and (n639,n640,n311);
not (n640,n633);
nand (n641,n642,n643);
or (n642,n332,n360);
or (n643,n333,n644);
nor (n644,n645,n649);
and (n645,n646,n346);
wire s0n646,s1n646,notn646;
or (n646,s0n646,s1n646);
not(notn646,n132);
and (s0n646,notn646,n647);
and (s1n646,n132,n648);
wire s0n647,s1n647,notn647;
or (n647,s0n647,s1n647);
not(notn647,n24);
and (s0n647,notn647,1'b0);
and (s1n647,n24,n296);
xor (n648,n295,n297);
and (n649,n650,n347);
not (n650,n646);
nand (n651,n652,n653);
or (n652,n17,n137);
or (n653,n18,n654);
nor (n654,n655,n656);
and (n655,n89,n263);
and (n656,n82,n270);
xor (n657,n658,n846);
xor (n658,n659,n785);
or (n659,n660,n784);
and (n660,n661,n702);
xor (n661,n662,n663);
xor (n662,n603,n616);
xor (n663,n664,n689);
xor (n664,n665,n668);
nand (n665,n666,n667);
or (n666,n392,n421);
or (n667,n393,n592);
nand (n668,n669,n685);
or (n669,n670,n682);
or (n670,n671,n679);
not (n671,n672);
and (n672,n673,n678);
nand (n673,n674,n405);
not (n674,n675);
wire s0n675,s1n675,notn675;
or (n675,s0n675,s1n675);
not(notn675,n71);
and (s0n675,notn675,n676);
and (s1n675,n71,n677);
wire s0n676,s1n676,notn676;
or (n676,s0n676,s1n676);
not(notn676,n24);
and (s0n676,notn676,1'b0);
and (s1n676,n24,n448);
xor (n677,n447,n449);
nand (n678,n675,n412);
nor (n679,n680,n681);
and (n680,n675,n454);
and (n681,n674,n450);
nor (n682,n683,n684);
and (n683,n450,n455);
and (n684,n454,n456);
or (n685,n672,n686);
nor (n686,n687,n688);
and (n687,n415,n454);
and (n688,n419,n450);
xor (n689,n690,n696);
nor (n690,n691,n454);
nor (n691,n692,n695);
and (n692,n693,n412);
not (n693,n694);
and (n694,n456,n675);
and (n695,n674,n455);
nand (n696,n697,n701);
or (n697,n459,n698);
nor (n698,n699,n700);
and (n699,n646,n336);
and (n700,n650,n337);
or (n701,n470,n460);
or (n702,n703,n783);
and (n703,n704,n752);
xor (n704,n705,n721);
and (n705,n706,n712);
nor (n706,n707,n412);
nor (n707,n708,n711);
and (n708,n709,n217);
not (n709,n710);
and (n710,n456,n395);
and (n711,n402,n455);
nand (n712,n713,n717);
or (n713,n459,n714);
nor (n714,n715,n716);
and (n715,n354,n336);
and (n716,n358,n337);
or (n717,n460,n718);
nor (n718,n719,n720);
and (n719,n362,n336);
and (n720,n366,n337);
or (n721,n722,n751);
and (n722,n723,n742);
xor (n723,n724,n733);
nand (n724,n725,n729);
or (n725,n245,n726);
nor (n726,n727,n728);
and (n727,n79,n92);
and (n728,n74,n135);
or (n729,n730,n253);
nor (n730,n731,n732);
and (n731,n79,n139);
and (n732,n74,n146);
nand (n733,n734,n738);
or (n734,n735,n316);
nor (n735,n736,n737);
and (n736,n646,n310);
and (n737,n650,n311);
or (n738,n739,n317);
nor (n739,n740,n741);
and (n740,n472,n310);
and (n741,n476,n311);
nand (n742,n743,n747);
or (n743,n332,n744);
nor (n744,n745,n746);
and (n745,n567,n346);
and (n746,n571,n347);
or (n747,n748,n333);
nor (n748,n749,n750);
and (n749,n496,n346);
and (n750,n500,n347);
and (n751,n724,n733);
or (n752,n753,n782);
and (n753,n754,n773);
xor (n754,n755,n764);
nand (n755,n756,n760);
or (n756,n483,n757);
nor (n757,n758,n759);
and (n758,n263,n260);
and (n759,n270,n256);
or (n760,n484,n761);
nor (n761,n762,n763);
and (n762,n274,n260);
and (n763,n281,n256);
nand (n764,n765,n769);
or (n765,n509,n766);
nor (n766,n767,n768);
and (n767,n519,n585);
and (n768,n520,n589);
or (n769,n770,n529);
nor (n770,n771,n772);
and (n771,n519,n549);
and (n772,n520,n553);
nand (n773,n774,n778);
or (n774,n535,n775);
nor (n775,n776,n777);
and (n776,n214,n227);
and (n777,n209,n231);
or (n778,n779,n537);
nor (n779,n780,n781);
and (n780,n214,n236);
and (n781,n209,n240);
and (n782,n755,n764);
and (n783,n705,n721);
and (n784,n662,n663);
xor (n785,n786,n802);
xor (n786,n787,n790);
or (n787,n788,n789);
and (n788,n664,n689);
and (n789,n665,n668);
xor (n790,n791,n799);
xor (n791,n792,n798);
nand (n792,n793,n794);
or (n793,n670,n686);
or (n794,n672,n795);
nor (n795,n796,n797);
and (n796,n423,n454);
and (n797,n427,n450);
and (n798,n690,n696);
or (n799,n800,n801);
and (n800,n242,n330);
and (n801,n243,n282);
or (n802,n803,n845);
and (n803,n804,n832);
xor (n804,n805,n821);
or (n805,n806,n820);
and (n806,n807,n814);
xor (n807,n808,n811);
nand (n808,n809,n810);
or (n809,n739,n316);
or (n810,n284,n317);
nand (n811,n812,n813);
or (n812,n332,n748);
or (n813,n352,n333);
nand (n814,n815,n819);
or (n815,n17,n816);
nor (n816,n817,n818);
and (n817,n89,n181);
and (n818,n82,n185);
or (n819,n18,n90);
and (n820,n808,n811);
or (n821,n822,n831);
and (n822,n823,n828);
xor (n823,n824,n825);
nor (n824,n672,n455);
nand (n825,n826,n827);
or (n826,n459,n718);
or (n827,n460,n698);
nand (n828,n829,n830);
or (n829,n483,n761);
or (n830,n484,n606);
and (n831,n824,n825);
or (n832,n833,n844);
and (n833,n834,n841);
xor (n834,n835,n838);
nand (n835,n836,n837);
or (n836,n509,n770);
or (n837,n529,n612);
nand (n838,n839,n840);
or (n839,n535,n779);
or (n840,n618,n537);
nand (n841,n842,n843);
or (n842,n245,n730);
or (n843,n261,n253);
and (n844,n835,n838);
and (n845,n805,n821);
or (n846,n847,n879);
and (n847,n848,n878);
xor (n848,n849,n877);
or (n849,n850,n876);
and (n850,n851,n875);
xor (n851,n852,n874);
or (n852,n853,n873);
and (n853,n854,n867);
xor (n854,n855,n861);
nand (n855,n856,n860);
or (n856,n17,n857);
nor (n857,n858,n859);
and (n858,n89,n172);
and (n859,n82,n176);
or (n860,n18,n816);
nand (n861,n862,n866);
or (n862,n149,n863);
nor (n863,n864,n865);
and (n864,n152,n557);
and (n865,n153,n561);
or (n866,n178,n372);
nand (n867,n868,n872);
or (n868,n188,n869);
nor (n869,n870,n871);
and (n870,n423,n217);
and (n871,n427,n218);
or (n872,n233,n382);
and (n873,n855,n861);
xor (n874,n807,n814);
xor (n875,n834,n841);
and (n876,n852,n874);
xor (n877,n804,n832);
xor (n878,n12,n367);
and (n879,n849,n877);
or (n880,n881,n1007);
and (n881,n882,n923);
xor (n882,n883,n884);
xor (n883,n661,n702);
or (n884,n885,n922);
and (n885,n886,n889);
xor (n886,n887,n888);
xor (n887,n823,n828);
xor (n888,n369,n390);
or (n889,n890,n921);
and (n890,n891,n899);
xor (n891,n892,n898);
nand (n892,n893,n897);
or (n893,n392,n894);
nor (n894,n895,n896);
and (n895,n405,n455);
and (n896,n412,n456);
or (n897,n393,n413);
xor (n898,n706,n712);
or (n899,n900,n920);
and (n900,n901,n914);
xor (n901,n902,n908);
nand (n902,n903,n907);
or (n903,n245,n904);
nor (n904,n905,n906);
and (n905,n79,n181);
and (n906,n74,n185);
or (n907,n726,n253);
nand (n908,n909,n913);
or (n909,n332,n910);
nor (n910,n911,n912);
and (n911,n274,n346);
and (n912,n281,n347);
or (n913,n333,n744);
nand (n914,n915,n919);
or (n915,n17,n916);
nor (n916,n917,n918);
and (n917,n89,n374);
and (n918,n82,n378);
or (n919,n18,n857);
and (n920,n902,n908);
and (n921,n892,n898);
and (n922,n887,n888);
or (n923,n924,n1006);
and (n924,n925,n971);
xor (n925,n926,n927);
xor (n926,n704,n752);
or (n927,n928,n970);
and (n928,n929,n969);
xor (n929,n930,n947);
or (n930,n931,n946);
and (n931,n932,n940);
xor (n932,n933,n934);
nor (n933,n393,n455);
nand (n934,n935,n939);
or (n935,n936,n316);
nor (n936,n937,n938);
and (n937,n362,n310);
and (n938,n366,n311);
or (n939,n735,n317);
nand (n940,n941,n945);
or (n941,n483,n942);
nor (n942,n943,n944);
and (n943,n139,n260);
and (n944,n146,n256);
or (n945,n484,n757);
and (n946,n933,n934);
or (n947,n948,n968);
and (n948,n949,n962);
xor (n949,n950,n956);
nand (n950,n951,n955);
or (n951,n509,n952);
nor (n952,n953,n954);
and (n953,n236,n519);
and (n954,n240,n520);
or (n955,n766,n529);
nand (n956,n957,n961);
or (n957,n535,n958);
nor (n958,n959,n960);
and (n959,n384,n214);
and (n960,n388,n209);
or (n961,n775,n537);
nand (n962,n963,n967);
or (n963,n459,n964);
nor (n964,n965,n966);
and (n965,n496,n336);
and (n966,n500,n337);
or (n967,n460,n714);
and (n968,n950,n956);
xor (n969,n723,n742);
and (n970,n930,n947);
or (n971,n972,n1005);
and (n972,n973,n976);
xor (n973,n974,n975);
xor (n974,n754,n773);
xor (n975,n854,n867);
or (n976,n977,n1004);
and (n977,n978,n991);
xor (n978,n979,n985);
nand (n979,n980,n984);
or (n980,n149,n981);
nor (n981,n982,n983);
and (n982,n152,n549);
and (n983,n153,n553);
or (n984,n178,n863);
nand (n985,n986,n990);
or (n986,n188,n987);
nor (n987,n988,n989);
and (n988,n415,n217);
and (n989,n419,n218);
or (n990,n233,n869);
and (n991,n992,n998);
nor (n992,n993,n217);
nor (n993,n994,n997);
and (n994,n995,n214);
not (n995,n996);
and (n996,n456,n191);
and (n997,n213,n455);
nand (n998,n999,n1003);
or (n999,n1000,n316);
nor (n1000,n1001,n1002);
and (n1001,n354,n310);
and (n1002,n358,n311);
or (n1003,n936,n317);
and (n1004,n979,n985);
and (n1005,n974,n975);
and (n1006,n926,n927);
and (n1007,n883,n884);
or (n1008,n1009,n1074);
and (n1009,n1010,n1073);
xor (n1010,n1011,n1012);
xor (n1011,n848,n878);
or (n1012,n1013,n1072);
and (n1013,n1014,n1017);
xor (n1014,n1015,n1016);
xor (n1015,n851,n875);
xor (n1016,n886,n889);
or (n1017,n1018,n1071);
and (n1018,n1019,n1070);
xor (n1019,n1020,n1021);
xor (n1020,n891,n899);
or (n1021,n1022,n1069);
and (n1022,n1023,n1068);
xor (n1023,n1024,n1046);
or (n1024,n1025,n1045);
and (n1025,n1026,n1039);
xor (n1026,n1027,n1033);
nand (n1027,n1028,n1032);
or (n1028,n483,n1029);
nor (n1029,n1030,n1031);
and (n1030,n92,n260);
and (n1031,n135,n256);
or (n1032,n484,n942);
nand (n1033,n1034,n1038);
or (n1034,n509,n1035);
nor (n1035,n1036,n1037);
and (n1036,n519,n227);
and (n1037,n231,n520);
or (n1038,n529,n952);
nand (n1039,n1040,n1044);
or (n1040,n535,n1041);
nor (n1041,n1042,n1043);
and (n1042,n423,n214);
and (n1043,n427,n209);
or (n1044,n958,n537);
and (n1045,n1027,n1033);
or (n1046,n1047,n1067);
and (n1047,n1048,n1061);
xor (n1048,n1049,n1055);
nand (n1049,n1050,n1054);
or (n1050,n459,n1051);
nor (n1051,n1052,n1053);
and (n1052,n336,n567);
and (n1053,n571,n337);
or (n1054,n964,n460);
nand (n1055,n1056,n1060);
or (n1056,n245,n1057);
nor (n1057,n1058,n1059);
and (n1058,n79,n172);
and (n1059,n74,n176);
or (n1060,n904,n253);
nand (n1061,n1062,n1066);
or (n1062,n332,n1063);
nor (n1063,n1064,n1065);
and (n1064,n263,n346);
and (n1065,n270,n347);
or (n1066,n333,n910);
and (n1067,n1049,n1055);
xor (n1068,n901,n914);
and (n1069,n1024,n1046);
xor (n1070,n929,n969);
and (n1071,n1020,n1021);
and (n1072,n1015,n1016);
xor (n1073,n882,n923);
and (n1074,n1011,n1012);
nor (n1075,n6,n1008);
not (n1076,n1077);
nor (n1077,n1078,n2218);
and (n1078,n1079,n2211);
or (n1079,n1080,n2210);
and (n1080,n1081,n1260);
xor (n1081,n1082,n1253);
or (n1082,n1083,n1252);
and (n1083,n1084,n1167);
xor (n1084,n1085,n1086);
xor (n1085,n1019,n1070);
xor (n1086,n1087,n1117);
xor (n1087,n1088,n1116);
or (n1088,n1089,n1115);
and (n1089,n1090,n1093);
xor (n1090,n1091,n1092);
xor (n1091,n932,n940);
xor (n1092,n949,n962);
or (n1093,n1094,n1114);
and (n1094,n1095,n1108);
xor (n1095,n1096,n1102);
nand (n1096,n1097,n1101);
or (n1097,n17,n1098);
nor (n1098,n1099,n1100);
and (n1099,n89,n557);
and (n1100,n82,n561);
or (n1101,n18,n916);
nand (n1102,n1103,n1107);
or (n1103,n149,n1104);
nor (n1104,n1105,n1106);
and (n1105,n152,n585);
and (n1106,n153,n589);
or (n1107,n981,n178);
nand (n1108,n1109,n1113);
or (n1109,n188,n1110);
nor (n1110,n1111,n1112);
and (n1111,n218,n455);
and (n1112,n217,n456);
or (n1113,n233,n987);
and (n1114,n1096,n1102);
and (n1115,n1091,n1092);
xor (n1116,n973,n976);
or (n1117,n1118,n1166);
and (n1118,n1119,n1165);
xor (n1119,n1120,n1121);
xor (n1120,n978,n991);
or (n1121,n1122,n1164);
and (n1122,n1123,n1142);
xor (n1123,n1124,n1125);
xor (n1124,n992,n998);
or (n1125,n1126,n1141);
and (n1126,n1127,n1135);
xor (n1127,n1128,n1129);
nor (n1128,n233,n455);
nand (n1129,n1130,n1134);
or (n1130,n1131,n316);
nor (n1131,n1132,n1133);
and (n1132,n496,n310);
and (n1133,n500,n311);
or (n1134,n1000,n317);
nand (n1135,n1136,n1137);
or (n1136,n1029,n484);
or (n1137,n483,n1138);
nor (n1138,n1139,n1140);
and (n1139,n181,n260);
and (n1140,n185,n256);
and (n1141,n1128,n1129);
or (n1142,n1143,n1163);
and (n1143,n1144,n1157);
xor (n1144,n1145,n1151);
nand (n1145,n1146,n1150);
or (n1146,n509,n1147);
nor (n1147,n1148,n1149);
and (n1148,n384,n519);
and (n1149,n388,n520);
or (n1150,n1035,n529);
nand (n1151,n1152,n1156);
or (n1152,n535,n1153);
nor (n1153,n1154,n1155);
and (n1154,n415,n214);
and (n1155,n419,n209);
or (n1156,n1041,n537);
nand (n1157,n1158,n1162);
or (n1158,n459,n1159);
nor (n1159,n1160,n1161);
and (n1160,n336,n274);
and (n1161,n281,n337);
or (n1162,n460,n1051);
and (n1163,n1145,n1151);
and (n1164,n1124,n1125);
xor (n1165,n1023,n1068);
and (n1166,n1120,n1121);
or (n1167,n1168,n1251);
and (n1168,n1169,n1199);
xor (n1169,n1170,n1198);
or (n1170,n1171,n1197);
and (n1171,n1172,n1196);
xor (n1172,n1173,n1195);
or (n1173,n1174,n1194);
and (n1174,n1175,n1188);
xor (n1175,n1176,n1182);
nand (n1176,n1177,n1181);
or (n1177,n245,n1178);
nor (n1178,n1179,n1180);
and (n1179,n79,n374);
and (n1180,n74,n378);
or (n1181,n1057,n253);
nand (n1182,n1183,n1187);
or (n1183,n332,n1184);
nor (n1184,n1185,n1186);
and (n1185,n139,n346);
and (n1186,n146,n347);
or (n1187,n333,n1063);
nand (n1188,n1189,n1193);
or (n1189,n17,n1190);
nor (n1190,n1191,n1192);
and (n1191,n89,n549);
and (n1192,n82,n553);
or (n1193,n18,n1098);
and (n1194,n1176,n1182);
xor (n1195,n1048,n1061);
xor (n1196,n1026,n1039);
and (n1197,n1173,n1195);
xor (n1198,n1090,n1093);
or (n1199,n1200,n1250);
and (n1200,n1201,n1249);
xor (n1201,n1202,n1203);
xor (n1202,n1095,n1108);
or (n1203,n1204,n1248);
and (n1204,n1205,n1225);
xor (n1205,n1206,n1212);
nand (n1206,n1207,n1211);
or (n1207,n149,n1208);
nor (n1208,n1209,n1210);
and (n1209,n152,n236);
and (n1210,n153,n240);
or (n1211,n1104,n178);
and (n1212,n1213,n1219);
nor (n1213,n1214,n214);
nor (n1214,n1215,n1218);
and (n1215,n519,n1216);
not (n1216,n1217);
and (n1217,n456,n540);
and (n1218,n539,n455);
nand (n1219,n1220,n1224);
or (n1220,n1221,n316);
nor (n1221,n1222,n1223);
and (n1222,n567,n310);
and (n1223,n571,n311);
or (n1224,n1131,n317);
or (n1225,n1226,n1247);
and (n1226,n1227,n1240);
xor (n1227,n1228,n1234);
nand (n1228,n1229,n1233);
or (n1229,n483,n1230);
nor (n1230,n1231,n1232);
and (n1231,n172,n260);
and (n1232,n176,n256);
or (n1233,n1138,n484);
nand (n1234,n1235,n1239);
or (n1235,n509,n1236);
nor (n1236,n1237,n1238);
and (n1237,n423,n519);
and (n1238,n427,n520);
or (n1239,n529,n1147);
nand (n1240,n1241,n1246);
or (n1241,n1242,n535);
not (n1242,n1243);
nand (n1243,n1244,n1245);
or (n1244,n214,n456);
or (n1245,n209,n455);
or (n1246,n1153,n537);
and (n1247,n1228,n1234);
and (n1248,n1206,n1212);
xor (n1249,n1123,n1142);
and (n1250,n1202,n1203);
and (n1251,n1170,n1198);
and (n1252,n1085,n1086);
xor (n1253,n1254,n1257);
xor (n1254,n1255,n1256);
xor (n1255,n925,n971);
xor (n1256,n1014,n1017);
or (n1257,n1258,n1259);
and (n1258,n1087,n1117);
and (n1259,n1088,n1116);
nand (n1260,n1261,n2204);
or (n1261,n1262,n2197);
nand (n1262,n1263,n2186);
not (n1263,n1264);
nor (n1264,n1265,n2175);
nor (n1265,n1266,n2124);
nand (n1266,n1267,n1998);
or (n1267,n1268,n1997);
and (n1268,n1269,n1587);
xor (n1269,n1270,n1501);
or (n1270,n1271,n1500);
and (n1271,n1272,n1449);
xor (n1272,n1273,n1356);
xor (n1273,n1274,n1325);
xor (n1274,n1275,n1296);
xor (n1275,n1276,n1287);
xor (n1276,n1277,n1278);
nor (n1277,n529,n455);
nand (n1278,n1279,n1283);
or (n1279,n1280,n316);
nor (n1280,n1281,n1282);
and (n1281,n310,n139);
and (n1282,n146,n311);
or (n1283,n1284,n317);
nor (n1284,n1285,n1286);
and (n1285,n263,n310);
and (n1286,n270,n311);
nand (n1287,n1288,n1292);
or (n1288,n459,n1289);
nor (n1289,n1290,n1291);
and (n1290,n336,n181);
and (n1291,n185,n337);
or (n1292,n460,n1293);
nor (n1293,n1294,n1295);
and (n1294,n92,n336);
and (n1295,n135,n337);
or (n1296,n1297,n1324);
and (n1297,n1298,n1314);
xor (n1298,n1299,n1305);
nand (n1299,n1300,n1304);
or (n1300,n459,n1301);
nor (n1301,n1302,n1303);
and (n1302,n336,n172);
and (n1303,n176,n337);
or (n1304,n460,n1289);
nand (n1305,n1306,n1310);
or (n1306,n483,n1307);
nor (n1307,n1308,n1309);
and (n1308,n585,n260);
and (n1309,n589,n256);
or (n1310,n484,n1311);
nor (n1311,n1312,n1313);
and (n1312,n549,n260);
and (n1313,n553,n256);
nand (n1314,n1315,n1320);
or (n1315,n1316,n245);
not (n1316,n1317);
nand (n1317,n1318,n1319);
or (n1318,n74,n231);
or (n1319,n79,n227);
or (n1320,n1321,n253);
nor (n1321,n1322,n1323);
and (n1322,n79,n236);
and (n1323,n74,n240);
and (n1324,n1299,n1305);
or (n1325,n1326,n1355);
and (n1326,n1327,n1346);
xor (n1327,n1328,n1337);
nand (n1328,n1329,n1333);
or (n1329,n332,n1330);
nor (n1330,n1331,n1332);
and (n1331,n557,n346);
and (n1332,n561,n347);
or (n1333,n1334,n333);
nor (n1334,n1335,n1336);
and (n1335,n374,n346);
and (n1336,n378,n347);
nand (n1337,n1338,n1342);
or (n1338,n17,n1339);
nor (n1339,n1340,n1341);
and (n1340,n423,n89);
and (n1341,n427,n82);
or (n1342,n1343,n18);
nor (n1343,n1344,n1345);
and (n1344,n384,n89);
and (n1345,n388,n82);
nand (n1346,n1347,n1351);
or (n1347,n178,n1348);
nor (n1348,n1349,n1350);
and (n1349,n415,n152);
and (n1350,n419,n153);
or (n1351,n149,n1352);
nor (n1352,n1353,n1354);
and (n1353,n153,n455);
and (n1354,n152,n456);
and (n1355,n1328,n1337);
xor (n1356,n1357,n1405);
xor (n1357,n1358,n1385);
xor (n1358,n1359,n1372);
xor (n1359,n1360,n1366);
nand (n1360,n1361,n1362);
or (n1361,n17,n1343);
or (n1362,n1363,n18);
nor (n1363,n1364,n1365);
and (n1364,n89,n227);
and (n1365,n82,n231);
nand (n1366,n1367,n1368);
or (n1367,n149,n1348);
or (n1368,n1369,n178);
nor (n1369,n1370,n1371);
and (n1370,n423,n152);
and (n1371,n427,n153);
and (n1372,n1373,n1379);
nand (n1373,n1374,n1378);
or (n1374,n1375,n316);
nor (n1375,n1376,n1377);
and (n1376,n310,n92);
and (n1377,n135,n311);
or (n1378,n1280,n317);
nor (n1379,n1380,n152);
nor (n1380,n1381,n1384);
and (n1381,n89,n1382);
not (n1382,n1383);
and (n1383,n456,n162);
and (n1384,n166,n455);
xor (n1385,n1386,n1399);
xor (n1386,n1387,n1393);
nand (n1387,n1388,n1389);
or (n1388,n483,n1311);
or (n1389,n1390,n484);
nor (n1390,n1391,n1392);
and (n1391,n557,n260);
and (n1392,n561,n256);
nand (n1393,n1394,n1395);
or (n1394,n245,n1321);
or (n1395,n1396,n253);
nor (n1396,n1397,n1398);
and (n1397,n79,n585);
and (n1398,n74,n589);
nand (n1399,n1400,n1404);
or (n1400,n333,n1401);
nor (n1401,n1402,n1403);
and (n1402,n172,n346);
and (n1403,n176,n347);
or (n1404,n332,n1334);
or (n1405,n1406,n1448);
and (n1406,n1407,n1426);
xor (n1407,n1408,n1409);
xor (n1408,n1373,n1379);
or (n1409,n1410,n1425);
and (n1410,n1411,n1419);
xor (n1411,n1412,n1413);
nor (n1412,n178,n455);
nand (n1413,n1414,n1418);
or (n1414,n1415,n316);
nor (n1415,n1416,n1417);
and (n1416,n310,n181);
and (n1417,n185,n311);
or (n1418,n1375,n317);
nand (n1419,n1420,n1421);
or (n1420,n460,n1301);
or (n1421,n459,n1422);
nor (n1422,n1423,n1424);
and (n1423,n374,n336);
and (n1424,n378,n337);
and (n1425,n1412,n1413);
or (n1426,n1427,n1447);
and (n1427,n1428,n1441);
xor (n1428,n1429,n1435);
nand (n1429,n1430,n1434);
or (n1430,n483,n1431);
nor (n1431,n1432,n1433);
and (n1432,n236,n260);
and (n1433,n240,n256);
or (n1434,n1307,n484);
nand (n1435,n1436,n1437);
or (n1436,n253,n1316);
or (n1437,n245,n1438);
nor (n1438,n1439,n1440);
and (n1439,n79,n384);
and (n1440,n74,n388);
nand (n1441,n1442,n1443);
or (n1442,n18,n1339);
or (n1443,n17,n1444);
nor (n1444,n1445,n1446);
and (n1445,n415,n89);
and (n1446,n419,n82);
and (n1447,n1429,n1435);
and (n1448,n1408,n1409);
or (n1449,n1450,n1499);
and (n1450,n1451,n1454);
xor (n1451,n1452,n1453);
xor (n1452,n1327,n1346);
xor (n1453,n1298,n1314);
or (n1454,n1455,n1498);
and (n1455,n1456,n1476);
xor (n1456,n1457,n1463);
nand (n1457,n1458,n1462);
or (n1458,n332,n1459);
nor (n1459,n1460,n1461);
and (n1460,n549,n346);
and (n1461,n553,n347);
or (n1462,n333,n1330);
and (n1463,n1464,n1470);
nand (n1464,n1465,n1469);
or (n1465,n1466,n316);
nor (n1466,n1467,n1468);
and (n1467,n172,n310);
and (n1468,n176,n311);
or (n1469,n1415,n317);
nor (n1470,n1471,n89);
nor (n1471,n1472,n1475);
and (n1472,n79,n1473);
not (n1473,n1474);
and (n1474,n456,n20);
and (n1475,n78,n455);
or (n1476,n1477,n1497);
and (n1477,n1478,n1491);
xor (n1478,n1479,n1485);
nand (n1479,n1480,n1484);
or (n1480,n459,n1481);
nor (n1481,n1482,n1483);
and (n1482,n557,n336);
and (n1483,n561,n337);
or (n1484,n460,n1422);
nand (n1485,n1486,n1490);
or (n1486,n483,n1487);
nor (n1487,n1488,n1489);
and (n1488,n227,n260);
and (n1489,n231,n256);
or (n1490,n1431,n484);
nand (n1491,n1492,n1496);
or (n1492,n245,n1493);
nor (n1493,n1494,n1495);
and (n1494,n423,n79);
and (n1495,n427,n74);
or (n1496,n1438,n253);
and (n1497,n1479,n1485);
and (n1498,n1457,n1463);
and (n1499,n1452,n1453);
and (n1500,n1273,n1356);
xor (n1501,n1502,n1535);
xor (n1502,n1503,n1532);
xor (n1503,n1504,n1511);
xor (n1504,n1505,n1508);
or (n1505,n1506,n1507);
and (n1506,n1386,n1399);
and (n1507,n1387,n1393);
or (n1508,n1509,n1510);
and (n1509,n1359,n1372);
and (n1510,n1360,n1366);
xor (n1511,n1512,n1525);
xor (n1512,n1513,n1519);
nand (n1513,n1514,n1515);
or (n1514,n245,n1396);
or (n1515,n1516,n253);
nor (n1516,n1517,n1518);
and (n1517,n79,n549);
and (n1518,n74,n553);
nand (n1519,n1520,n1521);
or (n1520,n332,n1401);
or (n1521,n333,n1522);
nor (n1522,n1523,n1524);
and (n1523,n181,n346);
and (n1524,n185,n347);
nand (n1525,n1526,n1531);
or (n1526,n18,n1527);
not (n1527,n1528);
nand (n1528,n1529,n1530);
or (n1529,n240,n82);
or (n1530,n89,n236);
or (n1531,n17,n1363);
or (n1532,n1533,n1534);
and (n1533,n1357,n1405);
and (n1534,n1358,n1385);
xor (n1535,n1536,n1563);
xor (n1536,n1537,n1560);
xor (n1537,n1538,n1554);
xor (n1538,n1539,n1545);
nand (n1539,n1540,n1541);
or (n1540,n459,n1293);
or (n1541,n460,n1542);
nor (n1542,n1543,n1544);
and (n1543,n336,n139);
and (n1544,n146,n337);
nand (n1545,n1546,n1550);
or (n1546,n509,n1547);
nor (n1547,n1548,n1549);
and (n1548,n520,n455);
and (n1549,n519,n456);
or (n1550,n1551,n529);
nor (n1551,n1552,n1553);
and (n1552,n415,n519);
and (n1553,n419,n520);
nand (n1554,n1555,n1559);
or (n1555,n1556,n484);
nor (n1556,n1557,n1558);
and (n1557,n374,n260);
and (n1558,n378,n256);
or (n1559,n483,n1390);
or (n1560,n1561,n1562);
and (n1561,n1274,n1325);
and (n1562,n1275,n1296);
xor (n1563,n1564,n1584);
xor (n1564,n1565,n1571);
nand (n1565,n1566,n1567);
or (n1566,n149,n1369);
or (n1567,n1568,n178);
nor (n1568,n1569,n1570);
and (n1569,n384,n152);
and (n1570,n388,n153);
xor (n1571,n1572,n1578);
nand (n1572,n1573,n1574);
or (n1573,n1284,n316);
or (n1574,n1575,n317);
nor (n1575,n1576,n1577);
and (n1576,n274,n310);
and (n1577,n281,n311);
nor (n1578,n1579,n519);
nor (n1579,n1580,n1583);
and (n1580,n152,n1581);
not (n1581,n1582);
and (n1582,n456,n513);
and (n1583,n524,n455);
or (n1584,n1585,n1586);
and (n1585,n1276,n1287);
and (n1586,n1277,n1278);
or (n1587,n1588,n1996);
and (n1588,n1589,n1620);
xor (n1589,n1590,n1619);
or (n1590,n1591,n1618);
and (n1591,n1592,n1617);
xor (n1592,n1593,n1616);
or (n1593,n1594,n1615);
and (n1594,n1595,n1598);
xor (n1595,n1596,n1597);
xor (n1596,n1411,n1419);
xor (n1597,n1428,n1441);
or (n1598,n1599,n1614);
and (n1599,n1600,n1613);
xor (n1600,n1601,n1607);
nand (n1601,n1602,n1606);
or (n1602,n17,n1603);
nor (n1603,n1604,n1605);
and (n1604,n82,n455);
and (n1605,n89,n456);
or (n1606,n1444,n18);
nand (n1607,n1608,n1612);
or (n1608,n332,n1609);
nor (n1609,n1610,n1611);
and (n1610,n585,n346);
and (n1611,n589,n347);
or (n1612,n1459,n333);
xor (n1613,n1464,n1470);
and (n1614,n1601,n1607);
and (n1615,n1596,n1597);
xor (n1616,n1407,n1426);
xor (n1617,n1451,n1454);
and (n1618,n1593,n1616);
xor (n1619,n1272,n1449);
nand (n1620,n1621,n1993,n1995);
or (n1621,n1622,n1988);
nand (n1622,n1623,n1977);
or (n1623,n1624,n1976);
and (n1624,n1625,n1746);
xor (n1625,n1626,n1731);
or (n1626,n1627,n1730);
and (n1627,n1628,n1696);
xor (n1628,n1629,n1651);
xor (n1629,n1630,n1645);
xor (n1630,n1631,n1638);
nand (n1631,n1632,n1637);
or (n1632,n483,n1633);
not (n1633,n1634);
nor (n1634,n1635,n1636);
and (n1635,n260,n388);
and (n1636,n384,n256);
or (n1637,n1487,n484);
nand (n1638,n1639,n1644);
or (n1639,n1640,n245);
not (n1640,n1641);
nand (n1641,n1642,n1643);
or (n1642,n419,n74);
or (n1643,n415,n79);
or (n1644,n1493,n253);
nand (n1645,n1646,n1650);
or (n1646,n332,n1647);
nor (n1647,n1648,n1649);
and (n1648,n236,n346);
and (n1649,n240,n347);
or (n1650,n333,n1609);
or (n1651,n1652,n1695);
and (n1652,n1653,n1675);
xor (n1653,n1654,n1660);
nand (n1654,n1655,n1659);
or (n1655,n332,n1656);
nor (n1656,n1657,n1658);
and (n1657,n227,n346);
and (n1658,n231,n347);
or (n1659,n1647,n333);
xor (n1660,n1661,n1667);
nor (n1661,n1662,n79);
nor (n1662,n1663,n1666);
and (n1663,n1664,n260);
not (n1664,n1665);
and (n1665,n456,n248);
and (n1666,n252,n455);
nand (n1667,n1668,n1671);
or (n1668,n316,n1669);
not (n1669,n1670);
xnor (n1670,n557,n310);
or (n1671,n1672,n317);
nor (n1672,n1673,n1674);
and (n1673,n310,n374);
and (n1674,n378,n311);
or (n1675,n1676,n1694);
and (n1676,n1677,n1685);
xor (n1677,n1678,n1679);
nor (n1678,n253,n455);
nand (n1679,n1680,n1681);
or (n1680,n317,n1669);
or (n1681,n1682,n316);
nor (n1682,n1683,n1684);
and (n1683,n310,n549);
and (n1684,n553,n311);
nand (n1685,n1686,n1690);
or (n1686,n483,n1687);
nor (n1687,n1688,n1689);
and (n1688,n415,n260);
and (n1689,n419,n256);
or (n1690,n1691,n484);
nor (n1691,n1692,n1693);
and (n1692,n423,n260);
and (n1693,n427,n256);
and (n1694,n1678,n1679);
and (n1695,n1654,n1660);
xor (n1696,n1697,n1711);
xor (n1697,n1698,n1699);
and (n1698,n1661,n1667);
xor (n1699,n1700,n1705);
xor (n1700,n1701,n1702);
nor (n1701,n18,n455);
nand (n1702,n1703,n1704);
or (n1703,n1672,n316);
or (n1704,n1466,n317);
nand (n1705,n1706,n1710);
or (n1706,n459,n1707);
nor (n1707,n1708,n1709);
and (n1708,n549,n336);
and (n1709,n553,n337);
or (n1710,n460,n1481);
or (n1711,n1712,n1729);
and (n1712,n1713,n1723);
xor (n1713,n1714,n1720);
nand (n1714,n1715,n1719);
or (n1715,n459,n1716);
nor (n1716,n1717,n1718);
and (n1717,n336,n585);
and (n1718,n589,n337);
or (n1719,n1707,n460);
nand (n1720,n1721,n1722);
or (n1721,n484,n1633);
or (n1722,n1691,n483);
nand (n1723,n1724,n1725);
or (n1724,n253,n1640);
or (n1725,n245,n1726);
nor (n1726,n1727,n1728);
and (n1727,n74,n455);
and (n1728,n79,n456);
and (n1729,n1714,n1720);
and (n1730,n1629,n1651);
xor (n1731,n1732,n1737);
xor (n1732,n1733,n1734);
xor (n1733,n1478,n1491);
or (n1734,n1735,n1736);
and (n1735,n1697,n1711);
and (n1736,n1698,n1699);
xor (n1737,n1738,n1745);
xor (n1738,n1739,n1742);
or (n1739,n1740,n1741);
and (n1740,n1700,n1705);
and (n1741,n1701,n1702);
or (n1742,n1743,n1744);
and (n1743,n1630,n1645);
and (n1744,n1631,n1638);
xor (n1745,n1600,n1613);
or (n1746,n1747,n1975);
and (n1747,n1748,n1785);
xor (n1748,n1749,n1784);
or (n1749,n1750,n1783);
and (n1750,n1751,n1782);
xor (n1751,n1752,n1781);
or (n1752,n1753,n1780);
and (n1753,n1754,n1767);
xor (n1754,n1755,n1761);
nand (n1755,n1756,n1760);
or (n1756,n459,n1757);
nor (n1757,n1758,n1759);
and (n1758,n236,n336);
and (n1759,n337,n240);
or (n1760,n1716,n460);
nand (n1761,n1762,n1766);
or (n1762,n332,n1763);
nor (n1763,n1764,n1765);
and (n1764,n384,n346);
and (n1765,n388,n347);
or (n1766,n1656,n333);
and (n1767,n1768,n1774);
nor (n1768,n1769,n260);
nor (n1769,n1770,n1773);
and (n1770,n1771,n346);
not (n1771,n1772);
and (n1772,n456,n486);
and (n1773,n490,n455);
nand (n1774,n1775,n1779);
or (n1775,n1776,n316);
nor (n1776,n1777,n1778);
and (n1777,n310,n585);
and (n1778,n589,n311);
or (n1779,n1682,n317);
and (n1780,n1755,n1761);
xor (n1781,n1713,n1723);
xor (n1782,n1653,n1675);
and (n1783,n1752,n1781);
xor (n1784,n1628,n1696);
nand (n1785,n1786,n1972,n1974);
or (n1786,n1787,n1845);
nand (n1787,n1788,n1840);
not (n1788,n1789);
nor (n1789,n1790,n1816);
xor (n1790,n1791,n1815);
xor (n1791,n1792,n1814);
or (n1792,n1793,n1813);
and (n1793,n1794,n1807);
xor (n1794,n1795,n1801);
nand (n1795,n1796,n1800);
or (n1796,n483,n1797);
nor (n1797,n1798,n1799);
and (n1798,n256,n455);
and (n1799,n260,n456);
or (n1800,n1687,n484);
nand (n1801,n1802,n1806);
or (n1802,n1803,n459);
nor (n1803,n1804,n1805);
and (n1804,n337,n231);
and (n1805,n336,n227);
or (n1806,n1757,n460);
nand (n1807,n1808,n1812);
or (n1808,n332,n1809);
nor (n1809,n1810,n1811);
and (n1810,n423,n346);
and (n1811,n427,n347);
or (n1812,n1763,n333);
and (n1813,n1795,n1801);
xor (n1814,n1677,n1685);
xor (n1815,n1754,n1767);
or (n1816,n1817,n1839);
and (n1817,n1818,n1838);
xor (n1818,n1819,n1820);
xor (n1819,n1768,n1774);
or (n1820,n1821,n1837);
and (n1821,n1822,n1831);
xor (n1822,n1823,n1824);
nor (n1823,n484,n455);
nand (n1824,n1825,n1830);
or (n1825,n1826,n316);
not (n1826,n1827);
nand (n1827,n1828,n1829);
or (n1828,n311,n240);
nand (n1829,n240,n311);
or (n1830,n1776,n317);
nand (n1831,n1832,n1836);
or (n1832,n459,n1833);
nor (n1833,n1834,n1835);
and (n1834,n336,n384);
and (n1835,n337,n388);
or (n1836,n1803,n460);
and (n1837,n1823,n1824);
xor (n1838,n1794,n1807);
and (n1839,n1819,n1820);
or (n1840,n1841,n1842);
xor (n1841,n1751,n1782);
or (n1842,n1843,n1844);
and (n1843,n1791,n1815);
and (n1844,n1792,n1814);
nor (n1845,n1846,n1971);
and (n1846,n1847,n1966);
or (n1847,n1848,n1965);
and (n1848,n1849,n1890);
xor (n1849,n1850,n1883);
or (n1850,n1851,n1882);
and (n1851,n1852,n1868);
xor (n1852,n1853,n1859);
nand (n1853,n1854,n1858);
or (n1854,n459,n1855);
nor (n1855,n1856,n1857);
and (n1856,n337,n427);
and (n1857,n336,n423);
or (n1858,n1833,n460);
or (n1859,n1860,n1864);
nor (n1860,n1861,n333);
nor (n1861,n1862,n1863);
and (n1862,n346,n415);
and (n1863,n347,n419);
nor (n1864,n332,n1865);
nor (n1865,n1866,n1867);
and (n1866,n347,n455);
and (n1867,n346,n456);
xor (n1868,n1869,n1875);
nor (n1869,n1870,n346);
nor (n1870,n1871,n1874);
and (n1871,n1872,n336);
not (n1872,n1873);
and (n1873,n456,n340);
and (n1874,n350,n455);
nand (n1875,n1876,n1881);
or (n1876,n316,n1877);
not (n1877,n1878);
nand (n1878,n1879,n1880);
or (n1879,n310,n227);
nand (n1880,n227,n310);
nand (n1881,n1827,n318);
and (n1882,n1853,n1859);
xor (n1883,n1884,n1889);
xor (n1884,n1885,n1888);
nand (n1885,n1886,n1887);
or (n1886,n332,n1861);
or (n1887,n1809,n333);
and (n1888,n1869,n1875);
xor (n1889,n1822,n1831);
or (n1890,n1891,n1964);
and (n1891,n1892,n1912);
xor (n1892,n1893,n1911);
or (n1893,n1894,n1910);
and (n1894,n1895,n1904);
xor (n1895,n1896,n1897);
and (n1896,n334,n456);
nand (n1897,n1898,n1903);
or (n1898,n316,n1899);
not (n1899,n1900);
nand (n1900,n1901,n1902);
or (n1901,n311,n388);
nand (n1902,n388,n311);
nand (n1903,n1878,n318);
nand (n1904,n1905,n1909);
or (n1905,n459,n1906);
nor (n1906,n1907,n1908);
and (n1907,n336,n415);
and (n1908,n337,n419);
or (n1909,n1855,n460);
and (n1910,n1896,n1897);
xor (n1911,n1852,n1868);
or (n1912,n1913,n1963);
and (n1913,n1914,n1931);
xor (n1914,n1915,n1930);
and (n1915,n1916,n1922);
and (n1916,n1917,n337);
nand (n1917,n1918,n1921);
nand (n1918,n1919,n310);
not (n1919,n1920);
and (n1920,n456,n462);
nand (n1921,n466,n455);
nand (n1922,n1923,n1924);
or (n1923,n317,n1899);
nand (n1924,n1925,n1929);
not (n1925,n1926);
nor (n1926,n1927,n1928);
and (n1927,n427,n311);
and (n1928,n423,n310);
not (n1929,n316);
xor (n1930,n1895,n1904);
or (n1931,n1932,n1962);
and (n1932,n1933,n1941);
xor (n1933,n1934,n1940);
nand (n1934,n1935,n1939);
or (n1935,n459,n1936);
nor (n1936,n1937,n1938);
and (n1937,n337,n455);
and (n1938,n336,n456);
or (n1939,n1906,n460);
xor (n1940,n1916,n1922);
or (n1941,n1942,n1961);
and (n1942,n1943,n1951);
xor (n1943,n1944,n1945);
nor (n1944,n460,n455);
nand (n1945,n1946,n1950);
or (n1946,n1947,n316);
or (n1947,n1948,n1949);
and (n1948,n310,n419);
and (n1949,n415,n311);
or (n1950,n1926,n317);
nor (n1951,n1952,n1959);
nor (n1952,n1953,n1955);
and (n1953,n1954,n318);
not (n1954,n1947);
and (n1955,n1956,n1929);
nand (n1956,n1957,n1958);
or (n1957,n310,n456);
or (n1958,n311,n455);
or (n1959,n310,n1960);
and (n1960,n456,n318);
and (n1961,n1944,n1945);
and (n1962,n1934,n1940);
and (n1963,n1915,n1930);
and (n1964,n1893,n1911);
and (n1965,n1850,n1883);
or (n1966,n1967,n1968);
xor (n1967,n1818,n1838);
or (n1968,n1969,n1970);
and (n1969,n1884,n1889);
and (n1970,n1885,n1888);
and (n1971,n1967,n1968);
nand (n1972,n1840,n1973);
and (n1973,n1790,n1816);
nand (n1974,n1841,n1842);
and (n1975,n1749,n1784);
and (n1976,n1626,n1731);
or (n1977,n1978,n1985);
xor (n1978,n1979,n1984);
xor (n1979,n1980,n1981);
xor (n1980,n1456,n1476);
or (n1981,n1982,n1983);
and (n1982,n1738,n1745);
and (n1983,n1739,n1742);
xor (n1984,n1595,n1598);
or (n1985,n1986,n1987);
and (n1986,n1732,n1737);
and (n1987,n1733,n1734);
nor (n1988,n1989,n1990);
xor (n1989,n1592,n1617);
or (n1990,n1991,n1992);
and (n1991,n1979,n1984);
and (n1992,n1980,n1981);
or (n1993,n1988,n1994);
nand (n1994,n1978,n1985);
nand (n1995,n1989,n1990);
and (n1996,n1590,n1619);
and (n1997,n1270,n1501);
nor (n1998,n1999,n2119);
nor (n1999,n2000,n2110);
xor (n2000,n2001,n2065);
xor (n2001,n2002,n2040);
xor (n2002,n2003,n2025);
xor (n2003,n2004,n2005);
xor (n2004,n1227,n1240);
xor (n2005,n2006,n2019);
xor (n2006,n2007,n2013);
nand (n2007,n2008,n2012);
or (n2008,n459,n2009);
nor (n2009,n2010,n2011);
and (n2010,n336,n263);
and (n2011,n270,n337);
or (n2012,n460,n1159);
nand (n2013,n2014,n2018);
or (n2014,n245,n2015);
nor (n2015,n2016,n2017);
and (n2016,n79,n557);
and (n2017,n74,n561);
or (n2018,n1178,n253);
nand (n2019,n2020,n2024);
or (n2020,n2021,n332);
nor (n2021,n2022,n2023);
and (n2022,n92,n346);
and (n2023,n135,n347);
or (n2024,n333,n1184);
xor (n2025,n2026,n2039);
xor (n2026,n2027,n2033);
nand (n2027,n2028,n2032);
or (n2028,n17,n2029);
nor (n2029,n2030,n2031);
and (n2030,n89,n585);
and (n2031,n82,n589);
or (n2032,n1190,n18);
nand (n2033,n2034,n2038);
or (n2034,n149,n2035);
nor (n2035,n2036,n2037);
and (n2036,n152,n227);
and (n2037,n231,n153);
or (n2038,n178,n1208);
xor (n2039,n1213,n1219);
or (n2040,n2041,n2064);
and (n2041,n2042,n2049);
xor (n2042,n2043,n2046);
or (n2043,n2044,n2045);
and (n2044,n1564,n1584);
and (n2045,n1565,n1571);
or (n2046,n2047,n2048);
and (n2047,n1504,n1511);
and (n2048,n1505,n1508);
xor (n2049,n2050,n2061);
xor (n2050,n2051,n2052);
and (n2051,n1572,n1578);
xor (n2052,n2053,n2058);
xor (n2053,n2054,n2055);
nor (n2054,n537,n455);
nand (n2055,n2056,n2057);
or (n2056,n1575,n316);
or (n2057,n1221,n317);
nand (n2058,n2059,n2060);
or (n2059,n459,n1542);
or (n2060,n460,n2009);
or (n2061,n2062,n2063);
and (n2062,n1538,n1554);
and (n2063,n1539,n1545);
and (n2064,n2043,n2046);
xor (n2065,n2066,n2101);
xor (n2066,n2067,n2070);
or (n2067,n2068,n2069);
and (n2068,n2050,n2061);
and (n2069,n2051,n2052);
xor (n2070,n2071,n2088);
xor (n2071,n2072,n2075);
or (n2072,n2073,n2074);
and (n2073,n2053,n2058);
and (n2074,n2054,n2055);
or (n2075,n2076,n2087);
and (n2076,n2077,n2084);
xor (n2077,n2078,n2081);
nand (n2078,n2079,n2080);
or (n2079,n332,n1522);
or (n2080,n333,n2021);
nand (n2081,n2082,n2083);
or (n2082,n1527,n17);
or (n2083,n2029,n18);
nand (n2084,n2085,n2086);
or (n2085,n149,n1568);
or (n2086,n2035,n178);
and (n2087,n2078,n2081);
or (n2088,n2089,n2100);
and (n2089,n2090,n2097);
xor (n2090,n2091,n2094);
nand (n2091,n2092,n2093);
or (n2092,n509,n1551);
or (n2093,n1236,n529);
nand (n2094,n2095,n2096);
or (n2095,n483,n1556);
or (n2096,n1230,n484);
nand (n2097,n2098,n2099);
or (n2098,n245,n1516);
or (n2099,n2015,n253);
and (n2100,n2091,n2094);
or (n2101,n2102,n2109);
and (n2102,n2103,n2108);
xor (n2103,n2104,n2107);
or (n2104,n2105,n2106);
and (n2105,n1512,n1525);
and (n2106,n1513,n1519);
xor (n2107,n2077,n2084);
xor (n2108,n2090,n2097);
and (n2109,n2104,n2107);
or (n2110,n2111,n2118);
and (n2111,n2112,n2117);
xor (n2112,n2113,n2114);
xor (n2113,n2103,n2108);
or (n2114,n2115,n2116);
and (n2115,n1536,n1563);
and (n2116,n1537,n1560);
xor (n2117,n2042,n2049);
and (n2118,n2113,n2114);
nor (n2119,n2120,n2121);
xor (n2120,n2112,n2117);
or (n2121,n2122,n2123);
and (n2122,n1502,n1535);
and (n2123,n1503,n1532);
or (n2124,n2125,n2170);
nor (n2125,n2126,n2161);
xor (n2126,n2127,n2146);
xor (n2127,n2128,n2129);
xor (n2128,n1201,n1249);
or (n2129,n2130,n2145);
and (n2130,n2131,n2138);
xor (n2131,n2132,n2135);
or (n2132,n2133,n2134);
and (n2133,n2071,n2088);
and (n2134,n2072,n2075);
or (n2135,n2136,n2137);
and (n2136,n2003,n2025);
and (n2137,n2004,n2005);
xor (n2138,n2139,n2144);
xor (n2139,n2140,n2143);
or (n2140,n2141,n2142);
and (n2141,n2006,n2019);
and (n2142,n2007,n2013);
xor (n2143,n1175,n1188);
xor (n2144,n1127,n1135);
and (n2145,n2132,n2135);
xor (n2146,n2147,n2152);
xor (n2147,n2148,n2151);
or (n2148,n2149,n2150);
and (n2149,n2139,n2144);
and (n2150,n2140,n2143);
xor (n2151,n1172,n1196);
or (n2152,n2153,n2160);
and (n2153,n2154,n2159);
xor (n2154,n2155,n2156);
xor (n2155,n1144,n1157);
or (n2156,n2157,n2158);
and (n2157,n2026,n2039);
and (n2158,n2027,n2033);
xor (n2159,n1205,n1225);
and (n2160,n2155,n2156);
or (n2161,n2162,n2169);
and (n2162,n2163,n2168);
xor (n2163,n2164,n2165);
xor (n2164,n2154,n2159);
or (n2165,n2166,n2167);
and (n2166,n2066,n2101);
and (n2167,n2067,n2070);
xor (n2168,n2131,n2138);
and (n2169,n2164,n2165);
nor (n2170,n2171,n2174);
or (n2171,n2172,n2173);
and (n2172,n2001,n2065);
and (n2173,n2002,n2040);
xor (n2174,n2163,n2168);
nand (n2175,n2176,n2185);
or (n2176,n2177,n2125);
nor (n2177,n2178,n2184);
and (n2178,n2179,n2183);
nand (n2179,n2180,n2182);
or (n2180,n1999,n2181);
nand (n2181,n2120,n2121);
nand (n2182,n2000,n2110);
not (n2183,n2170);
and (n2184,n2171,n2174);
nand (n2185,n2126,n2161);
or (n2186,n2187,n2194);
xor (n2187,n2188,n2193);
xor (n2188,n2189,n2190);
xor (n2189,n1119,n1165);
or (n2190,n2191,n2192);
and (n2191,n2147,n2152);
and (n2192,n2148,n2151);
xor (n2193,n1169,n1199);
or (n2194,n2195,n2196);
and (n2195,n2127,n2146);
and (n2196,n2128,n2129);
and (n2197,n2198,n2200);
not (n2198,n2199);
xor (n2199,n1084,n1167);
not (n2200,n2201);
or (n2201,n2202,n2203);
and (n2202,n2188,n2193);
and (n2203,n2189,n2190);
nor (n2204,n2205,n2209);
and (n2205,n2206,n2207);
not (n2206,n2197);
not (n2207,n2208);
nand (n2208,n2187,n2194);
nor (n2209,n2198,n2200);
and (n2210,n1082,n1253);
nand (n2211,n2212,n2216);
not (n2212,n2213);
or (n2213,n2214,n2215);
and (n2214,n1254,n1257);
and (n2215,n1255,n1256);
not (n2216,n2217);
xor (n2217,n1010,n1073);
nor (n2218,n2216,n2212);
or (n2219,n1077,n3);
xor (n2220,n2221,n3865);
xor (n2221,n2222,n3862);
xor (n2222,n2223,n3861);
xor (n2223,n2224,n3853);
xor (n2224,n2225,n3852);
xor (n2225,n2226,n3837);
xor (n2226,n2227,n3836);
xor (n2227,n2228,n3816);
xor (n2228,n2229,n3815);
xor (n2229,n2230,n3788);
xor (n2230,n2231,n3787);
xor (n2231,n2232,n3755);
xor (n2232,n2233,n3754);
xor (n2233,n2234,n3715);
xor (n2234,n2235,n3714);
xor (n2235,n2236,n3670);
xor (n2236,n2237,n3669);
xor (n2237,n2238,n3618);
xor (n2238,n2239,n3617);
xor (n2239,n2240,n3561);
xor (n2240,n2241,n3560);
xor (n2241,n2242,n3497);
xor (n2242,n2243,n3496);
xor (n2243,n2244,n3428);
xor (n2244,n2245,n3427);
xor (n2245,n2246,n3352);
xor (n2246,n2247,n3351);
xor (n2247,n2248,n3271);
xor (n2248,n2249,n3270);
xor (n2249,n2250,n3183);
xor (n2250,n2251,n3182);
xor (n2251,n2252,n3090);
xor (n2252,n2253,n3089);
xor (n2253,n2254,n2991);
xor (n2254,n2255,n2990);
xor (n2255,n2256,n2886);
xor (n2256,n2257,n2885);
xor (n2257,n2258,n2774);
xor (n2258,n2259,n2773);
xor (n2259,n2260,n2657);
xor (n2260,n2261,n2656);
xor (n2261,n2262,n2533);
xor (n2262,n2263,n2532);
xor (n2263,n2264,n2404);
xor (n2264,n2265,n2403);
xor (n2265,n2266,n2269);
xor (n2266,n2267,n2268);
and (n2267,n633,n318);
and (n2268,n322,n311);
or (n2269,n2270,n2273);
and (n2270,n2271,n2272);
and (n2271,n322,n318);
and (n2272,n286,n311);
and (n2273,n2274,n2275);
xor (n2274,n2271,n2272);
or (n2275,n2276,n2279);
and (n2276,n2277,n2278);
and (n2277,n286,n318);
and (n2278,n472,n311);
and (n2279,n2280,n2281);
xor (n2280,n2277,n2278);
or (n2281,n2282,n2285);
and (n2282,n2283,n2284);
and (n2283,n472,n318);
and (n2284,n646,n311);
and (n2285,n2286,n2287);
xor (n2286,n2283,n2284);
or (n2287,n2288,n2291);
and (n2288,n2289,n2290);
and (n2289,n646,n318);
and (n2290,n362,n311);
and (n2291,n2292,n2293);
xor (n2292,n2289,n2290);
or (n2293,n2294,n2297);
and (n2294,n2295,n2296);
and (n2295,n362,n318);
and (n2296,n354,n311);
and (n2297,n2298,n2299);
xor (n2298,n2295,n2296);
or (n2299,n2300,n2303);
and (n2300,n2301,n2302);
and (n2301,n354,n318);
and (n2302,n496,n311);
and (n2303,n2304,n2305);
xor (n2304,n2301,n2302);
or (n2305,n2306,n2309);
and (n2306,n2307,n2308);
and (n2307,n496,n318);
and (n2308,n567,n311);
and (n2309,n2310,n2311);
xor (n2310,n2307,n2308);
or (n2311,n2312,n2315);
and (n2312,n2313,n2314);
and (n2313,n567,n318);
and (n2314,n274,n311);
and (n2315,n2316,n2317);
xor (n2316,n2313,n2314);
or (n2317,n2318,n2321);
and (n2318,n2319,n2320);
and (n2319,n274,n318);
and (n2320,n263,n311);
and (n2321,n2322,n2323);
xor (n2322,n2319,n2320);
or (n2323,n2324,n2327);
and (n2324,n2325,n2326);
and (n2325,n263,n318);
and (n2326,n139,n311);
and (n2327,n2328,n2329);
xor (n2328,n2325,n2326);
or (n2329,n2330,n2333);
and (n2330,n2331,n2332);
and (n2331,n139,n318);
and (n2332,n92,n311);
and (n2333,n2334,n2335);
xor (n2334,n2331,n2332);
or (n2335,n2336,n2339);
and (n2336,n2337,n2338);
and (n2337,n92,n318);
and (n2338,n181,n311);
and (n2339,n2340,n2341);
xor (n2340,n2337,n2338);
or (n2341,n2342,n2345);
and (n2342,n2343,n2344);
and (n2343,n181,n318);
and (n2344,n172,n311);
and (n2345,n2346,n2347);
xor (n2346,n2343,n2344);
or (n2347,n2348,n2351);
and (n2348,n2349,n2350);
and (n2349,n172,n318);
and (n2350,n374,n311);
and (n2351,n2352,n2353);
xor (n2352,n2349,n2350);
or (n2353,n2354,n2357);
and (n2354,n2355,n2356);
and (n2355,n374,n318);
and (n2356,n557,n311);
and (n2357,n2358,n2359);
xor (n2358,n2355,n2356);
or (n2359,n2360,n2363);
and (n2360,n2361,n2362);
and (n2361,n557,n318);
and (n2362,n549,n311);
and (n2363,n2364,n2365);
xor (n2364,n2361,n2362);
or (n2365,n2366,n2369);
and (n2366,n2367,n2368);
and (n2367,n549,n318);
and (n2368,n585,n311);
and (n2369,n2370,n2371);
xor (n2370,n2367,n2368);
or (n2371,n2372,n2375);
and (n2372,n2373,n2374);
and (n2373,n585,n318);
and (n2374,n236,n311);
and (n2375,n2376,n2377);
xor (n2376,n2373,n2374);
or (n2377,n2378,n2381);
and (n2378,n2379,n2380);
and (n2379,n236,n318);
and (n2380,n227,n311);
and (n2381,n2382,n2383);
xor (n2382,n2379,n2380);
or (n2383,n2384,n2387);
and (n2384,n2385,n2386);
and (n2385,n227,n318);
and (n2386,n384,n311);
and (n2387,n2388,n2389);
xor (n2388,n2385,n2386);
or (n2389,n2390,n2393);
and (n2390,n2391,n2392);
and (n2391,n384,n318);
and (n2392,n423,n311);
and (n2393,n2394,n2395);
xor (n2394,n2391,n2392);
or (n2395,n2396,n2398);
and (n2396,n2397,n1949);
and (n2397,n423,n318);
and (n2398,n2399,n2400);
xor (n2399,n2397,n1949);
and (n2400,n2401,n2402);
and (n2401,n415,n318);
and (n2402,n456,n311);
and (n2403,n286,n462);
or (n2404,n2405,n2408);
and (n2405,n2406,n2407);
xor (n2406,n2274,n2275);
and (n2407,n472,n462);
and (n2408,n2409,n2410);
xor (n2409,n2406,n2407);
or (n2410,n2411,n2414);
and (n2411,n2412,n2413);
xor (n2412,n2280,n2281);
and (n2413,n646,n462);
and (n2414,n2415,n2416);
xor (n2415,n2412,n2413);
or (n2416,n2417,n2420);
and (n2417,n2418,n2419);
xor (n2418,n2286,n2287);
and (n2419,n362,n462);
and (n2420,n2421,n2422);
xor (n2421,n2418,n2419);
or (n2422,n2423,n2426);
and (n2423,n2424,n2425);
xor (n2424,n2292,n2293);
and (n2425,n354,n462);
and (n2426,n2427,n2428);
xor (n2427,n2424,n2425);
or (n2428,n2429,n2432);
and (n2429,n2430,n2431);
xor (n2430,n2298,n2299);
and (n2431,n496,n462);
and (n2432,n2433,n2434);
xor (n2433,n2430,n2431);
or (n2434,n2435,n2438);
and (n2435,n2436,n2437);
xor (n2436,n2304,n2305);
and (n2437,n567,n462);
and (n2438,n2439,n2440);
xor (n2439,n2436,n2437);
or (n2440,n2441,n2444);
and (n2441,n2442,n2443);
xor (n2442,n2310,n2311);
and (n2443,n274,n462);
and (n2444,n2445,n2446);
xor (n2445,n2442,n2443);
or (n2446,n2447,n2450);
and (n2447,n2448,n2449);
xor (n2448,n2316,n2317);
and (n2449,n263,n462);
and (n2450,n2451,n2452);
xor (n2451,n2448,n2449);
or (n2452,n2453,n2456);
and (n2453,n2454,n2455);
xor (n2454,n2322,n2323);
and (n2455,n139,n462);
and (n2456,n2457,n2458);
xor (n2457,n2454,n2455);
or (n2458,n2459,n2462);
and (n2459,n2460,n2461);
xor (n2460,n2328,n2329);
and (n2461,n92,n462);
and (n2462,n2463,n2464);
xor (n2463,n2460,n2461);
or (n2464,n2465,n2468);
and (n2465,n2466,n2467);
xor (n2466,n2334,n2335);
and (n2467,n181,n462);
and (n2468,n2469,n2470);
xor (n2469,n2466,n2467);
or (n2470,n2471,n2474);
and (n2471,n2472,n2473);
xor (n2472,n2340,n2341);
and (n2473,n172,n462);
and (n2474,n2475,n2476);
xor (n2475,n2472,n2473);
or (n2476,n2477,n2480);
and (n2477,n2478,n2479);
xor (n2478,n2346,n2347);
and (n2479,n374,n462);
and (n2480,n2481,n2482);
xor (n2481,n2478,n2479);
or (n2482,n2483,n2486);
and (n2483,n2484,n2485);
xor (n2484,n2352,n2353);
and (n2485,n557,n462);
and (n2486,n2487,n2488);
xor (n2487,n2484,n2485);
or (n2488,n2489,n2492);
and (n2489,n2490,n2491);
xor (n2490,n2358,n2359);
and (n2491,n549,n462);
and (n2492,n2493,n2494);
xor (n2493,n2490,n2491);
or (n2494,n2495,n2498);
and (n2495,n2496,n2497);
xor (n2496,n2364,n2365);
and (n2497,n585,n462);
and (n2498,n2499,n2500);
xor (n2499,n2496,n2497);
or (n2500,n2501,n2504);
and (n2501,n2502,n2503);
xor (n2502,n2370,n2371);
and (n2503,n236,n462);
and (n2504,n2505,n2506);
xor (n2505,n2502,n2503);
or (n2506,n2507,n2510);
and (n2507,n2508,n2509);
xor (n2508,n2376,n2377);
and (n2509,n227,n462);
and (n2510,n2511,n2512);
xor (n2511,n2508,n2509);
or (n2512,n2513,n2516);
and (n2513,n2514,n2515);
xor (n2514,n2382,n2383);
and (n2515,n384,n462);
and (n2516,n2517,n2518);
xor (n2517,n2514,n2515);
or (n2518,n2519,n2522);
and (n2519,n2520,n2521);
xor (n2520,n2388,n2389);
and (n2521,n423,n462);
and (n2522,n2523,n2524);
xor (n2523,n2520,n2521);
or (n2524,n2525,n2528);
and (n2525,n2526,n2527);
xor (n2526,n2394,n2395);
and (n2527,n415,n462);
and (n2528,n2529,n2530);
xor (n2529,n2526,n2527);
and (n2530,n2531,n1920);
xor (n2531,n2399,n2400);
and (n2532,n472,n337);
or (n2533,n2534,n2537);
and (n2534,n2535,n2536);
xor (n2535,n2409,n2410);
and (n2536,n646,n337);
and (n2537,n2538,n2539);
xor (n2538,n2535,n2536);
or (n2539,n2540,n2543);
and (n2540,n2541,n2542);
xor (n2541,n2415,n2416);
and (n2542,n362,n337);
and (n2543,n2544,n2545);
xor (n2544,n2541,n2542);
or (n2545,n2546,n2549);
and (n2546,n2547,n2548);
xor (n2547,n2421,n2422);
and (n2548,n354,n337);
and (n2549,n2550,n2551);
xor (n2550,n2547,n2548);
or (n2551,n2552,n2555);
and (n2552,n2553,n2554);
xor (n2553,n2427,n2428);
and (n2554,n496,n337);
and (n2555,n2556,n2557);
xor (n2556,n2553,n2554);
or (n2557,n2558,n2561);
and (n2558,n2559,n2560);
xor (n2559,n2433,n2434);
and (n2560,n567,n337);
and (n2561,n2562,n2563);
xor (n2562,n2559,n2560);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2439,n2440);
and (n2566,n274,n337);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2445,n2446);
and (n2572,n263,n337);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
or (n2575,n2576,n2579);
and (n2576,n2577,n2578);
xor (n2577,n2451,n2452);
and (n2578,n139,n337);
and (n2579,n2580,n2581);
xor (n2580,n2577,n2578);
or (n2581,n2582,n2585);
and (n2582,n2583,n2584);
xor (n2583,n2457,n2458);
and (n2584,n92,n337);
and (n2585,n2586,n2587);
xor (n2586,n2583,n2584);
or (n2587,n2588,n2591);
and (n2588,n2589,n2590);
xor (n2589,n2463,n2464);
and (n2590,n181,n337);
and (n2591,n2592,n2593);
xor (n2592,n2589,n2590);
or (n2593,n2594,n2597);
and (n2594,n2595,n2596);
xor (n2595,n2469,n2470);
and (n2596,n172,n337);
and (n2597,n2598,n2599);
xor (n2598,n2595,n2596);
or (n2599,n2600,n2603);
and (n2600,n2601,n2602);
xor (n2601,n2475,n2476);
and (n2602,n374,n337);
and (n2603,n2604,n2605);
xor (n2604,n2601,n2602);
or (n2605,n2606,n2609);
and (n2606,n2607,n2608);
xor (n2607,n2481,n2482);
and (n2608,n557,n337);
and (n2609,n2610,n2611);
xor (n2610,n2607,n2608);
or (n2611,n2612,n2615);
and (n2612,n2613,n2614);
xor (n2613,n2487,n2488);
and (n2614,n549,n337);
and (n2615,n2616,n2617);
xor (n2616,n2613,n2614);
or (n2617,n2618,n2621);
and (n2618,n2619,n2620);
xor (n2619,n2493,n2494);
and (n2620,n585,n337);
and (n2621,n2622,n2623);
xor (n2622,n2619,n2620);
or (n2623,n2624,n2627);
and (n2624,n2625,n2626);
xor (n2625,n2499,n2500);
and (n2626,n236,n337);
and (n2627,n2628,n2629);
xor (n2628,n2625,n2626);
or (n2629,n2630,n2633);
and (n2630,n2631,n2632);
xor (n2631,n2505,n2506);
and (n2632,n227,n337);
and (n2633,n2634,n2635);
xor (n2634,n2631,n2632);
or (n2635,n2636,n2639);
and (n2636,n2637,n2638);
xor (n2637,n2511,n2512);
and (n2638,n384,n337);
and (n2639,n2640,n2641);
xor (n2640,n2637,n2638);
or (n2641,n2642,n2645);
and (n2642,n2643,n2644);
xor (n2643,n2517,n2518);
and (n2644,n423,n337);
and (n2645,n2646,n2647);
xor (n2646,n2643,n2644);
or (n2647,n2648,n2651);
and (n2648,n2649,n2650);
xor (n2649,n2523,n2524);
and (n2650,n415,n337);
and (n2651,n2652,n2653);
xor (n2652,n2649,n2650);
and (n2653,n2654,n2655);
xor (n2654,n2529,n2530);
and (n2655,n456,n337);
and (n2656,n646,n340);
or (n2657,n2658,n2661);
and (n2658,n2659,n2660);
xor (n2659,n2538,n2539);
and (n2660,n362,n340);
and (n2661,n2662,n2663);
xor (n2662,n2659,n2660);
or (n2663,n2664,n2667);
and (n2664,n2665,n2666);
xor (n2665,n2544,n2545);
and (n2666,n354,n340);
and (n2667,n2668,n2669);
xor (n2668,n2665,n2666);
or (n2669,n2670,n2673);
and (n2670,n2671,n2672);
xor (n2671,n2550,n2551);
and (n2672,n496,n340);
and (n2673,n2674,n2675);
xor (n2674,n2671,n2672);
or (n2675,n2676,n2679);
and (n2676,n2677,n2678);
xor (n2677,n2556,n2557);
and (n2678,n567,n340);
and (n2679,n2680,n2681);
xor (n2680,n2677,n2678);
or (n2681,n2682,n2685);
and (n2682,n2683,n2684);
xor (n2683,n2562,n2563);
and (n2684,n274,n340);
and (n2685,n2686,n2687);
xor (n2686,n2683,n2684);
or (n2687,n2688,n2691);
and (n2688,n2689,n2690);
xor (n2689,n2568,n2569);
and (n2690,n263,n340);
and (n2691,n2692,n2693);
xor (n2692,n2689,n2690);
or (n2693,n2694,n2697);
and (n2694,n2695,n2696);
xor (n2695,n2574,n2575);
and (n2696,n139,n340);
and (n2697,n2698,n2699);
xor (n2698,n2695,n2696);
or (n2699,n2700,n2703);
and (n2700,n2701,n2702);
xor (n2701,n2580,n2581);
and (n2702,n92,n340);
and (n2703,n2704,n2705);
xor (n2704,n2701,n2702);
or (n2705,n2706,n2709);
and (n2706,n2707,n2708);
xor (n2707,n2586,n2587);
and (n2708,n181,n340);
and (n2709,n2710,n2711);
xor (n2710,n2707,n2708);
or (n2711,n2712,n2715);
and (n2712,n2713,n2714);
xor (n2713,n2592,n2593);
and (n2714,n172,n340);
and (n2715,n2716,n2717);
xor (n2716,n2713,n2714);
or (n2717,n2718,n2721);
and (n2718,n2719,n2720);
xor (n2719,n2598,n2599);
and (n2720,n374,n340);
and (n2721,n2722,n2723);
xor (n2722,n2719,n2720);
or (n2723,n2724,n2727);
and (n2724,n2725,n2726);
xor (n2725,n2604,n2605);
and (n2726,n557,n340);
and (n2727,n2728,n2729);
xor (n2728,n2725,n2726);
or (n2729,n2730,n2733);
and (n2730,n2731,n2732);
xor (n2731,n2610,n2611);
and (n2732,n549,n340);
and (n2733,n2734,n2735);
xor (n2734,n2731,n2732);
or (n2735,n2736,n2739);
and (n2736,n2737,n2738);
xor (n2737,n2616,n2617);
and (n2738,n585,n340);
and (n2739,n2740,n2741);
xor (n2740,n2737,n2738);
or (n2741,n2742,n2745);
and (n2742,n2743,n2744);
xor (n2743,n2622,n2623);
and (n2744,n236,n340);
and (n2745,n2746,n2747);
xor (n2746,n2743,n2744);
or (n2747,n2748,n2751);
and (n2748,n2749,n2750);
xor (n2749,n2628,n2629);
and (n2750,n227,n340);
and (n2751,n2752,n2753);
xor (n2752,n2749,n2750);
or (n2753,n2754,n2757);
and (n2754,n2755,n2756);
xor (n2755,n2634,n2635);
and (n2756,n384,n340);
and (n2757,n2758,n2759);
xor (n2758,n2755,n2756);
or (n2759,n2760,n2763);
and (n2760,n2761,n2762);
xor (n2761,n2640,n2641);
and (n2762,n423,n340);
and (n2763,n2764,n2765);
xor (n2764,n2761,n2762);
or (n2765,n2766,n2769);
and (n2766,n2767,n2768);
xor (n2767,n2646,n2647);
and (n2768,n415,n340);
and (n2769,n2770,n2771);
xor (n2770,n2767,n2768);
and (n2771,n2772,n1873);
xor (n2772,n2652,n2653);
and (n2773,n362,n347);
or (n2774,n2775,n2778);
and (n2775,n2776,n2777);
xor (n2776,n2662,n2663);
and (n2777,n354,n347);
and (n2778,n2779,n2780);
xor (n2779,n2776,n2777);
or (n2780,n2781,n2784);
and (n2781,n2782,n2783);
xor (n2782,n2668,n2669);
and (n2783,n496,n347);
and (n2784,n2785,n2786);
xor (n2785,n2782,n2783);
or (n2786,n2787,n2790);
and (n2787,n2788,n2789);
xor (n2788,n2674,n2675);
and (n2789,n567,n347);
and (n2790,n2791,n2792);
xor (n2791,n2788,n2789);
or (n2792,n2793,n2796);
and (n2793,n2794,n2795);
xor (n2794,n2680,n2681);
and (n2795,n274,n347);
and (n2796,n2797,n2798);
xor (n2797,n2794,n2795);
or (n2798,n2799,n2802);
and (n2799,n2800,n2801);
xor (n2800,n2686,n2687);
and (n2801,n263,n347);
and (n2802,n2803,n2804);
xor (n2803,n2800,n2801);
or (n2804,n2805,n2808);
and (n2805,n2806,n2807);
xor (n2806,n2692,n2693);
and (n2807,n139,n347);
and (n2808,n2809,n2810);
xor (n2809,n2806,n2807);
or (n2810,n2811,n2814);
and (n2811,n2812,n2813);
xor (n2812,n2698,n2699);
and (n2813,n92,n347);
and (n2814,n2815,n2816);
xor (n2815,n2812,n2813);
or (n2816,n2817,n2820);
and (n2817,n2818,n2819);
xor (n2818,n2704,n2705);
and (n2819,n181,n347);
and (n2820,n2821,n2822);
xor (n2821,n2818,n2819);
or (n2822,n2823,n2826);
and (n2823,n2824,n2825);
xor (n2824,n2710,n2711);
and (n2825,n172,n347);
and (n2826,n2827,n2828);
xor (n2827,n2824,n2825);
or (n2828,n2829,n2832);
and (n2829,n2830,n2831);
xor (n2830,n2716,n2717);
and (n2831,n374,n347);
and (n2832,n2833,n2834);
xor (n2833,n2830,n2831);
or (n2834,n2835,n2838);
and (n2835,n2836,n2837);
xor (n2836,n2722,n2723);
and (n2837,n557,n347);
and (n2838,n2839,n2840);
xor (n2839,n2836,n2837);
or (n2840,n2841,n2844);
and (n2841,n2842,n2843);
xor (n2842,n2728,n2729);
and (n2843,n549,n347);
and (n2844,n2845,n2846);
xor (n2845,n2842,n2843);
or (n2846,n2847,n2850);
and (n2847,n2848,n2849);
xor (n2848,n2734,n2735);
and (n2849,n585,n347);
and (n2850,n2851,n2852);
xor (n2851,n2848,n2849);
or (n2852,n2853,n2856);
and (n2853,n2854,n2855);
xor (n2854,n2740,n2741);
and (n2855,n236,n347);
and (n2856,n2857,n2858);
xor (n2857,n2854,n2855);
or (n2858,n2859,n2862);
and (n2859,n2860,n2861);
xor (n2860,n2746,n2747);
and (n2861,n227,n347);
and (n2862,n2863,n2864);
xor (n2863,n2860,n2861);
or (n2864,n2865,n2868);
and (n2865,n2866,n2867);
xor (n2866,n2752,n2753);
and (n2867,n384,n347);
and (n2868,n2869,n2870);
xor (n2869,n2866,n2867);
or (n2870,n2871,n2874);
and (n2871,n2872,n2873);
xor (n2872,n2758,n2759);
and (n2873,n423,n347);
and (n2874,n2875,n2876);
xor (n2875,n2872,n2873);
or (n2876,n2877,n2880);
and (n2877,n2878,n2879);
xor (n2878,n2764,n2765);
and (n2879,n415,n347);
and (n2880,n2881,n2882);
xor (n2881,n2878,n2879);
and (n2882,n2883,n2884);
xor (n2883,n2770,n2771);
and (n2884,n456,n347);
and (n2885,n354,n486);
or (n2886,n2887,n2890);
and (n2887,n2888,n2889);
xor (n2888,n2779,n2780);
and (n2889,n496,n486);
and (n2890,n2891,n2892);
xor (n2891,n2888,n2889);
or (n2892,n2893,n2896);
and (n2893,n2894,n2895);
xor (n2894,n2785,n2786);
and (n2895,n567,n486);
and (n2896,n2897,n2898);
xor (n2897,n2894,n2895);
or (n2898,n2899,n2902);
and (n2899,n2900,n2901);
xor (n2900,n2791,n2792);
and (n2901,n274,n486);
and (n2902,n2903,n2904);
xor (n2903,n2900,n2901);
or (n2904,n2905,n2908);
and (n2905,n2906,n2907);
xor (n2906,n2797,n2798);
and (n2907,n263,n486);
and (n2908,n2909,n2910);
xor (n2909,n2906,n2907);
or (n2910,n2911,n2914);
and (n2911,n2912,n2913);
xor (n2912,n2803,n2804);
and (n2913,n139,n486);
and (n2914,n2915,n2916);
xor (n2915,n2912,n2913);
or (n2916,n2917,n2920);
and (n2917,n2918,n2919);
xor (n2918,n2809,n2810);
and (n2919,n92,n486);
and (n2920,n2921,n2922);
xor (n2921,n2918,n2919);
or (n2922,n2923,n2926);
and (n2923,n2924,n2925);
xor (n2924,n2815,n2816);
and (n2925,n181,n486);
and (n2926,n2927,n2928);
xor (n2927,n2924,n2925);
or (n2928,n2929,n2932);
and (n2929,n2930,n2931);
xor (n2930,n2821,n2822);
and (n2931,n172,n486);
and (n2932,n2933,n2934);
xor (n2933,n2930,n2931);
or (n2934,n2935,n2938);
and (n2935,n2936,n2937);
xor (n2936,n2827,n2828);
and (n2937,n374,n486);
and (n2938,n2939,n2940);
xor (n2939,n2936,n2937);
or (n2940,n2941,n2944);
and (n2941,n2942,n2943);
xor (n2942,n2833,n2834);
and (n2943,n557,n486);
and (n2944,n2945,n2946);
xor (n2945,n2942,n2943);
or (n2946,n2947,n2950);
and (n2947,n2948,n2949);
xor (n2948,n2839,n2840);
and (n2949,n549,n486);
and (n2950,n2951,n2952);
xor (n2951,n2948,n2949);
or (n2952,n2953,n2956);
and (n2953,n2954,n2955);
xor (n2954,n2845,n2846);
and (n2955,n585,n486);
and (n2956,n2957,n2958);
xor (n2957,n2954,n2955);
or (n2958,n2959,n2962);
and (n2959,n2960,n2961);
xor (n2960,n2851,n2852);
and (n2961,n236,n486);
and (n2962,n2963,n2964);
xor (n2963,n2960,n2961);
or (n2964,n2965,n2968);
and (n2965,n2966,n2967);
xor (n2966,n2857,n2858);
and (n2967,n227,n486);
and (n2968,n2969,n2970);
xor (n2969,n2966,n2967);
or (n2970,n2971,n2974);
and (n2971,n2972,n2973);
xor (n2972,n2863,n2864);
and (n2973,n384,n486);
and (n2974,n2975,n2976);
xor (n2975,n2972,n2973);
or (n2976,n2977,n2980);
and (n2977,n2978,n2979);
xor (n2978,n2869,n2870);
and (n2979,n423,n486);
and (n2980,n2981,n2982);
xor (n2981,n2978,n2979);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
xor (n2984,n2875,n2876);
and (n2985,n415,n486);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
and (n2988,n2989,n1772);
xor (n2989,n2881,n2882);
and (n2990,n496,n256);
or (n2991,n2992,n2995);
and (n2992,n2993,n2994);
xor (n2993,n2891,n2892);
and (n2994,n567,n256);
and (n2995,n2996,n2997);
xor (n2996,n2993,n2994);
or (n2997,n2998,n3001);
and (n2998,n2999,n3000);
xor (n2999,n2897,n2898);
and (n3000,n274,n256);
and (n3001,n3002,n3003);
xor (n3002,n2999,n3000);
or (n3003,n3004,n3007);
and (n3004,n3005,n3006);
xor (n3005,n2903,n2904);
and (n3006,n263,n256);
and (n3007,n3008,n3009);
xor (n3008,n3005,n3006);
or (n3009,n3010,n3013);
and (n3010,n3011,n3012);
xor (n3011,n2909,n2910);
and (n3012,n139,n256);
and (n3013,n3014,n3015);
xor (n3014,n3011,n3012);
or (n3015,n3016,n3019);
and (n3016,n3017,n3018);
xor (n3017,n2915,n2916);
and (n3018,n92,n256);
and (n3019,n3020,n3021);
xor (n3020,n3017,n3018);
or (n3021,n3022,n3025);
and (n3022,n3023,n3024);
xor (n3023,n2921,n2922);
and (n3024,n181,n256);
and (n3025,n3026,n3027);
xor (n3026,n3023,n3024);
or (n3027,n3028,n3031);
and (n3028,n3029,n3030);
xor (n3029,n2927,n2928);
and (n3030,n172,n256);
and (n3031,n3032,n3033);
xor (n3032,n3029,n3030);
or (n3033,n3034,n3037);
and (n3034,n3035,n3036);
xor (n3035,n2933,n2934);
and (n3036,n374,n256);
and (n3037,n3038,n3039);
xor (n3038,n3035,n3036);
or (n3039,n3040,n3043);
and (n3040,n3041,n3042);
xor (n3041,n2939,n2940);
and (n3042,n557,n256);
and (n3043,n3044,n3045);
xor (n3044,n3041,n3042);
or (n3045,n3046,n3049);
and (n3046,n3047,n3048);
xor (n3047,n2945,n2946);
and (n3048,n549,n256);
and (n3049,n3050,n3051);
xor (n3050,n3047,n3048);
or (n3051,n3052,n3055);
and (n3052,n3053,n3054);
xor (n3053,n2951,n2952);
and (n3054,n585,n256);
and (n3055,n3056,n3057);
xor (n3056,n3053,n3054);
or (n3057,n3058,n3061);
and (n3058,n3059,n3060);
xor (n3059,n2957,n2958);
and (n3060,n236,n256);
and (n3061,n3062,n3063);
xor (n3062,n3059,n3060);
or (n3063,n3064,n3067);
and (n3064,n3065,n3066);
xor (n3065,n2963,n2964);
and (n3066,n227,n256);
and (n3067,n3068,n3069);
xor (n3068,n3065,n3066);
or (n3069,n3070,n3072);
and (n3070,n3071,n1636);
xor (n3071,n2969,n2970);
and (n3072,n3073,n3074);
xor (n3073,n3071,n1636);
or (n3074,n3075,n3078);
and (n3075,n3076,n3077);
xor (n3076,n2975,n2976);
and (n3077,n423,n256);
and (n3078,n3079,n3080);
xor (n3079,n3076,n3077);
or (n3080,n3081,n3084);
and (n3081,n3082,n3083);
xor (n3082,n2981,n2982);
and (n3083,n415,n256);
and (n3084,n3085,n3086);
xor (n3085,n3082,n3083);
and (n3086,n3087,n3088);
xor (n3087,n2987,n2988);
and (n3088,n456,n256);
and (n3089,n567,n248);
or (n3090,n3091,n3094);
and (n3091,n3092,n3093);
xor (n3092,n2996,n2997);
and (n3093,n274,n248);
and (n3094,n3095,n3096);
xor (n3095,n3092,n3093);
or (n3096,n3097,n3100);
and (n3097,n3098,n3099);
xor (n3098,n3002,n3003);
and (n3099,n263,n248);
and (n3100,n3101,n3102);
xor (n3101,n3098,n3099);
or (n3102,n3103,n3106);
and (n3103,n3104,n3105);
xor (n3104,n3008,n3009);
and (n3105,n139,n248);
and (n3106,n3107,n3108);
xor (n3107,n3104,n3105);
or (n3108,n3109,n3112);
and (n3109,n3110,n3111);
xor (n3110,n3014,n3015);
and (n3111,n92,n248);
and (n3112,n3113,n3114);
xor (n3113,n3110,n3111);
or (n3114,n3115,n3118);
and (n3115,n3116,n3117);
xor (n3116,n3020,n3021);
and (n3117,n181,n248);
and (n3118,n3119,n3120);
xor (n3119,n3116,n3117);
or (n3120,n3121,n3124);
and (n3121,n3122,n3123);
xor (n3122,n3026,n3027);
and (n3123,n172,n248);
and (n3124,n3125,n3126);
xor (n3125,n3122,n3123);
or (n3126,n3127,n3130);
and (n3127,n3128,n3129);
xor (n3128,n3032,n3033);
and (n3129,n374,n248);
and (n3130,n3131,n3132);
xor (n3131,n3128,n3129);
or (n3132,n3133,n3136);
and (n3133,n3134,n3135);
xor (n3134,n3038,n3039);
and (n3135,n557,n248);
and (n3136,n3137,n3138);
xor (n3137,n3134,n3135);
or (n3138,n3139,n3142);
and (n3139,n3140,n3141);
xor (n3140,n3044,n3045);
and (n3141,n549,n248);
and (n3142,n3143,n3144);
xor (n3143,n3140,n3141);
or (n3144,n3145,n3148);
and (n3145,n3146,n3147);
xor (n3146,n3050,n3051);
and (n3147,n585,n248);
and (n3148,n3149,n3150);
xor (n3149,n3146,n3147);
or (n3150,n3151,n3154);
and (n3151,n3152,n3153);
xor (n3152,n3056,n3057);
and (n3153,n236,n248);
and (n3154,n3155,n3156);
xor (n3155,n3152,n3153);
or (n3156,n3157,n3160);
and (n3157,n3158,n3159);
xor (n3158,n3062,n3063);
and (n3159,n227,n248);
and (n3160,n3161,n3162);
xor (n3161,n3158,n3159);
or (n3162,n3163,n3166);
and (n3163,n3164,n3165);
xor (n3164,n3068,n3069);
and (n3165,n384,n248);
and (n3166,n3167,n3168);
xor (n3167,n3164,n3165);
or (n3168,n3169,n3172);
and (n3169,n3170,n3171);
xor (n3170,n3073,n3074);
and (n3171,n423,n248);
and (n3172,n3173,n3174);
xor (n3173,n3170,n3171);
or (n3174,n3175,n3178);
and (n3175,n3176,n3177);
xor (n3176,n3079,n3080);
and (n3177,n415,n248);
and (n3178,n3179,n3180);
xor (n3179,n3176,n3177);
and (n3180,n3181,n1665);
xor (n3181,n3085,n3086);
and (n3182,n274,n74);
or (n3183,n3184,n3187);
and (n3184,n3185,n3186);
xor (n3185,n3095,n3096);
and (n3186,n263,n74);
and (n3187,n3188,n3189);
xor (n3188,n3185,n3186);
or (n3189,n3190,n3193);
and (n3190,n3191,n3192);
xor (n3191,n3101,n3102);
and (n3192,n139,n74);
and (n3193,n3194,n3195);
xor (n3194,n3191,n3192);
or (n3195,n3196,n3199);
and (n3196,n3197,n3198);
xor (n3197,n3107,n3108);
and (n3198,n92,n74);
and (n3199,n3200,n3201);
xor (n3200,n3197,n3198);
or (n3201,n3202,n3205);
and (n3202,n3203,n3204);
xor (n3203,n3113,n3114);
and (n3204,n181,n74);
and (n3205,n3206,n3207);
xor (n3206,n3203,n3204);
or (n3207,n3208,n3211);
and (n3208,n3209,n3210);
xor (n3209,n3119,n3120);
and (n3210,n172,n74);
and (n3211,n3212,n3213);
xor (n3212,n3209,n3210);
or (n3213,n3214,n3217);
and (n3214,n3215,n3216);
xor (n3215,n3125,n3126);
and (n3216,n374,n74);
and (n3217,n3218,n3219);
xor (n3218,n3215,n3216);
or (n3219,n3220,n3223);
and (n3220,n3221,n3222);
xor (n3221,n3131,n3132);
and (n3222,n557,n74);
and (n3223,n3224,n3225);
xor (n3224,n3221,n3222);
or (n3225,n3226,n3229);
and (n3226,n3227,n3228);
xor (n3227,n3137,n3138);
and (n3228,n549,n74);
and (n3229,n3230,n3231);
xor (n3230,n3227,n3228);
or (n3231,n3232,n3235);
and (n3232,n3233,n3234);
xor (n3233,n3143,n3144);
and (n3234,n585,n74);
and (n3235,n3236,n3237);
xor (n3236,n3233,n3234);
or (n3237,n3238,n3241);
and (n3238,n3239,n3240);
xor (n3239,n3149,n3150);
and (n3240,n236,n74);
and (n3241,n3242,n3243);
xor (n3242,n3239,n3240);
or (n3243,n3244,n3247);
and (n3244,n3245,n3246);
xor (n3245,n3155,n3156);
and (n3246,n227,n74);
and (n3247,n3248,n3249);
xor (n3248,n3245,n3246);
or (n3249,n3250,n3253);
and (n3250,n3251,n3252);
xor (n3251,n3161,n3162);
and (n3252,n384,n74);
and (n3253,n3254,n3255);
xor (n3254,n3251,n3252);
or (n3255,n3256,n3259);
and (n3256,n3257,n3258);
xor (n3257,n3167,n3168);
and (n3258,n423,n74);
and (n3259,n3260,n3261);
xor (n3260,n3257,n3258);
or (n3261,n3262,n3265);
and (n3262,n3263,n3264);
xor (n3263,n3173,n3174);
and (n3264,n415,n74);
and (n3265,n3266,n3267);
xor (n3266,n3263,n3264);
and (n3267,n3268,n3269);
xor (n3268,n3179,n3180);
and (n3269,n456,n74);
and (n3270,n263,n20);
or (n3271,n3272,n3275);
and (n3272,n3273,n3274);
xor (n3273,n3188,n3189);
and (n3274,n139,n20);
and (n3275,n3276,n3277);
xor (n3276,n3273,n3274);
or (n3277,n3278,n3281);
and (n3278,n3279,n3280);
xor (n3279,n3194,n3195);
and (n3280,n92,n20);
and (n3281,n3282,n3283);
xor (n3282,n3279,n3280);
or (n3283,n3284,n3287);
and (n3284,n3285,n3286);
xor (n3285,n3200,n3201);
and (n3286,n181,n20);
and (n3287,n3288,n3289);
xor (n3288,n3285,n3286);
or (n3289,n3290,n3293);
and (n3290,n3291,n3292);
xor (n3291,n3206,n3207);
and (n3292,n172,n20);
and (n3293,n3294,n3295);
xor (n3294,n3291,n3292);
or (n3295,n3296,n3299);
and (n3296,n3297,n3298);
xor (n3297,n3212,n3213);
and (n3298,n374,n20);
and (n3299,n3300,n3301);
xor (n3300,n3297,n3298);
or (n3301,n3302,n3305);
and (n3302,n3303,n3304);
xor (n3303,n3218,n3219);
and (n3304,n557,n20);
and (n3305,n3306,n3307);
xor (n3306,n3303,n3304);
or (n3307,n3308,n3311);
and (n3308,n3309,n3310);
xor (n3309,n3224,n3225);
and (n3310,n549,n20);
and (n3311,n3312,n3313);
xor (n3312,n3309,n3310);
or (n3313,n3314,n3317);
and (n3314,n3315,n3316);
xor (n3315,n3230,n3231);
and (n3316,n585,n20);
and (n3317,n3318,n3319);
xor (n3318,n3315,n3316);
or (n3319,n3320,n3323);
and (n3320,n3321,n3322);
xor (n3321,n3236,n3237);
and (n3322,n236,n20);
and (n3323,n3324,n3325);
xor (n3324,n3321,n3322);
or (n3325,n3326,n3329);
and (n3326,n3327,n3328);
xor (n3327,n3242,n3243);
and (n3328,n227,n20);
and (n3329,n3330,n3331);
xor (n3330,n3327,n3328);
or (n3331,n3332,n3335);
and (n3332,n3333,n3334);
xor (n3333,n3248,n3249);
and (n3334,n384,n20);
and (n3335,n3336,n3337);
xor (n3336,n3333,n3334);
or (n3337,n3338,n3341);
and (n3338,n3339,n3340);
xor (n3339,n3254,n3255);
and (n3340,n423,n20);
and (n3341,n3342,n3343);
xor (n3342,n3339,n3340);
or (n3343,n3344,n3347);
and (n3344,n3345,n3346);
xor (n3345,n3260,n3261);
and (n3346,n415,n20);
and (n3347,n3348,n3349);
xor (n3348,n3345,n3346);
and (n3349,n3350,n1474);
xor (n3350,n3266,n3267);
and (n3351,n139,n82);
or (n3352,n3353,n3356);
and (n3353,n3354,n3355);
xor (n3354,n3276,n3277);
and (n3355,n92,n82);
and (n3356,n3357,n3358);
xor (n3357,n3354,n3355);
or (n3358,n3359,n3362);
and (n3359,n3360,n3361);
xor (n3360,n3282,n3283);
and (n3361,n181,n82);
and (n3362,n3363,n3364);
xor (n3363,n3360,n3361);
or (n3364,n3365,n3368);
and (n3365,n3366,n3367);
xor (n3366,n3288,n3289);
and (n3367,n172,n82);
and (n3368,n3369,n3370);
xor (n3369,n3366,n3367);
or (n3370,n3371,n3374);
and (n3371,n3372,n3373);
xor (n3372,n3294,n3295);
and (n3373,n374,n82);
and (n3374,n3375,n3376);
xor (n3375,n3372,n3373);
or (n3376,n3377,n3380);
and (n3377,n3378,n3379);
xor (n3378,n3300,n3301);
and (n3379,n557,n82);
and (n3380,n3381,n3382);
xor (n3381,n3378,n3379);
or (n3382,n3383,n3386);
and (n3383,n3384,n3385);
xor (n3384,n3306,n3307);
and (n3385,n549,n82);
and (n3386,n3387,n3388);
xor (n3387,n3384,n3385);
or (n3388,n3389,n3392);
and (n3389,n3390,n3391);
xor (n3390,n3312,n3313);
and (n3391,n585,n82);
and (n3392,n3393,n3394);
xor (n3393,n3390,n3391);
or (n3394,n3395,n3398);
and (n3395,n3396,n3397);
xor (n3396,n3318,n3319);
and (n3397,n236,n82);
and (n3398,n3399,n3400);
xor (n3399,n3396,n3397);
or (n3400,n3401,n3404);
and (n3401,n3402,n3403);
xor (n3402,n3324,n3325);
and (n3403,n227,n82);
and (n3404,n3405,n3406);
xor (n3405,n3402,n3403);
or (n3406,n3407,n3410);
and (n3407,n3408,n3409);
xor (n3408,n3330,n3331);
and (n3409,n384,n82);
and (n3410,n3411,n3412);
xor (n3411,n3408,n3409);
or (n3412,n3413,n3416);
and (n3413,n3414,n3415);
xor (n3414,n3336,n3337);
and (n3415,n423,n82);
and (n3416,n3417,n3418);
xor (n3417,n3414,n3415);
or (n3418,n3419,n3422);
and (n3419,n3420,n3421);
xor (n3420,n3342,n3343);
and (n3421,n415,n82);
and (n3422,n3423,n3424);
xor (n3423,n3420,n3421);
and (n3424,n3425,n3426);
xor (n3425,n3348,n3349);
and (n3426,n456,n82);
and (n3427,n92,n162);
or (n3428,n3429,n3432);
and (n3429,n3430,n3431);
xor (n3430,n3357,n3358);
and (n3431,n181,n162);
and (n3432,n3433,n3434);
xor (n3433,n3430,n3431);
or (n3434,n3435,n3438);
and (n3435,n3436,n3437);
xor (n3436,n3363,n3364);
and (n3437,n172,n162);
and (n3438,n3439,n3440);
xor (n3439,n3436,n3437);
or (n3440,n3441,n3444);
and (n3441,n3442,n3443);
xor (n3442,n3369,n3370);
and (n3443,n374,n162);
and (n3444,n3445,n3446);
xor (n3445,n3442,n3443);
or (n3446,n3447,n3450);
and (n3447,n3448,n3449);
xor (n3448,n3375,n3376);
and (n3449,n557,n162);
and (n3450,n3451,n3452);
xor (n3451,n3448,n3449);
or (n3452,n3453,n3456);
and (n3453,n3454,n3455);
xor (n3454,n3381,n3382);
and (n3455,n549,n162);
and (n3456,n3457,n3458);
xor (n3457,n3454,n3455);
or (n3458,n3459,n3462);
and (n3459,n3460,n3461);
xor (n3460,n3387,n3388);
and (n3461,n585,n162);
and (n3462,n3463,n3464);
xor (n3463,n3460,n3461);
or (n3464,n3465,n3468);
and (n3465,n3466,n3467);
xor (n3466,n3393,n3394);
and (n3467,n236,n162);
and (n3468,n3469,n3470);
xor (n3469,n3466,n3467);
or (n3470,n3471,n3474);
and (n3471,n3472,n3473);
xor (n3472,n3399,n3400);
and (n3473,n227,n162);
and (n3474,n3475,n3476);
xor (n3475,n3472,n3473);
or (n3476,n3477,n3480);
and (n3477,n3478,n3479);
xor (n3478,n3405,n3406);
and (n3479,n384,n162);
and (n3480,n3481,n3482);
xor (n3481,n3478,n3479);
or (n3482,n3483,n3486);
and (n3483,n3484,n3485);
xor (n3484,n3411,n3412);
and (n3485,n423,n162);
and (n3486,n3487,n3488);
xor (n3487,n3484,n3485);
or (n3488,n3489,n3492);
and (n3489,n3490,n3491);
xor (n3490,n3417,n3418);
and (n3491,n415,n162);
and (n3492,n3493,n3494);
xor (n3493,n3490,n3491);
and (n3494,n3495,n1383);
xor (n3495,n3423,n3424);
and (n3496,n181,n153);
or (n3497,n3498,n3501);
and (n3498,n3499,n3500);
xor (n3499,n3433,n3434);
and (n3500,n172,n153);
and (n3501,n3502,n3503);
xor (n3502,n3499,n3500);
or (n3503,n3504,n3507);
and (n3504,n3505,n3506);
xor (n3505,n3439,n3440);
and (n3506,n374,n153);
and (n3507,n3508,n3509);
xor (n3508,n3505,n3506);
or (n3509,n3510,n3513);
and (n3510,n3511,n3512);
xor (n3511,n3445,n3446);
and (n3512,n557,n153);
and (n3513,n3514,n3515);
xor (n3514,n3511,n3512);
or (n3515,n3516,n3519);
and (n3516,n3517,n3518);
xor (n3517,n3451,n3452);
and (n3518,n549,n153);
and (n3519,n3520,n3521);
xor (n3520,n3517,n3518);
or (n3521,n3522,n3525);
and (n3522,n3523,n3524);
xor (n3523,n3457,n3458);
and (n3524,n585,n153);
and (n3525,n3526,n3527);
xor (n3526,n3523,n3524);
or (n3527,n3528,n3531);
and (n3528,n3529,n3530);
xor (n3529,n3463,n3464);
and (n3530,n236,n153);
and (n3531,n3532,n3533);
xor (n3532,n3529,n3530);
or (n3533,n3534,n3537);
and (n3534,n3535,n3536);
xor (n3535,n3469,n3470);
and (n3536,n227,n153);
and (n3537,n3538,n3539);
xor (n3538,n3535,n3536);
or (n3539,n3540,n3543);
and (n3540,n3541,n3542);
xor (n3541,n3475,n3476);
and (n3542,n384,n153);
and (n3543,n3544,n3545);
xor (n3544,n3541,n3542);
or (n3545,n3546,n3549);
and (n3546,n3547,n3548);
xor (n3547,n3481,n3482);
and (n3548,n423,n153);
and (n3549,n3550,n3551);
xor (n3550,n3547,n3548);
or (n3551,n3552,n3555);
and (n3552,n3553,n3554);
xor (n3553,n3487,n3488);
and (n3554,n415,n153);
and (n3555,n3556,n3557);
xor (n3556,n3553,n3554);
and (n3557,n3558,n3559);
xor (n3558,n3493,n3494);
and (n3559,n456,n153);
and (n3560,n172,n513);
or (n3561,n3562,n3565);
and (n3562,n3563,n3564);
xor (n3563,n3502,n3503);
and (n3564,n374,n513);
and (n3565,n3566,n3567);
xor (n3566,n3563,n3564);
or (n3567,n3568,n3571);
and (n3568,n3569,n3570);
xor (n3569,n3508,n3509);
and (n3570,n557,n513);
and (n3571,n3572,n3573);
xor (n3572,n3569,n3570);
or (n3573,n3574,n3577);
and (n3574,n3575,n3576);
xor (n3575,n3514,n3515);
and (n3576,n549,n513);
and (n3577,n3578,n3579);
xor (n3578,n3575,n3576);
or (n3579,n3580,n3583);
and (n3580,n3581,n3582);
xor (n3581,n3520,n3521);
and (n3582,n585,n513);
and (n3583,n3584,n3585);
xor (n3584,n3581,n3582);
or (n3585,n3586,n3589);
and (n3586,n3587,n3588);
xor (n3587,n3526,n3527);
and (n3588,n236,n513);
and (n3589,n3590,n3591);
xor (n3590,n3587,n3588);
or (n3591,n3592,n3595);
and (n3592,n3593,n3594);
xor (n3593,n3532,n3533);
and (n3594,n227,n513);
and (n3595,n3596,n3597);
xor (n3596,n3593,n3594);
or (n3597,n3598,n3601);
and (n3598,n3599,n3600);
xor (n3599,n3538,n3539);
and (n3600,n384,n513);
and (n3601,n3602,n3603);
xor (n3602,n3599,n3600);
or (n3603,n3604,n3607);
and (n3604,n3605,n3606);
xor (n3605,n3544,n3545);
and (n3606,n423,n513);
and (n3607,n3608,n3609);
xor (n3608,n3605,n3606);
or (n3609,n3610,n3613);
and (n3610,n3611,n3612);
xor (n3611,n3550,n3551);
and (n3612,n415,n513);
and (n3613,n3614,n3615);
xor (n3614,n3611,n3612);
and (n3615,n3616,n1582);
xor (n3616,n3556,n3557);
and (n3617,n374,n520);
or (n3618,n3619,n3622);
and (n3619,n3620,n3621);
xor (n3620,n3566,n3567);
and (n3621,n557,n520);
and (n3622,n3623,n3624);
xor (n3623,n3620,n3621);
or (n3624,n3625,n3628);
and (n3625,n3626,n3627);
xor (n3626,n3572,n3573);
and (n3627,n549,n520);
and (n3628,n3629,n3630);
xor (n3629,n3626,n3627);
or (n3630,n3631,n3634);
and (n3631,n3632,n3633);
xor (n3632,n3578,n3579);
and (n3633,n585,n520);
and (n3634,n3635,n3636);
xor (n3635,n3632,n3633);
or (n3636,n3637,n3640);
and (n3637,n3638,n3639);
xor (n3638,n3584,n3585);
and (n3639,n236,n520);
and (n3640,n3641,n3642);
xor (n3641,n3638,n3639);
or (n3642,n3643,n3646);
and (n3643,n3644,n3645);
xor (n3644,n3590,n3591);
and (n3645,n227,n520);
and (n3646,n3647,n3648);
xor (n3647,n3644,n3645);
or (n3648,n3649,n3652);
and (n3649,n3650,n3651);
xor (n3650,n3596,n3597);
and (n3651,n384,n520);
and (n3652,n3653,n3654);
xor (n3653,n3650,n3651);
or (n3654,n3655,n3658);
and (n3655,n3656,n3657);
xor (n3656,n3602,n3603);
and (n3657,n423,n520);
and (n3658,n3659,n3660);
xor (n3659,n3656,n3657);
or (n3660,n3661,n3664);
and (n3661,n3662,n3663);
xor (n3662,n3608,n3609);
and (n3663,n415,n520);
and (n3664,n3665,n3666);
xor (n3665,n3662,n3663);
and (n3666,n3667,n3668);
xor (n3667,n3614,n3615);
and (n3668,n456,n520);
and (n3669,n557,n540);
or (n3670,n3671,n3674);
and (n3671,n3672,n3673);
xor (n3672,n3623,n3624);
and (n3673,n549,n540);
and (n3674,n3675,n3676);
xor (n3675,n3672,n3673);
or (n3676,n3677,n3680);
and (n3677,n3678,n3679);
xor (n3678,n3629,n3630);
and (n3679,n585,n540);
and (n3680,n3681,n3682);
xor (n3681,n3678,n3679);
or (n3682,n3683,n3686);
and (n3683,n3684,n3685);
xor (n3684,n3635,n3636);
and (n3685,n236,n540);
and (n3686,n3687,n3688);
xor (n3687,n3684,n3685);
or (n3688,n3689,n3692);
and (n3689,n3690,n3691);
xor (n3690,n3641,n3642);
and (n3691,n227,n540);
and (n3692,n3693,n3694);
xor (n3693,n3690,n3691);
or (n3694,n3695,n3698);
and (n3695,n3696,n3697);
xor (n3696,n3647,n3648);
and (n3697,n384,n540);
and (n3698,n3699,n3700);
xor (n3699,n3696,n3697);
or (n3700,n3701,n3704);
and (n3701,n3702,n3703);
xor (n3702,n3653,n3654);
and (n3703,n423,n540);
and (n3704,n3705,n3706);
xor (n3705,n3702,n3703);
or (n3706,n3707,n3710);
and (n3707,n3708,n3709);
xor (n3708,n3659,n3660);
and (n3709,n415,n540);
and (n3710,n3711,n3712);
xor (n3711,n3708,n3709);
and (n3712,n3713,n1217);
xor (n3713,n3665,n3666);
and (n3714,n549,n209);
or (n3715,n3716,n3719);
and (n3716,n3717,n3718);
xor (n3717,n3675,n3676);
and (n3718,n585,n209);
and (n3719,n3720,n3721);
xor (n3720,n3717,n3718);
or (n3721,n3722,n3725);
and (n3722,n3723,n3724);
xor (n3723,n3681,n3682);
and (n3724,n236,n209);
and (n3725,n3726,n3727);
xor (n3726,n3723,n3724);
or (n3727,n3728,n3731);
and (n3728,n3729,n3730);
xor (n3729,n3687,n3688);
and (n3730,n227,n209);
and (n3731,n3732,n3733);
xor (n3732,n3729,n3730);
or (n3733,n3734,n3737);
and (n3734,n3735,n3736);
xor (n3735,n3693,n3694);
and (n3736,n384,n209);
and (n3737,n3738,n3739);
xor (n3738,n3735,n3736);
or (n3739,n3740,n3743);
and (n3740,n3741,n3742);
xor (n3741,n3699,n3700);
and (n3742,n423,n209);
and (n3743,n3744,n3745);
xor (n3744,n3741,n3742);
or (n3745,n3746,n3749);
and (n3746,n3747,n3748);
xor (n3747,n3705,n3706);
and (n3748,n415,n209);
and (n3749,n3750,n3751);
xor (n3750,n3747,n3748);
and (n3751,n3752,n3753);
xor (n3752,n3711,n3712);
and (n3753,n456,n209);
and (n3754,n585,n191);
or (n3755,n3756,n3759);
and (n3756,n3757,n3758);
xor (n3757,n3720,n3721);
and (n3758,n236,n191);
and (n3759,n3760,n3761);
xor (n3760,n3757,n3758);
or (n3761,n3762,n3765);
and (n3762,n3763,n3764);
xor (n3763,n3726,n3727);
and (n3764,n227,n191);
and (n3765,n3766,n3767);
xor (n3766,n3763,n3764);
or (n3767,n3768,n3771);
and (n3768,n3769,n3770);
xor (n3769,n3732,n3733);
and (n3770,n384,n191);
and (n3771,n3772,n3773);
xor (n3772,n3769,n3770);
or (n3773,n3774,n3777);
and (n3774,n3775,n3776);
xor (n3775,n3738,n3739);
and (n3776,n423,n191);
and (n3777,n3778,n3779);
xor (n3778,n3775,n3776);
or (n3779,n3780,n3783);
and (n3780,n3781,n3782);
xor (n3781,n3744,n3745);
and (n3782,n415,n191);
and (n3783,n3784,n3785);
xor (n3784,n3781,n3782);
and (n3785,n3786,n996);
xor (n3786,n3750,n3751);
and (n3787,n236,n218);
or (n3788,n3789,n3792);
and (n3789,n3790,n3791);
xor (n3790,n3760,n3761);
and (n3791,n227,n218);
and (n3792,n3793,n3794);
xor (n3793,n3790,n3791);
or (n3794,n3795,n3798);
and (n3795,n3796,n3797);
xor (n3796,n3766,n3767);
and (n3797,n384,n218);
and (n3798,n3799,n3800);
xor (n3799,n3796,n3797);
or (n3800,n3801,n3804);
and (n3801,n3802,n3803);
xor (n3802,n3772,n3773);
and (n3803,n423,n218);
and (n3804,n3805,n3806);
xor (n3805,n3802,n3803);
or (n3806,n3807,n3810);
and (n3807,n3808,n3809);
xor (n3808,n3778,n3779);
and (n3809,n415,n218);
and (n3810,n3811,n3812);
xor (n3811,n3808,n3809);
and (n3812,n3813,n3814);
xor (n3813,n3784,n3785);
and (n3814,n456,n218);
and (n3815,n227,n395);
or (n3816,n3817,n3820);
and (n3817,n3818,n3819);
xor (n3818,n3793,n3794);
and (n3819,n384,n395);
and (n3820,n3821,n3822);
xor (n3821,n3818,n3819);
or (n3822,n3823,n3826);
and (n3823,n3824,n3825);
xor (n3824,n3799,n3800);
and (n3825,n423,n395);
and (n3826,n3827,n3828);
xor (n3827,n3824,n3825);
or (n3828,n3829,n3832);
and (n3829,n3830,n3831);
xor (n3830,n3805,n3806);
and (n3831,n415,n395);
and (n3832,n3833,n3834);
xor (n3833,n3830,n3831);
and (n3834,n3835,n710);
xor (n3835,n3811,n3812);
and (n3836,n384,n405);
or (n3837,n3838,n3841);
and (n3838,n3839,n3840);
xor (n3839,n3821,n3822);
and (n3840,n423,n405);
and (n3841,n3842,n3843);
xor (n3842,n3839,n3840);
or (n3843,n3844,n3847);
and (n3844,n3845,n3846);
xor (n3845,n3827,n3828);
and (n3846,n415,n405);
and (n3847,n3848,n3849);
xor (n3848,n3845,n3846);
and (n3849,n3850,n3851);
xor (n3850,n3833,n3834);
and (n3851,n456,n405);
and (n3852,n423,n675);
or (n3853,n3854,n3857);
and (n3854,n3855,n3856);
xor (n3855,n3842,n3843);
and (n3856,n415,n675);
and (n3857,n3858,n3859);
xor (n3858,n3855,n3856);
and (n3859,n3860,n694);
xor (n3860,n3848,n3849);
and (n3861,n415,n450);
and (n3862,n3863,n3864);
xor (n3863,n3858,n3859);
and (n3864,n456,n450);
and (n3865,n456,n438);
endmodule
