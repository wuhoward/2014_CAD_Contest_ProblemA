module top (out,n14,n17,n18,n22,n25,n26,n36,n39,n40
        ,n44,n54,n57,n58,n62,n69,n72,n73,n77,n85
        ,n88,n89,n93,n103,n106,n107,n111,n116,n313,n374
        ,n470,n541,n627);
output out;
input n14;
input n17;
input n18;
input n22;
input n25;
input n26;
input n36;
input n39;
input n40;
input n44;
input n54;
input n57;
input n58;
input n62;
input n69;
input n72;
input n73;
input n77;
input n85;
input n88;
input n89;
input n93;
input n103;
input n106;
input n107;
input n111;
input n116;
input n313;
input n374;
input n470;
input n541;
input n627;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
xor (out,n0,n1311);
buf (n0,n1);
xor (n1,n2,n336);
xor (n2,n3,n271);
xor (n3,n4,n231);
or (n4,n5,n207,n230);
and (n5,n6,n178);
or (n6,n7,n150,n177);
and (n7,n8,n118);
or (n8,n9,n98,n117);
and (n9,n10,n49);
or (n10,n11,n32,n48);
and (n11,n12,n19);
not (n12,n13);
and (n13,n14,n15);
not (n15,n16);
and (n16,n17,n18);
xnor (n19,n20,n29);
not (n20,n21);
and (n21,n22,n23);
and (n23,n24,n27);
xor (n24,n25,n26);
not (n27,n28);
xor (n28,n26,n14);
and (n29,n25,n30);
not (n30,n31);
and (n31,n26,n14);
and (n32,n19,n33);
xnor (n33,n34,n45);
nor (n34,n35,n43);
and (n35,n36,n37);
and (n37,n38,n41);
xor (n38,n39,n40);
not (n41,n42);
xor (n42,n40,n25);
and (n43,n44,n42);
and (n45,n39,n46);
not (n46,n47);
and (n47,n40,n25);
and (n48,n12,n33);
or (n49,n50,n81,n97);
and (n50,n51,n66);
xnor (n51,n52,n63);
nor (n52,n53,n61);
and (n53,n54,n55);
and (n55,n56,n59);
xor (n56,n57,n58);
not (n59,n60);
xor (n60,n58,n39);
and (n61,n62,n60);
and (n63,n57,n64);
not (n64,n65);
and (n65,n58,n39);
xnor (n66,n67,n78);
nor (n67,n68,n76);
and (n68,n69,n70);
and (n70,n71,n74);
xor (n71,n72,n73);
not (n74,n75);
xor (n75,n73,n57);
and (n76,n77,n75);
and (n78,n72,n79);
not (n79,n80);
and (n80,n73,n57);
and (n81,n66,n82);
xnor (n82,n83,n94);
nor (n83,n84,n92);
and (n84,n85,n86);
and (n86,n87,n90);
xor (n87,n88,n89);
not (n90,n91);
xor (n91,n89,n72);
and (n92,n93,n91);
and (n94,n88,n95);
not (n95,n96);
and (n96,n89,n72);
and (n97,n51,n82);
and (n98,n49,n99);
and (n99,n100,n115);
xnor (n100,n101,n112);
nor (n101,n102,n110);
and (n102,n103,n104);
and (n104,n105,n108);
xor (n105,n106,n107);
not (n108,n109);
xor (n109,n107,n88);
and (n110,n111,n109);
and (n112,n106,n113);
not (n113,n114);
and (n114,n107,n88);
and (n115,n116,n106);
and (n117,n10,n99);
or (n118,n119,n146,n149);
and (n119,n120,n132);
not (n120,n121);
xor (n121,n122,n128);
xor (n122,n123,n124);
not (n123,n29);
xnor (n124,n125,n45);
nor (n125,n126,n127);
and (n126,n44,n37);
and (n127,n22,n42);
xnor (n128,n129,n63);
nor (n129,n130,n131);
and (n130,n62,n55);
and (n131,n36,n60);
xor (n132,n133,n142);
xor (n133,n134,n138);
xnor (n134,n135,n78);
nor (n135,n136,n137);
and (n136,n77,n70);
and (n137,n54,n75);
xnor (n138,n139,n94);
nor (n139,n140,n141);
and (n140,n93,n86);
and (n141,n69,n91);
xnor (n142,n143,n112);
nor (n143,n144,n145);
and (n144,n111,n104);
and (n145,n85,n109);
and (n146,n132,n147);
not (n147,n148);
and (n148,n103,n106);
and (n149,n120,n147);
and (n150,n118,n151);
xor (n151,n152,n168);
xor (n152,n153,n154);
and (n153,n111,n106);
xor (n154,n155,n164);
xor (n155,n156,n160);
xnor (n156,n157,n78);
nor (n157,n158,n159);
and (n158,n54,n70);
and (n159,n62,n75);
xnor (n160,n161,n94);
nor (n161,n162,n163);
and (n162,n69,n86);
and (n163,n77,n91);
xnor (n164,n165,n112);
nor (n165,n166,n167);
and (n166,n85,n104);
and (n167,n93,n109);
xor (n168,n169,n173);
xor (n169,n123,n170);
xnor (n170,n171,n45);
not (n171,n172);
and (n172,n22,n37);
xnor (n173,n174,n63);
nor (n174,n175,n176);
and (n175,n36,n55);
and (n176,n44,n60);
and (n177,n8,n151);
xor (n178,n179,n196);
xor (n179,n180,n192);
or (n180,n181,n190,n191);
and (n181,n182,n186);
or (n182,n183,n184,n185);
and (n183,n29,n124);
and (n184,n124,n128);
and (n185,n29,n128);
or (n186,n187,n188,n189);
and (n187,n134,n138);
and (n188,n138,n142);
and (n189,n134,n142);
and (n190,n186,n148);
and (n191,n182,n148);
or (n192,n193,n194,n195);
and (n193,n153,n154);
and (n194,n154,n168);
and (n195,n153,n168);
xor (n196,n197,n206);
xor (n197,n198,n202);
xnor (n198,n199,n94);
nor (n199,n200,n201);
and (n200,n77,n86);
and (n201,n54,n91);
xnor (n202,n203,n112);
nor (n203,n204,n205);
and (n204,n93,n104);
and (n205,n69,n109);
and (n206,n85,n106);
and (n207,n178,n208);
xor (n208,n209,n221);
not (n209,n210);
xor (n210,n211,n217);
xor (n211,n212,n213);
not (n212,n45);
xnor (n213,n214,n63);
nor (n214,n215,n216);
and (n215,n44,n55);
and (n216,n22,n60);
xnor (n217,n218,n78);
nor (n218,n219,n220);
and (n219,n62,n70);
and (n220,n36,n75);
xnor (n221,n222,n226);
or (n222,n223,n224,n225);
and (n223,n156,n160);
and (n224,n160,n164);
and (n225,n156,n164);
or (n226,n227,n228,n229);
and (n227,n123,n170);
and (n228,n170,n173);
and (n229,n123,n173);
and (n230,n6,n208);
xor (n231,n232,n238);
xor (n232,n233,n237);
or (n233,n234,n235,n236);
and (n234,n180,n192);
and (n235,n192,n196);
and (n236,n180,n196);
and (n237,n209,n221);
xor (n238,n239,n250);
xor (n239,n240,n241);
or (n240,n222,n226);
xor (n241,n242,n246);
xor (n242,n212,n243);
xnor (n243,n244,n63);
not (n244,n245);
and (n245,n22,n55);
xnor (n246,n247,n78);
nor (n247,n248,n249);
and (n248,n36,n70);
and (n249,n44,n75);
xor (n250,n251,n260);
xor (n251,n252,n256);
or (n252,n253,n254,n255);
and (n253,n198,n202);
and (n254,n202,n206);
and (n255,n198,n206);
or (n256,n257,n258,n259);
and (n257,n45,n213);
and (n258,n213,n217);
and (n259,n45,n217);
xor (n260,n261,n270);
xor (n261,n262,n266);
xnor (n262,n263,n94);
nor (n263,n264,n265);
and (n264,n54,n86);
and (n265,n62,n91);
xnor (n266,n267,n112);
nor (n267,n268,n269);
and (n268,n69,n104);
and (n269,n77,n109);
and (n270,n93,n106);
and (n271,n272,n334);
or (n272,n273,n330,n333);
and (n273,n274,n328);
or (n274,n275,n324,n327);
and (n275,n276,n315);
or (n276,n277,n306,n314);
and (n277,n278,n290);
or (n278,n279,n284,n289);
and (n279,n13,n280);
xnor (n280,n281,n29);
nor (n281,n282,n283);
and (n282,n44,n23);
and (n283,n22,n28);
and (n284,n280,n285);
xnor (n285,n286,n45);
nor (n286,n287,n288);
and (n287,n62,n37);
and (n288,n36,n42);
and (n289,n13,n285);
or (n290,n291,n300,n305);
and (n291,n292,n296);
xnor (n292,n293,n63);
nor (n293,n294,n295);
and (n294,n77,n55);
and (n295,n54,n60);
xnor (n296,n297,n78);
nor (n297,n298,n299);
and (n298,n93,n70);
and (n299,n69,n75);
and (n300,n296,n301);
xnor (n301,n302,n94);
nor (n302,n303,n304);
and (n303,n111,n86);
and (n304,n85,n91);
and (n305,n292,n301);
and (n306,n290,n307);
or (n307,n308,n312);
xnor (n308,n309,n112);
nor (n309,n310,n311);
and (n310,n116,n104);
and (n311,n103,n109);
and (n312,n313,n106);
and (n314,n278,n307);
or (n315,n316,n321,n323);
and (n316,n317,n319);
xor (n317,n318,n33);
xor (n318,n12,n19);
xor (n319,n320,n82);
xor (n320,n51,n66);
and (n321,n319,n322);
xor (n322,n100,n115);
and (n323,n317,n322);
and (n324,n315,n325);
xor (n325,n326,n132);
xor (n326,n148,n121);
and (n327,n276,n325);
xor (n328,n329,n148);
xor (n329,n182,n186);
and (n330,n328,n331);
xor (n331,n332,n151);
xor (n332,n8,n118);
and (n333,n274,n331);
xor (n334,n335,n208);
xor (n335,n6,n178);
or (n336,n337,n417);
and (n337,n338,n339);
xor (n338,n272,n334);
and (n339,n340,n415);
or (n340,n341,n411,n414);
and (n341,n342,n409);
or (n342,n343,n405,n408);
and (n343,n344,n394);
or (n344,n345,n376,n393);
and (n345,n346,n362);
or (n346,n347,n356,n361);
and (n347,n348,n349);
not (n348,n18);
xnor (n349,n350,n13);
not (n350,n351);
and (n351,n22,n352);
and (n352,n353,n354);
xor (n353,n14,n17);
not (n354,n355);
xor (n355,n17,n18);
and (n356,n349,n357);
xnor (n357,n358,n29);
nor (n358,n359,n360);
and (n359,n36,n23);
and (n360,n44,n28);
and (n361,n348,n357);
or (n362,n363,n372,n375);
and (n363,n364,n368);
xnor (n364,n365,n94);
nor (n365,n366,n367);
and (n366,n103,n86);
and (n367,n111,n91);
xnor (n368,n369,n112);
nor (n369,n370,n371);
and (n370,n313,n104);
and (n371,n116,n109);
and (n372,n368,n373);
and (n373,n374,n106);
and (n375,n364,n373);
and (n376,n362,n377);
or (n377,n378,n387,n392);
and (n378,n379,n383);
xnor (n379,n380,n45);
nor (n380,n381,n382);
and (n381,n54,n37);
and (n382,n62,n42);
xnor (n383,n384,n63);
nor (n384,n385,n386);
and (n385,n69,n55);
and (n386,n77,n60);
and (n387,n383,n388);
xnor (n388,n389,n78);
nor (n389,n390,n391);
and (n390,n85,n70);
and (n391,n93,n75);
and (n392,n379,n388);
and (n393,n346,n377);
or (n394,n395,n401,n404);
and (n395,n396,n399);
not (n396,n397);
xor (n397,n398,n285);
xor (n398,n12,n280);
xor (n399,n400,n301);
xor (n400,n292,n296);
and (n401,n399,n402);
not (n402,n403);
xor (n403,n308,n312);
and (n404,n396,n402);
and (n405,n394,n406);
xor (n406,n407,n322);
xor (n407,n317,n319);
and (n408,n344,n406);
xor (n409,n410,n99);
xor (n410,n10,n49);
and (n411,n409,n412);
xor (n412,n413,n325);
xor (n413,n276,n315);
and (n414,n342,n412);
xor (n415,n416,n331);
xor (n416,n274,n328);
and (n417,n418,n419);
xor (n418,n338,n339);
or (n419,n420,n490);
and (n420,n421,n422);
xor (n421,n340,n415);
and (n422,n423,n488);
or (n423,n424,n484,n487);
and (n424,n425,n482);
or (n425,n426,n478,n481);
and (n426,n427,n473);
or (n427,n428,n457,n472);
and (n428,n429,n445);
or (n429,n430,n439,n444);
and (n430,n431,n435);
xnor (n431,n432,n45);
nor (n432,n433,n434);
and (n433,n77,n37);
and (n434,n54,n42);
xnor (n435,n436,n63);
nor (n436,n437,n438);
and (n437,n93,n55);
and (n438,n69,n60);
and (n439,n435,n440);
xnor (n440,n441,n78);
nor (n441,n442,n443);
and (n442,n111,n70);
and (n443,n85,n75);
and (n444,n431,n440);
or (n445,n446,n451,n456);
and (n446,n18,n447);
xnor (n447,n448,n13);
nor (n448,n449,n450);
and (n449,n44,n352);
and (n450,n22,n355);
and (n451,n447,n452);
xnor (n452,n453,n29);
nor (n453,n454,n455);
and (n454,n62,n23);
and (n455,n36,n28);
and (n456,n18,n452);
and (n457,n445,n458);
or (n458,n459,n468,n471);
and (n459,n460,n464);
xnor (n460,n461,n94);
nor (n461,n462,n463);
and (n462,n116,n86);
and (n463,n103,n91);
xnor (n464,n465,n112);
nor (n465,n466,n467);
and (n466,n374,n104);
and (n467,n313,n109);
and (n468,n464,n469);
and (n469,n470,n106);
and (n471,n460,n469);
and (n472,n429,n458);
or (n473,n474,n476);
xor (n474,n475,n373);
xor (n475,n364,n368);
xor (n476,n477,n388);
xor (n477,n379,n383);
and (n478,n473,n479);
xor (n479,n480,n403);
xor (n480,n397,n399);
and (n481,n427,n479);
xor (n482,n483,n307);
xor (n483,n278,n290);
and (n484,n482,n485);
xor (n485,n486,n406);
xor (n486,n344,n394);
and (n487,n425,n485);
xor (n488,n489,n412);
xor (n489,n342,n409);
and (n490,n491,n492);
xor (n491,n421,n422);
or (n492,n493,n573);
and (n493,n494,n495);
xor (n494,n423,n488);
and (n495,n496,n571);
or (n496,n497,n567,n570);
and (n497,n498,n563);
or (n498,n499,n559,n562);
and (n499,n500,n548);
or (n500,n501,n534,n547);
and (n501,n502,n518);
or (n502,n503,n512,n517);
and (n503,n504,n508);
xnor (n504,n505,n29);
nor (n505,n506,n507);
and (n506,n54,n23);
and (n507,n62,n28);
xnor (n508,n509,n45);
nor (n509,n510,n511);
and (n510,n69,n37);
and (n511,n77,n42);
and (n512,n508,n513);
xnor (n513,n514,n63);
nor (n514,n515,n516);
and (n515,n85,n55);
and (n516,n93,n60);
and (n517,n504,n513);
or (n518,n519,n528,n533);
and (n519,n520,n524);
xnor (n520,n521,n78);
nor (n521,n522,n523);
and (n522,n103,n70);
and (n523,n111,n75);
xnor (n524,n525,n94);
nor (n525,n526,n527);
and (n526,n313,n86);
and (n527,n116,n91);
and (n528,n524,n529);
xnor (n529,n530,n112);
nor (n530,n531,n532);
and (n531,n470,n104);
and (n532,n374,n109);
and (n533,n520,n529);
and (n534,n518,n535);
and (n535,n536,n543);
xnor (n536,n537,n18);
not (n537,n538);
and (n538,n22,n539);
and (n539,n540,n542);
xor (n540,n18,n541);
not (n542,n541);
xnor (n543,n544,n13);
nor (n544,n545,n546);
and (n545,n36,n352);
and (n546,n44,n355);
and (n547,n502,n535);
or (n548,n549,n555,n558);
and (n549,n550,n552);
xor (n550,n551,n440);
xor (n551,n431,n435);
not (n552,n553);
xor (n553,n554,n452);
xor (n554,n348,n447);
and (n555,n552,n556);
xor (n556,n557,n469);
xor (n557,n460,n464);
and (n558,n550,n556);
and (n559,n548,n560);
xor (n560,n561,n357);
xor (n561,n348,n349);
and (n562,n500,n560);
and (n563,n564,n566);
xor (n564,n565,n458);
xor (n565,n429,n445);
xnor (n566,n474,n476);
and (n567,n563,n568);
xor (n568,n569,n377);
xor (n569,n346,n362);
and (n570,n498,n568);
xor (n571,n572,n485);
xor (n572,n425,n482);
and (n573,n574,n575);
xor (n574,n494,n495);
or (n575,n576,n655);
and (n576,n577,n578);
xor (n577,n496,n571);
or (n578,n579,n651,n654);
and (n579,n580,n649);
or (n580,n581,n646,n648);
and (n581,n582,n644);
or (n582,n583,n640,n643);
and (n583,n584,n630);
or (n584,n585,n618,n629);
and (n585,n586,n602);
or (n586,n587,n596,n601);
and (n587,n588,n592);
xnor (n588,n589,n18);
nor (n589,n590,n591);
and (n590,n44,n539);
and (n591,n22,n541);
xnor (n592,n593,n13);
nor (n593,n594,n595);
and (n594,n62,n352);
and (n595,n36,n355);
and (n596,n592,n597);
xnor (n597,n598,n29);
nor (n598,n599,n600);
and (n599,n77,n23);
and (n600,n54,n28);
and (n601,n588,n597);
or (n602,n603,n612,n617);
and (n603,n604,n608);
xnor (n604,n605,n45);
nor (n605,n606,n607);
and (n606,n93,n37);
and (n607,n69,n42);
xnor (n608,n609,n63);
nor (n609,n610,n611);
and (n610,n111,n55);
and (n611,n85,n60);
and (n612,n608,n613);
xnor (n613,n614,n78);
nor (n614,n615,n616);
and (n615,n116,n70);
and (n616,n103,n75);
and (n617,n604,n613);
and (n618,n602,n619);
and (n619,n620,n624);
xnor (n620,n621,n94);
nor (n621,n622,n623);
and (n622,n374,n86);
and (n623,n313,n91);
xnor (n624,n625,n112);
nor (n625,n626,n628);
and (n626,n627,n104);
and (n628,n470,n109);
and (n629,n586,n619);
or (n630,n631,n636,n639);
and (n631,n632,n634);
not (n632,n633);
nand (n633,n627,n106);
xor (n634,n635,n513);
xor (n635,n504,n508);
and (n636,n634,n637);
xor (n637,n638,n529);
xor (n638,n520,n524);
and (n639,n632,n637);
and (n640,n630,n641);
xor (n641,n642,n556);
xor (n642,n550,n552);
and (n643,n584,n641);
xor (n644,n645,n560);
xor (n645,n500,n548);
and (n646,n644,n647);
xor (n647,n564,n566);
and (n648,n582,n647);
xor (n649,n650,n568);
xor (n650,n498,n563);
and (n651,n649,n652);
xor (n652,n653,n479);
xor (n653,n427,n473);
and (n654,n580,n652);
and (n655,n656,n657);
xor (n656,n577,n578);
or (n657,n658,n735);
and (n658,n659,n661);
xor (n659,n660,n652);
xor (n660,n580,n649);
and (n661,n662,n733);
or (n662,n663,n729,n732);
and (n663,n664,n724);
or (n664,n665,n721,n723);
and (n665,n666,n712);
or (n666,n667,n694,n711);
and (n667,n668,n682);
or (n668,n669,n678,n681);
and (n669,n670,n674);
xnor (n670,n671,n78);
nor (n671,n672,n673);
and (n672,n313,n70);
and (n673,n116,n75);
xnor (n674,n675,n94);
nor (n675,n676,n677);
and (n676,n470,n86);
and (n677,n374,n91);
and (n678,n674,n679);
xnor (n679,n680,n112);
nand (n680,n627,n109);
and (n681,n670,n679);
or (n682,n683,n692,n693);
and (n683,n684,n688);
xnor (n684,n685,n18);
nor (n685,n686,n687);
and (n686,n36,n539);
and (n687,n44,n541);
xnor (n688,n689,n13);
nor (n689,n690,n691);
and (n690,n54,n352);
and (n691,n62,n355);
and (n692,n688,n112);
and (n693,n684,n112);
and (n694,n682,n695);
or (n695,n696,n705,n710);
and (n696,n697,n701);
xnor (n697,n698,n29);
nor (n698,n699,n700);
and (n699,n69,n23);
and (n700,n77,n28);
xnor (n701,n702,n45);
nor (n702,n703,n704);
and (n703,n85,n37);
and (n704,n93,n42);
and (n705,n701,n706);
xnor (n706,n707,n63);
nor (n707,n708,n709);
and (n708,n103,n55);
and (n709,n111,n60);
and (n710,n697,n706);
and (n711,n668,n695);
or (n712,n713,n718,n720);
and (n713,n714,n716);
xor (n714,n715,n597);
xor (n715,n588,n592);
xor (n716,n717,n613);
xor (n717,n604,n608);
and (n718,n716,n719);
xor (n719,n620,n624);
and (n720,n714,n719);
and (n721,n712,n722);
xor (n722,n536,n543);
and (n723,n666,n722);
and (n724,n725,n727);
xor (n725,n726,n619);
xor (n726,n586,n602);
xor (n727,n728,n637);
xor (n728,n632,n634);
and (n729,n724,n730);
xor (n730,n731,n535);
xor (n731,n502,n518);
and (n732,n664,n730);
xor (n733,n734,n647);
xor (n734,n582,n644);
and (n735,n736,n737);
xor (n736,n659,n661);
or (n737,n738,n745);
and (n738,n739,n740);
xor (n739,n662,n733);
and (n740,n741,n743);
xor (n741,n742,n730);
xor (n742,n664,n724);
xor (n743,n744,n641);
xor (n744,n584,n630);
and (n745,n746,n778);
xor (n746,n747,n772);
xor (n747,n748,n752);
or (n748,n663,n749,n751);
and (n749,n724,n750);
xnor (n750,n550,n556);
and (n751,n664,n750);
xor (n752,n753,n762);
xor (n753,n754,n757);
or (n754,n583,n755,n756);
and (n755,n630,n553);
and (n756,n584,n553);
xor (n757,n758,n458);
xor (n758,n429,n759);
or (n759,n760,n451,n761);
and (n760,n348,n447);
and (n761,n348,n452);
xor (n762,n763,n765);
xor (n763,n500,n764);
or (n764,n550,n556);
xor (n765,n766,n771);
xor (n766,n767,n769);
xor (n767,n768,n379);
xor (n768,n349,n357);
xor (n769,n770,n364);
xor (n770,n383,n388);
xnor (n771,n368,n373);
or (n772,n773,n775,n777);
and (n773,n730,n774);
xor (n774,n744,n553);
and (n775,n774,n776);
xor (n776,n742,n750);
and (n777,n730,n776);
or (n778,n779,n838);
and (n779,n780,n782);
xor (n780,n781,n776);
xor (n781,n730,n774);
or (n782,n783,n835,n837);
and (n783,n784,n833);
or (n784,n785,n829,n832);
and (n785,n786,n824);
or (n786,n787,n820,n823);
and (n787,n788,n804);
or (n788,n789,n798,n803);
and (n789,n790,n794);
xnor (n790,n791,n18);
nor (n791,n792,n793);
and (n792,n62,n539);
and (n793,n36,n541);
xnor (n794,n795,n13);
nor (n795,n796,n797);
and (n796,n77,n352);
and (n797,n54,n355);
and (n798,n794,n799);
xnor (n799,n800,n29);
nor (n800,n801,n802);
and (n801,n93,n23);
and (n802,n69,n28);
and (n803,n790,n799);
or (n804,n805,n814,n819);
and (n805,n806,n810);
xnor (n806,n807,n45);
nor (n807,n808,n809);
and (n808,n111,n37);
and (n809,n85,n42);
xnor (n810,n811,n63);
nor (n811,n812,n813);
and (n812,n116,n55);
and (n813,n103,n60);
and (n814,n810,n815);
xnor (n815,n816,n78);
nor (n816,n817,n818);
and (n817,n374,n70);
and (n818,n313,n75);
and (n819,n806,n815);
and (n820,n804,n821);
xor (n821,n822,n679);
xor (n822,n670,n674);
and (n823,n788,n821);
and (n824,n825,n827);
xor (n825,n826,n112);
xor (n826,n684,n688);
xor (n827,n828,n706);
xor (n828,n697,n701);
and (n829,n824,n830);
xor (n830,n831,n719);
xor (n831,n714,n716);
and (n832,n786,n830);
xor (n833,n834,n722);
xor (n834,n666,n712);
and (n835,n833,n836);
xor (n836,n725,n727);
and (n837,n784,n836);
and (n838,n839,n840);
xor (n839,n780,n782);
or (n840,n841,n895);
and (n841,n842,n844);
xor (n842,n843,n836);
xor (n843,n784,n833);
or (n844,n845,n891,n894);
and (n845,n846,n889);
or (n846,n847,n886,n888);
and (n847,n848,n884);
or (n848,n849,n878,n883);
and (n849,n850,n862);
or (n850,n851,n860,n861);
and (n851,n852,n856);
xnor (n852,n853,n18);
nor (n853,n854,n855);
and (n854,n54,n539);
and (n855,n62,n541);
xnor (n856,n857,n13);
nor (n857,n858,n859);
and (n858,n69,n352);
and (n859,n77,n355);
and (n860,n856,n94);
and (n861,n852,n94);
or (n862,n863,n872,n877);
and (n863,n864,n868);
xnor (n864,n865,n29);
nor (n865,n866,n867);
and (n866,n85,n23);
and (n867,n93,n28);
xnor (n868,n869,n45);
nor (n869,n870,n871);
and (n870,n103,n37);
and (n871,n111,n42);
and (n872,n868,n873);
xnor (n873,n874,n63);
nor (n874,n875,n876);
and (n875,n313,n55);
and (n876,n116,n60);
and (n877,n864,n873);
and (n878,n862,n879);
xnor (n879,n880,n94);
nor (n880,n881,n882);
and (n881,n627,n86);
and (n882,n470,n91);
and (n883,n850,n879);
xor (n884,n885,n821);
xor (n885,n788,n804);
and (n886,n884,n887);
xor (n887,n825,n827);
and (n888,n848,n887);
xor (n889,n890,n695);
xor (n890,n668,n682);
and (n891,n889,n892);
xor (n892,n893,n830);
xor (n893,n786,n824);
and (n894,n846,n892);
and (n895,n896,n897);
xor (n896,n842,n844);
or (n897,n898,n968);
and (n898,n899,n901);
xor (n899,n900,n892);
xor (n900,n846,n889);
or (n901,n902,n964,n967);
and (n902,n903,n959);
or (n903,n904,n955,n958);
and (n904,n905,n945);
or (n905,n906,n939,n944);
and (n906,n907,n923);
or (n907,n908,n917,n922);
and (n908,n909,n913);
xnor (n909,n910,n45);
nor (n910,n911,n912);
and (n911,n116,n37);
and (n912,n103,n42);
xnor (n913,n914,n63);
nor (n914,n915,n916);
and (n915,n374,n55);
and (n916,n313,n60);
and (n917,n913,n918);
xnor (n918,n919,n78);
nor (n919,n920,n921);
and (n920,n627,n70);
and (n921,n470,n75);
and (n922,n909,n918);
or (n923,n924,n933,n938);
and (n924,n925,n929);
xnor (n925,n926,n18);
nor (n926,n927,n928);
and (n927,n77,n539);
and (n928,n54,n541);
xnor (n929,n930,n13);
nor (n930,n931,n932);
and (n931,n93,n352);
and (n932,n69,n355);
and (n933,n929,n934);
xnor (n934,n935,n29);
nor (n935,n936,n937);
and (n936,n111,n23);
and (n937,n85,n28);
and (n938,n925,n934);
and (n939,n923,n940);
xnor (n940,n941,n78);
nor (n941,n942,n943);
and (n942,n470,n70);
and (n943,n374,n75);
and (n944,n907,n940);
or (n945,n946,n951,n954);
and (n946,n947,n949);
xnor (n947,n948,n94);
nand (n948,n627,n91);
xor (n949,n950,n94);
xor (n950,n852,n856);
and (n951,n949,n952);
xor (n952,n953,n873);
xor (n953,n864,n868);
and (n954,n947,n952);
and (n955,n945,n956);
xor (n956,n957,n815);
xor (n957,n806,n810);
and (n958,n905,n956);
and (n959,n960,n962);
xor (n960,n961,n799);
xor (n961,n790,n794);
xor (n962,n963,n879);
xor (n963,n850,n862);
and (n964,n959,n965);
xor (n965,n966,n887);
xor (n966,n848,n884);
and (n967,n903,n965);
and (n968,n969,n970);
xor (n969,n899,n901);
or (n970,n971,n1023);
and (n971,n972,n974);
xor (n972,n973,n965);
xor (n973,n903,n959);
or (n974,n975,n1020,n1022);
and (n975,n976,n1018);
or (n976,n977,n1014,n1017);
and (n977,n978,n1012);
or (n978,n979,n1008,n1011);
and (n979,n980,n996);
or (n980,n981,n990,n995);
and (n981,n982,n986);
xnor (n982,n983,n29);
nor (n983,n984,n985);
and (n984,n103,n23);
and (n985,n111,n28);
xnor (n986,n987,n45);
nor (n987,n988,n989);
and (n988,n313,n37);
and (n989,n116,n42);
and (n990,n986,n991);
xnor (n991,n992,n63);
nor (n992,n993,n994);
and (n993,n470,n55);
and (n994,n374,n60);
and (n995,n982,n991);
or (n996,n997,n1006,n1007);
and (n997,n998,n1002);
xnor (n998,n999,n18);
nor (n999,n1000,n1001);
and (n1000,n69,n539);
and (n1001,n77,n541);
xnor (n1002,n1003,n13);
nor (n1003,n1004,n1005);
and (n1004,n85,n352);
and (n1005,n93,n355);
and (n1006,n1002,n78);
and (n1007,n998,n78);
and (n1008,n996,n1009);
xor (n1009,n1010,n918);
xor (n1010,n909,n913);
and (n1011,n980,n1009);
xor (n1012,n1013,n940);
xor (n1013,n907,n923);
and (n1014,n1012,n1015);
xor (n1015,n1016,n952);
xor (n1016,n947,n949);
and (n1017,n978,n1015);
xor (n1018,n1019,n956);
xor (n1019,n905,n945);
and (n1020,n1018,n1021);
xor (n1021,n960,n962);
and (n1022,n976,n1021);
and (n1023,n1024,n1025);
xor (n1024,n972,n974);
or (n1025,n1026,n1064);
and (n1026,n1027,n1029);
xor (n1027,n1028,n1021);
xor (n1028,n976,n1018);
and (n1029,n1030,n1062);
or (n1030,n1031,n1058,n1061);
and (n1031,n1032,n1056);
or (n1032,n1033,n1052,n1055);
and (n1033,n1034,n1050);
or (n1034,n1035,n1044,n1049);
and (n1035,n1036,n1040);
xnor (n1036,n1037,n18);
nor (n1037,n1038,n1039);
and (n1038,n93,n539);
and (n1039,n69,n541);
xnor (n1040,n1041,n13);
nor (n1041,n1042,n1043);
and (n1042,n111,n352);
and (n1043,n85,n355);
and (n1044,n1040,n1045);
xnor (n1045,n1046,n29);
nor (n1046,n1047,n1048);
and (n1047,n116,n23);
and (n1048,n103,n28);
and (n1049,n1036,n1045);
xnor (n1050,n1051,n78);
nand (n1051,n627,n75);
and (n1052,n1050,n1053);
xor (n1053,n1054,n991);
xor (n1054,n982,n986);
and (n1055,n1034,n1053);
xor (n1056,n1057,n934);
xor (n1057,n925,n929);
and (n1058,n1056,n1059);
xor (n1059,n1060,n1009);
xor (n1060,n980,n996);
and (n1061,n1032,n1059);
xor (n1062,n1063,n1015);
xor (n1063,n978,n1012);
and (n1064,n1065,n1066);
xor (n1065,n1027,n1029);
or (n1066,n1067,n1119);
and (n1067,n1068,n1069);
xor (n1068,n1030,n1062);
and (n1069,n1070,n1117);
or (n1070,n1071,n1113,n1116);
and (n1071,n1072,n1106);
or (n1072,n1073,n1100,n1105);
and (n1073,n1074,n1088);
or (n1074,n1075,n1084,n1087);
and (n1075,n1076,n1080);
xnor (n1076,n1077,n29);
nor (n1077,n1078,n1079);
and (n1078,n313,n23);
and (n1079,n116,n28);
xnor (n1080,n1081,n45);
nor (n1081,n1082,n1083);
and (n1082,n470,n37);
and (n1083,n374,n42);
and (n1084,n1080,n1085);
xnor (n1085,n1086,n63);
nand (n1086,n627,n60);
and (n1087,n1076,n1085);
or (n1088,n1089,n1098,n1099);
and (n1089,n1090,n1094);
xnor (n1090,n1091,n18);
nor (n1091,n1092,n1093);
and (n1092,n85,n539);
and (n1093,n93,n541);
xnor (n1094,n1095,n13);
nor (n1095,n1096,n1097);
and (n1096,n103,n352);
and (n1097,n111,n355);
and (n1098,n1094,n63);
and (n1099,n1090,n63);
and (n1100,n1088,n1101);
xnor (n1101,n1102,n45);
nor (n1102,n1103,n1104);
and (n1103,n374,n37);
and (n1104,n313,n42);
and (n1105,n1074,n1101);
and (n1106,n1107,n1111);
xnor (n1107,n1108,n63);
nor (n1108,n1109,n1110);
and (n1109,n627,n55);
and (n1110,n470,n60);
xor (n1111,n1112,n1045);
xor (n1112,n1036,n1040);
and (n1113,n1106,n1114);
xor (n1114,n1115,n78);
xor (n1115,n998,n1002);
and (n1116,n1072,n1114);
xor (n1117,n1118,n1059);
xor (n1118,n1032,n1056);
and (n1119,n1120,n1121);
xor (n1120,n1068,n1069);
or (n1121,n1122,n1129);
and (n1122,n1123,n1124);
xor (n1123,n1070,n1117);
and (n1124,n1125,n1127);
xor (n1125,n1126,n1053);
xor (n1126,n1034,n1050);
xor (n1127,n1128,n1114);
xor (n1128,n1072,n1106);
and (n1129,n1130,n1131);
xor (n1130,n1123,n1124);
or (n1131,n1132,n1165);
and (n1132,n1133,n1134);
xor (n1133,n1125,n1127);
or (n1134,n1135,n1162,n1164);
and (n1135,n1136,n1160);
or (n1136,n1137,n1156,n1159);
and (n1137,n1138,n1154);
or (n1138,n1139,n1148,n1153);
and (n1139,n1140,n1144);
xnor (n1140,n1141,n18);
nor (n1141,n1142,n1143);
and (n1142,n111,n539);
and (n1143,n85,n541);
xnor (n1144,n1145,n13);
nor (n1145,n1146,n1147);
and (n1146,n116,n352);
and (n1147,n103,n355);
and (n1148,n1144,n1149);
xnor (n1149,n1150,n29);
nor (n1150,n1151,n1152);
and (n1151,n374,n23);
and (n1152,n313,n28);
and (n1153,n1140,n1149);
xor (n1154,n1155,n1085);
xor (n1155,n1076,n1080);
and (n1156,n1154,n1157);
xor (n1157,n1158,n63);
xor (n1158,n1090,n1094);
and (n1159,n1138,n1157);
xor (n1160,n1161,n1101);
xor (n1161,n1074,n1088);
and (n1162,n1160,n1163);
xor (n1163,n1107,n1111);
and (n1164,n1136,n1163);
and (n1165,n1166,n1167);
xor (n1166,n1133,n1134);
or (n1167,n1168,n1201);
and (n1168,n1169,n1171);
xor (n1169,n1170,n1163);
xor (n1170,n1136,n1160);
and (n1171,n1172,n1199);
or (n1172,n1173,n1193,n1198);
and (n1173,n1174,n1186);
or (n1174,n1175,n1184,n1185);
and (n1175,n1176,n1180);
xnor (n1176,n1177,n18);
nor (n1177,n1178,n1179);
and (n1178,n103,n539);
and (n1179,n111,n541);
xnor (n1180,n1181,n13);
nor (n1181,n1182,n1183);
and (n1182,n313,n352);
and (n1183,n116,n355);
and (n1184,n1180,n45);
and (n1185,n1176,n45);
and (n1186,n1187,n1191);
xnor (n1187,n1188,n29);
nor (n1188,n1189,n1190);
and (n1189,n470,n23);
and (n1190,n374,n28);
xnor (n1191,n1192,n45);
nand (n1192,n627,n42);
and (n1193,n1186,n1194);
xnor (n1194,n1195,n45);
nor (n1195,n1196,n1197);
and (n1196,n627,n37);
and (n1197,n470,n42);
and (n1198,n1174,n1194);
xor (n1199,n1200,n1157);
xor (n1200,n1138,n1154);
and (n1201,n1202,n1203);
xor (n1202,n1169,n1171);
or (n1203,n1204,n1211);
and (n1204,n1205,n1206);
xor (n1205,n1172,n1199);
and (n1206,n1207,n1209);
xor (n1207,n1208,n1149);
xor (n1208,n1140,n1144);
xor (n1209,n1210,n1194);
xor (n1210,n1174,n1186);
and (n1211,n1212,n1213);
xor (n1212,n1205,n1206);
or (n1213,n1214,n1239);
and (n1214,n1215,n1216);
xor (n1215,n1207,n1209);
or (n1216,n1217,n1236,n1238);
and (n1217,n1218,n1234);
or (n1218,n1219,n1228,n1233);
and (n1219,n1220,n1224);
xnor (n1220,n1221,n18);
nor (n1221,n1222,n1223);
and (n1222,n116,n539);
and (n1223,n103,n541);
xnor (n1224,n1225,n13);
nor (n1225,n1226,n1227);
and (n1226,n374,n352);
and (n1227,n313,n355);
and (n1228,n1224,n1229);
xnor (n1229,n1230,n29);
nor (n1230,n1231,n1232);
and (n1231,n627,n23);
and (n1232,n470,n28);
and (n1233,n1220,n1229);
xor (n1234,n1235,n45);
xor (n1235,n1176,n1180);
and (n1236,n1234,n1237);
xor (n1237,n1187,n1191);
and (n1238,n1218,n1237);
and (n1239,n1240,n1241);
xor (n1240,n1215,n1216);
or (n1241,n1242,n1260);
and (n1242,n1243,n1245);
xor (n1243,n1244,n1237);
xor (n1244,n1218,n1234);
and (n1245,n1246,n1258);
or (n1246,n1247,n1256,n1257);
and (n1247,n1248,n1252);
xnor (n1248,n1249,n18);
nor (n1249,n1250,n1251);
and (n1250,n313,n539);
and (n1251,n116,n541);
xnor (n1252,n1253,n13);
nor (n1253,n1254,n1255);
and (n1254,n470,n352);
and (n1255,n374,n355);
and (n1256,n1252,n29);
and (n1257,n1248,n29);
xor (n1258,n1259,n1229);
xor (n1259,n1220,n1224);
and (n1260,n1261,n1262);
xor (n1261,n1243,n1245);
or (n1262,n1263,n1270);
and (n1263,n1264,n1265);
xor (n1264,n1246,n1258);
and (n1265,n1266,n1268);
xnor (n1266,n1267,n29);
nand (n1267,n627,n28);
xor (n1268,n1269,n29);
xor (n1269,n1248,n1252);
and (n1270,n1271,n1272);
xor (n1271,n1264,n1265);
or (n1272,n1273,n1284);
and (n1273,n1274,n1275);
xor (n1274,n1266,n1268);
and (n1275,n1276,n1280);
xnor (n1276,n1277,n18);
nor (n1277,n1278,n1279);
and (n1278,n374,n539);
and (n1279,n313,n541);
xnor (n1280,n1281,n13);
nor (n1281,n1282,n1283);
and (n1282,n627,n352);
and (n1283,n470,n355);
and (n1284,n1285,n1286);
xor (n1285,n1274,n1275);
or (n1286,n1287,n1294);
and (n1287,n1288,n1289);
xor (n1288,n1276,n1280);
and (n1289,n1290,n13);
xnor (n1290,n1291,n18);
nor (n1291,n1292,n1293);
and (n1292,n470,n539);
and (n1293,n374,n541);
and (n1294,n1295,n1296);
xor (n1295,n1288,n1289);
or (n1296,n1297,n1301);
and (n1297,n1298,n1300);
xnor (n1298,n1299,n13);
nand (n1299,n627,n355);
xor (n1300,n1290,n13);
and (n1301,n1302,n1303);
xor (n1302,n1298,n1300);
and (n1303,n1304,n1308);
xnor (n1304,n1305,n18);
nor (n1305,n1306,n1307);
and (n1306,n627,n539);
and (n1307,n470,n541);
and (n1308,n1309,n18);
xnor (n1309,n1310,n18);
nand (n1310,n627,n541);
buf (n1311,n1312);
xor (n1312,n1313,n1408);
xor (n1313,n1314,n1377);
xor (n1314,n1315,n1363);
xor (n1315,n1316,n1332);
or (n1316,n1317,n1322,n1331);
and (n1317,n1318,n210);
or (n1318,n1319,n186);
or (n1319,n1320,n184,n1321);
and (n1320,n123,n124);
and (n1321,n123,n128);
and (n1322,n210,n1323);
xor (n1323,n1324,n196);
xor (n1324,n1325,n1328);
or (n1325,n224,n1326,n1327);
and (n1326,n164,n153);
and (n1327,n160,n153);
or (n1328,n228,n1329,n1330);
and (n1329,n173,n156);
and (n1330,n170,n156);
and (n1331,n1318,n1323);
or (n1332,n1333,n1359,n1362);
and (n1333,n1334,n1355);
or (n1334,n1335,n1351,n1354);
and (n1335,n1336,n1347);
or (n1336,n1337,n1344,n1346);
and (n1337,n1338,n1341);
or (n1338,n32,n1339,n1340);
and (n1339,n33,n51);
and (n1340,n19,n51);
or (n1341,n81,n1342,n1343);
and (n1342,n82,n100);
and (n1343,n66,n100);
and (n1344,n1341,n1345);
buf (n1345,n115);
and (n1346,n1338,n1345);
or (n1347,n1348,n1349,n1350);
and (n1348,n148,n121);
and (n1349,n121,n132);
and (n1350,n148,n132);
and (n1351,n1347,n1352);
xor (n1352,n1353,n153);
xor (n1353,n160,n164);
and (n1354,n1336,n1352);
and (n1355,n1356,n1358);
xor (n1356,n1357,n156);
xor (n1357,n170,n173);
xnor (n1358,n1319,n186);
and (n1359,n1355,n1360);
xor (n1360,n1361,n1323);
xor (n1361,n1318,n210);
and (n1362,n1334,n1360);
xor (n1363,n1364,n1371);
xor (n1364,n1365,n1369);
or (n1365,n1366,n1367,n1368);
and (n1366,n1325,n1328);
and (n1367,n1328,n196);
and (n1368,n1325,n196);
xor (n1369,n1370,n262);
xor (n1370,n243,n246);
xor (n1371,n1372,n1376);
xor (n1372,n252,n1373);
or (n1373,n1374,n258,n1375);
and (n1374,n212,n213);
and (n1375,n212,n217);
xnor (n1376,n266,n270);
and (n1377,n1378,n1406);
or (n1378,n1379,n1403,n1405);
and (n1379,n1380,n1401);
or (n1380,n1381,n1399,n1400);
and (n1381,n1382,n1390);
or (n1382,n1383,n1387,n1389);
and (n1383,n1384,n290);
or (n1384,n1385,n284,n1386);
and (n1385,n12,n280);
and (n1386,n12,n285);
and (n1387,n290,n1388);
and (n1388,n308,n312);
and (n1389,n1384,n1388);
or (n1390,n1391,n1396,n1398);
and (n1391,n1392,n1394);
xor (n1392,n1393,n51);
xor (n1393,n19,n33);
xor (n1394,n1395,n100);
xor (n1395,n66,n82);
and (n1396,n1394,n1397);
not (n1397,n115);
and (n1398,n1392,n1397);
and (n1399,n1390,n325);
and (n1400,n1382,n325);
xor (n1401,n1402,n1352);
xor (n1402,n1336,n1347);
and (n1403,n1401,n1404);
xor (n1404,n1356,n1358);
and (n1405,n1380,n1404);
xor (n1406,n1407,n1360);
xor (n1407,n1334,n1355);
or (n1408,n1409,n1443);
and (n1409,n1410,n1411);
xor (n1410,n1378,n1406);
and (n1411,n1412,n1441);
or (n1412,n1413,n1437,n1440);
and (n1413,n1414,n1435);
or (n1414,n1415,n1431,n1434);
and (n1415,n1416,n1427);
or (n1416,n1417,n1424,n1426);
and (n1417,n1418,n1421);
or (n1418,n356,n1419,n1420);
and (n1419,n357,n379);
and (n1420,n349,n379);
or (n1421,n387,n1422,n1423);
and (n1422,n388,n364);
and (n1423,n383,n364);
and (n1424,n1421,n1425);
or (n1425,n368,n373);
and (n1426,n1418,n1425);
or (n1427,n1428,n1429,n1430);
and (n1428,n397,n399);
and (n1429,n399,n403);
and (n1430,n397,n403);
and (n1431,n1427,n1432);
xor (n1432,n1433,n1397);
xor (n1433,n1392,n1394);
and (n1434,n1416,n1432);
xor (n1435,n1436,n1345);
xor (n1436,n1338,n1341);
and (n1437,n1435,n1438);
xor (n1438,n1439,n325);
xor (n1439,n1382,n1390);
and (n1440,n1414,n1438);
xor (n1441,n1442,n1404);
xor (n1442,n1380,n1401);
and (n1443,n1444,n1445);
xor (n1444,n1410,n1411);
or (n1445,n1446,n1470);
and (n1446,n1447,n1448);
xor (n1447,n1412,n1441);
and (n1448,n1449,n1468);
or (n1449,n1450,n1464,n1467);
and (n1450,n1451,n1462);
or (n1451,n1452,n1460,n1461);
and (n1452,n1453,n1456);
or (n1453,n1454,n1455,n472);
and (n1454,n429,n759);
and (n1455,n759,n458);
or (n1456,n1457,n1458,n1459);
and (n1457,n767,n769);
and (n1458,n769,n771);
and (n1459,n767,n771);
and (n1460,n1456,n479);
and (n1461,n1453,n479);
xor (n1462,n1463,n1388);
xor (n1463,n1384,n290);
and (n1464,n1462,n1465);
xor (n1465,n1466,n1432);
xor (n1466,n1416,n1427);
and (n1467,n1451,n1465);
xor (n1468,n1469,n1438);
xor (n1469,n1414,n1435);
and (n1470,n1471,n1472);
xor (n1471,n1447,n1448);
or (n1472,n1473,n1490);
and (n1473,n1474,n1475);
xor (n1474,n1449,n1468);
and (n1475,n1476,n1488);
or (n1476,n1477,n1484,n1487);
and (n1477,n1478,n1482);
or (n1478,n1479,n1480,n1481);
and (n1479,n500,n764);
and (n1480,n764,n765);
and (n1481,n500,n765);
xor (n1482,n1483,n1425);
xor (n1483,n1418,n1421);
and (n1484,n1482,n1485);
xor (n1485,n1486,n479);
xor (n1486,n1453,n1456);
and (n1487,n1478,n1485);
xor (n1488,n1489,n1465);
xor (n1489,n1451,n1462);
and (n1490,n1491,n1492);
xor (n1491,n1474,n1475);
or (n1492,n1493,n1502);
and (n1493,n1494,n1495);
xor (n1494,n1476,n1488);
and (n1495,n1496,n1500);
or (n1496,n1497,n1498,n1499);
and (n1497,n754,n757);
and (n1498,n757,n762);
and (n1499,n754,n762);
xor (n1500,n1501,n1485);
xor (n1501,n1478,n1482);
and (n1502,n1503,n1504);
xor (n1503,n1494,n1495);
or (n1504,n1505,n1508);
and (n1505,n1506,n1507);
xor (n1506,n1496,n1500);
and (n1507,n748,n752);
and (n1508,n1509,n1510);
xor (n1509,n1506,n1507);
or (n1510,n1511,n745);
and (n1511,n747,n772);
endmodule
