module top (out,n14,n18,n21,n23,n29,n31,n42,n44,n47
        ,n51,n53,n59,n67,n116,n172,n286,n290,n296,n306
        ,n309,n313,n371,n425);
output out;
input n14;
input n18;
input n21;
input n23;
input n29;
input n31;
input n42;
input n44;
input n47;
input n51;
input n53;
input n59;
input n67;
input n116;
input n172;
input n286;
input n290;
input n296;
input n306;
input n309;
input n313;
input n371;
input n425;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n16;
wire n17;
wire n19;
wire n20;
wire n22;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n287;
wire n288;
wire n289;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n307;
wire n308;
wire n310;
wire n311;
wire n312;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
xor (out,n0,n620);
buf (n0,n1);
xor (n1,n2,n528);
xor (n2,n3,n275);
buf (n3,n4);
buf (n4,n5);
xor (n5,n6,n154);
xor (n6,n7,n108);
xor (n7,n8,n85);
xor (n8,n9,n34);
or (n9,n10,n24,n33);
and (n10,n11,n19);
nor (n11,n12,n15);
not (n12,n13);
buf (n13,n14);
and (n15,n16,n13);
not (n16,n17);
buf (n17,n18);
and (n19,n20,n22);
buf (n20,n21);
buf (n22,n23);
and (n24,n19,n25);
nor (n25,n26,n32);
and (n26,n27,n30);
not (n27,n28);
buf (n28,n29);
buf (n30,n31);
not (n32,n30);
and (n33,n11,n25);
or (n34,n35,n71,n84);
and (n35,n36,n69);
or (n36,n37,n62,n68);
and (n37,n38,n55);
or (n38,n39,n48,n54);
and (n39,n40,n45);
and (n40,n41,n43);
buf (n41,n42);
buf (n43,n44);
and (n45,n46,n30);
buf (n46,n47);
and (n48,n45,n49);
and (n49,n50,n52);
buf (n50,n51);
buf (n52,n53);
and (n54,n40,n49);
xor (n55,n56,n61);
xor (n56,n57,n60);
and (n57,n41,n58);
buf (n58,n59);
and (n60,n46,n43);
and (n61,n50,n30);
and (n62,n55,n63);
xor (n63,n64,n65);
and (n64,n13,n22);
and (n65,n20,n66);
buf (n66,n67);
and (n68,n38,n63);
xor (n69,n70,n25);
xor (n70,n11,n19);
and (n71,n69,n72);
xor (n72,n73,n79);
xor (n73,n74,n78);
or (n74,n75,n76,n77);
and (n75,n57,n60);
and (n76,n60,n61);
and (n77,n57,n61);
and (n78,n64,n65);
xor (n79,n80,n83);
xor (n80,n81,n82);
and (n81,n41,n66);
and (n82,n46,n58);
and (n83,n50,n43);
and (n84,n36,n72);
xor (n85,n86,n100);
xor (n86,n87,n91);
or (n87,n88,n89,n90);
and (n88,n74,n78);
and (n89,n78,n79);
and (n90,n74,n79);
xor (n91,n92,n97);
xor (n92,n93,n96);
nor (n93,n94,n95);
not (n94,n20);
and (n95,n16,n20);
and (n96,n41,n22);
nor (n97,n98,n99);
and (n98,n27,n43);
not (n99,n43);
xor (n100,n101,n107);
xor (n101,n102,n106);
or (n102,n103,n104,n105);
and (n103,n81,n82);
and (n104,n82,n83);
and (n105,n81,n83);
and (n106,n46,n66);
and (n107,n50,n58);
or (n108,n109,n150,n153);
and (n109,n110,n129);
or (n110,n111,n124,n128);
and (n111,n112,n121);
or (n112,n113,n118,n120);
and (n113,n114,n117);
and (n114,n115,n22);
buf (n115,n116);
and (n117,n13,n66);
and (n118,n117,n119);
and (n119,n20,n58);
and (n120,n114,n119);
nor (n121,n122,n123);
not (n122,n115);
and (n123,n16,n115);
and (n124,n121,n125);
nor (n125,n126,n127);
and (n126,n27,n52);
not (n127,n52);
and (n128,n112,n125);
or (n129,n130,n146,n149);
and (n130,n131,n144);
or (n131,n132,n140,n143);
and (n132,n133,n138);
or (n133,n134,1'b0,1'b0);
and (n134,n135,n136);
and (n135,n41,n30);
and (n136,n46,n52);
xor (n138,n139,n119);
xor (n139,n114,n117);
and (n140,n138,n141);
xor (n141,n142,n49);
xor (n142,n40,n45);
and (n143,n133,n141);
xor (n144,n145,n125);
xor (n145,n112,n121);
and (n146,n144,n147);
xor (n147,n148,n63);
xor (n148,n38,n55);
and (n149,n131,n147);
and (n150,n129,n151);
xor (n151,n152,n72);
xor (n152,n36,n69);
and (n153,n110,n151);
or (n154,n155,n177);
and (n155,n156,n158);
xor (n156,n157,n151);
xor (n157,n110,n129);
or (n158,1'b0,n159,1'b0);
and (n159,n160,n175);
or (n160,n161,n168,n174);
and (n161,n162,n166);
or (n162,1'b0,n163,1'b0);
and (n163,n164,n165);
and (n164,n20,n43);
xor (n165,n135,n136);
xor (n166,n167,n141);
xor (n167,n133,n138);
and (n168,n166,n169);
nor (n169,n170,n173);
not (n170,n171);
buf (n171,n172);
and (n173,n16,n171);
and (n174,n162,n169);
xor (n175,n176,n147);
xor (n176,n131,n144);
and (n177,n178,n179);
xor (n178,n156,n158);
or (n179,n180,n212);
and (n180,n181,n182);
xor (n181,n160,n175);
or (n182,n183,n208,n211);
and (n183,n184,n191);
or (n184,n185,n188,n190);
and (n185,n186,n187);
and (n186,n171,n22);
and (n187,n115,n66);
and (n188,n187,n189);
and (n189,n13,n58);
and (n190,n186,n189);
or (n191,n192,n205,n207);
and (n192,n193,n203);
or (n193,n194,n200,n202);
and (n194,n195,n199);
or (n195,n196,1'b0,1'b0);
and (n196,n197,n198);
and (n197,n13,n30);
and (n198,n20,n52);
and (n199,n20,n30);
and (n200,n199,n201);
and (n201,n41,n52);
and (n202,n195,n201);
xor (n203,n204,n189);
xor (n204,n186,n187);
and (n205,n203,n206);
xor (n206,n164,n165);
and (n207,n193,n206);
and (n208,n191,n209);
xor (n209,n210,n169);
xor (n210,n162,n166);
and (n211,n184,n209);
and (n212,n213,n214);
xor (n213,n181,n182);
or (n214,n215,n244);
and (n215,n216,n218);
xor (n216,n217,n209);
xor (n217,n184,n191);
or (n218,n219,n240,n243);
and (n219,n220,n223);
and (n220,n221,n222);
and (n221,n115,n58);
and (n222,n13,n43);
or (n223,n224,n236,n239);
and (n224,n225,n235);
or (n225,n226,n232,n234);
and (n226,n227,n231);
or (n227,n228,1'b0,1'b0);
and (n228,n229,n230);
and (n229,n115,n30);
and (n230,n13,n52);
and (n231,n115,n43);
and (n232,n231,n233);
xor (n233,n197,n198);
and (n234,n227,n233);
xor (n235,n221,n222);
and (n236,n235,n237);
xor (n237,n238,n201);
xor (n238,n195,n199);
and (n239,n225,n237);
and (n240,n223,n241);
xor (n241,n242,n206);
xor (n242,n193,n203);
and (n243,n220,n241);
and (n244,n245,n246);
xor (n245,n216,n218);
or (n246,n247,n270);
and (n247,n248,n250);
xor (n248,n249,n241);
xor (n249,n220,n223);
and (n250,n251,n268);
or (n251,n252,n264,n267);
and (n252,n253,n263);
or (n253,n254,n260,n262);
and (n254,n255,n259);
or (n255,n256,1'b0,1'b0);
and (n256,n257,n258);
and (n257,n171,n30);
and (n258,n115,n52);
and (n259,n171,n43);
and (n260,n259,n261);
xor (n261,n229,n230);
and (n262,n255,n261);
and (n263,n171,n58);
and (n264,n263,n265);
xor (n265,n266,n233);
xor (n266,n227,n231);
and (n267,n253,n265);
xor (n268,n269,n237);
xor (n269,n225,n235);
and (n270,n271,n272);
xor (n271,n248,n250);
and (n272,n273,n274);
and (n273,n171,n66);
xor (n274,n251,n268);
buf (n275,n276);
buf (n276,n277);
xor (n277,n278,n407);
xor (n278,n279,n363);
xor (n279,n280,n341);
xor (n280,n281,n298);
or (n281,n282,n291,n297);
and (n282,n283,n288);
nor (n283,n284,n287);
not (n284,n285);
buf (n285,n286);
and (n287,n16,n285);
and (n288,n289,n22);
buf (n289,n290);
and (n291,n288,n292);
nor (n292,n293,n32);
and (n293,n294,n30);
not (n294,n295);
buf (n295,n296);
and (n297,n283,n292);
or (n298,n299,n327,n340);
and (n299,n300,n325);
or (n300,n301,n320,n324);
and (n301,n302,n315);
or (n302,n303,n310,n314);
and (n303,n304,n307);
and (n304,n305,n43);
buf (n305,n306);
and (n307,n308,n30);
buf (n308,n309);
and (n310,n307,n311);
and (n311,n312,n52);
buf (n312,n313);
and (n314,n304,n311);
xor (n315,n316,n319);
xor (n316,n317,n318);
and (n317,n305,n58);
and (n318,n308,n43);
and (n319,n312,n30);
and (n320,n315,n321);
xor (n321,n322,n323);
and (n322,n285,n22);
and (n323,n289,n66);
and (n324,n302,n321);
xor (n325,n326,n292);
xor (n326,n283,n288);
and (n327,n325,n328);
xor (n328,n329,n335);
xor (n329,n330,n334);
or (n330,n331,n332,n333);
and (n331,n317,n318);
and (n332,n318,n319);
and (n333,n317,n319);
and (n334,n322,n323);
xor (n335,n336,n339);
xor (n336,n337,n338);
and (n337,n305,n66);
and (n338,n308,n58);
and (n339,n312,n43);
and (n340,n300,n328);
xor (n341,n342,n355);
xor (n342,n343,n347);
or (n343,n344,n345,n346);
and (n344,n330,n334);
and (n345,n334,n335);
and (n346,n330,n335);
xor (n347,n348,n353);
xor (n348,n349,n352);
nor (n349,n350,n351);
not (n350,n289);
and (n351,n16,n289);
and (n352,n305,n22);
nor (n353,n354,n99);
and (n354,n294,n43);
xor (n355,n356,n362);
xor (n356,n357,n361);
or (n357,n358,n359,n360);
and (n358,n337,n338);
and (n359,n338,n339);
and (n360,n337,n339);
and (n361,n308,n66);
and (n362,n312,n58);
or (n363,n364,n403,n406);
and (n364,n365,n383);
or (n365,n366,n379,n382);
and (n366,n367,n376);
or (n367,n368,n373,n375);
and (n368,n369,n372);
and (n369,n370,n22);
buf (n370,n371);
and (n372,n285,n66);
and (n373,n372,n374);
and (n374,n289,n58);
and (n375,n369,n374);
nor (n376,n377,n378);
not (n377,n370);
and (n378,n16,n370);
and (n379,n376,n380);
nor (n380,n381,n127);
and (n381,n294,n52);
and (n382,n367,n380);
or (n383,n384,n399,n402);
and (n384,n385,n397);
or (n385,n386,n393,n396);
and (n386,n387,n391);
or (n387,n388,1'b0,1'b0);
and (n388,n389,n390);
and (n389,n305,n30);
and (n390,n308,n52);
xor (n391,n392,n374);
xor (n392,n369,n372);
and (n393,n391,n394);
xor (n394,n395,n311);
xor (n395,n304,n307);
and (n396,n387,n394);
xor (n397,n398,n380);
xor (n398,n367,n376);
and (n399,n397,n400);
xor (n400,n401,n321);
xor (n401,n302,n315);
and (n402,n385,n400);
and (n403,n383,n404);
xor (n404,n405,n328);
xor (n405,n300,n325);
and (n406,n365,n404);
or (n407,n408,n430);
and (n408,n409,n411);
xor (n409,n410,n404);
xor (n410,n365,n383);
or (n411,1'b0,n412,1'b0);
and (n412,n413,n428);
or (n413,n414,n421,n427);
and (n414,n415,n419);
or (n415,1'b0,n416,1'b0);
and (n416,n417,n418);
and (n417,n289,n43);
xor (n418,n389,n390);
xor (n419,n420,n394);
xor (n420,n387,n391);
and (n421,n419,n422);
nor (n422,n423,n426);
not (n423,n424);
buf (n424,n425);
and (n426,n16,n424);
and (n427,n415,n422);
xor (n428,n429,n400);
xor (n429,n385,n397);
and (n430,n431,n432);
xor (n431,n409,n411);
or (n432,n433,n465);
and (n433,n434,n435);
xor (n434,n413,n428);
or (n435,n436,n461,n464);
and (n436,n437,n444);
or (n437,n438,n441,n443);
and (n438,n439,n440);
and (n439,n424,n22);
and (n440,n370,n66);
and (n441,n440,n442);
and (n442,n285,n58);
and (n443,n439,n442);
or (n444,n445,n458,n460);
and (n445,n446,n456);
or (n446,n447,n453,n455);
and (n447,n448,n452);
or (n448,n449,1'b0,1'b0);
and (n449,n450,n451);
and (n450,n285,n30);
and (n451,n289,n52);
and (n452,n289,n30);
and (n453,n452,n454);
and (n454,n305,n52);
and (n455,n448,n454);
xor (n456,n457,n442);
xor (n457,n439,n440);
and (n458,n456,n459);
xor (n459,n417,n418);
and (n460,n446,n459);
and (n461,n444,n462);
xor (n462,n463,n422);
xor (n463,n415,n419);
and (n464,n437,n462);
and (n465,n466,n467);
xor (n466,n434,n435);
or (n467,n468,n497);
and (n468,n469,n471);
xor (n469,n470,n462);
xor (n470,n437,n444);
or (n471,n472,n493,n496);
and (n472,n473,n476);
and (n473,n474,n475);
and (n474,n370,n58);
and (n475,n285,n43);
or (n476,n477,n489,n492);
and (n477,n478,n488);
or (n478,n479,n485,n487);
and (n479,n480,n484);
or (n480,n481,1'b0,1'b0);
and (n481,n482,n483);
and (n482,n370,n30);
and (n483,n285,n52);
and (n484,n370,n43);
and (n485,n484,n486);
xor (n486,n450,n451);
and (n487,n480,n486);
xor (n488,n474,n475);
and (n489,n488,n490);
xor (n490,n491,n454);
xor (n491,n448,n452);
and (n492,n478,n490);
and (n493,n476,n494);
xor (n494,n495,n459);
xor (n495,n446,n456);
and (n496,n473,n494);
and (n497,n498,n499);
xor (n498,n469,n471);
or (n499,n500,n523);
and (n500,n501,n503);
xor (n501,n502,n494);
xor (n502,n473,n476);
and (n503,n504,n521);
or (n504,n505,n517,n520);
and (n505,n506,n516);
or (n506,n507,n513,n515);
and (n507,n508,n512);
or (n508,n509,1'b0,1'b0);
and (n509,n510,n511);
and (n510,n424,n30);
and (n511,n370,n52);
and (n512,n424,n43);
and (n513,n512,n514);
xor (n514,n482,n483);
and (n515,n508,n514);
and (n516,n424,n58);
and (n517,n516,n518);
xor (n518,n519,n486);
xor (n519,n480,n484);
and (n520,n506,n518);
xor (n521,n522,n490);
xor (n522,n478,n488);
and (n523,n524,n525);
xor (n524,n501,n503);
and (n525,n526,n527);
and (n526,n424,n66);
xor (n527,n504,n521);
or (n528,n529,n536,n619);
and (n529,n530,n533);
buf (n530,n531);
buf (n531,n532);
xor (n532,n178,n179);
buf (n533,n534);
buf (n534,n535);
xor (n535,n431,n432);
and (n536,n533,n537);
or (n537,n538,n545,n618);
and (n538,n539,n542);
buf (n539,n540);
buf (n540,n541);
xor (n541,n213,n214);
buf (n542,n543);
buf (n543,n544);
xor (n544,n466,n467);
and (n545,n542,n546);
or (n546,n547,n554,n617);
and (n547,n548,n551);
buf (n548,n549);
buf (n549,n550);
xor (n550,n245,n246);
buf (n551,n552);
buf (n552,n553);
xor (n553,n498,n499);
and (n554,n551,n555);
or (n555,n556,n563,n616);
and (n556,n557,n560);
buf (n557,n558);
buf (n558,n559);
xor (n559,n271,n272);
buf (n560,n561);
buf (n561,n562);
xor (n562,n524,n525);
and (n563,n560,n564);
or (n564,n565,n572,n615);
and (n565,n566,n569);
buf (n566,n567);
buf (n567,n568);
xor (n568,n273,n274);
buf (n569,n570);
buf (n570,n571);
xor (n571,n526,n527);
and (n572,n569,n573);
or (n573,n574,n583,n614);
and (n574,n575,n579);
buf (n575,n576);
buf (n576,n577);
xor (n577,n578,n265);
xor (n578,n253,n263);
buf (n579,n580);
buf (n580,n581);
xor (n581,n582,n518);
xor (n582,n506,n516);
and (n583,n579,n584);
or (n584,n585,n594,n613);
and (n585,n586,n590);
buf (n586,n587);
buf (n587,n588);
xor (n588,n589,n261);
xor (n589,n255,n259);
buf (n590,n591);
buf (n591,n592);
xor (n592,n593,n514);
xor (n593,n508,n512);
and (n594,n590,n595);
or (n595,n596,n603,n612);
and (n596,n597,n600);
buf (n597,n598);
buf (n598,n599);
xor (n599,n257,n258);
buf (n600,n601);
buf (n601,n602);
xor (n602,n510,n511);
and (n603,n600,n604);
or (n604,n605,1'b0,1'b0);
and (n605,n606,n609);
buf (n606,n607);
buf (n607,n608);
and (n608,n171,n52);
buf (n609,n610);
buf (n610,n611);
and (n611,n424,n52);
and (n612,n597,n604);
and (n613,n586,n595);
and (n614,n575,n584);
and (n615,n566,n573);
and (n616,n557,n564);
and (n617,n548,n555);
and (n618,n539,n546);
and (n619,n530,n537);
buf (n620,n621);
xor (n621,n622,n779);
xor (n622,n623,n745);
xor (n623,n624,n716);
xor (n624,n625,n671);
and (n625,n626,n652);
or (n626,n627,n643,n651);
and (n627,n628,n636);
and (n628,n629,n22);
xor (n629,n630,n631);
xor (n630,n13,n285);
or (n631,n632,n633,n635);
and (n632,n115,n370);
and (n633,n370,n634);
and (n634,n171,n424);
and (n635,n115,n634);
and (n636,n637,n66);
xor (n637,n638,n639);
xor (n638,n20,n289);
or (n639,n640,n641,n642);
and (n640,n13,n285);
and (n641,n285,n631);
and (n642,n13,n631);
and (n643,n636,n644);
and (n644,n645,n58);
xor (n645,n646,n647);
xor (n646,n41,n305);
or (n647,n648,n649,n650);
and (n648,n20,n289);
and (n649,n289,n639);
and (n650,n20,n639);
and (n651,n628,n644);
nor (n652,n653,n127);
and (n653,n654,n52);
not (n654,n655);
or (n655,n656,n657,n670);
and (n656,n28,n295);
and (n657,n295,n658);
or (n658,n659,n660,n669);
and (n659,n50,n312);
and (n660,n312,n661);
or (n661,n662,n663,n668);
and (n662,n46,n308);
and (n663,n308,n664);
or (n664,n665,n666,n667);
and (n665,n41,n305);
and (n666,n305,n647);
and (n667,n41,n647);
and (n668,n46,n664);
and (n669,n50,n661);
and (n670,n28,n658);
or (n671,n672,n713,n715);
and (n672,n673,n695);
or (n673,n674,n691,n694);
and (n674,n675,n680);
nor (n675,n676,n679);
not (n676,n677);
xor (n677,n678,n634);
xor (n678,n115,n370);
and (n679,n16,n677);
xor (n680,n681,n688);
xor (n681,n682,n685);
and (n682,n683,n43);
xor (n683,n684,n664);
xor (n684,n46,n308);
and (n685,n686,n30);
xor (n686,n687,n661);
xor (n687,n50,n312);
and (n688,n689,n52);
xor (n689,n690,n658);
xor (n690,n28,n295);
and (n691,n680,n692);
xor (n692,n693,n644);
xor (n693,n628,n636);
and (n694,n675,n692);
xor (n695,n696,n706);
xor (n696,n697,n701);
or (n697,n698,n699,n700);
and (n698,n682,n685);
and (n699,n685,n688);
and (n700,n682,n688);
xor (n701,n702,n705);
xor (n702,n703,n704);
and (n703,n683,n58);
and (n704,n686,n43);
and (n705,n689,n30);
xor (n706,n707,n712);
xor (n707,n708,n711);
nor (n708,n709,n710);
not (n709,n629);
and (n710,n16,n629);
and (n711,n637,n22);
and (n712,n645,n66);
and (n713,n695,n714);
xor (n714,n626,n652);
and (n715,n673,n714);
xor (n716,n717,n730);
xor (n717,n718,n722);
or (n718,n719,n720,n721);
and (n719,n697,n701);
and (n720,n701,n706);
and (n721,n697,n706);
xor (n722,n723,n728);
xor (n723,n724,n727);
nor (n724,n725,n726);
not (n725,n637);
and (n726,n16,n637);
and (n727,n645,n22);
nor (n728,n729,n32);
and (n729,n654,n30);
xor (n730,n731,n740);
xor (n731,n732,n736);
or (n732,n733,n734,n735);
and (n733,n703,n704);
and (n734,n704,n705);
and (n735,n703,n705);
or (n736,n737,n738,n739);
and (n737,n708,n711);
and (n738,n711,n712);
and (n739,n708,n712);
xor (n740,n741,n744);
xor (n741,n742,n743);
and (n742,n683,n66);
and (n743,n686,n58);
and (n744,n689,n43);
or (n745,n746,n775,n778);
and (n746,n747,n758);
and (n747,n748,n755);
or (n748,n749,n752,n754);
and (n749,n750,n751);
and (n750,n629,n66);
and (n751,n637,n58);
and (n752,n751,n753);
and (n753,n645,n43);
and (n754,n750,n753);
and (n755,n756,n757);
and (n756,n683,n30);
and (n757,n686,n52);
or (n758,n759,n771,n774);
and (n759,n760,n770);
or (n760,n761,n767,n769);
and (n761,n762,n765);
and (n762,n763,n764);
and (n763,n645,n30);
and (n764,n683,n52);
xor (n765,n766,n753);
xor (n766,n750,n751);
and (n767,n765,n768);
xor (n768,n756,n757);
and (n769,n762,n768);
xor (n770,n748,n755);
and (n771,n770,n772);
xor (n772,n773,n692);
xor (n773,n675,n680);
and (n774,n760,n772);
and (n775,n758,n776);
xor (n776,n777,n714);
xor (n777,n673,n695);
and (n778,n747,n776);
or (n779,n780,n805);
and (n780,n781,n783);
xor (n781,n782,n776);
xor (n782,n747,n758);
or (n783,n784,n801,n804);
and (n784,n785,n791);
and (n785,n786,n790);
nor (n786,n787,n789);
not (n787,n788);
xor (n788,n171,n424);
and (n789,n16,n788);
and (n790,n677,n22);
or (n791,n792,n798,n800);
and (n792,n793,n796);
and (n793,n794,n795);
and (n794,n637,n43);
xor (n795,n763,n764);
xor (n796,n797,n768);
xor (n797,n762,n765);
and (n798,n796,n799);
xor (n799,n786,n790);
and (n800,n793,n799);
and (n801,n791,n802);
xor (n802,n803,n772);
xor (n803,n760,n770);
and (n804,n785,n802);
and (n805,n806,n807);
xor (n806,n781,n783);
or (n807,n808,n840);
and (n808,n809,n811);
xor (n809,n810,n802);
xor (n810,n785,n791);
or (n811,n812,n836,n839);
and (n812,n813,n820);
or (n813,n814,n817,n819);
and (n814,n815,n816);
and (n815,n788,n22);
and (n816,n677,n66);
and (n817,n816,n818);
and (n818,n629,n58);
and (n819,n815,n818);
or (n820,n821,n833,n835);
and (n821,n822,n831);
or (n822,n823,n828,n830);
and (n823,n824,n827);
and (n824,n825,n826);
and (n825,n629,n30);
and (n826,n637,n52);
and (n827,n637,n30);
and (n828,n827,n829);
and (n829,n645,n52);
and (n830,n824,n829);
xor (n831,n832,n818);
xor (n832,n815,n816);
and (n833,n831,n834);
xor (n834,n794,n795);
and (n835,n822,n834);
and (n836,n820,n837);
xor (n837,n838,n799);
xor (n838,n793,n796);
and (n839,n813,n837);
and (n840,n841,n842);
xor (n841,n809,n811);
or (n842,n843,n871);
and (n843,n844,n846);
xor (n844,n845,n837);
xor (n845,n813,n820);
or (n846,n847,n867,n870);
and (n847,n848,n851);
and (n848,n849,n850);
and (n849,n677,n58);
and (n850,n629,n43);
or (n851,n852,n863,n866);
and (n852,n853,n862);
or (n853,n854,n859,n861);
and (n854,n855,n858);
and (n855,n856,n857);
and (n856,n677,n30);
and (n857,n629,n52);
and (n858,n677,n43);
and (n859,n858,n860);
xor (n860,n825,n826);
and (n861,n855,n860);
xor (n862,n849,n850);
and (n863,n862,n864);
xor (n864,n865,n829);
xor (n865,n824,n827);
and (n866,n853,n864);
and (n867,n851,n868);
xor (n868,n869,n834);
xor (n869,n822,n831);
and (n870,n848,n868);
and (n871,n872,n873);
xor (n872,n844,n846);
or (n873,n874,n896);
and (n874,n875,n877);
xor (n875,n876,n868);
xor (n876,n848,n851);
and (n877,n878,n894);
or (n878,n879,n890,n893);
and (n879,n880,n889);
or (n880,n881,n886,n888);
and (n881,n882,n885);
and (n882,n883,n884);
and (n883,n788,n30);
and (n884,n677,n52);
and (n885,n788,n43);
and (n886,n885,n887);
xor (n887,n856,n857);
and (n888,n882,n887);
and (n889,n788,n58);
and (n890,n889,n891);
xor (n891,n892,n860);
xor (n892,n855,n858);
and (n893,n880,n891);
xor (n894,n895,n864);
xor (n895,n853,n862);
and (n896,n897,n898);
xor (n897,n875,n877);
and (n898,n899,n900);
and (n899,n788,n66);
xor (n900,n878,n894);
endmodule
