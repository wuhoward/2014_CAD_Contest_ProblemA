module top (out,n3,n4,n5,n24,n26,n34,n35,n45,n52
        ,n53,n61,n62,n71,n78,n80,n86,n93,n102,n103
        ,n105,n109,n114,n116,n121,n132,n141,n147,n157,n163
        ,n172,n179,n181,n190,n196,n204,n214,n222);
output out;
input n3;
input n4;
input n5;
input n24;
input n26;
input n34;
input n35;
input n45;
input n52;
input n53;
input n61;
input n62;
input n71;
input n78;
input n80;
input n86;
input n93;
input n102;
input n103;
input n105;
input n109;
input n114;
input n116;
input n121;
input n132;
input n141;
input n147;
input n157;
input n163;
input n172;
input n179;
input n181;
input n190;
input n196;
input n204;
input n214;
input n222;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n104;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
xnor (out,n0,n1017);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n1014);
nand (n7,n8,n1013);
or (n8,n9,n496);
not (n9,n10);
nand (n10,n11,n495);
not (n11,n12);
nor (n12,n13,n437);
xor (n13,n14,n368);
xor (n14,n15,n224);
xor (n15,n16,n149);
xor (n16,n17,n96);
xor (n17,n18,n73);
xor (n18,n19,n47);
nand (n19,n20,n41);
or (n20,n21,n29);
not (n21,n22);
nand (n22,n23,n27);
or (n23,n24,n25);
not (n25,n26);
or (n27,n28,n26);
not (n28,n24);
not (n29,n30);
nor (n30,n31,n37);
nand (n31,n32,n36);
or (n32,n33,n35);
not (n33,n34);
nand (n36,n35,n33);
nor (n37,n38,n40);
and (n38,n39,n24);
not (n39,n35);
and (n40,n35,n28);
nand (n41,n42,n31);
nor (n42,n43,n46);
and (n43,n28,n44);
not (n44,n45);
and (n46,n45,n24);
nand (n47,n48,n67);
or (n48,n49,n56);
nor (n49,n50,n54);
and (n50,n51,n53);
not (n51,n52);
and (n54,n52,n55);
not (n55,n53);
nand (n56,n57,n64);
not (n57,n58);
nand (n58,n59,n63);
or (n59,n60,n62);
not (n60,n61);
nand (n63,n62,n60);
nand (n64,n65,n66);
nand (n65,n60,n53);
nand (n66,n61,n55);
nand (n67,n68,n58);
nor (n68,n69,n72);
and (n69,n70,n55);
not (n70,n71);
and (n72,n71,n53);
nand (n73,n74,n88);
or (n74,n75,n83);
not (n75,n76);
nand (n76,n77,n81);
or (n77,n78,n79);
not (n79,n80);
or (n81,n82,n80);
not (n82,n78);
nor (n83,n84,n87);
and (n84,n85,n53);
not (n85,n86);
and (n87,n86,n55);
or (n88,n89,n91);
nand (n89,n83,n90);
xor (n90,n85,n82);
nor (n91,n92,n94);
and (n92,n93,n82);
and (n94,n78,n95);
not (n95,n93);
xor (n96,n97,n125);
xor (n97,n98,n106);
and (n98,n99,n105);
nand (n99,n100,n104);
or (n100,n101,n103);
not (n101,n102);
nand (n104,n103,n101);
nand (n106,n107,n118);
or (n107,n108,n110);
not (n108,n109);
not (n110,n111);
nor (n111,n112,n117);
and (n112,n113,n115);
not (n113,n114);
not (n115,n116);
and (n117,n114,n116);
or (n118,n119,n124);
nor (n119,n120,n122);
and (n120,n115,n121);
and (n122,n116,n123);
not (n123,n121);
nand (n124,n108,n116);
nand (n125,n126,n143);
or (n126,n127,n137);
nand (n127,n128,n134);
not (n128,n129);
nand (n129,n130,n133);
or (n130,n131,n116);
not (n131,n132);
nand (n133,n131,n116);
nand (n134,n135,n136);
or (n135,n34,n131);
nand (n136,n131,n34);
not (n137,n138);
nor (n138,n139,n142);
and (n139,n140,n33);
not (n140,n141);
and (n142,n141,n34);
nand (n143,n129,n144);
nor (n144,n145,n148);
and (n145,n146,n33);
not (n146,n147);
and (n148,n147,n34);
xor (n149,n150,n198);
xor (n150,n151,n174);
nand (n151,n152,n168);
or (n152,n153,n159);
not (n153,n154);
nand (n154,n155,n158);
or (n155,n102,n156);
not (n156,n157);
or (n158,n101,n157);
nand (n159,n160,n165);
not (n160,n161);
nand (n161,n162,n164);
or (n162,n82,n163);
nand (n164,n82,n163);
nand (n165,n166,n167);
or (n166,n163,n101);
nand (n167,n101,n163);
nand (n168,n169,n161);
nand (n169,n170,n173);
or (n170,n102,n171);
not (n171,n172);
or (n173,n101,n172);
nand (n174,n175,n192);
or (n175,n176,n187);
nand (n176,n177,n183);
nand (n177,n178,n182);
or (n178,n179,n180);
not (n180,n181);
nand (n182,n180,n179);
not (n183,n184);
nand (n184,n185,n186);
or (n185,n28,n179);
nand (n186,n179,n28);
nor (n187,n188,n191);
and (n188,n189,n181);
not (n189,n190);
and (n191,n190,n180);
or (n192,n183,n193);
nor (n193,n194,n197);
and (n194,n195,n181);
not (n195,n196);
and (n197,n196,n180);
nand (n198,n199,n216);
or (n199,n200,n211);
not (n200,n201);
nor (n201,n202,n208);
nor (n202,n203,n206);
and (n203,n204,n205);
not (n205,n62);
and (n206,n62,n207);
not (n207,n204);
nand (n208,n209,n210);
or (n209,n180,n204);
nand (n210,n204,n180);
nor (n211,n212,n215);
and (n212,n213,n62);
not (n213,n214);
and (n215,n214,n205);
or (n216,n217,n218);
not (n217,n208);
not (n218,n219);
nand (n219,n220,n223);
or (n220,n62,n221);
not (n221,n222);
or (n223,n205,n222);
or (n224,n225,n367);
and (n225,n226,n305);
xor (n226,n227,n267);
or (n227,n228,n266);
and (n228,n229,n249);
xor (n229,n230,n240);
nand (n230,n231,n235);
or (n231,n232,n56);
nor (n232,n233,n234);
and (n233,n95,n53);
and (n234,n93,n55);
nand (n235,n236,n58);
not (n236,n237);
nor (n237,n238,n239);
and (n238,n55,n80);
and (n239,n53,n79);
nand (n240,n241,n245);
or (n241,n242,n89);
nor (n242,n243,n244);
and (n243,n82,n157);
and (n244,n78,n156);
or (n245,n83,n246);
nor (n246,n247,n248);
and (n247,n82,n172);
and (n248,n78,n171);
and (n249,n250,n256);
nor (n250,n251,n82);
nor (n251,n252,n254);
and (n252,n253,n55);
nand (n253,n105,n86);
and (n254,n255,n85);
not (n255,n105);
nand (n256,n257,n262);
or (n257,n108,n258);
not (n258,n259);
nor (n259,n260,n261);
and (n260,n140,n115);
and (n261,n141,n116);
or (n262,n263,n124);
nor (n263,n264,n265);
and (n264,n44,n116);
and (n265,n45,n115);
and (n266,n230,n240);
xor (n267,n268,n285);
xor (n268,n269,n272);
nand (n269,n270,n271);
or (n270,n89,n246);
or (n271,n83,n91);
xor (n272,n273,n279);
nor (n273,n274,n101);
nor (n274,n275,n277);
and (n275,n276,n82);
nand (n276,n105,n163);
and (n277,n255,n278);
not (n278,n163);
nand (n279,n280,n284);
or (n280,n281,n124);
nor (n281,n282,n283);
and (n282,n146,n116);
and (n283,n147,n115);
or (n284,n119,n108);
or (n285,n286,n304);
and (n286,n287,n293);
xor (n287,n288,n289);
nor (n288,n160,n255);
nand (n289,n290,n291);
or (n290,n124,n258);
nand (n291,n292,n109);
not (n292,n281);
nand (n293,n294,n299);
or (n294,n127,n295);
not (n295,n296);
nand (n296,n297,n298);
or (n297,n34,n25);
or (n298,n33,n26);
or (n299,n128,n300);
not (n300,n301);
nand (n301,n302,n303);
or (n302,n34,n44);
or (n303,n33,n45);
and (n304,n288,n289);
or (n305,n306,n366);
and (n306,n307,n365);
xor (n307,n308,n339);
or (n308,n309,n338);
and (n309,n310,n328);
xor (n310,n311,n318);
nand (n311,n312,n317);
or (n312,n313,n127);
not (n313,n314);
nor (n314,n315,n316);
and (n315,n195,n33);
and (n316,n196,n34);
nand (n317,n296,n129);
nand (n318,n319,n324);
or (n319,n320,n176);
not (n320,n321);
nand (n321,n322,n323);
or (n322,n181,n70);
or (n323,n180,n71);
nand (n324,n184,n325);
nand (n325,n326,n327);
or (n326,n181,n213);
or (n327,n180,n214);
nand (n328,n329,n334);
or (n329,n200,n330);
not (n330,n331);
nand (n331,n332,n333);
or (n332,n62,n79);
or (n333,n205,n80);
or (n334,n217,n335);
nor (n335,n336,n337);
and (n336,n205,n52);
and (n337,n62,n51);
and (n338,n311,n318);
or (n339,n340,n364);
and (n340,n341,n358);
xor (n341,n342,n352);
nand (n342,n343,n347);
or (n343,n29,n344);
nor (n344,n345,n346);
and (n345,n28,n222);
and (n346,n24,n221);
or (n347,n348,n351);
nor (n348,n349,n350);
and (n349,n28,n190);
and (n350,n24,n189);
not (n351,n31);
nand (n352,n353,n357);
or (n353,n56,n354);
nor (n354,n355,n356);
and (n355,n55,n172);
and (n356,n53,n171);
or (n357,n232,n57);
nand (n358,n359,n363);
or (n359,n89,n360);
nor (n360,n361,n362);
and (n361,n255,n78);
and (n362,n105,n82);
or (n363,n242,n83);
and (n364,n342,n352);
xor (n365,n287,n293);
and (n366,n308,n339);
and (n367,n227,n267);
xor (n368,n369,n417);
xor (n369,n370,n373);
or (n370,n371,n372);
and (n371,n268,n285);
and (n372,n269,n272);
xor (n373,n374,n397);
xor (n374,n375,n376);
and (n375,n273,n279);
or (n376,n377,n396);
and (n377,n378,n389);
xor (n378,n379,n382);
nand (n379,n380,n381);
or (n380,n300,n127);
nand (n381,n129,n138);
nand (n382,n383,n388);
or (n383,n384,n159);
not (n384,n385);
nand (n385,n386,n387);
or (n386,n101,n105);
or (n387,n102,n255);
nand (n388,n154,n161);
nand (n389,n390,n395);
or (n390,n176,n391);
not (n391,n392);
nor (n392,n393,n394);
and (n393,n221,n180);
and (n394,n222,n181);
or (n395,n183,n187);
and (n396,n379,n382);
or (n397,n398,n416);
and (n398,n399,n413);
xor (n399,n400,n407);
nand (n400,n401,n406);
or (n401,n402,n200);
not (n402,n403);
nor (n403,n404,n405);
and (n404,n70,n205);
and (n405,n71,n62);
or (n406,n211,n217);
nand (n407,n408,n412);
or (n408,n409,n29);
nor (n409,n410,n411);
and (n410,n28,n196);
and (n411,n24,n195);
nand (n412,n31,n22);
nand (n413,n414,n415);
or (n414,n56,n237);
or (n415,n57,n49);
and (n416,n400,n407);
or (n417,n418,n436);
and (n418,n419,n435);
xor (n419,n420,n434);
or (n420,n421,n433);
and (n421,n422,n430);
xor (n422,n423,n427);
nand (n423,n424,n426);
or (n424,n425,n176);
not (n425,n325);
nand (n426,n184,n392);
nand (n427,n428,n429);
or (n428,n200,n335);
nand (n429,n208,n403);
nand (n430,n431,n432);
or (n431,n29,n348);
or (n432,n409,n351);
and (n433,n423,n427);
xor (n434,n399,n413);
xor (n435,n378,n389);
and (n436,n420,n434);
or (n437,n438,n494);
and (n438,n439,n493);
xor (n439,n440,n441);
xor (n440,n419,n435);
or (n441,n442,n492);
and (n442,n443,n446);
xor (n443,n444,n445);
xor (n444,n422,n430);
xor (n445,n229,n249);
or (n446,n447,n491);
and (n447,n448,n469);
xor (n448,n449,n450);
xor (n449,n250,n256);
or (n450,n451,n468);
and (n451,n452,n462);
xor (n452,n453,n455);
and (n453,n454,n105);
not (n454,n83);
nand (n455,n456,n461);
or (n456,n457,n127);
not (n457,n458);
nand (n458,n459,n460);
or (n459,n34,n189);
or (n460,n33,n190);
nand (n461,n129,n314);
nand (n462,n463,n464);
or (n463,n320,n183);
or (n464,n176,n465);
nor (n465,n466,n467);
and (n466,n51,n181);
and (n467,n52,n180);
and (n468,n453,n455);
or (n469,n470,n490);
and (n470,n471,n484);
xor (n471,n472,n478);
nand (n472,n473,n477);
or (n473,n474,n200);
nor (n474,n475,n476);
and (n475,n95,n62);
and (n476,n93,n205);
nand (n477,n331,n208);
nand (n478,n479,n483);
or (n479,n480,n124);
nor (n480,n481,n482);
and (n481,n115,n26);
and (n482,n116,n25);
or (n483,n263,n108);
nand (n484,n485,n489);
or (n485,n486,n56);
nor (n486,n487,n488);
and (n487,n55,n157);
and (n488,n53,n156);
or (n489,n354,n57);
and (n490,n472,n478);
and (n491,n449,n450);
and (n492,n444,n445);
xor (n493,n226,n305);
and (n494,n440,n441);
nand (n495,n13,n437);
not (n496,n497);
nand (n497,n498,n1000);
or (n498,n499,n936);
not (n499,n500);
nand (n500,n501,n925,n935);
nand (n501,n502,n680,n784);
nand (n502,n503,n644);
not (n503,n504);
xor (n504,n505,n603);
xor (n505,n506,n541);
xor (n506,n507,n523);
xor (n507,n508,n514);
nand (n508,n509,n513);
or (n509,n56,n510);
nor (n510,n511,n512);
and (n511,n255,n53);
and (n512,n55,n105);
or (n513,n57,n486);
nand (n514,n515,n519);
or (n515,n29,n516);
nor (n516,n517,n518);
and (n517,n28,n71);
and (n518,n24,n70);
or (n519,n520,n351);
nor (n520,n521,n522);
and (n521,n28,n214);
and (n522,n24,n213);
nand (n523,n524,n540);
or (n524,n525,n532);
not (n525,n526);
nand (n526,n527,n53);
nand (n527,n528,n529);
or (n528,n105,n61);
nand (n529,n530,n205);
not (n530,n531);
and (n531,n105,n61);
not (n532,n533);
nand (n533,n534,n539);
or (n534,n535,n127);
not (n535,n536);
nand (n536,n537,n538);
or (n537,n34,n221);
or (n538,n33,n222);
nand (n539,n129,n458);
or (n540,n533,n526);
xor (n541,n542,n592);
xor (n542,n543,n564);
or (n543,n544,n563);
and (n544,n545,n553);
xor (n545,n546,n547);
and (n546,n58,n105);
nand (n547,n548,n552);
or (n548,n549,n127);
nor (n549,n550,n551);
and (n550,n213,n34);
and (n551,n214,n33);
nand (n552,n129,n536);
nand (n553,n554,n559);
or (n554,n176,n555);
not (n555,n556);
nor (n556,n557,n558);
and (n557,n95,n180);
and (n558,n93,n181);
or (n559,n183,n560);
nor (n560,n561,n562);
and (n561,n80,n180);
and (n562,n79,n181);
and (n563,n546,n547);
or (n564,n565,n591);
and (n565,n566,n585);
xor (n566,n567,n576);
nand (n567,n568,n572);
or (n568,n200,n569);
nor (n569,n570,n571);
and (n570,n156,n62);
and (n571,n157,n205);
or (n572,n217,n573);
nor (n573,n574,n575);
and (n574,n172,n205);
and (n575,n171,n62);
nand (n576,n577,n581);
or (n577,n578,n124);
nor (n578,n579,n580);
and (n579,n115,n190);
and (n580,n116,n189);
or (n581,n582,n108);
nor (n582,n583,n584);
and (n583,n115,n196);
and (n584,n116,n195);
nand (n585,n586,n590);
or (n586,n29,n587);
nor (n587,n588,n589);
and (n588,n28,n52);
and (n589,n24,n51);
or (n590,n516,n351);
and (n591,n567,n576);
xor (n592,n593,n600);
xor (n593,n594,n597);
nand (n594,n595,n596);
or (n595,n176,n560);
or (n596,n465,n183);
nand (n597,n598,n599);
or (n598,n200,n573);
or (n599,n217,n474);
nand (n600,n601,n602);
or (n601,n582,n124);
or (n602,n480,n108);
or (n603,n604,n643);
and (n604,n605,n642);
xor (n605,n606,n619);
and (n606,n607,n613);
and (n607,n608,n62);
nand (n608,n609,n610);
or (n609,n105,n204);
nand (n610,n611,n180);
not (n611,n612);
and (n612,n105,n204);
nand (n613,n614,n618);
or (n614,n127,n615);
nor (n615,n616,n617);
and (n616,n33,n71);
and (n617,n34,n70);
or (n618,n128,n549);
or (n619,n620,n641);
and (n620,n621,n635);
xor (n621,n622,n629);
nand (n622,n623,n628);
or (n623,n624,n176);
not (n624,n625);
nor (n625,n626,n627);
and (n626,n172,n181);
and (n627,n171,n180);
nand (n628,n184,n556);
nand (n629,n630,n634);
or (n630,n200,n631);
nor (n631,n632,n633);
and (n632,n62,n255);
and (n633,n205,n105);
or (n634,n217,n569);
nand (n635,n636,n640);
or (n636,n124,n637);
nor (n637,n638,n639);
and (n638,n115,n222);
and (n639,n116,n221);
or (n640,n578,n108);
and (n641,n622,n629);
xor (n642,n545,n553);
and (n643,n606,n619);
not (n644,n645);
or (n645,n646,n679);
and (n646,n647,n678);
xor (n647,n648,n649);
xor (n648,n566,n585);
or (n649,n650,n677);
and (n650,n651,n659);
xor (n651,n652,n658);
nand (n652,n653,n657);
or (n653,n29,n654);
nor (n654,n655,n656);
and (n655,n28,n80);
and (n656,n24,n79);
or (n657,n587,n351);
xor (n658,n607,n613);
or (n659,n660,n676);
and (n660,n661,n669);
xor (n661,n662,n663);
and (n662,n208,n105);
nand (n663,n664,n668);
or (n664,n665,n124);
nor (n665,n666,n667);
and (n666,n115,n214);
and (n667,n116,n213);
or (n668,n637,n108);
nand (n669,n670,n675);
or (n670,n176,n671);
not (n671,n672);
nand (n672,n673,n674);
or (n673,n181,n156);
or (n674,n180,n157);
or (n675,n183,n624);
and (n676,n662,n663);
and (n677,n652,n658);
xor (n678,n605,n642);
and (n679,n648,n649);
nor (n680,n681,n721);
not (n681,n682);
or (n682,n683,n684);
xor (n683,n647,n678);
or (n684,n685,n720);
and (n685,n686,n719);
xor (n686,n687,n688);
xor (n687,n621,n635);
or (n688,n689,n718);
and (n689,n690,n703);
xor (n690,n691,n697);
nand (n691,n692,n696);
or (n692,n127,n693);
nor (n693,n694,n695);
and (n694,n33,n52);
and (n695,n34,n51);
or (n696,n128,n615);
nand (n697,n698,n702);
or (n698,n29,n699);
nor (n699,n700,n701);
and (n700,n28,n93);
and (n701,n24,n95);
or (n702,n654,n351);
and (n703,n704,n711);
nor (n704,n705,n180);
nor (n705,n706,n709);
and (n706,n707,n28);
not (n707,n708);
and (n708,n105,n179);
and (n709,n255,n710);
not (n710,n179);
nand (n711,n712,n717);
or (n712,n124,n713);
not (n713,n714);
nor (n714,n715,n716);
and (n715,n71,n116);
and (n716,n70,n115);
or (n717,n665,n108);
and (n718,n691,n697);
xor (n719,n651,n659);
and (n720,n687,n688);
nand (n721,n722,n778);
not (n722,n723);
nor (n723,n724,n753);
xor (n724,n725,n752);
xor (n725,n726,n751);
or (n726,n727,n750);
and (n727,n728,n744);
xor (n728,n729,n736);
nand (n729,n730,n735);
or (n730,n731,n176);
not (n731,n732);
nand (n732,n733,n734);
or (n733,n180,n105);
or (n734,n181,n255);
nand (n735,n184,n672);
nand (n736,n737,n742);
or (n737,n738,n127);
not (n738,n739);
nand (n739,n740,n741);
or (n740,n34,n79);
or (n741,n33,n80);
nand (n742,n743,n129);
not (n743,n693);
nand (n744,n745,n749);
or (n745,n29,n746);
nor (n746,n747,n748);
and (n747,n28,n172);
and (n748,n24,n171);
or (n749,n699,n351);
and (n750,n729,n736);
xor (n751,n661,n669);
xor (n752,n690,n703);
or (n753,n754,n777);
and (n754,n755,n776);
xor (n755,n756,n757);
xor (n756,n704,n711);
or (n757,n758,n775);
and (n758,n759,n768);
xor (n759,n760,n761);
and (n760,n184,n105);
nand (n761,n762,n763);
or (n762,n108,n713);
or (n763,n764,n124);
not (n764,n765);
nand (n765,n766,n767);
or (n766,n52,n115);
nand (n767,n115,n52);
nand (n768,n769,n774);
or (n769,n770,n127);
not (n770,n771);
nand (n771,n772,n773);
or (n772,n34,n95);
or (n773,n33,n93);
nand (n774,n129,n739);
and (n775,n760,n761);
xor (n776,n728,n744);
and (n777,n756,n757);
not (n778,n779);
nor (n779,n780,n781);
xor (n780,n686,n719);
or (n781,n782,n783);
and (n782,n725,n752);
and (n783,n726,n751);
or (n784,n785,n924);
and (n785,n786,n813);
xor (n786,n787,n812);
or (n787,n788,n811);
and (n788,n789,n810);
xor (n789,n790,n796);
nand (n790,n791,n795);
or (n791,n29,n792);
nor (n792,n793,n794);
and (n793,n28,n157);
and (n794,n24,n156);
or (n795,n746,n351);
nor (n796,n797,n805);
not (n797,n798);
nand (n798,n799,n804);
or (n799,n124,n800);
not (n800,n801);
nor (n801,n802,n803);
and (n802,n80,n116);
and (n803,n79,n115);
nand (n804,n765,n109);
nand (n805,n806,n24);
nand (n806,n807,n809);
or (n807,n808,n34);
and (n808,n105,n35);
or (n809,n105,n35);
xor (n810,n759,n768);
and (n811,n790,n796);
xor (n812,n755,n776);
or (n813,n814,n923);
and (n814,n815,n839);
xor (n815,n816,n838);
or (n816,n817,n837);
and (n817,n818,n833);
xor (n818,n819,n826);
nand (n819,n820,n825);
or (n820,n821,n127);
not (n821,n822);
nor (n822,n823,n824);
and (n823,n171,n33);
and (n824,n172,n34);
nand (n825,n129,n771);
nand (n826,n827,n832);
or (n827,n828,n29);
not (n828,n829);
nand (n829,n830,n831);
or (n830,n28,n105);
or (n831,n255,n24);
or (n832,n792,n351);
nand (n833,n834,n836);
or (n834,n835,n797);
not (n835,n805);
or (n836,n798,n805);
and (n837,n819,n826);
xor (n838,n789,n810);
or (n839,n840,n922);
and (n840,n841,n862);
xor (n841,n842,n861);
or (n842,n843,n860);
and (n843,n844,n853);
xor (n844,n845,n846);
and (n845,n31,n105);
nand (n846,n847,n852);
or (n847,n848,n127);
not (n848,n849);
nor (n849,n850,n851);
and (n850,n156,n33);
and (n851,n157,n34);
nand (n852,n129,n822);
nand (n853,n854,n855);
or (n854,n108,n800);
or (n855,n124,n856);
not (n856,n857);
nor (n857,n858,n859);
and (n858,n95,n115);
and (n859,n93,n116);
and (n860,n845,n846);
xor (n861,n818,n833);
nand (n862,n863,n921);
or (n863,n864,n880);
nor (n864,n865,n866);
xor (n865,n844,n853);
and (n866,n867,n874);
nand (n867,n868,n869);
nand (n868,n857,n109);
nand (n869,n870,n873);
nor (n870,n871,n872);
and (n871,n171,n115);
and (n872,n172,n116);
not (n873,n124);
not (n874,n875);
nand (n875,n876,n34);
nand (n876,n877,n879);
or (n877,n878,n116);
and (n878,n105,n132);
or (n879,n105,n132);
nor (n880,n881,n920);
and (n881,n882,n894);
nand (n882,n883,n887);
nor (n883,n884,n886);
and (n884,n885,n874);
not (n885,n867);
and (n886,n867,n875);
nor (n887,n888,n889);
and (n888,n129,n849);
and (n889,n890,n891);
not (n890,n127);
nand (n891,n892,n893);
or (n892,n33,n105);
or (n893,n255,n34);
nand (n894,n895,n918);
or (n895,n896,n910);
not (n896,n897);
and (n897,n898,n908);
nand (n898,n899,n904);
or (n899,n108,n900);
not (n900,n901);
nor (n901,n902,n903);
and (n902,n156,n115);
and (n903,n157,n116);
nand (n904,n905,n873);
nand (n905,n906,n907);
or (n906,n115,n105);
or (n907,n116,n255);
nor (n908,n909,n115);
and (n909,n105,n109);
not (n910,n911);
nand (n911,n912,n917);
not (n912,n913);
nand (n913,n914,n916);
or (n914,n108,n915);
not (n915,n870);
nand (n916,n901,n873);
nand (n917,n129,n105);
nand (n918,n919,n913);
not (n919,n917);
nor (n920,n883,n887);
nand (n921,n865,n866);
and (n922,n842,n861);
and (n923,n816,n838);
and (n924,n787,n812);
nand (n925,n926,n502);
or (n926,n927,n929);
not (n927,n928);
nand (n928,n683,n684);
not (n929,n930);
nand (n930,n682,n931);
nand (n931,n932,n934);
or (n932,n779,n933);
nand (n933,n724,n753);
nand (n934,n780,n781);
nand (n935,n504,n645);
not (n936,n937);
nor (n937,n938,n963);
nor (n938,n939,n940);
xor (n939,n439,n493);
or (n940,n941,n962);
and (n941,n942,n945);
xor (n942,n943,n944);
xor (n943,n307,n365);
xor (n944,n443,n446);
or (n945,n946,n961);
and (n946,n947,n950);
xor (n947,n948,n949);
xor (n948,n341,n358);
xor (n949,n310,n328);
or (n950,n951,n960);
and (n951,n952,n957);
xor (n952,n953,n956);
nand (n953,n954,n955);
or (n954,n29,n520);
or (n955,n344,n351);
and (n956,n533,n525);
or (n957,n958,n959);
and (n958,n593,n600);
and (n959,n594,n597);
and (n960,n953,n956);
and (n961,n948,n949);
and (n962,n943,n944);
nand (n963,n964,n993);
nor (n964,n965,n988);
nor (n965,n966,n979);
xor (n966,n967,n978);
xor (n967,n968,n969);
xor (n968,n448,n469);
or (n969,n970,n977);
and (n970,n971,n974);
xor (n971,n972,n973);
xor (n972,n471,n484);
xor (n973,n452,n462);
or (n974,n975,n976);
and (n975,n507,n523);
and (n976,n508,n514);
and (n977,n972,n973);
xor (n978,n947,n950);
or (n979,n980,n987);
and (n980,n981,n986);
xor (n981,n982,n983);
xor (n982,n952,n957);
or (n983,n984,n985);
and (n984,n542,n592);
and (n985,n543,n564);
xor (n986,n971,n974);
and (n987,n982,n983);
nor (n988,n989,n992);
or (n989,n990,n991);
and (n990,n505,n603);
and (n991,n506,n541);
xor (n992,n981,n986);
nand (n993,n994,n996);
not (n994,n995);
xor (n995,n942,n945);
not (n996,n997);
or (n997,n998,n999);
and (n998,n967,n978);
and (n999,n968,n969);
nor (n1000,n1001,n1012);
and (n1001,n1002,n1003);
not (n1002,n938);
nand (n1003,n1004,n1011);
or (n1004,n1005,n1006);
not (n1005,n993);
not (n1006,n1007);
nand (n1007,n1008,n1010);
or (n1008,n965,n1009);
nand (n1009,n989,n992);
nand (n1010,n966,n979);
nand (n1011,n995,n997);
and (n1012,n939,n940);
or (n1013,n497,n10);
not (n1014,n1015);
nand (n1015,n1016,n3);
not (n1016,n4);
wire s0n1017,s1n1017,notn1017;
or (n1017,s0n1017,s1n1017);
not(notn1017,n4);
and (s0n1017,notn1017,n1018);
and (s1n1017,n4,1'b0);
wire s0n1018,s1n1018,notn1018;
or (n1018,s0n1018,s1n1018);
not(notn1018,n3);
and (s0n1018,notn1018,n5);
and (s1n1018,n3,n1019);
xor (n1019,n1020,n1722);
xor (n1020,n1021,n1719);
xor (n1021,n1022,n1718);
xor (n1022,n1023,n1709);
xor (n1023,n1024,n1708);
xor (n1024,n1025,n1693);
xor (n1025,n1026,n1692);
xor (n1026,n1027,n1671);
xor (n1027,n1028,n1670);
xor (n1028,n1029,n1643);
xor (n1029,n1030,n1642);
xor (n1030,n1031,n1610);
xor (n1031,n1032,n1609);
xor (n1032,n1033,n1571);
xor (n1033,n1034,n1570);
xor (n1034,n1035,n1526);
xor (n1035,n1036,n1525);
xor (n1036,n1037,n1477);
xor (n1037,n1038,n1476);
xor (n1038,n1039,n1420);
xor (n1039,n1040,n1419);
xor (n1040,n1041,n1356);
xor (n1041,n1042,n1355);
xor (n1042,n1043,n1287);
xor (n1043,n1044,n1286);
xor (n1044,n1045,n1214);
xor (n1045,n1046,n142);
xor (n1046,n1047,n1134);
xor (n1047,n1048,n1133);
xor (n1048,n1049,n1052);
xor (n1049,n1050,n1051);
and (n1050,n114,n109);
and (n1051,n121,n116);
or (n1052,n1053,n1056);
and (n1053,n1054,n1055);
and (n1054,n121,n109);
and (n1055,n147,n116);
and (n1056,n1057,n1058);
xor (n1057,n1054,n1055);
or (n1058,n1059,n1061);
and (n1059,n1060,n261);
and (n1060,n147,n109);
and (n1061,n1062,n1063);
xor (n1062,n1060,n261);
or (n1063,n1064,n1067);
and (n1064,n1065,n1066);
and (n1065,n141,n109);
and (n1066,n45,n116);
and (n1067,n1068,n1069);
xor (n1068,n1065,n1066);
or (n1069,n1070,n1073);
and (n1070,n1071,n1072);
and (n1071,n45,n109);
and (n1072,n26,n116);
and (n1073,n1074,n1075);
xor (n1074,n1071,n1072);
or (n1075,n1076,n1079);
and (n1076,n1077,n1078);
and (n1077,n26,n109);
and (n1078,n196,n116);
and (n1079,n1080,n1081);
xor (n1080,n1077,n1078);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
and (n1083,n196,n109);
and (n1084,n190,n116);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
and (n1089,n190,n109);
and (n1090,n222,n116);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
and (n1095,n222,n109);
and (n1096,n214,n116);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
or (n1099,n1100,n1102);
and (n1100,n1101,n715);
and (n1101,n214,n109);
and (n1102,n1103,n1104);
xor (n1103,n1101,n715);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
and (n1106,n71,n109);
and (n1107,n52,n116);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1113);
and (n1111,n1112,n802);
and (n1112,n52,n109);
and (n1113,n1114,n1115);
xor (n1114,n1112,n802);
or (n1115,n1116,n1118);
and (n1116,n1117,n859);
and (n1117,n80,n109);
and (n1118,n1119,n1120);
xor (n1119,n1117,n859);
or (n1120,n1121,n1123);
and (n1121,n1122,n872);
and (n1122,n93,n109);
and (n1123,n1124,n1125);
xor (n1124,n1122,n872);
or (n1125,n1126,n1128);
and (n1126,n1127,n903);
and (n1127,n172,n109);
and (n1128,n1129,n1130);
xor (n1129,n1127,n903);
and (n1130,n1131,n1132);
and (n1131,n157,n109);
and (n1132,n105,n116);
and (n1133,n147,n132);
or (n1134,n1135,n1138);
and (n1135,n1136,n1137);
xor (n1136,n1057,n1058);
and (n1137,n141,n132);
and (n1138,n1139,n1140);
xor (n1139,n1136,n1137);
or (n1140,n1141,n1144);
and (n1141,n1142,n1143);
xor (n1142,n1062,n1063);
and (n1143,n45,n132);
and (n1144,n1145,n1146);
xor (n1145,n1142,n1143);
or (n1146,n1147,n1150);
and (n1147,n1148,n1149);
xor (n1148,n1068,n1069);
and (n1149,n26,n132);
and (n1150,n1151,n1152);
xor (n1151,n1148,n1149);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
xor (n1154,n1074,n1075);
and (n1155,n196,n132);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
xor (n1160,n1080,n1081);
and (n1161,n190,n132);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
xor (n1166,n1086,n1087);
and (n1167,n222,n132);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1092,n1093);
and (n1173,n214,n132);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1098,n1099);
and (n1179,n71,n132);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1103,n1104);
and (n1185,n52,n132);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1109,n1110);
and (n1191,n80,n132);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1114,n1115);
and (n1197,n93,n132);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1119,n1120);
and (n1203,n172,n132);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1124,n1125);
and (n1209,n157,n132);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
and (n1212,n1213,n878);
xor (n1213,n1129,n1130);
or (n1214,n1215,n1218);
and (n1215,n1216,n1217);
xor (n1216,n1139,n1140);
and (n1217,n45,n34);
and (n1218,n1219,n1220);
xor (n1219,n1216,n1217);
or (n1220,n1221,n1224);
and (n1221,n1222,n1223);
xor (n1222,n1145,n1146);
and (n1223,n26,n34);
and (n1224,n1225,n1226);
xor (n1225,n1222,n1223);
or (n1226,n1227,n1229);
and (n1227,n1228,n316);
xor (n1228,n1151,n1152);
and (n1229,n1230,n1231);
xor (n1230,n1228,n316);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1157,n1158);
and (n1234,n190,n34);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1163,n1164);
and (n1240,n222,n34);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1169,n1170);
and (n1246,n214,n34);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1175,n1176);
and (n1252,n71,n34);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
or (n1255,n1256,n1259);
and (n1256,n1257,n1258);
xor (n1257,n1181,n1182);
and (n1258,n52,n34);
and (n1259,n1260,n1261);
xor (n1260,n1257,n1258);
or (n1261,n1262,n1265);
and (n1262,n1263,n1264);
xor (n1263,n1187,n1188);
and (n1264,n80,n34);
and (n1265,n1266,n1267);
xor (n1266,n1263,n1264);
or (n1267,n1268,n1271);
and (n1268,n1269,n1270);
xor (n1269,n1193,n1194);
and (n1270,n93,n34);
and (n1271,n1272,n1273);
xor (n1272,n1269,n1270);
or (n1273,n1274,n1276);
and (n1274,n1275,n824);
xor (n1275,n1199,n1200);
and (n1276,n1277,n1278);
xor (n1277,n1275,n824);
or (n1278,n1279,n1281);
and (n1279,n1280,n851);
xor (n1280,n1205,n1206);
and (n1281,n1282,n1283);
xor (n1282,n1280,n851);
and (n1283,n1284,n1285);
xor (n1284,n1211,n1212);
and (n1285,n105,n34);
and (n1286,n45,n35);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1219,n1220);
and (n1290,n26,n35);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1225,n1226);
and (n1296,n196,n35);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1230,n1231);
and (n1302,n190,n35);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1236,n1237);
and (n1308,n222,n35);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1242,n1243);
and (n1314,n214,n35);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1248,n1249);
and (n1320,n71,n35);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1254,n1255);
and (n1326,n52,n35);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1260,n1261);
and (n1332,n80,n35);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
or (n1335,n1336,n1339);
and (n1336,n1337,n1338);
xor (n1337,n1266,n1267);
and (n1338,n93,n35);
and (n1339,n1340,n1341);
xor (n1340,n1337,n1338);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1272,n1273);
and (n1344,n172,n35);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1351);
and (n1348,n1349,n1350);
xor (n1349,n1277,n1278);
and (n1350,n157,n35);
and (n1351,n1352,n1353);
xor (n1352,n1349,n1350);
and (n1353,n1354,n808);
xor (n1354,n1282,n1283);
and (n1355,n26,n24);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1292,n1293);
and (n1359,n196,n24);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1298,n1299);
and (n1365,n190,n24);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1304,n1305);
and (n1371,n222,n24);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1310,n1311);
and (n1377,n214,n24);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1316,n1317);
and (n1383,n71,n24);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1322,n1323);
and (n1389,n52,n24);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
or (n1392,n1393,n1396);
and (n1393,n1394,n1395);
xor (n1394,n1328,n1329);
and (n1395,n80,n24);
and (n1396,n1397,n1398);
xor (n1397,n1394,n1395);
or (n1398,n1399,n1402);
and (n1399,n1400,n1401);
xor (n1400,n1334,n1335);
and (n1401,n93,n24);
and (n1402,n1403,n1404);
xor (n1403,n1400,n1401);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1340,n1341);
and (n1407,n172,n24);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1414);
and (n1411,n1412,n1413);
xor (n1412,n1346,n1347);
and (n1413,n157,n24);
and (n1414,n1415,n1416);
xor (n1415,n1412,n1413);
and (n1416,n1417,n1418);
xor (n1417,n1352,n1353);
and (n1418,n105,n24);
and (n1419,n196,n179);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1361,n1362);
and (n1423,n190,n179);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1367,n1368);
and (n1429,n222,n179);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
or (n1432,n1433,n1436);
and (n1433,n1434,n1435);
xor (n1434,n1373,n1374);
and (n1435,n214,n179);
and (n1436,n1437,n1438);
xor (n1437,n1434,n1435);
or (n1438,n1439,n1442);
and (n1439,n1440,n1441);
xor (n1440,n1379,n1380);
and (n1441,n71,n179);
and (n1442,n1443,n1444);
xor (n1443,n1440,n1441);
or (n1444,n1445,n1448);
and (n1445,n1446,n1447);
xor (n1446,n1385,n1386);
and (n1447,n52,n179);
and (n1448,n1449,n1450);
xor (n1449,n1446,n1447);
or (n1450,n1451,n1454);
and (n1451,n1452,n1453);
xor (n1452,n1391,n1392);
and (n1453,n80,n179);
and (n1454,n1455,n1456);
xor (n1455,n1452,n1453);
or (n1456,n1457,n1460);
and (n1457,n1458,n1459);
xor (n1458,n1397,n1398);
and (n1459,n93,n179);
and (n1460,n1461,n1462);
xor (n1461,n1458,n1459);
or (n1462,n1463,n1466);
and (n1463,n1464,n1465);
xor (n1464,n1403,n1404);
and (n1465,n172,n179);
and (n1466,n1467,n1468);
xor (n1467,n1464,n1465);
or (n1468,n1469,n1472);
and (n1469,n1470,n1471);
xor (n1470,n1409,n1410);
and (n1471,n157,n179);
and (n1472,n1473,n1474);
xor (n1473,n1470,n1471);
and (n1474,n1475,n708);
xor (n1475,n1415,n1416);
and (n1476,n190,n181);
or (n1477,n1478,n1480);
and (n1478,n1479,n394);
xor (n1479,n1425,n1426);
and (n1480,n1481,n1482);
xor (n1481,n1479,n394);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1431,n1432);
and (n1485,n214,n181);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1437,n1438);
and (n1491,n71,n181);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1443,n1444);
and (n1497,n52,n181);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1449,n1450);
and (n1503,n80,n181);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1509);
and (n1507,n1508,n558);
xor (n1508,n1455,n1456);
and (n1509,n1510,n1511);
xor (n1510,n1508,n558);
or (n1511,n1512,n1514);
and (n1512,n1513,n626);
xor (n1513,n1461,n1462);
and (n1514,n1515,n1516);
xor (n1515,n1513,n626);
or (n1516,n1517,n1520);
and (n1517,n1518,n1519);
xor (n1518,n1467,n1468);
and (n1519,n157,n181);
and (n1520,n1521,n1522);
xor (n1521,n1518,n1519);
and (n1522,n1523,n1524);
xor (n1523,n1473,n1474);
and (n1524,n105,n181);
and (n1525,n222,n204);
or (n1526,n1527,n1530);
and (n1527,n1528,n1529);
xor (n1528,n1481,n1482);
and (n1529,n214,n204);
and (n1530,n1531,n1532);
xor (n1531,n1528,n1529);
or (n1532,n1533,n1536);
and (n1533,n1534,n1535);
xor (n1534,n1487,n1488);
and (n1535,n71,n204);
and (n1536,n1537,n1538);
xor (n1537,n1534,n1535);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1493,n1494);
and (n1541,n52,n204);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
or (n1544,n1545,n1548);
and (n1545,n1546,n1547);
xor (n1546,n1499,n1500);
and (n1547,n80,n204);
and (n1548,n1549,n1550);
xor (n1549,n1546,n1547);
or (n1550,n1551,n1554);
and (n1551,n1552,n1553);
xor (n1552,n1505,n1506);
and (n1553,n93,n204);
and (n1554,n1555,n1556);
xor (n1555,n1552,n1553);
or (n1556,n1557,n1560);
and (n1557,n1558,n1559);
xor (n1558,n1510,n1511);
and (n1559,n172,n204);
and (n1560,n1561,n1562);
xor (n1561,n1558,n1559);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
xor (n1564,n1515,n1516);
and (n1565,n157,n204);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
and (n1568,n1569,n612);
xor (n1569,n1521,n1522);
and (n1570,n214,n62);
or (n1571,n1572,n1574);
and (n1572,n1573,n405);
xor (n1573,n1531,n1532);
and (n1574,n1575,n1576);
xor (n1575,n1573,n405);
or (n1576,n1577,n1580);
and (n1577,n1578,n1579);
xor (n1578,n1537,n1538);
and (n1579,n52,n62);
and (n1580,n1581,n1582);
xor (n1581,n1578,n1579);
or (n1582,n1583,n1586);
and (n1583,n1584,n1585);
xor (n1584,n1543,n1544);
and (n1585,n80,n62);
and (n1586,n1587,n1588);
xor (n1587,n1584,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n1549,n1550);
and (n1591,n93,n62);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1555,n1556);
and (n1597,n172,n62);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1561,n1562);
and (n1603,n157,n62);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
and (n1606,n1607,n1608);
xor (n1607,n1567,n1568);
and (n1608,n105,n62);
and (n1609,n71,n61);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1575,n1576);
and (n1613,n52,n61);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
xor (n1618,n1581,n1582);
and (n1619,n80,n61);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
xor (n1624,n1587,n1588);
and (n1625,n93,n61);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1593,n1594);
and (n1631,n172,n61);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1599,n1600);
and (n1637,n157,n61);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
and (n1640,n1641,n531);
xor (n1641,n1605,n1606);
and (n1642,n52,n53);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1615,n1616);
and (n1646,n80,n53);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1621,n1622);
and (n1652,n93,n53);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1627,n1628);
and (n1658,n172,n53);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1633,n1634);
and (n1664,n157,n53);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
and (n1667,n1668,n1669);
xor (n1668,n1639,n1640);
and (n1669,n105,n53);
and (n1670,n80,n86);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1648,n1649);
and (n1674,n93,n86);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1654,n1655);
and (n1680,n172,n86);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1660,n1661);
and (n1686,n157,n86);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
and (n1689,n1690,n1691);
xor (n1690,n1666,n1667);
not (n1691,n253);
and (n1692,n93,n78);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1676,n1677);
and (n1696,n172,n78);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1682,n1683);
and (n1702,n157,n78);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
and (n1705,n1706,n1707);
xor (n1706,n1688,n1689);
and (n1707,n105,n78);
and (n1708,n172,n163);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1698,n1699);
and (n1712,n157,n163);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
and (n1715,n1716,n1717);
xor (n1716,n1704,n1705);
not (n1717,n276);
and (n1718,n157,n102);
and (n1719,n1720,n1721);
xor (n1720,n1714,n1715);
and (n1721,n105,n102);
and (n1722,n105,n103);
endmodule
