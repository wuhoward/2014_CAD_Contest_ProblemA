module top (out,n17,n22,n23,n24,n26,n27,n38,n41,n44
        ,n47,n50,n53,n56,n59,n62,n65,n68,n70,n73
        ,n82,n93,n98,n101,n104,n107,n110,n113,n116,n119
        ,n122,n125,n128,n139,n336,n351,n460,n472);
output out;
input n17;
input n22;
input n23;
input n24;
input n26;
input n27;
input n38;
input n41;
input n44;
input n47;
input n50;
input n53;
input n56;
input n59;
input n62;
input n65;
input n68;
input n70;
input n73;
input n82;
input n93;
input n98;
input n101;
input n104;
input n107;
input n110;
input n113;
input n116;
input n119;
input n122;
input n125;
input n128;
input n139;
input n336;
input n351;
input n460;
input n472;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n25;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n63;
wire n64;
wire n66;
wire n67;
wire n69;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n102;
wire n103;
wire n105;
wire n106;
wire n108;
wire n109;
wire n111;
wire n112;
wire n114;
wire n115;
wire n117;
wire n118;
wire n120;
wire n121;
wire n123;
wire n124;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
xor (out,n0,n909);
xor (n0,n1,n533);
xor (n1,n2,n448);
or (n2,n3,n447);
and (n3,n4,n361);
xor (n4,n5,n326);
or (n5,n6,n325);
and (n6,n7,n277);
xor (n7,n8,n177);
xor (n8,n9,n145);
xor (n9,n10,n83);
nor (n10,n11,n80);
not (n11,n12);
nor (n12,n13,n77);
and (n13,n14,n74);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n71);
and (s0n14,notn14,n15);
and (s1n14,n71,n34);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n18);
and (s0n15,notn15,1'b0);
and (s1n15,n18,n17);
or (n18,n19,n30);
or (n19,n20,n28);
nor (n20,n21,n23,n24,n25,n27);
not (n21,n22);
not (n25,n26);
nor (n28,n22,n29,n24,n25,n27);
not (n29,n23);
or (n30,n31,n33);
and (n31,n21,n23,n24,n25,n32);
not (n32,n27);
nor (n33,n21,n29,n24,n25,n27);
xor (n34,n35,n36);
not (n35,n17);
and (n36,n37,n39);
not (n37,n38);
and (n39,n40,n42);
not (n40,n41);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n57);
not (n55,n56);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n66);
not (n64,n65);
and (n66,n67,n69);
not (n67,n68);
not (n69,n70);
and (n71,n72,n73);
or (n72,n20,n31);
wire s0n74,s1n74,notn74;
or (n74,s0n74,s1n74);
not(notn74,n71);
and (s0n74,notn74,n75);
and (s1n74,n71,n76);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n18);
and (s0n75,notn75,1'b0);
and (s1n75,n18,n38);
xor (n76,n37,n39);
and (n77,n78,n79);
not (n78,n14);
not (n79,n74);
not (n80,n81);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n18);
and (s0n81,notn81,1'b0);
and (s1n81,n18,n82);
nand (n83,n84,n134);
or (n84,n85,n131);
nor (n85,n86,n129);
and (n86,n87,n91);
not (n87,n88);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n71);
and (s0n88,notn88,n89);
and (s1n88,n71,n90);
wire s0n89,s1n89,notn89;
or (n89,s0n89,s1n89);
not(notn89,n18);
and (s0n89,notn89,1'b0);
and (s1n89,n18,n68);
xor (n90,n67,n69);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n127);
and (s0n91,notn91,n92);
and (s1n91,n127,n94);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n18);
and (s0n92,notn92,1'b0);
and (s1n92,n18,n93);
xor (n94,n95,n96);
not (n95,n93);
and (n96,n97,n99);
not (n97,n98);
and (n99,n100,n102);
not (n100,n101);
and (n102,n103,n105);
not (n103,n104);
and (n105,n106,n108);
not (n106,n107);
and (n108,n109,n111);
not (n109,n110);
and (n111,n112,n114);
not (n112,n113);
and (n114,n115,n117);
not (n115,n116);
and (n117,n118,n120);
not (n118,n119);
and (n120,n121,n123);
not (n121,n122);
and (n123,n124,n126);
not (n124,n125);
not (n126,n82);
and (n127,n72,n128);
and (n129,n130,n88);
not (n130,n91);
nand (n131,n88,n132);
not (n132,n133);
wire s0n133,s1n133,notn133;
or (n133,s0n133,s1n133);
not(notn133,n18);
and (s0n133,notn133,1'b0);
and (s1n133,n18,n70);
or (n134,n135,n132);
nor (n135,n136,n143);
and (n136,n87,n137);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n127);
and (s0n137,notn137,n138);
and (s1n137,n127,n140);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n18);
and (s0n138,notn138,1'b0);
and (s1n138,n18,n139);
xor (n140,n141,n142);
not (n141,n139);
and (n142,n95,n96);
and (n143,n144,n88);
not (n144,n137);
nand (n145,n146,n165);
or (n146,n147,n154);
nor (n147,n148,n152);
and (n148,n87,n149);
wire s0n149,s1n149,notn149;
or (n149,s0n149,s1n149);
not(notn149,n71);
and (s0n149,notn149,n150);
and (s1n149,n71,n151);
wire s0n150,s1n150,notn150;
or (n150,s0n150,s1n150);
not(notn150,n18);
and (s0n150,notn150,1'b0);
and (s1n150,n18,n65);
xor (n151,n64,n66);
and (n152,n88,n153);
not (n153,n149);
nor (n154,n155,n163);
and (n155,n156,n160);
not (n156,n157);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n71);
and (s0n157,notn157,n158);
and (s1n157,n71,n159);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n18);
and (s0n158,notn158,1'b0);
and (s1n158,n18,n62);
xor (n159,n61,n63);
wire s0n160,s1n160,notn160;
or (n160,s0n160,s1n160);
not(notn160,n127);
and (s0n160,notn160,n161);
and (s1n160,n127,n162);
wire s0n161,s1n161,notn161;
or (n161,s0n161,s1n161);
not(notn161,n18);
and (s0n161,notn161,1'b0);
and (s1n161,n18,n98);
xor (n162,n97,n99);
and (n163,n164,n157);
not (n164,n160);
or (n165,n166,n170);
nand (n166,n147,n167);
nand (n167,n168,n169);
or (n168,n156,n149);
nand (n169,n156,n149);
nor (n170,n171,n175);
and (n171,n172,n156);
wire s0n172,s1n172,notn172;
or (n172,s0n172,s1n172);
not(notn172,n127);
and (s0n172,notn172,n173);
and (s1n172,n127,n174);
wire s0n173,s1n173,notn173;
or (n173,s0n173,s1n173);
not(notn173,n18);
and (s0n173,notn173,1'b0);
and (s1n173,n18,n101);
xor (n174,n100,n102);
and (n175,n176,n157);
not (n176,n172);
xor (n177,n178,n249);
xor (n178,n179,n215);
nand (n179,n180,n207);
or (n180,n181,n200);
nand (n181,n182,n193);
or (n182,n183,n190);
and (n183,n184,n187);
wire s0n184,s1n184,notn184;
or (n184,s0n184,s1n184);
not(notn184,n71);
and (s0n184,notn184,n185);
and (s1n184,n71,n186);
wire s0n185,s1n185,notn185;
or (n185,s0n185,s1n185);
not(notn185,n18);
and (s0n185,notn185,1'b0);
and (s1n185,n18,n56);
xor (n186,n55,n57);
wire s0n187,s1n187,notn187;
or (n187,s0n187,s1n187);
not(notn187,n71);
and (s0n187,notn187,n188);
and (s1n187,n71,n189);
wire s0n188,s1n188,notn188;
or (n188,s0n188,s1n188);
not(notn188,n18);
and (s0n188,notn188,1'b0);
and (s1n188,n18,n53);
xor (n189,n52,n54);
and (n190,n191,n192);
not (n191,n184);
not (n192,n187);
nor (n193,n194,n198);
and (n194,n195,n187);
wire s0n195,s1n195,notn195;
or (n195,s0n195,s1n195);
not(notn195,n71);
and (s0n195,notn195,n196);
and (s1n195,n71,n197);
wire s0n196,s1n196,notn196;
or (n196,s0n196,s1n196);
not(notn196,n18);
and (s0n196,notn196,1'b0);
and (s1n196,n18,n50);
xor (n197,n49,n51);
and (n198,n199,n192);
not (n199,n195);
nor (n200,n201,n205);
and (n201,n202,n199);
wire s0n202,s1n202,notn202;
or (n202,s0n202,s1n202);
not(notn202,n127);
and (s0n202,notn202,n203);
and (s1n202,n127,n204);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n18);
and (s0n203,notn203,1'b0);
and (s1n203,n18,n113);
xor (n204,n112,n114);
and (n205,n206,n195);
not (n206,n202);
or (n207,n208,n182);
nor (n208,n209,n213);
and (n209,n210,n199);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n127);
and (s0n210,notn210,n211);
and (s1n210,n127,n212);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n18);
and (s0n211,notn211,1'b0);
and (s1n211,n18,n110);
xor (n212,n109,n111);
and (n213,n214,n195);
not (n214,n210);
nand (n215,n216,n237);
or (n216,n217,n225);
not (n217,n218);
nor (n218,n219,n223);
and (n219,n195,n220);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n71);
and (s0n220,notn220,n221);
and (s1n220,n71,n222);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n18);
and (s0n221,notn221,1'b0);
and (s1n221,n18,n47);
xor (n222,n46,n48);
and (n223,n199,n224);
not (n224,n220);
not (n225,n226);
nand (n226,n227,n235);
or (n227,n228,n231);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n71);
and (s0n228,notn228,n229);
and (s1n228,n71,n230);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n18);
and (s0n229,notn229,1'b0);
and (s1n229,n18,n44);
xor (n230,n43,n45);
not (n231,n232);
wire s0n232,s1n232,notn232;
or (n232,s0n232,s1n232);
not(notn232,n127);
and (s0n232,notn232,n233);
and (s1n232,n127,n234);
wire s0n233,s1n233,notn233;
or (n233,s0n233,s1n233);
not(notn233,n18);
and (s0n233,notn233,1'b0);
and (s1n233,n18,n116);
xor (n234,n115,n117);
or (n235,n236,n232);
not (n236,n228);
or (n237,n238,n242);
nand (n238,n239,n217);
nor (n239,n240,n241);
and (n240,n220,n228);
and (n241,n224,n236);
nor (n242,n243,n247);
and (n243,n236,n244);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n127);
and (s0n244,notn244,n245);
and (s1n244,n127,n246);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n18);
and (s0n245,notn245,1'b0);
and (s1n245,n18,n119);
xor (n246,n118,n120);
and (n247,n228,n248);
not (n248,n244);
nand (n249,n250,n265);
or (n250,n251,n258);
or (n251,n252,n256);
and (n252,n253,n228);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n71);
and (s0n253,notn253,n254);
and (s1n253,n71,n255);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n18);
and (s0n254,notn254,1'b0);
and (s1n254,n18,n41);
xor (n255,n40,n42);
and (n256,n257,n236);
not (n257,n253);
nor (n258,n259,n263);
and (n259,n260,n79);
wire s0n260,s1n260,notn260;
or (n260,s0n260,s1n260);
not(notn260,n127);
and (s0n260,notn260,n261);
and (s1n260,n127,n262);
wire s0n261,s1n261,notn261;
or (n261,s0n261,s1n261);
not(notn261,n18);
and (s0n261,notn261,1'b0);
and (s1n261,n18,n122);
xor (n262,n121,n123);
and (n263,n264,n74);
not (n264,n260);
or (n265,n266,n270);
nand (n266,n251,n267);
nand (n267,n268,n269);
or (n268,n257,n74);
or (n269,n79,n253);
nor (n270,n271,n275);
and (n271,n272,n79);
wire s0n272,s1n272,notn272;
or (n272,s0n272,s1n272);
not(notn272,n127);
and (s0n272,notn272,n273);
and (s1n272,n127,n274);
wire s0n273,s1n273,notn273;
or (n273,s0n273,s1n273);
not(notn273,n18);
and (s0n273,notn273,1'b0);
and (s1n273,n18,n125);
xor (n274,n124,n126);
and (n275,n276,n74);
not (n276,n272);
or (n277,n278,n324);
and (n278,n279,n311);
xor (n279,n280,n286);
nand (n280,n281,n285);
or (n281,n266,n282);
nor (n282,n283,n284);
and (n283,n74,n80);
and (n284,n79,n81);
or (n285,n270,n251);
nand (n286,n287,n303);
or (n287,n288,n300);
nand (n288,n289,n296);
not (n289,n290);
nand (n290,n291,n295);
or (n291,n156,n292);
wire s0n292,s1n292,notn292;
or (n292,s0n292,s1n292);
not(notn292,n71);
and (s0n292,notn292,n293);
and (s1n292,n71,n294);
wire s0n293,s1n293,notn293;
or (n293,s0n293,s1n293);
not(notn293,n18);
and (s0n293,notn293,1'b0);
and (s1n293,n18,n59);
xor (n294,n58,n60);
nand (n295,n292,n156);
nor (n296,n297,n299);
and (n297,n191,n298);
not (n298,n292);
and (n299,n184,n292);
nor (n300,n301,n302);
and (n301,n210,n191);
and (n302,n214,n184);
or (n303,n304,n289);
nor (n304,n305,n309);
and (n305,n306,n191);
wire s0n306,s1n306,notn306;
or (n306,s0n306,s1n306);
not(notn306,n127);
and (s0n306,notn306,n307);
and (s1n306,n127,n308);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n18);
and (s0n307,notn307,1'b0);
and (s1n307,n18,n107);
xor (n308,n106,n108);
and (n309,n310,n184);
not (n310,n306);
xor (n311,n312,n318);
nand (n312,n313,n317);
or (n313,n314,n131);
nor (n314,n315,n316);
and (n315,n160,n87);
and (n316,n164,n88);
or (n317,n85,n132);
nor (n318,n319,n79);
nor (n319,n320,n323);
and (n320,n236,n321);
not (n321,n322);
and (n322,n81,n253);
and (n323,n257,n80);
and (n324,n280,n286);
and (n325,n8,n177);
xor (n326,n327,n358);
xor (n327,n328,n355);
xor (n328,n329,n342);
nand (n329,n330,n331);
or (n330,n135,n131);
or (n331,n332,n132);
nor (n332,n333,n340);
and (n333,n87,n334);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n127);
and (s0n334,notn334,n335);
and (s1n334,n127,n337);
wire s0n335,s1n335,notn335;
or (n335,s0n335,s1n335);
not(notn335,n18);
and (s0n335,notn335,1'b0);
and (s1n335,n18,n336);
xor (n337,n338,n339);
not (n338,n336);
and (n339,n141,n142);
and (n340,n341,n88);
not (n341,n334);
nor (n342,n343,n348);
nor (n343,n344,n347);
and (n344,n79,n345);
not (n345,n346);
and (n346,n81,n14);
and (n347,n78,n80);
not (n348,n349);
wire s0n349,s1n349,notn349;
or (n349,s0n349,s1n349);
not(notn349,n71);
and (s0n349,notn349,n350);
and (s1n349,n71,n352);
wire s0n350,s1n350,notn350;
or (n350,s0n350,s1n350);
not(notn350,n18);
and (s0n350,notn350,1'b0);
and (s1n350,n18,n351);
xor (n352,n353,n354);
not (n353,n351);
and (n354,n35,n36);
or (n355,n356,n357);
and (n356,n9,n145);
and (n357,n10,n83);
or (n358,n359,n360);
and (n359,n178,n249);
and (n360,n179,n215);
xor (n361,n362,n417);
xor (n362,n363,n397);
xor (n363,n364,n384);
xor (n364,n365,n378);
nand (n365,n366,n374);
or (n366,n288,n367);
nor (n367,n368,n372);
and (n368,n369,n191);
wire s0n369,s1n369,notn369;
or (n369,s0n369,s1n369);
not(notn369,n127);
and (s0n369,notn369,n370);
and (s1n369,n127,n371);
wire s0n370,s1n370,notn370;
or (n370,s0n370,s1n370);
not(notn370,n18);
and (s0n370,notn370,1'b0);
and (s1n370,n18,n104);
xor (n371,n103,n105);
and (n372,n373,n184);
not (n373,n369);
or (n374,n375,n289);
nor (n375,n376,n377);
and (n376,n172,n191);
and (n377,n176,n184);
nand (n378,n379,n380);
or (n379,n266,n258);
or (n380,n381,n251);
nor (n381,n382,n383);
and (n382,n244,n79);
and (n383,n248,n74);
nand (n384,n385,n389);
or (n385,n11,n386);
nor (n386,n387,n388);
and (n387,n272,n348);
and (n388,n276,n349);
or (n389,n390,n394);
or (n390,n391,n12);
nor (n391,n392,n393);
and (n392,n348,n14);
and (n393,n78,n349);
nor (n394,n395,n396);
and (n395,n349,n80);
and (n396,n348,n81);
xor (n397,n398,n411);
xor (n398,n399,n405);
nand (n399,n400,n401);
or (n400,n166,n154);
or (n401,n147,n402);
nor (n402,n403,n404);
and (n403,n156,n91);
and (n404,n130,n157);
nand (n405,n406,n407);
or (n406,n181,n208);
or (n407,n182,n408);
nor (n408,n409,n410);
and (n409,n306,n199);
and (n410,n310,n195);
nand (n411,n412,n413);
or (n412,n225,n238);
or (n413,n414,n217);
nor (n414,n415,n416);
and (n415,n236,n202);
and (n416,n228,n206);
or (n417,n418,n446);
and (n418,n419,n424);
xor (n419,n420,n423);
nand (n420,n421,n422);
or (n421,n288,n304);
or (n422,n289,n367);
and (n423,n312,n318);
or (n424,n425,n445);
and (n425,n426,n439);
xor (n426,n427,n433);
nand (n427,n428,n432);
or (n428,n166,n429);
nor (n429,n430,n431);
and (n430,n369,n156);
and (n431,n373,n157);
or (n432,n147,n170);
nand (n433,n434,n438);
or (n434,n181,n435);
nor (n435,n436,n437);
and (n436,n232,n199);
and (n437,n231,n195);
or (n438,n200,n182);
nand (n439,n440,n444);
or (n440,n238,n441);
nor (n441,n442,n443);
and (n442,n260,n236);
and (n443,n264,n228);
or (n444,n242,n217);
and (n445,n427,n433);
and (n446,n420,n423);
and (n447,n5,n326);
xor (n448,n449,n530);
xor (n449,n450,n490);
xor (n450,n451,n487);
xor (n451,n452,n484);
xor (n452,n453,n478);
xor (n453,n454,n465);
nor (n454,n455,n80);
not (n455,n456);
nand (n456,n457,n464);
or (n457,n348,n458);
wire s0n458,s1n458,notn458;
or (n458,s0n458,s1n458);
not(notn458,n71);
and (s0n458,notn458,n459);
and (s1n458,n71,n461);
wire s0n459,s1n459,notn459;
or (n459,s0n459,s1n459);
not(notn459,n18);
and (s0n459,notn459,1'b0);
and (s1n459,n18,n460);
xor (n461,n462,n463);
not (n462,n460);
and (n463,n353,n354);
nand (n464,n348,n458);
nand (n465,n466,n467);
or (n466,n332,n131);
or (n467,n468,n132);
nor (n468,n469,n476);
and (n469,n470,n87);
wire s0n470,s1n470,notn470;
or (n470,s0n470,s1n470);
not(notn470,n127);
and (s0n470,notn470,n471);
and (s1n470,n127,n473);
wire s0n471,s1n471,notn471;
or (n471,s0n471,s1n471);
not(notn471,n18);
and (s0n471,notn471,1'b0);
and (s1n471,n18,n472);
xor (n473,n474,n475);
not (n474,n472);
and (n475,n338,n339);
and (n476,n477,n88);
not (n477,n470);
nand (n478,n479,n480);
or (n479,n166,n402);
or (n480,n147,n481);
nor (n481,n482,n483);
and (n482,n137,n156);
and (n483,n144,n157);
or (n484,n485,n486);
and (n485,n398,n411);
and (n486,n399,n405);
or (n487,n488,n489);
and (n488,n364,n384);
and (n489,n365,n378);
xor (n490,n491,n527);
xor (n491,n492,n507);
xor (n492,n493,n506);
xor (n493,n494,n500);
nand (n494,n495,n496);
or (n495,n266,n381);
or (n496,n497,n251);
nor (n497,n498,n499);
and (n498,n79,n232);
and (n499,n74,n231);
nand (n500,n501,n502);
or (n501,n390,n386);
or (n502,n503,n11);
nor (n503,n504,n505);
and (n504,n260,n348);
and (n505,n264,n349);
and (n506,n329,n342);
xor (n507,n508,n521);
xor (n508,n509,n515);
nand (n509,n510,n511);
or (n510,n181,n408);
or (n511,n512,n182);
nor (n512,n513,n514);
and (n513,n369,n199);
and (n514,n373,n195);
nand (n515,n516,n517);
or (n516,n238,n414);
or (n517,n518,n217);
nor (n518,n519,n520);
and (n519,n236,n210);
and (n520,n228,n214);
nand (n521,n522,n526);
or (n522,n289,n523);
nor (n523,n524,n525);
and (n524,n160,n191);
and (n525,n164,n184);
or (n526,n288,n375);
or (n527,n528,n529);
and (n528,n327,n358);
and (n529,n328,n355);
or (n530,n531,n532);
and (n531,n362,n417);
and (n532,n363,n397);
nand (n533,n534,n906,n908);
or (n534,n535,n901);
nand (n535,n536,n890);
or (n536,n537,n889);
and (n537,n538,n659);
xor (n538,n539,n644);
or (n539,n540,n643);
and (n540,n541,n609);
xor (n541,n542,n564);
xor (n542,n543,n558);
xor (n543,n544,n551);
nand (n544,n545,n550);
or (n545,n181,n546);
not (n546,n547);
nor (n547,n548,n549);
and (n548,n199,n248);
and (n549,n244,n195);
or (n550,n435,n182);
nand (n551,n552,n557);
or (n552,n553,n238);
not (n553,n554);
nand (n554,n555,n556);
or (n555,n276,n228);
or (n556,n272,n236);
or (n557,n441,n217);
nand (n558,n559,n563);
or (n559,n288,n560);
nor (n560,n561,n562);
and (n561,n202,n191);
and (n562,n206,n184);
or (n563,n289,n300);
or (n564,n565,n608);
and (n565,n566,n588);
xor (n566,n567,n573);
nand (n567,n568,n572);
or (n568,n288,n569);
nor (n569,n570,n571);
and (n570,n232,n191);
and (n571,n231,n184);
or (n572,n560,n289);
xor (n573,n574,n580);
nor (n574,n575,n236);
nor (n575,n576,n579);
and (n576,n577,n199);
not (n577,n578);
and (n578,n81,n220);
and (n579,n224,n80);
nand (n580,n581,n584);
or (n581,n131,n582);
not (n582,n583);
xnor (n583,n369,n87);
or (n584,n585,n132);
nor (n585,n586,n587);
and (n586,n87,n172);
and (n587,n176,n88);
or (n588,n589,n607);
and (n589,n590,n598);
xor (n590,n591,n592);
nor (n591,n217,n80);
nand (n592,n593,n594);
or (n593,n132,n582);
or (n594,n595,n131);
nor (n595,n596,n597);
and (n596,n87,n306);
and (n597,n310,n88);
nand (n598,n599,n603);
or (n599,n181,n600);
nor (n600,n601,n602);
and (n601,n272,n199);
and (n602,n276,n195);
or (n603,n604,n182);
nor (n604,n605,n606);
and (n605,n260,n199);
and (n606,n264,n195);
and (n607,n591,n592);
and (n608,n567,n573);
xor (n609,n610,n624);
xor (n610,n611,n612);
and (n611,n574,n580);
xor (n612,n613,n618);
xor (n613,n614,n615);
nor (n614,n251,n80);
nand (n615,n616,n617);
or (n616,n585,n131);
or (n617,n314,n132);
nand (n618,n619,n623);
or (n619,n166,n620);
nor (n620,n621,n622);
and (n621,n306,n156);
and (n622,n310,n157);
or (n623,n147,n429);
or (n624,n625,n642);
and (n625,n626,n636);
xor (n626,n627,n633);
nand (n627,n628,n632);
or (n628,n166,n629);
nor (n629,n630,n631);
and (n630,n156,n210);
and (n631,n214,n157);
or (n632,n620,n147);
nand (n633,n634,n635);
or (n634,n182,n546);
or (n635,n604,n181);
nand (n636,n637,n638);
or (n637,n217,n553);
or (n638,n238,n639);
nor (n639,n640,n641);
and (n640,n228,n80);
and (n641,n236,n81);
and (n642,n627,n633);
and (n643,n542,n564);
xor (n644,n645,n650);
xor (n645,n646,n647);
xor (n646,n426,n439);
or (n647,n648,n649);
and (n648,n610,n624);
and (n649,n611,n612);
xor (n650,n651,n658);
xor (n651,n652,n655);
or (n652,n653,n654);
and (n653,n613,n618);
and (n654,n614,n615);
or (n655,n656,n657);
and (n656,n543,n558);
and (n657,n544,n551);
xor (n658,n279,n311);
or (n659,n660,n888);
and (n660,n661,n698);
xor (n661,n662,n697);
or (n662,n663,n696);
and (n663,n664,n695);
xor (n664,n665,n694);
or (n665,n666,n693);
and (n666,n667,n680);
xor (n667,n668,n674);
nand (n668,n669,n673);
or (n669,n166,n670);
nor (n670,n671,n672);
and (n671,n202,n156);
and (n672,n157,n206);
or (n673,n629,n147);
nand (n674,n675,n679);
or (n675,n288,n676);
nor (n676,n677,n678);
and (n677,n244,n191);
and (n678,n248,n184);
or (n679,n569,n289);
and (n680,n681,n687);
nor (n681,n682,n199);
nor (n682,n683,n686);
and (n683,n684,n191);
not (n684,n685);
and (n685,n81,n187);
and (n686,n192,n80);
nand (n687,n688,n692);
or (n688,n689,n131);
nor (n689,n690,n691);
and (n690,n87,n210);
and (n691,n214,n88);
or (n692,n595,n132);
and (n693,n668,n674);
xor (n694,n626,n636);
xor (n695,n566,n588);
and (n696,n665,n694);
xor (n697,n541,n609);
nand (n698,n699,n885,n887);
or (n699,n700,n758);
nand (n700,n701,n753);
not (n701,n702);
nor (n702,n703,n729);
xor (n703,n704,n728);
xor (n704,n705,n727);
or (n705,n706,n726);
and (n706,n707,n720);
xor (n707,n708,n714);
nand (n708,n709,n713);
or (n709,n181,n710);
nor (n710,n711,n712);
and (n711,n195,n80);
and (n712,n199,n81);
or (n713,n600,n182);
nand (n714,n715,n719);
or (n715,n716,n166);
nor (n716,n717,n718);
and (n717,n157,n231);
and (n718,n156,n232);
or (n719,n670,n147);
nand (n720,n721,n725);
or (n721,n288,n722);
nor (n722,n723,n724);
and (n723,n260,n191);
and (n724,n264,n184);
or (n725,n676,n289);
and (n726,n708,n714);
xor (n727,n590,n598);
xor (n728,n667,n680);
or (n729,n730,n752);
and (n730,n731,n751);
xor (n731,n732,n733);
xor (n732,n681,n687);
or (n733,n734,n750);
and (n734,n735,n744);
xor (n735,n736,n737);
nor (n736,n182,n80);
nand (n737,n738,n743);
or (n738,n739,n131);
not (n739,n740);
nand (n740,n741,n742);
or (n741,n88,n206);
nand (n742,n206,n88);
or (n743,n689,n132);
nand (n744,n745,n749);
or (n745,n166,n746);
nor (n746,n747,n748);
and (n747,n156,n244);
and (n748,n157,n248);
or (n749,n716,n147);
and (n750,n736,n737);
xor (n751,n707,n720);
and (n752,n732,n733);
or (n753,n754,n755);
xor (n754,n664,n695);
or (n755,n756,n757);
and (n756,n704,n728);
and (n757,n705,n727);
nor (n758,n759,n884);
and (n759,n760,n879);
or (n760,n761,n878);
and (n761,n762,n803);
xor (n762,n763,n796);
or (n763,n764,n795);
and (n764,n765,n781);
xor (n765,n766,n772);
nand (n766,n767,n771);
or (n767,n166,n768);
nor (n768,n769,n770);
and (n769,n157,n264);
and (n770,n156,n260);
or (n771,n746,n147);
or (n772,n773,n777);
nor (n773,n774,n289);
nor (n774,n775,n776);
and (n775,n191,n272);
and (n776,n184,n276);
nor (n777,n288,n778);
nor (n778,n779,n780);
and (n779,n184,n80);
and (n780,n191,n81);
xor (n781,n782,n788);
nor (n782,n783,n191);
nor (n783,n784,n787);
and (n784,n785,n156);
not (n785,n786);
and (n786,n81,n292);
and (n787,n298,n80);
nand (n788,n789,n794);
or (n789,n131,n790);
not (n790,n791);
nand (n791,n792,n793);
or (n792,n87,n232);
nand (n793,n232,n87);
nand (n794,n740,n133);
and (n795,n766,n772);
xor (n796,n797,n802);
xor (n797,n798,n801);
nand (n798,n799,n800);
or (n799,n288,n774);
or (n800,n722,n289);
and (n801,n782,n788);
xor (n802,n735,n744);
or (n803,n804,n877);
and (n804,n805,n825);
xor (n805,n806,n824);
or (n806,n807,n823);
and (n807,n808,n817);
xor (n808,n809,n810);
and (n809,n290,n81);
nand (n810,n811,n816);
or (n811,n131,n812);
not (n812,n813);
nand (n813,n814,n815);
or (n814,n88,n248);
nand (n815,n248,n88);
nand (n816,n791,n133);
nand (n817,n818,n822);
or (n818,n166,n819);
nor (n819,n820,n821);
and (n820,n156,n272);
and (n821,n157,n276);
or (n822,n768,n147);
and (n823,n809,n810);
xor (n824,n765,n781);
or (n825,n826,n876);
and (n826,n827,n844);
xor (n827,n828,n843);
and (n828,n829,n835);
and (n829,n830,n157);
nand (n830,n831,n834);
nand (n831,n832,n87);
not (n832,n833);
and (n833,n81,n149);
nand (n834,n153,n80);
nand (n835,n836,n837);
or (n836,n132,n812);
nand (n837,n838,n842);
not (n838,n839);
nor (n839,n840,n841);
and (n840,n264,n88);
and (n841,n260,n87);
not (n842,n131);
xor (n843,n808,n817);
or (n844,n845,n875);
and (n845,n846,n854);
xor (n846,n847,n853);
nand (n847,n848,n852);
or (n848,n166,n849);
nor (n849,n850,n851);
and (n850,n157,n80);
and (n851,n156,n81);
or (n852,n819,n147);
xor (n853,n829,n835);
or (n854,n855,n874);
and (n855,n856,n864);
xor (n856,n857,n858);
nor (n857,n147,n80);
nand (n858,n859,n863);
or (n859,n860,n131);
or (n860,n861,n862);
and (n861,n87,n276);
and (n862,n272,n88);
or (n863,n839,n132);
nor (n864,n865,n872);
nor (n865,n866,n868);
and (n866,n867,n133);
not (n867,n860);
and (n868,n869,n842);
nand (n869,n870,n871);
or (n870,n87,n81);
or (n871,n88,n80);
or (n872,n87,n873);
and (n873,n81,n133);
and (n874,n857,n858);
and (n875,n847,n853);
and (n876,n828,n843);
and (n877,n806,n824);
and (n878,n763,n796);
or (n879,n880,n881);
xor (n880,n731,n751);
or (n881,n882,n883);
and (n882,n797,n802);
and (n883,n798,n801);
and (n884,n880,n881);
nand (n885,n753,n886);
and (n886,n703,n729);
nand (n887,n754,n755);
and (n888,n662,n697);
and (n889,n539,n644);
or (n890,n891,n898);
xor (n891,n892,n897);
xor (n892,n893,n894);
xor (n893,n419,n424);
or (n894,n895,n896);
and (n895,n651,n658);
and (n896,n652,n655);
xor (n897,n7,n277);
or (n898,n899,n900);
and (n899,n645,n650);
and (n900,n646,n647);
nor (n901,n902,n903);
xor (n902,n4,n361);
or (n903,n904,n905);
and (n904,n892,n897);
and (n905,n893,n894);
or (n906,n901,n907);
nand (n907,n891,n898);
nand (n908,n902,n903);
xor (n909,n910,n1449);
xor (n910,n911,n1446);
xor (n911,n912,n1445);
xor (n912,n913,n1437);
xor (n913,n914,n1436);
xor (n914,n915,n1421);
xor (n915,n916,n1420);
xor (n916,n917,n1400);
xor (n917,n918,n1399);
xor (n918,n919,n1372);
xor (n919,n920,n1371);
xor (n920,n921,n1339);
xor (n921,n922,n1338);
xor (n922,n923,n1300);
xor (n923,n924,n1299);
xor (n924,n925,n1255);
xor (n925,n926,n1254);
xor (n926,n927,n1203);
xor (n927,n928,n1202);
xor (n928,n929,n1146);
xor (n929,n930,n1145);
xor (n930,n931,n1082);
xor (n931,n932,n1081);
xor (n932,n933,n1013);
xor (n933,n934,n1012);
xor (n934,n935,n938);
xor (n935,n936,n937);
and (n936,n470,n133);
and (n937,n334,n88);
or (n938,n939,n942);
and (n939,n940,n941);
and (n940,n334,n133);
and (n941,n137,n88);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
and (n946,n137,n133);
and (n947,n91,n88);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
and (n952,n91,n133);
and (n953,n160,n88);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n960);
and (n957,n958,n959);
and (n958,n160,n133);
and (n959,n172,n88);
and (n960,n961,n962);
xor (n961,n958,n959);
or (n962,n963,n966);
and (n963,n964,n965);
and (n964,n172,n133);
and (n965,n369,n88);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n972);
and (n969,n970,n971);
and (n970,n369,n133);
and (n971,n306,n88);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
and (n976,n306,n133);
and (n977,n210,n88);
and (n978,n979,n980);
xor (n979,n976,n977);
or (n980,n981,n984);
and (n981,n982,n983);
and (n982,n210,n133);
and (n983,n202,n88);
and (n984,n985,n986);
xor (n985,n982,n983);
or (n986,n987,n990);
and (n987,n988,n989);
and (n988,n202,n133);
and (n989,n232,n88);
and (n990,n991,n992);
xor (n991,n988,n989);
or (n992,n993,n996);
and (n993,n994,n995);
and (n994,n232,n133);
and (n995,n244,n88);
and (n996,n997,n998);
xor (n997,n994,n995);
or (n998,n999,n1002);
and (n999,n1000,n1001);
and (n1000,n244,n133);
and (n1001,n260,n88);
and (n1002,n1003,n1004);
xor (n1003,n1000,n1001);
or (n1004,n1005,n1007);
and (n1005,n1006,n862);
and (n1006,n260,n133);
and (n1007,n1008,n1009);
xor (n1008,n1006,n862);
and (n1009,n1010,n1011);
and (n1010,n272,n133);
and (n1011,n81,n88);
and (n1012,n137,n149);
or (n1013,n1014,n1017);
and (n1014,n1015,n1016);
xor (n1015,n943,n944);
and (n1016,n91,n149);
and (n1017,n1018,n1019);
xor (n1018,n1015,n1016);
or (n1019,n1020,n1023);
and (n1020,n1021,n1022);
xor (n1021,n949,n950);
and (n1022,n160,n149);
and (n1023,n1024,n1025);
xor (n1024,n1021,n1022);
or (n1025,n1026,n1029);
and (n1026,n1027,n1028);
xor (n1027,n955,n956);
and (n1028,n172,n149);
and (n1029,n1030,n1031);
xor (n1030,n1027,n1028);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
xor (n1033,n961,n962);
and (n1034,n369,n149);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
xor (n1039,n967,n968);
and (n1040,n306,n149);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1047);
and (n1044,n1045,n1046);
xor (n1045,n973,n974);
and (n1046,n210,n149);
and (n1047,n1048,n1049);
xor (n1048,n1045,n1046);
or (n1049,n1050,n1053);
and (n1050,n1051,n1052);
xor (n1051,n979,n980);
and (n1052,n202,n149);
and (n1053,n1054,n1055);
xor (n1054,n1051,n1052);
or (n1055,n1056,n1059);
and (n1056,n1057,n1058);
xor (n1057,n985,n986);
and (n1058,n232,n149);
and (n1059,n1060,n1061);
xor (n1060,n1057,n1058);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n991,n992);
and (n1064,n244,n149);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n997,n998);
and (n1070,n260,n149);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n1003,n1004);
and (n1076,n272,n149);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
and (n1079,n1080,n833);
xor (n1080,n1008,n1009);
and (n1081,n91,n157);
or (n1082,n1083,n1086);
and (n1083,n1084,n1085);
xor (n1084,n1018,n1019);
and (n1085,n160,n157);
and (n1086,n1087,n1088);
xor (n1087,n1084,n1085);
or (n1088,n1089,n1092);
and (n1089,n1090,n1091);
xor (n1090,n1024,n1025);
and (n1091,n172,n157);
and (n1092,n1093,n1094);
xor (n1093,n1090,n1091);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
xor (n1096,n1030,n1031);
and (n1097,n369,n157);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
xor (n1102,n1036,n1037);
and (n1103,n306,n157);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1042,n1043);
and (n1109,n210,n157);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1048,n1049);
and (n1115,n202,n157);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1054,n1055);
and (n1121,n232,n157);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1060,n1061);
and (n1127,n244,n157);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1066,n1067);
and (n1133,n260,n157);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1072,n1073);
and (n1139,n272,n157);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
and (n1142,n1143,n1144);
xor (n1143,n1078,n1079);
and (n1144,n81,n157);
and (n1145,n160,n292);
or (n1146,n1147,n1150);
and (n1147,n1148,n1149);
xor (n1148,n1087,n1088);
and (n1149,n172,n292);
and (n1150,n1151,n1152);
xor (n1151,n1148,n1149);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
xor (n1154,n1093,n1094);
and (n1155,n369,n292);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
xor (n1160,n1099,n1100);
and (n1161,n306,n292);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
xor (n1166,n1105,n1106);
and (n1167,n210,n292);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1111,n1112);
and (n1173,n202,n292);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1117,n1118);
and (n1179,n232,n292);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1123,n1124);
and (n1185,n244,n292);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1129,n1130);
and (n1191,n260,n292);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1135,n1136);
and (n1197,n272,n292);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
and (n1200,n1201,n786);
xor (n1201,n1141,n1142);
and (n1202,n172,n184);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1151,n1152);
and (n1206,n369,n184);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1157,n1158);
and (n1212,n306,n184);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1163,n1164);
and (n1218,n210,n184);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1169,n1170);
and (n1224,n202,n184);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1175,n1176);
and (n1230,n232,n184);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1181,n1182);
and (n1236,n244,n184);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1187,n1188);
and (n1242,n260,n184);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1193,n1194);
and (n1248,n272,n184);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
and (n1251,n1252,n1253);
xor (n1252,n1199,n1200);
and (n1253,n81,n184);
and (n1254,n369,n187);
or (n1255,n1256,n1259);
and (n1256,n1257,n1258);
xor (n1257,n1208,n1209);
and (n1258,n306,n187);
and (n1259,n1260,n1261);
xor (n1260,n1257,n1258);
or (n1261,n1262,n1265);
and (n1262,n1263,n1264);
xor (n1263,n1214,n1215);
and (n1264,n210,n187);
and (n1265,n1266,n1267);
xor (n1266,n1263,n1264);
or (n1267,n1268,n1271);
and (n1268,n1269,n1270);
xor (n1269,n1220,n1221);
and (n1270,n202,n187);
and (n1271,n1272,n1273);
xor (n1272,n1269,n1270);
or (n1273,n1274,n1277);
and (n1274,n1275,n1276);
xor (n1275,n1226,n1227);
and (n1276,n232,n187);
and (n1277,n1278,n1279);
xor (n1278,n1275,n1276);
or (n1279,n1280,n1283);
and (n1280,n1281,n1282);
xor (n1281,n1232,n1233);
and (n1282,n244,n187);
and (n1283,n1284,n1285);
xor (n1284,n1281,n1282);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1238,n1239);
and (n1288,n260,n187);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1244,n1245);
and (n1294,n272,n187);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
and (n1297,n1298,n685);
xor (n1298,n1250,n1251);
and (n1299,n306,n195);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1260,n1261);
and (n1303,n210,n195);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1266,n1267);
and (n1309,n202,n195);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1272,n1273);
and (n1315,n232,n195);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1321);
and (n1319,n1320,n549);
xor (n1320,n1278,n1279);
and (n1321,n1322,n1323);
xor (n1322,n1320,n549);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1284,n1285);
and (n1326,n260,n195);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1290,n1291);
and (n1332,n272,n195);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
and (n1335,n1336,n1337);
xor (n1336,n1296,n1297);
and (n1337,n81,n195);
and (n1338,n210,n220);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1305,n1306);
and (n1342,n202,n220);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
xor (n1347,n1311,n1312);
and (n1348,n232,n220);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
xor (n1353,n1317,n1318);
and (n1354,n244,n220);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1322,n1323);
and (n1360,n260,n220);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1328,n1329);
and (n1366,n272,n220);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
and (n1369,n1370,n578);
xor (n1370,n1334,n1335);
and (n1371,n202,n228);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1344,n1345);
and (n1375,n232,n228);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1350,n1351);
and (n1381,n244,n228);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1356,n1357);
and (n1387,n260,n228);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1362,n1363);
and (n1393,n272,n228);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
and (n1396,n1397,n1398);
xor (n1397,n1368,n1369);
and (n1398,n81,n228);
and (n1399,n232,n253);
or (n1400,n1401,n1404);
and (n1401,n1402,n1403);
xor (n1402,n1377,n1378);
and (n1403,n244,n253);
and (n1404,n1405,n1406);
xor (n1405,n1402,n1403);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1383,n1384);
and (n1409,n260,n253);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1389,n1390);
and (n1415,n272,n253);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
and (n1418,n1419,n322);
xor (n1419,n1395,n1396);
and (n1420,n244,n74);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1405,n1406);
and (n1424,n260,n74);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1411,n1412);
and (n1430,n272,n74);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
and (n1433,n1434,n1435);
xor (n1434,n1417,n1418);
and (n1435,n81,n74);
and (n1436,n260,n14);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1426,n1427);
and (n1440,n272,n14);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
and (n1443,n1444,n346);
xor (n1444,n1432,n1433);
and (n1445,n272,n349);
and (n1446,n1447,n1448);
xor (n1447,n1442,n1443);
and (n1448,n81,n349);
and (n1449,n81,n458);
endmodule
