module top (out,n20,n21,n22,n24,n25,n31,n32,n38,n39
        ,n50,n51,n56,n57,n62,n73,n74,n82,n94,n95
        ,n103,n114,n148,n221,n226,n227,n261,n273,n331,n370
        ,n476,n482,n491,n501,n507);
output out;
input n20;
input n21;
input n22;
input n24;
input n25;
input n31;
input n32;
input n38;
input n39;
input n50;
input n51;
input n56;
input n57;
input n62;
input n73;
input n74;
input n82;
input n94;
input n95;
input n103;
input n114;
input n148;
input n221;
input n226;
input n227;
input n261;
input n273;
input n331;
input n370;
input n476;
input n482;
input n491;
input n501;
input n507;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
xor (out,n0,n1031);
nand (n0,n1,n973);
nand (n1,n2,n22);
nor (n2,n3,n970);
and (n3,n4,n187);
nor (n4,n5,n186);
and (n5,n6,n165);
not (n6,n7);
or (n7,n8,n164);
and (n8,n9,n124);
xor (n9,n10,n85);
or (n10,n11,n84);
and (n11,n12,n70);
xor (n12,n13,n42);
nand (n13,n14,n34);
or (n14,n15,n28);
and (n15,n16,n27);
nand (n16,n17,n26);
or (n17,n18,n23);
not (n18,n19);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,n20);
and (s1n19,n22,n21);
wire s0n23,s1n23,notn23;
or (n23,s0n23,s1n23);
not(notn23,n22);
and (s0n23,notn23,n24);
and (s1n23,n22,n25);
nand (n26,n23,n18);
not (n27,n28);
nand (n28,n29,n33);
or (n29,n18,n30);
wire s0n30,s1n30,notn30;
or (n30,s0n30,s1n30);
not(notn30,n22);
and (s0n30,notn30,n31);
and (s1n30,n22,n32);
nand (n33,n30,n18);
nand (n34,n35,n40);
or (n35,n23,n36);
not (n36,n37);
and (n37,n38,n39);
or (n40,n41,n37);
not (n41,n23);
nand (n42,n43,n65);
or (n43,n44,n59);
nand (n44,n45,n53);
not (n45,n46);
nand (n46,n47,n52);
or (n47,n48,n23);
not (n48,n49);
wire s0n49,s1n49,notn49;
or (n49,s0n49,s1n49);
not(notn49,n22);
and (s0n49,notn49,n50);
and (s1n49,n22,n51);
nand (n52,n23,n48);
nand (n53,n54,n58);
or (n54,n48,n55);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n22);
and (s0n55,notn55,n56);
and (s1n55,n22,n57);
nand (n58,n55,n48);
nor (n59,n60,n63);
and (n60,n61,n62);
not (n61,n55);
and (n63,n55,n64);
not (n64,n62);
or (n65,n45,n66);
nor (n66,n67,n68);
and (n67,n61,n39);
and (n68,n55,n69);
not (n69,n39);
nor (n70,n71,n79);
nand (n71,n72,n75);
wire s0n72,s1n72,notn72;
or (n72,s0n72,s1n72);
not(notn72,n22);
and (s0n72,notn72,n73);
and (s1n72,n22,n74);
not (n75,n76);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n22);
and (s0n76,notn76,1'b0);
and (s1n76,n22,n78);
and (n78,n38,n74);
nor (n79,n80,n83);
and (n80,n76,n81);
not (n81,n82);
and (n83,n75,n82);
and (n84,n13,n42);
xor (n85,n86,n116);
xor (n86,n87,n110);
nand (n87,n88,n106);
or (n88,n89,n100);
nand (n89,n90,n97);
nor (n90,n91,n96);
and (n91,n92,n55);
not (n92,n93);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n22);
and (s0n93,notn93,n94);
and (s1n93,n22,n95);
and (n96,n93,n61);
nand (n97,n98,n99);
or (n98,n92,n72);
nand (n99,n72,n92);
nor (n100,n101,n104);
and (n101,n102,n103);
not (n102,n72);
and (n104,n72,n105);
not (n105,n103);
or (n106,n90,n107);
nor (n107,n108,n109);
and (n108,n102,n62);
and (n109,n72,n64);
nor (n110,n71,n111);
nor (n111,n112,n115);
and (n112,n76,n113);
not (n113,n114);
and (n115,n75,n114);
nor (n116,n117,n120);
and (n117,n118,n119);
not (n118,n44);
not (n119,n66);
and (n120,n46,n121);
nand (n121,n122,n123);
or (n122,n55,n36);
or (n123,n61,n37);
or (n124,n125,n163);
and (n125,n126,n141);
xor (n126,n127,n133);
nand (n127,n128,n132);
or (n128,n89,n129);
nor (n129,n130,n131);
and (n130,n102,n114);
and (n131,n72,n113);
or (n132,n90,n100);
nand (n133,n134,n136);
or (n134,n135,n27);
not (n135,n34);
nand (n136,n137,n15);
not (n137,n138);
nor (n138,n139,n140);
and (n139,n41,n39);
and (n140,n23,n69);
or (n141,n142,n162);
and (n142,n143,n156);
xor (n143,n144,n150);
nor (n144,n71,n145);
nor (n145,n146,n149);
and (n146,n76,n147);
not (n147,n148);
and (n149,n75,n148);
nand (n150,n151,n155);
or (n151,n44,n152);
nor (n152,n153,n154);
and (n153,n103,n61);
and (n154,n105,n55);
or (n155,n45,n59);
nand (n156,n157,n161);
or (n157,n89,n158);
nor (n158,n159,n160);
and (n159,n102,n82);
and (n160,n72,n81);
or (n161,n90,n129);
and (n162,n144,n150);
and (n163,n127,n133);
and (n164,n10,n85);
not (n165,n166);
xor (n166,n167,n183);
xor (n167,n168,n169);
not (n168,n116);
xor (n169,n170,n179);
xor (n170,n171,n173);
nand (n171,n172,n121);
or (n172,n118,n46);
nand (n173,n174,n175);
or (n174,n89,n107);
or (n175,n90,n176);
nor (n176,n177,n178);
and (n177,n102,n39);
and (n178,n72,n69);
nor (n179,n71,n180);
nor (n180,n181,n182);
and (n181,n76,n105);
and (n182,n75,n103);
or (n183,n184,n185);
and (n184,n86,n116);
and (n185,n87,n110);
nor (n186,n6,n165);
nand (n187,n188,n969);
or (n188,n189,n244);
nor (n189,n190,n243);
or (n190,n191,n242);
and (n191,n192,n195);
xor (n192,n193,n194);
xor (n193,n12,n70);
xor (n194,n126,n141);
or (n195,n196,n241);
and (n196,n197,n214);
xor (n197,n198,n199);
not (n198,n133);
or (n199,n200,n206);
nand (n200,n201,n205);
or (n201,n89,n202);
nor (n202,n203,n204);
and (n203,n102,n148);
and (n204,n72,n147);
or (n205,n90,n158);
nand (n206,n207,n213);
or (n207,n208,n209);
not (n208,n15);
not (n209,n210);
nand (n210,n211,n212);
or (n211,n23,n64);
or (n212,n41,n62);
or (n213,n27,n138);
or (n214,n215,n240);
and (n215,n216,n234);
xor (n216,n217,n223);
nor (n217,n71,n218);
nor (n218,n219,n222);
and (n219,n76,n220);
not (n220,n221);
and (n222,n75,n221);
nand (n223,n224,n230);
or (n224,n225,n228);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n22);
and (s0n225,notn225,n226);
and (s1n225,n22,n227);
nor (n228,n229,n225);
not (n229,n30);
not (n230,n231);
nor (n231,n232,n233);
and (n232,n229,n37);
and (n233,n30,n36);
nand (n234,n235,n236);
or (n235,n152,n45);
or (n236,n44,n237);
nor (n237,n238,n239);
and (n238,n61,n114);
and (n239,n55,n113);
and (n240,n217,n223);
and (n241,n198,n199);
and (n242,n193,n194);
xor (n243,n9,n124);
not (n244,n245);
nand (n245,n246,n956);
or (n246,n247,n454);
not (n247,n248);
and (n248,n249,n435,n448);
nor (n249,n250,n412);
nor (n250,n251,n381);
or (n251,n252,n380);
and (n252,n253,n340);
xor (n253,n254,n284);
xor (n254,n255,n275);
xor (n255,n256,n269);
nand (n256,n257,n264);
or (n257,n258,n89);
not (n258,n259);
nor (n259,n260,n262);
and (n260,n261,n72);
and (n262,n263,n102);
not (n263,n261);
nand (n264,n265,n266);
not (n265,n90);
nor (n266,n267,n268);
and (n267,n221,n72);
and (n268,n220,n102);
nor (n269,n71,n270);
nor (n270,n271,n274);
and (n271,n76,n272);
not (n272,n273);
and (n274,n75,n273);
nand (n275,n276,n280);
or (n276,n44,n277);
nor (n277,n278,n279);
and (n278,n61,n148);
and (n279,n55,n147);
or (n280,n45,n281);
nor (n281,n282,n283);
and (n282,n61,n82);
and (n283,n55,n81);
xor (n284,n285,n318);
xor (n285,n286,n305);
xor (n286,n287,n298);
nand (n287,n288,n293);
or (n288,n289,n290);
not (n289,n228);
nor (n290,n291,n292);
and (n291,n229,n62);
and (n292,n30,n64);
or (n293,n294,n297);
nor (n294,n295,n296);
and (n295,n229,n39);
and (n296,n30,n69);
not (n297,n225);
nand (n298,n299,n303);
or (n299,n208,n300);
nor (n300,n301,n302);
and (n301,n41,n114);
and (n302,n23,n113);
or (n303,n304,n27);
xor (n304,n103,n41);
and (n305,n306,n312);
nand (n306,n307,n311);
or (n307,n289,n308);
nor (n308,n309,n310);
and (n309,n229,n103);
and (n310,n30,n105);
or (n311,n290,n297);
nand (n312,n313,n317);
or (n313,n208,n314);
nor (n314,n315,n316);
and (n315,n41,n82);
and (n316,n23,n81);
or (n317,n27,n300);
or (n318,n319,n339);
and (n319,n320,n333);
xor (n320,n321,n327);
nand (n321,n322,n326);
or (n322,n323,n89);
nor (n323,n324,n325);
and (n324,n273,n102);
and (n325,n272,n72);
nand (n326,n265,n259);
nor (n327,n71,n328);
nor (n328,n329,n332);
and (n329,n76,n330);
not (n330,n331);
and (n332,n75,n331);
nand (n333,n334,n338);
or (n334,n44,n335);
nor (n335,n336,n337);
and (n336,n61,n221);
and (n337,n55,n220);
or (n338,n45,n277);
and (n339,n321,n327);
or (n340,n341,n379);
and (n341,n342,n357);
xor (n342,n343,n344);
xor (n343,n306,n312);
and (n344,n345,n351);
nand (n345,n346,n350);
or (n346,n289,n347);
nor (n347,n348,n349);
and (n348,n229,n114);
and (n349,n30,n113);
or (n350,n308,n297);
nand (n351,n352,n356);
or (n352,n208,n353);
nor (n353,n354,n355);
and (n354,n41,n148);
and (n355,n23,n147);
or (n356,n314,n27);
or (n357,n358,n378);
and (n358,n359,n372);
xor (n359,n360,n366);
nand (n360,n361,n365);
or (n361,n89,n362);
nor (n362,n363,n364);
and (n363,n102,n331);
and (n364,n72,n330);
or (n365,n90,n323);
nor (n366,n71,n367);
nor (n367,n368,n371);
and (n368,n76,n369);
not (n369,n370);
and (n371,n75,n370);
nand (n372,n373,n374);
or (n373,n335,n45);
or (n374,n44,n375);
nor (n375,n376,n377);
and (n376,n61,n261);
and (n377,n55,n263);
and (n378,n360,n366);
and (n379,n343,n344);
and (n380,n254,n284);
xor (n381,n382,n409);
xor (n382,n383,n396);
xor (n383,n384,n393);
xor (n384,n385,n389);
nand (n385,n386,n388);
or (n386,n387,n89);
not (n387,n266);
or (n388,n90,n202);
nor (n389,n71,n390);
nor (n390,n391,n392);
and (n391,n76,n263);
and (n392,n75,n261);
nand (n393,n394,n395);
or (n394,n44,n281);
or (n395,n45,n237);
xor (n396,n397,n406);
xor (n397,n398,n405);
xor (n398,n399,n402);
nand (n399,n400,n401);
or (n400,n289,n294);
or (n401,n231,n297);
nand (n402,n403,n404);
or (n403,n304,n208);
nand (n404,n28,n210);
and (n405,n287,n298);
or (n406,n407,n408);
and (n407,n255,n275);
and (n408,n256,n269);
or (n409,n410,n411);
and (n410,n285,n318);
and (n411,n286,n305);
not (n412,n413);
nand (n413,n414,n431);
not (n414,n415);
xor (n415,n416,n421);
xor (n416,n417,n418);
xor (n417,n216,n234);
or (n418,n419,n420);
and (n419,n397,n406);
and (n420,n398,n405);
xor (n421,n422,n427);
xor (n422,n423,n424);
and (n423,n399,n402);
or (n424,n425,n426);
and (n425,n384,n393);
and (n426,n385,n389);
nand (n427,n428,n199);
or (n428,n429,n430);
not (n429,n206);
not (n430,n200);
not (n431,n432);
or (n432,n433,n434);
and (n433,n382,n409);
and (n434,n383,n396);
nand (n435,n436,n438);
not (n436,n437);
xor (n437,n192,n195);
not (n438,n439);
or (n439,n440,n447);
and (n440,n441,n444);
xor (n441,n442,n443);
xor (n442,n143,n156);
xor (n443,n197,n214);
or (n444,n445,n446);
and (n445,n422,n427);
and (n446,n423,n424);
and (n447,n442,n443);
not (n448,n449);
nor (n449,n450,n451);
xor (n450,n441,n444);
or (n451,n452,n453);
and (n452,n416,n421);
and (n453,n417,n418);
not (n454,n455);
nand (n455,n456,n945,n955);
nand (n456,n457,n866);
nand (n457,n458,n722,n865);
nand (n458,n459,n675);
nand (n459,n460,n674);
or (n460,n461,n629);
nor (n461,n462,n628);
and (n462,n463,n600);
not (n463,n464);
nor (n464,n465,n560);
or (n465,n466,n559);
and (n466,n467,n530);
xor (n467,n468,n511);
or (n468,n469,n510);
and (n469,n470,n497);
xor (n470,n471,n485);
nand (n471,n472,n479);
or (n472,n473,n89);
not (n473,n474);
nand (n474,n475,n477);
or (n475,n102,n476);
or (n477,n72,n478);
not (n478,n476);
or (n479,n90,n480);
nor (n480,n481,n483);
and (n481,n482,n102);
and (n483,n484,n72);
not (n484,n482);
nand (n485,n486,n493);
or (n486,n487,n208);
not (n487,n488);
nand (n488,n489,n492);
or (n489,n23,n490);
not (n490,n491);
or (n492,n41,n491);
nand (n493,n28,n494);
nor (n494,n495,n496);
and (n495,n370,n23);
and (n496,n369,n41);
nand (n497,n498,n504);
or (n498,n44,n499);
nor (n499,n500,n502);
and (n500,n61,n501);
and (n502,n55,n503);
not (n503,n501);
or (n504,n45,n505);
nor (n505,n506,n508);
and (n506,n61,n507);
and (n508,n55,n509);
not (n509,n507);
and (n510,n471,n485);
xor (n511,n512,n524);
xor (n512,n513,n515);
and (n513,n514,n476);
not (n514,n71);
nand (n515,n516,n520);
or (n516,n289,n517);
nor (n517,n518,n519);
and (n518,n272,n30);
and (n519,n273,n229);
or (n520,n521,n297);
nor (n521,n522,n523);
and (n522,n229,n261);
and (n523,n30,n263);
nand (n524,n525,n526);
or (n525,n89,n480);
or (n526,n90,n527);
nor (n527,n528,n529);
and (n528,n501,n102);
and (n529,n503,n72);
xor (n530,n531,n545);
xor (n531,n532,n539);
nand (n532,n533,n535);
or (n533,n208,n534);
not (n534,n494);
or (n535,n27,n536);
nor (n536,n537,n538);
and (n537,n41,n331);
and (n538,n23,n330);
nand (n539,n540,n541);
or (n540,n44,n505);
or (n541,n45,n542);
nor (n542,n543,n544);
and (n543,n61,n491);
and (n544,n55,n490);
and (n545,n546,n551);
nor (n546,n547,n102);
nor (n547,n548,n550);
and (n548,n61,n549);
nand (n549,n93,n476);
and (n550,n92,n478);
nand (n551,n552,n557);
or (n552,n553,n289);
not (n553,n554);
nor (n554,n555,n556);
and (n555,n331,n30);
and (n556,n330,n229);
nand (n557,n558,n225);
not (n558,n517);
and (n559,n468,n511);
xor (n560,n561,n583);
xor (n561,n562,n580);
xor (n562,n563,n574);
xor (n563,n564,n570);
nand (n564,n565,n566);
or (n565,n527,n89);
nand (n566,n567,n265);
nor (n567,n568,n569);
and (n568,n507,n72);
and (n569,n509,n102);
nor (n570,n71,n571);
nor (n571,n572,n573);
and (n572,n76,n484);
and (n573,n75,n482);
nand (n574,n575,n576);
or (n575,n289,n521);
or (n576,n577,n297);
nor (n577,n578,n579);
and (n578,n229,n221);
and (n579,n30,n220);
or (n580,n581,n582);
and (n581,n531,n545);
and (n582,n532,n539);
xor (n583,n584,n597);
xor (n584,n585,n591);
nand (n585,n586,n587);
or (n586,n44,n542);
or (n587,n45,n588);
nor (n588,n589,n590);
and (n589,n61,n370);
and (n590,n55,n369);
nand (n591,n592,n593);
or (n592,n208,n536);
or (n593,n594,n27);
nor (n594,n595,n596);
and (n595,n41,n273);
and (n596,n23,n272);
or (n597,n598,n599);
and (n598,n512,n524);
and (n599,n513,n515);
not (n600,n601);
nand (n601,n602,n603);
xor (n602,n467,n530);
or (n603,n604,n627);
and (n604,n605,n626);
xor (n605,n606,n607);
xor (n606,n546,n551);
or (n607,n608,n625);
and (n608,n609,n618);
xor (n609,n610,n611);
and (n610,n265,n476);
nand (n611,n612,n613);
or (n612,n297,n553);
nand (n613,n614,n228);
not (n614,n615);
nor (n615,n616,n617);
and (n616,n370,n229);
and (n617,n369,n30);
nand (n618,n619,n624);
or (n619,n620,n208);
not (n620,n621);
nor (n621,n622,n623);
and (n622,n507,n23);
and (n623,n41,n509);
nand (n624,n28,n488);
and (n625,n610,n611);
xor (n626,n470,n497);
and (n627,n606,n607);
and (n628,n465,n560);
nor (n629,n630,n671);
xor (n630,n631,n668);
xor (n631,n632,n651);
xor (n632,n633,n645);
xor (n633,n634,n641);
nand (n634,n635,n637);
or (n635,n636,n89);
not (n636,n567);
nand (n637,n265,n638);
nor (n638,n639,n640);
and (n639,n491,n72);
and (n640,n490,n102);
nor (n641,n71,n642);
nor (n642,n643,n644);
and (n643,n76,n503);
and (n644,n75,n501);
nand (n645,n646,n647);
or (n646,n44,n588);
or (n647,n45,n648);
nor (n648,n649,n650);
and (n649,n61,n331);
and (n650,n55,n330);
xor (n651,n652,n665);
xor (n652,n653,n659);
nand (n653,n654,n655);
or (n654,n289,n577);
or (n655,n656,n297);
nor (n656,n657,n658);
and (n657,n229,n148);
and (n658,n30,n147);
nand (n659,n660,n661);
or (n660,n208,n594);
or (n661,n662,n27);
nor (n662,n663,n664);
and (n663,n41,n261);
and (n664,n23,n263);
or (n665,n666,n667);
and (n666,n563,n574);
and (n667,n564,n570);
or (n668,n669,n670);
and (n669,n584,n597);
and (n670,n585,n591);
or (n671,n672,n673);
and (n672,n561,n583);
and (n673,n562,n580);
nand (n674,n630,n671);
nand (n675,n676,n718);
not (n676,n677);
xor (n677,n678,n717);
xor (n678,n679,n698);
xor (n679,n680,n692);
xor (n680,n681,n688);
nand (n681,n682,n684);
or (n682,n683,n89);
not (n683,n638);
nand (n684,n265,n685);
nor (n685,n686,n687);
and (n686,n370,n72);
and (n687,n369,n102);
nor (n688,n71,n689);
nor (n689,n690,n691);
and (n690,n76,n509);
and (n691,n75,n507);
nand (n692,n693,n694);
or (n693,n44,n648);
or (n694,n45,n695);
nor (n695,n696,n697);
and (n696,n61,n273);
and (n697,n55,n272);
xor (n698,n699,n714);
xor (n699,n700,n713);
xor (n700,n701,n707);
nand (n701,n702,n703);
or (n702,n289,n656);
or (n703,n704,n297);
nor (n704,n705,n706);
and (n705,n229,n82);
and (n706,n30,n81);
nand (n707,n708,n709);
or (n708,n208,n662);
or (n709,n27,n710);
nor (n710,n711,n712);
and (n711,n41,n221);
and (n712,n23,n220);
and (n713,n653,n659);
or (n714,n715,n716);
and (n715,n633,n645);
and (n716,n634,n641);
and (n717,n652,n665);
not (n718,n719);
or (n719,n720,n721);
and (n720,n631,n668);
and (n721,n632,n651);
nand (n722,n675,n723,n864);
nor (n723,n724,n861);
nor (n724,n725,n859);
and (n725,n726,n854);
or (n726,n727,n853);
and (n727,n728,n769);
xor (n728,n729,n762);
or (n729,n730,n761);
and (n730,n731,n749);
xor (n731,n732,n739);
nand (n732,n733,n738);
or (n733,n734,n208);
not (n734,n735);
nor (n735,n736,n737);
and (n736,n503,n41);
and (n737,n501,n23);
nand (n738,n28,n621);
nand (n739,n740,n745);
or (n740,n741,n45);
not (n741,n742);
nor (n742,n743,n744);
and (n743,n482,n55);
and (n744,n484,n61);
nand (n745,n118,n746);
nand (n746,n747,n748);
or (n747,n61,n476);
or (n748,n55,n478);
xor (n749,n750,n755);
and (n750,n751,n55);
nand (n751,n752,n754);
or (n752,n23,n753);
and (n753,n476,n49);
or (n754,n49,n476);
nand (n755,n756,n760);
or (n756,n289,n757);
nor (n757,n758,n759);
and (n758,n229,n491);
and (n759,n30,n490);
or (n760,n615,n297);
and (n761,n732,n739);
xor (n762,n763,n768);
xor (n763,n764,n767);
nand (n764,n765,n766);
or (n765,n741,n44);
or (n766,n45,n499);
and (n767,n750,n755);
xor (n768,n609,n618);
or (n769,n770,n852);
and (n770,n771,n792);
xor (n771,n772,n791);
or (n772,n773,n790);
and (n773,n774,n783);
xor (n774,n775,n776);
and (n775,n46,n476);
nand (n776,n777,n782);
or (n777,n778,n208);
not (n778,n779);
nor (n779,n780,n781);
and (n780,n482,n23);
and (n781,n484,n41);
nand (n782,n735,n28);
nand (n783,n784,n789);
or (n784,n289,n785);
not (n785,n786);
nor (n786,n787,n788);
and (n787,n509,n229);
and (n788,n507,n30);
or (n789,n757,n297);
and (n790,n775,n776);
xor (n791,n731,n749);
or (n792,n793,n851);
and (n793,n794,n850);
xor (n794,n795,n809);
nor (n795,n796,n804);
not (n796,n797);
nand (n797,n798,n803);
or (n798,n799,n289);
not (n799,n800);
nand (n800,n801,n802);
or (n801,n503,n30);
nand (n802,n30,n503);
nand (n803,n786,n225);
nand (n804,n805,n23);
nand (n805,n806,n808);
or (n806,n30,n807);
and (n807,n476,n19);
or (n808,n19,n476);
nand (n809,n810,n848);
or (n810,n811,n834);
not (n811,n812);
nand (n812,n813,n833);
or (n813,n814,n823);
nor (n814,n815,n822);
nand (n815,n816,n821);
or (n816,n817,n289);
not (n817,n818);
nand (n818,n819,n820);
or (n819,n484,n30);
nand (n820,n30,n484);
nand (n821,n800,n225);
nor (n822,n27,n478);
nand (n823,n824,n831);
nand (n824,n825,n830);
or (n825,n826,n289);
not (n826,n827);
nand (n827,n828,n829);
or (n828,n229,n476);
or (n829,n30,n478);
nand (n830,n818,n225);
nor (n831,n832,n229);
and (n832,n476,n225);
nand (n833,n815,n822);
not (n834,n835);
nand (n835,n836,n844);
not (n836,n837);
nand (n837,n838,n843);
or (n838,n839,n208);
not (n839,n840);
nand (n840,n841,n842);
or (n841,n41,n476);
or (n842,n23,n478);
nand (n843,n28,n779);
nor (n844,n845,n847);
and (n845,n796,n846);
not (n846,n804);
and (n847,n797,n804);
nand (n848,n849,n837);
not (n849,n844);
xor (n850,n774,n783);
and (n851,n795,n809);
and (n852,n772,n791);
and (n853,n729,n762);
or (n854,n855,n856);
xor (n855,n605,n626);
or (n856,n857,n858);
and (n857,n763,n768);
and (n858,n764,n767);
not (n859,n860);
nand (n860,n855,n856);
nand (n861,n862,n463);
not (n862,n863);
nor (n863,n602,n603);
not (n864,n629);
nand (n865,n677,n719);
nor (n866,n867,n924);
nand (n867,n868,n917);
not (n868,n869);
nor (n869,n870,n908);
xor (n870,n871,n899);
xor (n871,n872,n873);
xor (n872,n359,n372);
xor (n873,n874,n883);
xor (n874,n875,n876);
xor (n875,n345,n351);
and (n876,n877,n880);
nand (n877,n878,n879);
or (n878,n289,n704);
or (n879,n347,n297);
nand (n880,n881,n882);
or (n881,n208,n710);
or (n882,n353,n27);
or (n883,n884,n898);
and (n884,n885,n895);
xor (n885,n886,n891);
nand (n886,n887,n889);
or (n887,n888,n89);
not (n888,n685);
nand (n889,n890,n265);
not (n890,n362);
nor (n891,n71,n892);
nor (n892,n893,n894);
and (n893,n76,n490);
and (n894,n75,n491);
nand (n895,n896,n897);
or (n896,n44,n695);
or (n897,n45,n375);
and (n898,n886,n891);
or (n899,n900,n907);
and (n900,n901,n904);
xor (n901,n902,n903);
xor (n902,n877,n880);
and (n903,n701,n707);
or (n904,n905,n906);
and (n905,n680,n692);
and (n906,n681,n688);
and (n907,n902,n903);
or (n908,n909,n916);
and (n909,n910,n913);
xor (n910,n911,n912);
xor (n911,n885,n895);
xor (n912,n901,n904);
or (n913,n914,n915);
and (n914,n699,n714);
and (n915,n700,n713);
and (n916,n911,n912);
nand (n917,n918,n920);
not (n918,n919);
xor (n919,n910,n913);
not (n920,n921);
or (n921,n922,n923);
and (n922,n678,n717);
and (n923,n679,n698);
nand (n924,n925,n938);
nand (n925,n926,n934);
not (n926,n927);
xor (n927,n928,n931);
xor (n928,n929,n930);
xor (n929,n320,n333);
xor (n930,n342,n357);
or (n931,n932,n933);
and (n932,n874,n883);
and (n933,n875,n876);
not (n934,n935);
or (n935,n936,n937);
and (n936,n871,n899);
and (n937,n872,n873);
nand (n938,n939,n941);
not (n939,n940);
xor (n940,n253,n340);
not (n941,n942);
or (n942,n943,n944);
and (n943,n928,n931);
and (n944,n929,n930);
nand (n945,n946,n938);
nand (n946,n947,n954);
or (n947,n948,n949);
not (n948,n925);
not (n949,n950);
nand (n950,n951,n953);
or (n951,n869,n952);
nand (n952,n919,n921);
nand (n953,n870,n908);
nand (n954,n927,n935);
nand (n955,n942,n940);
not (n956,n957);
nand (n957,n958,n968);
or (n958,n959,n960);
not (n959,n435);
not (n960,n961);
nand (n961,n962,n967);
or (n962,n963,n449);
nor (n963,n964,n966);
and (n964,n965,n413);
and (n965,n251,n381);
nor (n966,n414,n431);
nand (n967,n450,n451);
or (n968,n436,n438);
nand (n969,n190,n243);
and (n970,n971,n972);
not (n971,n4);
not (n972,n187);
not (n973,n974);
and (n974,n975,n1030,n38);
nand (n975,n976,n1029);
or (n976,n977,n1011);
not (n977,n978);
nor (n978,n979,n1010);
and (n979,n980,n999);
not (n980,n981);
or (n981,n982,n998);
and (n982,n983,n995);
xor (n983,n984,n991);
nand (n984,n985,n990);
or (n985,n986,n90);
not (n986,n987);
nand (n987,n988,n989);
or (n988,n72,n36);
or (n989,n102,n37);
or (n990,n89,n176);
nand (n991,n992,n993,n514);
or (n992,n76,n62);
not (n993,n994);
and (n994,n62,n76);
or (n995,n996,n997);
and (n996,n170,n179);
and (n997,n171,n173);
and (n998,n984,n991);
not (n999,n1000);
xor (n1000,n1001,n1009);
xor (n1001,n1002,n1005);
nand (n1002,n1003,n987);
or (n1003,n1004,n265);
not (n1004,n89);
nor (n1005,n71,n1006);
nor (n1006,n1007,n1008);
and (n1007,n76,n69);
and (n1008,n75,n39);
not (n1009,n991);
and (n1010,n981,n1000);
nand (n1011,n1012,n1020,n1028);
nand (n1012,n455,n1013);
and (n1013,n248,n1014,n1015);
nor (n1014,n189,n5);
or (n1015,n1016,n1019);
or (n1016,n1017,n1018);
and (n1017,n167,n183);
and (n1018,n168,n169);
xor (n1019,n983,n995);
nand (n1020,n1021,n1015);
nand (n1021,n1022,n1024);
or (n1022,n1023,n956);
not (n1023,n1014);
nor (n1024,n1025,n186);
and (n1025,n1026,n1027);
not (n1026,n969);
not (n1027,n5);
nand (n1028,n1016,n1019);
nand (n1029,n977,n1011);
not (n1030,n22);
wire s0n1031,s1n1031,notn1031;
or (n1031,s0n1031,s1n1031);
not(notn1031,n22);
and (s0n1031,notn1031,n1032);
and (s1n1031,n22,n2332);
and (n1032,n38,n1033);
xor (n1033,n1034,n1848);
xor (n1034,n1035,n2330);
xor (n1035,n1036,n1843);
xor (n1036,n1037,n2323);
xor (n1037,n1038,n1837);
xor (n1038,n1039,n2311);
xor (n1039,n1040,n1831);
xor (n1040,n1041,n2294);
xor (n1041,n1042,n1825);
xor (n1042,n1043,n2272);
xor (n1043,n1044,n1819);
xor (n1044,n1045,n2245);
xor (n1045,n1046,n1813);
xor (n1046,n1047,n2213);
xor (n1047,n1048,n1807);
xor (n1048,n1049,n2176);
xor (n1049,n1050,n1801);
xor (n1050,n1051,n2134);
xor (n1051,n1052,n1795);
xor (n1052,n1053,n2087);
xor (n1053,n1054,n1789);
xor (n1054,n1055,n2035);
xor (n1055,n1056,n1783);
xor (n1056,n1057,n1978);
xor (n1057,n1058,n1777);
xor (n1058,n1059,n1916);
xor (n1059,n1060,n1771);
xor (n1060,n1061,n1849);
xor (n1061,n1062,n994);
xor (n1062,n1063,n1763);
xor (n1063,n1064,n1762);
xor (n1064,n1065,n1674);
xor (n1065,n1066,n1673);
xor (n1066,n1067,n1575);
xor (n1067,n1068,n1574);
xor (n1068,n1069,n1472);
xor (n1069,n1070,n1471);
xor (n1070,n1071,n1364);
xor (n1071,n1072,n1363);
xor (n1072,n1073,n1084);
xor (n1073,n1074,n1083);
xor (n1074,n1075,n1082);
xor (n1075,n1076,n1081);
xor (n1076,n1077,n1080);
xor (n1077,n1078,n1079);
and (n1078,n37,n225);
and (n1079,n37,n30);
and (n1080,n1078,n1079);
and (n1081,n37,n19);
and (n1082,n1076,n1081);
and (n1083,n37,n23);
or (n1084,n1085,n1086);
and (n1085,n1074,n1083);
and (n1086,n1073,n1087);
or (n1087,n1085,n1088);
and (n1088,n1073,n1089);
or (n1089,n1085,n1090);
and (n1090,n1073,n1091);
or (n1091,n1085,n1092);
and (n1092,n1073,n1093);
or (n1093,n1094,n1278);
and (n1094,n1095,n1277);
xor (n1095,n1075,n1096);
or (n1096,n1097,n1189);
and (n1097,n1098,n1188);
xor (n1098,n1077,n1099);
or (n1099,n1080,n1100);
and (n1100,n1101,n1103);
xor (n1101,n1078,n1102);
and (n1102,n39,n30);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n39,n225);
and (n1106,n62,n30);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n62,n225);
and (n1112,n103,n30);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n103,n225);
and (n1118,n114,n30);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n114,n225);
and (n1124,n82,n30);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
and (n1129,n82,n225);
and (n1130,n148,n30);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
and (n1135,n148,n225);
and (n1136,n221,n30);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
and (n1141,n221,n225);
and (n1142,n261,n30);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
and (n1147,n261,n225);
and (n1148,n273,n30);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1154);
and (n1152,n1153,n555);
and (n1153,n273,n225);
and (n1154,n1155,n1156);
xor (n1155,n1153,n555);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
and (n1158,n331,n225);
and (n1159,n370,n30);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
and (n1164,n370,n225);
and (n1165,n491,n30);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1171);
and (n1169,n1170,n788);
and (n1170,n491,n225);
and (n1171,n1172,n1173);
xor (n1172,n1170,n788);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
and (n1175,n507,n225);
and (n1176,n501,n30);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
and (n1181,n501,n225);
and (n1182,n482,n30);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
and (n1185,n1186,n1187);
and (n1186,n482,n225);
and (n1187,n476,n30);
and (n1188,n39,n19);
and (n1189,n1190,n1191);
xor (n1190,n1098,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1101,n1103);
and (n1194,n62,n19);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1108,n1109);
and (n1200,n103,n19);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1114,n1115);
and (n1206,n114,n19);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1120,n1121);
and (n1212,n82,n19);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1126,n1127);
and (n1218,n148,n19);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1132,n1133);
and (n1224,n221,n19);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1138,n1139);
and (n1230,n261,n19);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1144,n1145);
and (n1236,n273,n19);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1150,n1151);
and (n1242,n331,n19);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1155,n1156);
and (n1248,n370,n19);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1161,n1162);
and (n1254,n491,n19);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1167,n1168);
and (n1260,n507,n19);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1172,n1173);
and (n1266,n501,n19);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1178,n1179);
and (n1272,n482,n19);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
and (n1275,n1276,n807);
xor (n1276,n1184,n1185);
and (n1277,n39,n23);
and (n1278,n1279,n1280);
xor (n1279,n1095,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1190,n1191);
and (n1283,n62,n23);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1196,n1197);
and (n1289,n103,n23);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1202,n1203);
and (n1295,n114,n23);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1208,n1209);
and (n1301,n82,n23);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1214,n1215);
and (n1307,n148,n23);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1220,n1221);
and (n1313,n221,n23);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1226,n1227);
and (n1319,n261,n23);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1232,n1233);
and (n1325,n273,n23);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1238,n1239);
and (n1331,n331,n23);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1337);
and (n1335,n1336,n495);
xor (n1336,n1244,n1245);
and (n1337,n1338,n1339);
xor (n1338,n1336,n495);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1250,n1251);
and (n1342,n491,n23);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1348);
and (n1346,n1347,n622);
xor (n1347,n1256,n1257);
and (n1348,n1349,n1350);
xor (n1349,n1347,n622);
or (n1350,n1351,n1353);
and (n1351,n1352,n737);
xor (n1352,n1262,n1263);
and (n1353,n1354,n1355);
xor (n1354,n1352,n737);
or (n1355,n1356,n1358);
and (n1356,n1357,n780);
xor (n1357,n1268,n1269);
and (n1358,n1359,n1360);
xor (n1359,n1357,n780);
and (n1360,n1361,n1362);
xor (n1361,n1274,n1275);
and (n1362,n476,n23);
and (n1363,n37,n49);
or (n1364,n1365,n1367);
and (n1365,n1366,n1363);
xor (n1366,n1073,n1087);
and (n1367,n1368,n1369);
xor (n1368,n1366,n1363);
or (n1369,n1370,n1372);
and (n1370,n1371,n1363);
xor (n1371,n1073,n1089);
and (n1372,n1373,n1374);
xor (n1373,n1371,n1363);
or (n1374,n1375,n1377);
and (n1375,n1376,n1363);
xor (n1376,n1073,n1091);
and (n1377,n1378,n1379);
xor (n1378,n1376,n1363);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1073,n1093);
and (n1382,n39,n49);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
or (n1385,n1386,n1389);
and (n1386,n1387,n1388);
xor (n1387,n1279,n1280);
and (n1388,n62,n49);
and (n1389,n1390,n1391);
xor (n1390,n1387,n1388);
or (n1391,n1392,n1395);
and (n1392,n1393,n1394);
xor (n1393,n1285,n1286);
and (n1394,n103,n49);
and (n1395,n1396,n1397);
xor (n1396,n1393,n1394);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1291,n1292);
and (n1400,n114,n49);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
or (n1403,n1404,n1407);
and (n1404,n1405,n1406);
xor (n1405,n1297,n1298);
and (n1406,n82,n49);
and (n1407,n1408,n1409);
xor (n1408,n1405,n1406);
or (n1409,n1410,n1413);
and (n1410,n1411,n1412);
xor (n1411,n1303,n1304);
and (n1412,n148,n49);
and (n1413,n1414,n1415);
xor (n1414,n1411,n1412);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1309,n1310);
and (n1418,n221,n49);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1315,n1316);
and (n1424,n261,n49);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1321,n1322);
and (n1430,n273,n49);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
or (n1433,n1434,n1437);
and (n1434,n1435,n1436);
xor (n1435,n1327,n1328);
and (n1436,n331,n49);
and (n1437,n1438,n1439);
xor (n1438,n1435,n1436);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1333,n1334);
and (n1442,n370,n49);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1338,n1339);
and (n1448,n491,n49);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1344,n1345);
and (n1454,n507,n49);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
or (n1457,n1458,n1461);
and (n1458,n1459,n1460);
xor (n1459,n1349,n1350);
and (n1460,n501,n49);
and (n1461,n1462,n1463);
xor (n1462,n1459,n1460);
or (n1463,n1464,n1467);
and (n1464,n1465,n1466);
xor (n1465,n1354,n1355);
and (n1466,n482,n49);
and (n1467,n1468,n1469);
xor (n1468,n1465,n1466);
and (n1469,n1470,n753);
xor (n1470,n1359,n1360);
and (n1471,n37,n55);
or (n1472,n1473,n1475);
and (n1473,n1474,n1471);
xor (n1474,n1368,n1369);
and (n1475,n1476,n1477);
xor (n1476,n1474,n1471);
or (n1477,n1478,n1480);
and (n1478,n1479,n1471);
xor (n1479,n1373,n1374);
and (n1480,n1481,n1482);
xor (n1481,n1479,n1471);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1378,n1379);
and (n1485,n39,n55);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1384,n1385);
and (n1491,n62,n55);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1390,n1391);
and (n1497,n103,n55);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1396,n1397);
and (n1503,n114,n55);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1402,n1403);
and (n1509,n82,n55);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1408,n1409);
and (n1515,n148,n55);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1414,n1415);
and (n1521,n221,n55);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1420,n1421);
and (n1527,n261,n55);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1426,n1427);
and (n1533,n273,n55);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1432,n1433);
and (n1539,n331,n55);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1438,n1439);
and (n1545,n370,n55);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1444,n1445);
and (n1551,n491,n55);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
xor (n1556,n1450,n1451);
and (n1557,n507,n55);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1456,n1457);
and (n1563,n501,n55);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
or (n1566,n1567,n1569);
and (n1567,n1568,n743);
xor (n1568,n1462,n1463);
and (n1569,n1570,n1571);
xor (n1570,n1568,n743);
and (n1571,n1572,n1573);
xor (n1572,n1468,n1469);
and (n1573,n476,n55);
and (n1574,n37,n93);
or (n1575,n1576,n1578);
and (n1576,n1577,n1574);
xor (n1577,n1476,n1477);
and (n1578,n1579,n1580);
xor (n1579,n1577,n1574);
or (n1580,n1581,n1584);
and (n1581,n1582,n1583);
xor (n1582,n1481,n1482);
and (n1583,n39,n93);
and (n1584,n1585,n1586);
xor (n1585,n1582,n1583);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
xor (n1588,n1487,n1488);
and (n1589,n62,n93);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1493,n1494);
and (n1595,n103,n93);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1499,n1500);
and (n1601,n114,n93);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
xor (n1606,n1505,n1506);
and (n1607,n82,n93);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1511,n1512);
and (n1613,n148,n93);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
xor (n1618,n1517,n1518);
and (n1619,n221,n93);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
xor (n1624,n1523,n1524);
and (n1625,n261,n93);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1529,n1530);
and (n1631,n273,n93);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1535,n1536);
and (n1637,n331,n93);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1541,n1542);
and (n1643,n370,n93);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1547,n1548);
and (n1649,n491,n93);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1553,n1554);
and (n1655,n507,n93);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1559,n1560);
and (n1661,n501,n93);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1565,n1566);
and (n1667,n482,n93);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
and (n1670,n1671,n1672);
xor (n1671,n1570,n1571);
not (n1672,n549);
and (n1673,n37,n72);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1579,n1580);
and (n1677,n39,n72);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
or (n1680,n1681,n1684);
and (n1681,n1682,n1683);
xor (n1682,n1585,n1586);
and (n1683,n62,n72);
and (n1684,n1685,n1686);
xor (n1685,n1682,n1683);
or (n1686,n1687,n1690);
and (n1687,n1688,n1689);
xor (n1688,n1591,n1592);
and (n1689,n103,n72);
and (n1690,n1691,n1692);
xor (n1691,n1688,n1689);
or (n1692,n1693,n1696);
and (n1693,n1694,n1695);
xor (n1694,n1597,n1598);
and (n1695,n114,n72);
and (n1696,n1697,n1698);
xor (n1697,n1694,n1695);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
xor (n1700,n1603,n1604);
and (n1701,n82,n72);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1609,n1610);
and (n1707,n148,n72);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
or (n1710,n1711,n1713);
and (n1711,n1712,n267);
xor (n1712,n1615,n1616);
and (n1713,n1714,n1715);
xor (n1714,n1712,n267);
or (n1715,n1716,n1718);
and (n1716,n1717,n260);
xor (n1717,n1621,n1622);
and (n1718,n1719,n1720);
xor (n1719,n1717,n260);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
xor (n1722,n1627,n1628);
and (n1723,n273,n72);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
xor (n1728,n1633,n1634);
and (n1729,n331,n72);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1735);
and (n1733,n1734,n686);
xor (n1734,n1639,n1640);
and (n1735,n1736,n1737);
xor (n1736,n1734,n686);
or (n1737,n1738,n1740);
and (n1738,n1739,n639);
xor (n1739,n1645,n1646);
and (n1740,n1741,n1742);
xor (n1741,n1739,n639);
or (n1742,n1743,n1745);
and (n1743,n1744,n568);
xor (n1744,n1651,n1652);
and (n1745,n1746,n1747);
xor (n1746,n1744,n568);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1657,n1658);
and (n1750,n501,n72);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1663,n1664);
and (n1756,n482,n72);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
and (n1759,n1760,n1761);
xor (n1760,n1669,n1670);
and (n1761,n476,n72);
and (n1762,n39,n76);
or (n1763,n1764,n1766);
and (n1764,n1765,n994);
xor (n1765,n1679,n1680);
and (n1766,n1767,n1768);
xor (n1767,n1765,n994);
or (n1768,n1769,n1772);
and (n1769,n1770,n1771);
xor (n1770,n1685,n1686);
and (n1771,n103,n76);
and (n1772,n1773,n1774);
xor (n1773,n1770,n1771);
or (n1774,n1775,n1778);
and (n1775,n1776,n1777);
xor (n1776,n1691,n1692);
and (n1777,n114,n76);
and (n1778,n1779,n1780);
xor (n1779,n1776,n1777);
or (n1780,n1781,n1784);
and (n1781,n1782,n1783);
xor (n1782,n1697,n1698);
and (n1783,n82,n76);
and (n1784,n1785,n1786);
xor (n1785,n1782,n1783);
or (n1786,n1787,n1790);
and (n1787,n1788,n1789);
xor (n1788,n1703,n1704);
and (n1789,n148,n76);
and (n1790,n1791,n1792);
xor (n1791,n1788,n1789);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1709,n1710);
and (n1795,n221,n76);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1714,n1715);
and (n1801,n261,n76);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1719,n1720);
and (n1807,n273,n76);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1725,n1726);
and (n1813,n331,n76);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1731,n1732);
and (n1819,n370,n76);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
or (n1822,n1823,n1826);
and (n1823,n1824,n1825);
xor (n1824,n1736,n1737);
and (n1825,n491,n76);
and (n1826,n1827,n1828);
xor (n1827,n1824,n1825);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1741,n1742);
and (n1831,n507,n76);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1838);
and (n1835,n1836,n1837);
xor (n1836,n1746,n1747);
and (n1837,n501,n76);
and (n1838,n1839,n1840);
xor (n1839,n1836,n1837);
or (n1840,n1841,n1844);
and (n1841,n1842,n1843);
xor (n1842,n1752,n1753);
and (n1843,n482,n76);
and (n1844,n1845,n1846);
xor (n1845,n1842,n1843);
and (n1846,n1847,n1848);
xor (n1847,n1758,n1759);
and (n1848,n476,n76);
or (n1849,n1850,n1852);
and (n1850,n1851,n1771);
xor (n1851,n1767,n1768);
and (n1852,n1853,n1854);
xor (n1853,n1851,n1771);
or (n1854,n1855,n1857);
and (n1855,n1856,n1777);
xor (n1856,n1773,n1774);
and (n1857,n1858,n1859);
xor (n1858,n1856,n1777);
or (n1859,n1860,n1862);
and (n1860,n1861,n1783);
xor (n1861,n1779,n1780);
and (n1862,n1863,n1864);
xor (n1863,n1861,n1783);
or (n1864,n1865,n1867);
and (n1865,n1866,n1789);
xor (n1866,n1785,n1786);
and (n1867,n1868,n1869);
xor (n1868,n1866,n1789);
or (n1869,n1870,n1872);
and (n1870,n1871,n1795);
xor (n1871,n1791,n1792);
and (n1872,n1873,n1874);
xor (n1873,n1871,n1795);
or (n1874,n1875,n1877);
and (n1875,n1876,n1801);
xor (n1876,n1797,n1798);
and (n1877,n1878,n1879);
xor (n1878,n1876,n1801);
or (n1879,n1880,n1882);
and (n1880,n1881,n1807);
xor (n1881,n1803,n1804);
and (n1882,n1883,n1884);
xor (n1883,n1881,n1807);
or (n1884,n1885,n1887);
and (n1885,n1886,n1813);
xor (n1886,n1809,n1810);
and (n1887,n1888,n1889);
xor (n1888,n1886,n1813);
or (n1889,n1890,n1892);
and (n1890,n1891,n1819);
xor (n1891,n1815,n1816);
and (n1892,n1893,n1894);
xor (n1893,n1891,n1819);
or (n1894,n1895,n1897);
and (n1895,n1896,n1825);
xor (n1896,n1821,n1822);
and (n1897,n1898,n1899);
xor (n1898,n1896,n1825);
or (n1899,n1900,n1902);
and (n1900,n1901,n1831);
xor (n1901,n1827,n1828);
and (n1902,n1903,n1904);
xor (n1903,n1901,n1831);
or (n1904,n1905,n1907);
and (n1905,n1906,n1837);
xor (n1906,n1833,n1834);
and (n1907,n1908,n1909);
xor (n1908,n1906,n1837);
or (n1909,n1910,n1912);
and (n1910,n1911,n1843);
xor (n1911,n1839,n1840);
and (n1912,n1913,n1914);
xor (n1913,n1911,n1843);
and (n1914,n1915,n1848);
xor (n1915,n1845,n1846);
or (n1916,n1917,n1919);
and (n1917,n1918,n1777);
xor (n1918,n1853,n1854);
and (n1919,n1920,n1921);
xor (n1920,n1918,n1777);
or (n1921,n1922,n1924);
and (n1922,n1923,n1783);
xor (n1923,n1858,n1859);
and (n1924,n1925,n1926);
xor (n1925,n1923,n1783);
or (n1926,n1927,n1929);
and (n1927,n1928,n1789);
xor (n1928,n1863,n1864);
and (n1929,n1930,n1931);
xor (n1930,n1928,n1789);
or (n1931,n1932,n1934);
and (n1932,n1933,n1795);
xor (n1933,n1868,n1869);
and (n1934,n1935,n1936);
xor (n1935,n1933,n1795);
or (n1936,n1937,n1939);
and (n1937,n1938,n1801);
xor (n1938,n1873,n1874);
and (n1939,n1940,n1941);
xor (n1940,n1938,n1801);
or (n1941,n1942,n1944);
and (n1942,n1943,n1807);
xor (n1943,n1878,n1879);
and (n1944,n1945,n1946);
xor (n1945,n1943,n1807);
or (n1946,n1947,n1949);
and (n1947,n1948,n1813);
xor (n1948,n1883,n1884);
and (n1949,n1950,n1951);
xor (n1950,n1948,n1813);
or (n1951,n1952,n1954);
and (n1952,n1953,n1819);
xor (n1953,n1888,n1889);
and (n1954,n1955,n1956);
xor (n1955,n1953,n1819);
or (n1956,n1957,n1959);
and (n1957,n1958,n1825);
xor (n1958,n1893,n1894);
and (n1959,n1960,n1961);
xor (n1960,n1958,n1825);
or (n1961,n1962,n1964);
and (n1962,n1963,n1831);
xor (n1963,n1898,n1899);
and (n1964,n1965,n1966);
xor (n1965,n1963,n1831);
or (n1966,n1967,n1969);
and (n1967,n1968,n1837);
xor (n1968,n1903,n1904);
and (n1969,n1970,n1971);
xor (n1970,n1968,n1837);
or (n1971,n1972,n1974);
and (n1972,n1973,n1843);
xor (n1973,n1908,n1909);
and (n1974,n1975,n1976);
xor (n1975,n1973,n1843);
and (n1976,n1977,n1848);
xor (n1977,n1913,n1914);
or (n1978,n1979,n1981);
and (n1979,n1980,n1783);
xor (n1980,n1920,n1921);
and (n1981,n1982,n1983);
xor (n1982,n1980,n1783);
or (n1983,n1984,n1986);
and (n1984,n1985,n1789);
xor (n1985,n1925,n1926);
and (n1986,n1987,n1988);
xor (n1987,n1985,n1789);
or (n1988,n1989,n1991);
and (n1989,n1990,n1795);
xor (n1990,n1930,n1931);
and (n1991,n1992,n1993);
xor (n1992,n1990,n1795);
or (n1993,n1994,n1996);
and (n1994,n1995,n1801);
xor (n1995,n1935,n1936);
and (n1996,n1997,n1998);
xor (n1997,n1995,n1801);
or (n1998,n1999,n2001);
and (n1999,n2000,n1807);
xor (n2000,n1940,n1941);
and (n2001,n2002,n2003);
xor (n2002,n2000,n1807);
or (n2003,n2004,n2006);
and (n2004,n2005,n1813);
xor (n2005,n1945,n1946);
and (n2006,n2007,n2008);
xor (n2007,n2005,n1813);
or (n2008,n2009,n2011);
and (n2009,n2010,n1819);
xor (n2010,n1950,n1951);
and (n2011,n2012,n2013);
xor (n2012,n2010,n1819);
or (n2013,n2014,n2016);
and (n2014,n2015,n1825);
xor (n2015,n1955,n1956);
and (n2016,n2017,n2018);
xor (n2017,n2015,n1825);
or (n2018,n2019,n2021);
and (n2019,n2020,n1831);
xor (n2020,n1960,n1961);
and (n2021,n2022,n2023);
xor (n2022,n2020,n1831);
or (n2023,n2024,n2026);
and (n2024,n2025,n1837);
xor (n2025,n1965,n1966);
and (n2026,n2027,n2028);
xor (n2027,n2025,n1837);
or (n2028,n2029,n2031);
and (n2029,n2030,n1843);
xor (n2030,n1970,n1971);
and (n2031,n2032,n2033);
xor (n2032,n2030,n1843);
and (n2033,n2034,n1848);
xor (n2034,n1975,n1976);
or (n2035,n2036,n2038);
and (n2036,n2037,n1789);
xor (n2037,n1982,n1983);
and (n2038,n2039,n2040);
xor (n2039,n2037,n1789);
or (n2040,n2041,n2043);
and (n2041,n2042,n1795);
xor (n2042,n1987,n1988);
and (n2043,n2044,n2045);
xor (n2044,n2042,n1795);
or (n2045,n2046,n2048);
and (n2046,n2047,n1801);
xor (n2047,n1992,n1993);
and (n2048,n2049,n2050);
xor (n2049,n2047,n1801);
or (n2050,n2051,n2053);
and (n2051,n2052,n1807);
xor (n2052,n1997,n1998);
and (n2053,n2054,n2055);
xor (n2054,n2052,n1807);
or (n2055,n2056,n2058);
and (n2056,n2057,n1813);
xor (n2057,n2002,n2003);
and (n2058,n2059,n2060);
xor (n2059,n2057,n1813);
or (n2060,n2061,n2063);
and (n2061,n2062,n1819);
xor (n2062,n2007,n2008);
and (n2063,n2064,n2065);
xor (n2064,n2062,n1819);
or (n2065,n2066,n2068);
and (n2066,n2067,n1825);
xor (n2067,n2012,n2013);
and (n2068,n2069,n2070);
xor (n2069,n2067,n1825);
or (n2070,n2071,n2073);
and (n2071,n2072,n1831);
xor (n2072,n2017,n2018);
and (n2073,n2074,n2075);
xor (n2074,n2072,n1831);
or (n2075,n2076,n2078);
and (n2076,n2077,n1837);
xor (n2077,n2022,n2023);
and (n2078,n2079,n2080);
xor (n2079,n2077,n1837);
or (n2080,n2081,n2083);
and (n2081,n2082,n1843);
xor (n2082,n2027,n2028);
and (n2083,n2084,n2085);
xor (n2084,n2082,n1843);
and (n2085,n2086,n1848);
xor (n2086,n2032,n2033);
or (n2087,n2088,n2090);
and (n2088,n2089,n1795);
xor (n2089,n2039,n2040);
and (n2090,n2091,n2092);
xor (n2091,n2089,n1795);
or (n2092,n2093,n2095);
and (n2093,n2094,n1801);
xor (n2094,n2044,n2045);
and (n2095,n2096,n2097);
xor (n2096,n2094,n1801);
or (n2097,n2098,n2100);
and (n2098,n2099,n1807);
xor (n2099,n2049,n2050);
and (n2100,n2101,n2102);
xor (n2101,n2099,n1807);
or (n2102,n2103,n2105);
and (n2103,n2104,n1813);
xor (n2104,n2054,n2055);
and (n2105,n2106,n2107);
xor (n2106,n2104,n1813);
or (n2107,n2108,n2110);
and (n2108,n2109,n1819);
xor (n2109,n2059,n2060);
and (n2110,n2111,n2112);
xor (n2111,n2109,n1819);
or (n2112,n2113,n2115);
and (n2113,n2114,n1825);
xor (n2114,n2064,n2065);
and (n2115,n2116,n2117);
xor (n2116,n2114,n1825);
or (n2117,n2118,n2120);
and (n2118,n2119,n1831);
xor (n2119,n2069,n2070);
and (n2120,n2121,n2122);
xor (n2121,n2119,n1831);
or (n2122,n2123,n2125);
and (n2123,n2124,n1837);
xor (n2124,n2074,n2075);
and (n2125,n2126,n2127);
xor (n2126,n2124,n1837);
or (n2127,n2128,n2130);
and (n2128,n2129,n1843);
xor (n2129,n2079,n2080);
and (n2130,n2131,n2132);
xor (n2131,n2129,n1843);
and (n2132,n2133,n1848);
xor (n2133,n2084,n2085);
or (n2134,n2135,n2137);
and (n2135,n2136,n1801);
xor (n2136,n2091,n2092);
and (n2137,n2138,n2139);
xor (n2138,n2136,n1801);
or (n2139,n2140,n2142);
and (n2140,n2141,n1807);
xor (n2141,n2096,n2097);
and (n2142,n2143,n2144);
xor (n2143,n2141,n1807);
or (n2144,n2145,n2147);
and (n2145,n2146,n1813);
xor (n2146,n2101,n2102);
and (n2147,n2148,n2149);
xor (n2148,n2146,n1813);
or (n2149,n2150,n2152);
and (n2150,n2151,n1819);
xor (n2151,n2106,n2107);
and (n2152,n2153,n2154);
xor (n2153,n2151,n1819);
or (n2154,n2155,n2157);
and (n2155,n2156,n1825);
xor (n2156,n2111,n2112);
and (n2157,n2158,n2159);
xor (n2158,n2156,n1825);
or (n2159,n2160,n2162);
and (n2160,n2161,n1831);
xor (n2161,n2116,n2117);
and (n2162,n2163,n2164);
xor (n2163,n2161,n1831);
or (n2164,n2165,n2167);
and (n2165,n2166,n1837);
xor (n2166,n2121,n2122);
and (n2167,n2168,n2169);
xor (n2168,n2166,n1837);
or (n2169,n2170,n2172);
and (n2170,n2171,n1843);
xor (n2171,n2126,n2127);
and (n2172,n2173,n2174);
xor (n2173,n2171,n1843);
and (n2174,n2175,n1848);
xor (n2175,n2131,n2132);
or (n2176,n2177,n2179);
and (n2177,n2178,n1807);
xor (n2178,n2138,n2139);
and (n2179,n2180,n2181);
xor (n2180,n2178,n1807);
or (n2181,n2182,n2184);
and (n2182,n2183,n1813);
xor (n2183,n2143,n2144);
and (n2184,n2185,n2186);
xor (n2185,n2183,n1813);
or (n2186,n2187,n2189);
and (n2187,n2188,n1819);
xor (n2188,n2148,n2149);
and (n2189,n2190,n2191);
xor (n2190,n2188,n1819);
or (n2191,n2192,n2194);
and (n2192,n2193,n1825);
xor (n2193,n2153,n2154);
and (n2194,n2195,n2196);
xor (n2195,n2193,n1825);
or (n2196,n2197,n2199);
and (n2197,n2198,n1831);
xor (n2198,n2158,n2159);
and (n2199,n2200,n2201);
xor (n2200,n2198,n1831);
or (n2201,n2202,n2204);
and (n2202,n2203,n1837);
xor (n2203,n2163,n2164);
and (n2204,n2205,n2206);
xor (n2205,n2203,n1837);
or (n2206,n2207,n2209);
and (n2207,n2208,n1843);
xor (n2208,n2168,n2169);
and (n2209,n2210,n2211);
xor (n2210,n2208,n1843);
and (n2211,n2212,n1848);
xor (n2212,n2173,n2174);
or (n2213,n2214,n2216);
and (n2214,n2215,n1813);
xor (n2215,n2180,n2181);
and (n2216,n2217,n2218);
xor (n2217,n2215,n1813);
or (n2218,n2219,n2221);
and (n2219,n2220,n1819);
xor (n2220,n2185,n2186);
and (n2221,n2222,n2223);
xor (n2222,n2220,n1819);
or (n2223,n2224,n2226);
and (n2224,n2225,n1825);
xor (n2225,n2190,n2191);
and (n2226,n2227,n2228);
xor (n2227,n2225,n1825);
or (n2228,n2229,n2231);
and (n2229,n2230,n1831);
xor (n2230,n2195,n2196);
and (n2231,n2232,n2233);
xor (n2232,n2230,n1831);
or (n2233,n2234,n2236);
and (n2234,n2235,n1837);
xor (n2235,n2200,n2201);
and (n2236,n2237,n2238);
xor (n2237,n2235,n1837);
or (n2238,n2239,n2241);
and (n2239,n2240,n1843);
xor (n2240,n2205,n2206);
and (n2241,n2242,n2243);
xor (n2242,n2240,n1843);
and (n2243,n2244,n1848);
xor (n2244,n2210,n2211);
or (n2245,n2246,n2248);
and (n2246,n2247,n1819);
xor (n2247,n2217,n2218);
and (n2248,n2249,n2250);
xor (n2249,n2247,n1819);
or (n2250,n2251,n2253);
and (n2251,n2252,n1825);
xor (n2252,n2222,n2223);
and (n2253,n2254,n2255);
xor (n2254,n2252,n1825);
or (n2255,n2256,n2258);
and (n2256,n2257,n1831);
xor (n2257,n2227,n2228);
and (n2258,n2259,n2260);
xor (n2259,n2257,n1831);
or (n2260,n2261,n2263);
and (n2261,n2262,n1837);
xor (n2262,n2232,n2233);
and (n2263,n2264,n2265);
xor (n2264,n2262,n1837);
or (n2265,n2266,n2268);
and (n2266,n2267,n1843);
xor (n2267,n2237,n2238);
and (n2268,n2269,n2270);
xor (n2269,n2267,n1843);
and (n2270,n2271,n1848);
xor (n2271,n2242,n2243);
or (n2272,n2273,n2275);
and (n2273,n2274,n1825);
xor (n2274,n2249,n2250);
and (n2275,n2276,n2277);
xor (n2276,n2274,n1825);
or (n2277,n2278,n2280);
and (n2278,n2279,n1831);
xor (n2279,n2254,n2255);
and (n2280,n2281,n2282);
xor (n2281,n2279,n1831);
or (n2282,n2283,n2285);
and (n2283,n2284,n1837);
xor (n2284,n2259,n2260);
and (n2285,n2286,n2287);
xor (n2286,n2284,n1837);
or (n2287,n2288,n2290);
and (n2288,n2289,n1843);
xor (n2289,n2264,n2265);
and (n2290,n2291,n2292);
xor (n2291,n2289,n1843);
and (n2292,n2293,n1848);
xor (n2293,n2269,n2270);
or (n2294,n2295,n2297);
and (n2295,n2296,n1831);
xor (n2296,n2276,n2277);
and (n2297,n2298,n2299);
xor (n2298,n2296,n1831);
or (n2299,n2300,n2302);
and (n2300,n2301,n1837);
xor (n2301,n2281,n2282);
and (n2302,n2303,n2304);
xor (n2303,n2301,n1837);
or (n2304,n2305,n2307);
and (n2305,n2306,n1843);
xor (n2306,n2286,n2287);
and (n2307,n2308,n2309);
xor (n2308,n2306,n1843);
and (n2309,n2310,n1848);
xor (n2310,n2291,n2292);
or (n2311,n2312,n2314);
and (n2312,n2313,n1837);
xor (n2313,n2298,n2299);
and (n2314,n2315,n2316);
xor (n2315,n2313,n1837);
or (n2316,n2317,n2319);
and (n2317,n2318,n1843);
xor (n2318,n2303,n2304);
and (n2319,n2320,n2321);
xor (n2320,n2318,n1843);
and (n2321,n2322,n1848);
xor (n2322,n2308,n2309);
or (n2323,n2324,n2326);
and (n2324,n2325,n1843);
xor (n2325,n2315,n2316);
and (n2326,n2327,n2328);
xor (n2327,n2325,n1843);
and (n2328,n2329,n1848);
xor (n2329,n2320,n2321);
and (n2330,n2331,n1848);
xor (n2331,n2327,n2328);
xor (n2332,n2329,n1848);
endmodule
