module top (out,n17,n22,n24,n25,n27,n31,n34,n40,n58
        ,n72,n73,n74,n75,n76,n77,n78,n79,n83,n84
        ,n85,n89,n91,n93,n130,n132,n133,n134,n145,n146
        ,n147,n148,n160,n161,n162,n163,n176,n177,n178,n179
        ,n185,n187,n188,n191,n193,n196,n198,n199,n200,n280
        ,n386,n389,n391,n545,n547,n548,n551,n554,n555,n556
        ,n557,n560,n562,n566,n577,n578,n595,n598,n600,n601
        ,n603,n607,n613,n616,n618,n620,n624,n627,n629,n631
        ,n635,n638,n640,n642,n644,n652,n655,n657,n659,n663
        ,n666,n668,n670,n674,n677,n679,n681,n685,n688,n690
        ,n692,n700,n703,n705,n707,n711,n714,n716,n718,n722
        ,n725,n727,n729,n733,n736,n738,n740,n749,n752,n754
        ,n756,n770,n773,n775,n777,n796,n799,n801,n803,n812
        ,n815,n817,n819,n833,n836,n838,n840,n863,n866,n868
        ,n870,n886,n889,n891,n893,n938,n941,n943,n945,n949
        ,n952,n954,n956,n960,n963,n965,n967,n971,n974,n976
        ,n978,n986,n989,n991,n993,n997,n1000,n1002,n1004,n1008
        ,n1011,n1013,n1015,n1019,n1022,n1024,n1026,n1035,n1038,n1040
        ,n1042,n1047,n1050,n1052,n1054,n1064,n1067,n1069,n1071,n1089
        ,n1092,n1094,n1096,n1116,n1119,n1121,n1123,n1142,n1145,n1147
        ,n1149,n1171,n1174,n1176,n1178,n1190,n1193,n1195,n1197,n1229
        ,n1232,n1234,n1236,n1240,n1243,n1245,n1247,n1251,n1254,n1256
        ,n1258,n1262,n1265,n1267,n1269,n1290,n1293,n1295,n1297,n1304
        ,n1307,n1309,n1311,n1316,n1319,n1321,n1323,n1335,n1338,n1340
        ,n1342,n1351,n1354,n1356,n1358,n1368,n1371,n1373,n1375,n1383
        ,n1386,n1388,n1390,n1434,n1437,n1439,n1441,n1447,n1450,n1452
        ,n1454,n1464,n1467,n1469,n1471,n1500,n1503,n1505,n1507,n1619
        ,n1622,n1624,n1626,n1634,n1637,n1639,n1641,n1650,n1653,n1655
        ,n1657,n1666,n1669,n1671,n1673,n1681,n1684,n1686,n1688);
output out;
input n17;
input n22;
input n24;
input n25;
input n27;
input n31;
input n34;
input n40;
input n58;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n83;
input n84;
input n85;
input n89;
input n91;
input n93;
input n130;
input n132;
input n133;
input n134;
input n145;
input n146;
input n147;
input n148;
input n160;
input n161;
input n162;
input n163;
input n176;
input n177;
input n178;
input n179;
input n185;
input n187;
input n188;
input n191;
input n193;
input n196;
input n198;
input n199;
input n200;
input n280;
input n386;
input n389;
input n391;
input n545;
input n547;
input n548;
input n551;
input n554;
input n555;
input n556;
input n557;
input n560;
input n562;
input n566;
input n577;
input n578;
input n595;
input n598;
input n600;
input n601;
input n603;
input n607;
input n613;
input n616;
input n618;
input n620;
input n624;
input n627;
input n629;
input n631;
input n635;
input n638;
input n640;
input n642;
input n644;
input n652;
input n655;
input n657;
input n659;
input n663;
input n666;
input n668;
input n670;
input n674;
input n677;
input n679;
input n681;
input n685;
input n688;
input n690;
input n692;
input n700;
input n703;
input n705;
input n707;
input n711;
input n714;
input n716;
input n718;
input n722;
input n725;
input n727;
input n729;
input n733;
input n736;
input n738;
input n740;
input n749;
input n752;
input n754;
input n756;
input n770;
input n773;
input n775;
input n777;
input n796;
input n799;
input n801;
input n803;
input n812;
input n815;
input n817;
input n819;
input n833;
input n836;
input n838;
input n840;
input n863;
input n866;
input n868;
input n870;
input n886;
input n889;
input n891;
input n893;
input n938;
input n941;
input n943;
input n945;
input n949;
input n952;
input n954;
input n956;
input n960;
input n963;
input n965;
input n967;
input n971;
input n974;
input n976;
input n978;
input n986;
input n989;
input n991;
input n993;
input n997;
input n1000;
input n1002;
input n1004;
input n1008;
input n1011;
input n1013;
input n1015;
input n1019;
input n1022;
input n1024;
input n1026;
input n1035;
input n1038;
input n1040;
input n1042;
input n1047;
input n1050;
input n1052;
input n1054;
input n1064;
input n1067;
input n1069;
input n1071;
input n1089;
input n1092;
input n1094;
input n1096;
input n1116;
input n1119;
input n1121;
input n1123;
input n1142;
input n1145;
input n1147;
input n1149;
input n1171;
input n1174;
input n1176;
input n1178;
input n1190;
input n1193;
input n1195;
input n1197;
input n1229;
input n1232;
input n1234;
input n1236;
input n1240;
input n1243;
input n1245;
input n1247;
input n1251;
input n1254;
input n1256;
input n1258;
input n1262;
input n1265;
input n1267;
input n1269;
input n1290;
input n1293;
input n1295;
input n1297;
input n1304;
input n1307;
input n1309;
input n1311;
input n1316;
input n1319;
input n1321;
input n1323;
input n1335;
input n1338;
input n1340;
input n1342;
input n1351;
input n1354;
input n1356;
input n1358;
input n1368;
input n1371;
input n1373;
input n1375;
input n1383;
input n1386;
input n1388;
input n1390;
input n1434;
input n1437;
input n1439;
input n1441;
input n1447;
input n1450;
input n1452;
input n1454;
input n1464;
input n1467;
input n1469;
input n1471;
input n1500;
input n1503;
input n1505;
input n1507;
input n1619;
input n1622;
input n1624;
input n1626;
input n1634;
input n1637;
input n1639;
input n1641;
input n1650;
input n1653;
input n1655;
input n1657;
input n1666;
input n1669;
input n1671;
input n1673;
input n1681;
input n1684;
input n1686;
input n1688;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n26;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n80;
wire n81;
wire n82;
wire n86;
wire n87;
wire n88;
wire n90;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n189;
wire n190;
wire n192;
wire n194;
wire n195;
wire n197;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n387;
wire n388;
wire n390;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n546;
wire n549;
wire n550;
wire n552;
wire n553;
wire n558;
wire n559;
wire n561;
wire n563;
wire n564;
wire n565;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n596;
wire n597;
wire n599;
wire n602;
wire n604;
wire n605;
wire n606;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n614;
wire n615;
wire n617;
wire n619;
wire n621;
wire n622;
wire n623;
wire n625;
wire n626;
wire n628;
wire n630;
wire n632;
wire n633;
wire n634;
wire n636;
wire n637;
wire n639;
wire n641;
wire n643;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n653;
wire n654;
wire n656;
wire n658;
wire n660;
wire n661;
wire n662;
wire n664;
wire n665;
wire n667;
wire n669;
wire n671;
wire n672;
wire n673;
wire n675;
wire n676;
wire n678;
wire n680;
wire n682;
wire n683;
wire n684;
wire n686;
wire n687;
wire n689;
wire n691;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n701;
wire n702;
wire n704;
wire n706;
wire n708;
wire n709;
wire n710;
wire n712;
wire n713;
wire n715;
wire n717;
wire n719;
wire n720;
wire n721;
wire n723;
wire n724;
wire n726;
wire n728;
wire n730;
wire n731;
wire n732;
wire n734;
wire n735;
wire n737;
wire n739;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n750;
wire n751;
wire n753;
wire n755;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n771;
wire n772;
wire n774;
wire n776;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n797;
wire n798;
wire n800;
wire n802;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n813;
wire n814;
wire n816;
wire n818;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n834;
wire n835;
wire n837;
wire n839;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n864;
wire n865;
wire n867;
wire n869;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n887;
wire n888;
wire n890;
wire n892;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n939;
wire n940;
wire n942;
wire n944;
wire n946;
wire n947;
wire n948;
wire n950;
wire n951;
wire n953;
wire n955;
wire n957;
wire n958;
wire n959;
wire n961;
wire n962;
wire n964;
wire n966;
wire n968;
wire n969;
wire n970;
wire n972;
wire n973;
wire n975;
wire n977;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n987;
wire n988;
wire n990;
wire n992;
wire n994;
wire n995;
wire n996;
wire n998;
wire n999;
wire n1001;
wire n1003;
wire n1005;
wire n1006;
wire n1007;
wire n1009;
wire n1010;
wire n1012;
wire n1014;
wire n1016;
wire n1017;
wire n1018;
wire n1020;
wire n1021;
wire n1023;
wire n1025;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1036;
wire n1037;
wire n1039;
wire n1041;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1048;
wire n1049;
wire n1051;
wire n1053;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1065;
wire n1066;
wire n1068;
wire n1070;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1090;
wire n1091;
wire n1093;
wire n1095;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1117;
wire n1118;
wire n1120;
wire n1122;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1143;
wire n1144;
wire n1146;
wire n1148;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1172;
wire n1173;
wire n1175;
wire n1177;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1191;
wire n1192;
wire n1194;
wire n1196;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1230;
wire n1231;
wire n1233;
wire n1235;
wire n1237;
wire n1238;
wire n1239;
wire n1241;
wire n1242;
wire n1244;
wire n1246;
wire n1248;
wire n1249;
wire n1250;
wire n1252;
wire n1253;
wire n1255;
wire n1257;
wire n1259;
wire n1260;
wire n1261;
wire n1263;
wire n1264;
wire n1266;
wire n1268;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1291;
wire n1292;
wire n1294;
wire n1296;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1305;
wire n1306;
wire n1308;
wire n1310;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1317;
wire n1318;
wire n1320;
wire n1322;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1336;
wire n1337;
wire n1339;
wire n1341;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1352;
wire n1353;
wire n1355;
wire n1357;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1369;
wire n1370;
wire n1372;
wire n1374;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1384;
wire n1385;
wire n1387;
wire n1389;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1435;
wire n1436;
wire n1438;
wire n1440;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1448;
wire n1449;
wire n1451;
wire n1453;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1465;
wire n1466;
wire n1468;
wire n1470;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1501;
wire n1502;
wire n1504;
wire n1506;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1620;
wire n1621;
wire n1623;
wire n1625;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1635;
wire n1636;
wire n1638;
wire n1640;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1651;
wire n1652;
wire n1654;
wire n1656;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1667;
wire n1668;
wire n1670;
wire n1672;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1682;
wire n1683;
wire n1685;
wire n1687;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
xnor (out,n0,n2237);
or (n0,n1,n2215);
or (n1,n2,n2214);
and (n2,n3,n2152);
xor (n3,n4,n2121);
or (n4,n5,n2120);
and (n5,n6,n1945);
xor (n6,n7,n1901);
xor (n7,n8,n1778);
xor (n8,n9,n1276);
xor (n9,n10,n1271);
xor (n10,n11,n1028);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n931);
and (s0n11,notn11,1'b0);
and (s1n11,n931,n13);
xor (n13,n14,n742);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n588);
and (s0n14,notn14,1'b0);
and (s1n14,n588,n15);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n571);
and (s0n15,notn15,n16);
and (s1n15,n571,n558);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n18);
and (s0n16,notn16,1'b0);
and (s1n16,n18,n17);
and (n18,n19,n552);
and (n19,n20,n36);
or (n20,n21,n26,n30,n33);
and (n21,n22,n23);
and (n23,n24,n25);
and (n26,n27,n28);
and (n28,n29,n25);
not (n29,n24);
and (n30,n31,n32);
nor (n32,n29,n25);
and (n33,n34,n35);
nor (n35,n24,n25);
and (n36,n37,n551);
not (n37,n38);
wire s0n38,s1n38,notn38;
or (n38,s0n38,s1n38);
not(notn38,n550);
and (s0n38,notn38,n39);
and (s1n38,n550,1'b0);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n180);
and (s0n39,notn39,n40);
and (s1n39,n180,n41);
wire s0n41,s1n41,notn41;
or (n41,s0n41,s1n41);
not(notn41,n543);
and (s0n41,notn41,n42);
and (s1n41,n543,n517);
or (n42,n43,n485,n516,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n43,n44,n484);
or (n44,n45,n483);
or (n45,n46,n482);
or (n46,n47,n480);
or (n47,n48,n479);
or (n48,n49,n477);
or (n49,n50,n475);
nor (n50,n51,n400,n409,n421,n433,n444,n455,n466);
or (n51,1'b0,n52,n394,n398);
and (n52,n53,n393);
wire s0n53,s1n53,notn53;
or (n53,s0n53,s1n53);
not(notn53,n384);
and (s0n53,notn53,n54);
and (s1n53,n384,n292);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n251);
and (s0n54,notn54,1'b0);
and (s1n54,n251,n55);
or (n55,n56,n232,n236,n240,n243,n246,n248,1'b0);
and (n56,n57,n59);
not (n57,n58);
and (n59,n60,n205,n216,n226);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n94);
and (s0n60,notn60,n61);
and (s1n60,n94,1'b0);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n92);
and (s0n61,notn61,n62);
and (s1n61,n92,n90);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n86);
and (s0n62,notn62,n63);
and (s1n62,n86,n80);
wire s0n63,s1n63,notn63;
or (n63,s0n63,s1n63);
not(notn63,n79);
and (s0n63,notn63,n64);
and (s1n63,n79,1'b0);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n78);
and (s0n64,notn64,n65);
and (s1n64,n78,1'b1);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n77);
and (s0n65,notn65,n66);
and (s1n65,n77,1'b0);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n76);
and (s0n66,notn66,n67);
and (s1n66,n76,1'b1);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n75);
and (s0n67,notn67,n68);
and (s1n67,n75,1'b0);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n74);
and (s0n68,notn68,n69);
and (s1n68,n74,1'b1);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n73);
and (s0n69,notn69,n70);
and (s1n69,n73,1'b0);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n72);
and (s0n70,notn70,n57);
and (s1n70,n72,1'b1);
wire s0n80,s1n80,notn80;
or (n80,s0n80,s1n80);
not(notn80,n85);
and (s0n80,notn80,n81);
and (s1n80,n85,1'b0);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n84);
and (s0n81,notn81,n82);
and (s1n81,n84,1'b1);
not (n82,n83);
or (n86,n87,n89);
or (n87,n88,n83);
or (n88,n85,n84);
not (n90,n91);
or (n92,n91,n93);
not (n94,n95);
or (n95,n96,n203);
or (n96,n97,n201);
or (n97,n98,n195);
or (n98,n99,n194);
or (n99,n100,n190);
or (n100,n101,n189);
or (n101,n102,n184);
or (n102,n103,n183);
or (n103,n104,n182);
or (n104,n105,n180);
or (n105,n106,n174);
or (n106,n107,n173);
or (n107,n108,n172);
or (n108,n109,n171);
or (n109,n110,n170);
or (n110,n111,n169);
or (n111,n112,n168);
or (n112,n113,n167);
or (n113,n114,n164);
or (n114,n115,n158);
or (n115,n116,n157);
or (n116,n117,n156);
or (n117,n118,n155);
or (n118,n119,n154);
or (n119,n120,n153);
or (n120,n121,n151);
or (n121,n122,n149);
or (n122,n123,n143);
or (n123,n124,n142);
or (n124,n125,n141);
or (n125,n126,n140);
or (n126,n127,n139);
or (n127,n128,n137);
or (n128,n129,n135);
nor (n129,n130,n131,n133,n134);
not (n131,n132);
nor (n135,n130,n131,n136,n134);
not (n136,n133);
and (n137,n130,n132,n133,n138);
not (n138,n134);
and (n139,n130,n131,n133,n138);
nor (n140,n130,n132,n136,n134);
and (n141,n130,n131,n133,n134);
and (n142,n130,n132,n133,n134);
nor (n143,n144,n146,n147,n148);
not (n144,n145);
nor (n149,n144,n150,n147,n148);
not (n150,n146);
and (n151,n144,n146,n147,n152);
not (n152,n148);
and (n153,n145,n146,n147,n152);
and (n154,n145,n150,n147,n152);
and (n155,n144,n150,n147,n148);
and (n156,n145,n150,n147,n148);
and (n157,n145,n146,n147,n148);
nor (n158,n159,n161,n162,n163);
not (n159,n160);
and (n164,n160,n161,n165,n166);
not (n165,n162);
not (n166,n163);
and (n167,n159,n161,n165,n166);
and (n168,n160,n161,n162,n166);
nor (n169,n160,n161,n165,n166);
and (n170,n159,n161,n162,n163);
and (n171,n159,n161,n165,n163);
and (n172,n160,n161,n165,n163);
nor (n173,n159,n161,n162,n166);
nor (n174,n175,n177,n178,n179);
not (n175,n176);
nor (n180,n176,n181,n178,n179);
not (n181,n177);
and (n182,n175,n181,n178,n179);
and (n183,n176,n181,n178,n179);
nor (n184,n185,n186,n188);
not (n186,n187);
and (n189,n185,n187,n188);
and (n190,n191,n192);
not (n192,n193);
nor (n194,n191,n192);
nor (n195,n196,n197,n199,n200);
not (n197,n198);
and (n201,n196,n198,n199,n202);
not (n202,n200);
and (n203,n204,n197,n199,n202);
not (n204,n196);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n94);
and (s0n205,notn205,n206);
and (s1n205,n94,1'b0);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n92);
and (s0n206,notn206,n207);
and (s1n206,n92,1'b0);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n86);
and (s0n207,notn207,n208);
and (s1n207,n86,n88);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n79);
and (s0n208,notn208,n209);
and (s1n208,n79,1'b1);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n78);
and (s0n209,notn209,n210);
and (s1n209,n78,1'b1);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n77);
and (s0n210,notn210,n211);
and (s1n210,n77,1'b0);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n76);
and (s0n211,notn211,n212);
and (s1n211,n76,1'b0);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n75);
and (s0n212,notn212,n213);
and (s1n212,n75,1'b1);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n74);
and (s0n213,notn213,n214);
and (s1n213,n74,1'b1);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n73);
and (s0n214,notn214,n215);
and (s1n214,n73,1'b0);
not (n215,n72);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n94);
and (s0n216,notn216,n217);
and (s1n216,n94,1'b0);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n92);
and (s0n217,notn217,n218);
and (s1n217,n92,1'b0);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n86);
and (s0n218,notn218,n219);
and (s1n218,n86,n225);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n79);
and (s0n219,notn219,n220);
and (s1n219,n79,1'b1);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n78);
and (s0n220,notn220,n221);
and (s1n220,n78,1'b1);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n77);
and (s0n221,notn221,n222);
and (s1n221,n77,1'b0);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n76);
and (s0n222,notn222,n223);
and (s1n222,n76,1'b0);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n75);
and (s0n223,notn223,n224);
and (s1n223,n75,1'b0);
not (n224,n74);
not (n225,n88);
not (n226,n227);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n94);
and (s0n227,notn227,n228);
and (s1n227,n94,1'b0);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n92);
and (s0n228,notn228,n229);
and (s1n228,n92,1'b0);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n86);
and (s0n229,notn229,n230);
and (s1n229,n86,1'b0);
wire s0n230,s1n230,notn230;
or (n230,s0n230,s1n230);
not(notn230,n79);
and (s0n230,notn230,n231);
and (s1n230,n79,1'b0);
not (n231,n78);
and (n232,n233,n234);
not (n233,n73);
and (n234,n235,n205,n216,n226);
not (n235,n60);
and (n236,n237,n238);
not (n237,n75);
and (n238,n60,n239,n216,n226);
not (n239,n205);
and (n240,n241,n242);
not (n241,n77);
and (n242,n235,n239,n216,n226);
and (n243,n244,n245);
not (n244,n79);
nor (n245,n235,n239,n216,n227);
and (n246,n82,n247);
nor (n247,n60,n239,n216,n227);
and (n248,n249,n250);
not (n249,n85);
nor (n250,n235,n205,n216,n227);
or (n251,n252,n281);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n279);
and (s0n252,notn252,n253);
and (s1n252,n279,1'b0);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n278);
and (s0n253,notn253,n254);
and (s1n253,n278,n273);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n272);
and (s0n254,notn254,n255);
and (s1n254,n272,n261);
wire s0n255,s1n255,notn255;
or (n255,s0n255,s1n255);
not(notn255,n260);
and (s0n255,notn255,n256);
and (s1n255,n260,n123);
or (n256,n257,n154);
or (n257,n258,n153);
or (n258,n259,n151);
or (n259,n143,n149);
or (n260,n130,n132,n133,n134);
or (n261,1'b0,1'b0,n262,n268,n270);
and (n262,n263,n266);
or (n263,1'b0,1'b0,n264,n184);
and (n264,n265,n187,n188);
not (n265,n185);
and (n266,n175,n181,n178,n267);
not (n267,n179);
and (n268,n191,n269);
and (n269,n176,n181,n178,n267);
or (n270,n271,n182);
or (n271,n174,n180);
or (n272,n176,n177,n178,n179);
or (n273,n274,n173);
or (n274,n275,n171);
or (n275,n276,n168);
or (n276,n277,n167);
or (n277,n158,n164);
or (n278,n160,n161,n162,n163);
not (n279,n280);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n279);
and (s0n281,notn281,n282);
and (s1n281,n279,1'b0);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n278);
and (s0n282,notn282,n283);
and (s1n282,n278,n291);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n272);
and (s0n283,notn283,n284);
and (s1n283,n272,n287);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n260);
and (s0n284,notn284,n285);
and (s1n284,n260,1'b0);
or (n285,n286,n157);
or (n286,n155,n156);
or (n287,1'b0,n183,n288,n290,1'b0);
and (n288,n289,n266);
or (n289,1'b0,n189,n264,1'b0);
and (n290,n193,n269);
or (n291,n170,n172);
not (n292,n293);
nor (n293,n54,n294,n310,n330,n347,n361,n372,n380);
wire s0n294,s1n294,notn294;
or (n294,s0n294,s1n294);
not(notn294,n251);
and (s0n294,notn294,1'b0);
and (s1n294,n251,n295);
or (n295,n296,n298,n300,n302,n304,n306,n308,1'b0);
and (n296,n297,n59);
xnor (n297,n72,n58);
and (n298,n299,n234);
xnor (n299,n74,n73);
and (n300,n301,n238);
xnor (n301,n76,n75);
and (n302,n303,n242);
xnor (n303,n78,n77);
and (n304,n305,n245);
xnor (n305,n89,n79);
and (n306,n307,n247);
xnor (n307,n84,n83);
and (n308,n309,n250);
xnor (n309,n93,n85);
wire s0n310,s1n310,notn310;
or (n310,s0n310,s1n310);
not(notn310,n251);
and (s0n310,notn310,1'b0);
and (s1n310,n251,n311);
or (n311,n312,n315,n318,n321,n324,n327,1'b0,1'b0);
and (n312,n313,n59);
xnor (n313,n73,n314);
or (n314,n72,n58);
and (n315,n316,n234);
xnor (n316,n75,n317);
or (n317,n74,n73);
and (n318,n319,n238);
xnor (n319,n77,n320);
or (n320,n76,n75);
and (n321,n322,n242);
xnor (n322,n79,n323);
or (n323,n78,n77);
and (n324,n325,n245);
xnor (n325,n83,n326);
or (n326,n89,n79);
and (n327,n328,n247);
xnor (n328,n85,n329);
or (n329,n84,n83);
wire s0n330,s1n330,notn330;
or (n330,s0n330,s1n330);
not(notn330,n251);
and (s0n330,notn330,1'b0);
and (s1n330,n251,n331);
or (n331,n332,n335,n338,n341,n344,1'b0,1'b0,1'b0);
and (n332,n333,n59);
xnor (n333,n74,n334);
or (n334,n73,n314);
and (n335,n336,n234);
xnor (n336,n76,n337);
or (n337,n75,n317);
and (n338,n339,n238);
xnor (n339,n78,n340);
or (n340,n77,n320);
and (n341,n342,n242);
xnor (n342,n89,n343);
or (n343,n79,n323);
and (n344,n345,n245);
xnor (n345,n84,n346);
or (n346,n83,n326);
wire s0n347,s1n347,notn347;
or (n347,s0n347,s1n347);
not(notn347,n251);
and (s0n347,notn347,1'b0);
and (s1n347,n251,n348);
or (n348,n349,n352,n355,n358,1'b0,1'b0,1'b0,1'b0);
and (n349,n350,n59);
xnor (n350,n75,n351);
or (n351,n74,n334);
and (n352,n353,n234);
xnor (n353,n77,n354);
or (n354,n76,n337);
and (n355,n356,n238);
xnor (n356,n79,n357);
or (n357,n78,n340);
and (n358,n359,n242);
xnor (n359,n83,n360);
or (n360,n89,n343);
wire s0n361,s1n361,notn361;
or (n361,s0n361,s1n361);
not(notn361,n251);
and (s0n361,notn361,1'b0);
and (s1n361,n251,n362);
or (n362,n363,n366,n369,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n363,n364,n59);
xnor (n364,n76,n365);
or (n365,n75,n351);
and (n366,n367,n234);
xnor (n367,n78,n368);
or (n368,n77,n354);
and (n369,n370,n238);
xnor (n370,n89,n371);
or (n371,n79,n357);
wire s0n372,s1n372,notn372;
or (n372,s0n372,s1n372);
not(notn372,n251);
and (s0n372,notn372,1'b0);
and (s1n372,n251,n373);
or (n373,n374,n377,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n374,n375,n59);
xnor (n375,n77,n376);
or (n376,n76,n365);
and (n377,n378,n234);
xnor (n378,n79,n379);
or (n379,n78,n368);
wire s0n380,s1n380,notn380;
or (n380,s0n380,s1n380);
not(notn380,n251);
and (s0n380,notn380,1'b0);
and (s1n380,n251,n381);
and (n381,n382,n59);
xnor (n382,n78,n383);
or (n383,n77,n376);
nor (n384,n385,n387,n390);
not (n385,n386);
not (n387,n388);
xor (n388,n389,n386);
xor (n390,n391,n392);
and (n392,n389,n386);
and (n393,n252,n281);
and (n394,n395,n396);
xor (n395,n294,n54);
nor (n396,n252,n397);
not (n397,n281);
and (n398,n54,n399);
and (n399,n252,n397);
not (n400,n401);
or (n401,1'b0,n402,n404,n408);
and (n402,n403,n393);
wire s0n403,s1n403,notn403;
or (n403,s0n403,s1n403);
not(notn403,n384);
and (s0n403,notn403,n294);
and (s1n403,n384,1'b0);
and (n404,n405,n396);
xor (n405,n406,n407);
not (n406,n310);
not (n407,n294);
and (n408,n294,n399);
or (n409,1'b0,n410,n412,n420);
and (n410,n411,n393);
wire s0n411,s1n411,notn411;
or (n411,s0n411,s1n411);
not(notn411,n384);
and (s0n411,notn411,n310);
and (s1n411,n384,1'b0);
and (n412,n413,n396);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n54);
and (s0n413,notn413,n414);
and (s1n413,n54,n417);
xor (n414,n415,n416);
not (n415,n330);
and (n416,n406,n407);
xor (n417,n330,n418);
and (n418,n310,n419);
and (n419,n294,n54);
and (n420,n310,n399);
not (n421,n422);
or (n422,1'b0,n423,n425,n432);
and (n423,n424,n393);
wire s0n424,s1n424,notn424;
or (n424,s0n424,s1n424);
not(notn424,n384);
and (s0n424,notn424,n330);
and (s1n424,n384,1'b0);
and (n425,n426,n396);
wire s0n426,s1n426,notn426;
or (n426,s0n426,s1n426);
not(notn426,n54);
and (s0n426,notn426,n427);
and (s1n426,n54,n430);
xor (n427,n428,n429);
not (n428,n347);
and (n429,n415,n416);
xor (n430,n347,n431);
and (n431,n330,n418);
and (n432,n330,n399);
or (n433,1'b0,n434,n436,n443);
and (n434,n435,n393);
wire s0n435,s1n435,notn435;
or (n435,s0n435,s1n435);
not(notn435,n384);
and (s0n435,notn435,n347);
and (s1n435,n384,1'b0);
and (n436,n437,n396);
wire s0n437,s1n437,notn437;
or (n437,s0n437,s1n437);
not(notn437,n54);
and (s0n437,notn437,n438);
and (s1n437,n54,n441);
xor (n438,n439,n440);
not (n439,n361);
and (n440,n428,n429);
xor (n441,n361,n442);
and (n442,n347,n431);
and (n443,n347,n399);
or (n444,1'b0,n445,n447,n454);
and (n445,n446,n393);
wire s0n446,s1n446,notn446;
or (n446,s0n446,s1n446);
not(notn446,n384);
and (s0n446,notn446,n361);
and (s1n446,n384,1'b0);
and (n447,n448,n396);
wire s0n448,s1n448,notn448;
or (n448,s0n448,s1n448);
not(notn448,n54);
and (s0n448,notn448,n449);
and (s1n448,n54,n452);
xor (n449,n450,n451);
not (n450,n372);
and (n451,n439,n440);
xor (n452,n372,n453);
and (n453,n361,n442);
and (n454,n361,n399);
or (n455,1'b0,n456,n458,n465);
and (n456,n457,n393);
wire s0n457,s1n457,notn457;
or (n457,s0n457,s1n457);
not(notn457,n384);
and (s0n457,notn457,n372);
and (s1n457,n384,1'b0);
and (n458,n459,n396);
wire s0n459,s1n459,notn459;
or (n459,s0n459,s1n459);
not(notn459,n54);
and (s0n459,notn459,n460);
and (s1n459,n54,n463);
xor (n460,n461,n462);
not (n461,n380);
and (n462,n450,n451);
xor (n463,n380,n464);
and (n464,n372,n453);
and (n465,n372,n399);
or (n466,1'b0,n467,n469,n474);
and (n467,n468,n393);
wire s0n468,s1n468,notn468;
or (n468,s0n468,s1n468);
not(notn468,n384);
and (s0n468,notn468,n380);
and (s1n468,n384,1'b0);
and (n469,n470,n396);
wire s0n470,s1n470,notn470;
or (n470,s0n470,s1n470);
not(notn470,n54);
and (s0n470,notn470,n471);
and (s1n470,n54,n473);
not (n471,n472);
and (n472,n461,n462);
and (n473,n380,n464);
and (n474,n380,n399);
nor (n475,n476,n400,n409,n421,n433,n444,n455,n466);
not (n476,n51);
nor (n477,n51,n401,n478,n421,n433,n444,n455,n466);
not (n478,n409);
nor (n479,n476,n401,n478,n421,n433,n444,n455,n466);
nor (n480,n51,n400,n478,n422,n481,n444,n455,n466);
not (n481,n433);
nor (n482,n476,n400,n478,n422,n481,n444,n455,n466);
nor (n483,n51,n401,n409,n421,n481,n444,n455,n466);
nor (n484,n476,n401,n409,n421,n481,n444,n455,n466);
or (n485,n486,n501);
or (n486,n487,n500);
or (n487,n488,n499);
or (n488,n489,n498);
or (n489,n490,n497);
or (n490,n491,n496);
or (n491,n492,n495);
or (n492,n493,n494);
nor (n493,n51,n400,n478,n422,n433,n444,n455,n466);
nor (n494,n476,n400,n478,n422,n433,n444,n455,n466);
nor (n495,n51,n401,n409,n421,n433,n444,n455,n466);
nor (n496,n476,n401,n409,n421,n433,n444,n455,n466);
nor (n497,n51,n400,n409,n422,n481,n444,n455,n466);
nor (n498,n476,n400,n409,n422,n481,n444,n455,n466);
nor (n499,n51,n401,n478,n422,n481,n444,n455,n466);
nor (n500,n476,n401,n478,n422,n481,n444,n455,n466);
or (n501,n502,n515);
or (n502,n503,n514);
or (n503,n504,n513);
or (n504,n505,n512);
or (n505,n506,n511);
or (n506,n507,n510);
or (n507,n508,n509);
nor (n508,n51,n400,n478,n421,n433,n444,n455,n466);
nor (n509,n476,n400,n478,n421,n433,n444,n455,n466);
nor (n510,n51,n401,n409,n422,n481,n444,n455,n466);
nor (n511,n476,n401,n409,n422,n481,n444,n455,n466);
nor (n512,n51,n400,n409,n421,n481,n444,n455,n466);
nor (n513,n476,n400,n409,n421,n481,n444,n455,n466);
nor (n514,n51,n401,n478,n421,n481,n444,n455,n466);
nor (n515,n476,n401,n478,n421,n481,n444,n455,n466);
nor (n516,n476,n401,n478,n422,n433,n444,n455,n466);
or (n517,1'b0,n518,n525,n532,n293);
or (n518,n519,n483);
or (n519,n520,n482);
or (n520,n521,n480);
or (n521,n522,n500);
or (n522,n523,n477);
or (n523,n524,n475);
or (n524,n496,n50);
or (n525,n526,n499);
or (n526,n527,n498);
or (n527,n528,n497);
or (n528,n529,n511);
or (n529,n530,n495);
or (n530,n531,n494);
or (n531,n516,n493);
or (n532,n533,n510);
or (n533,n534,n509);
or (n534,n535,n508);
or (n535,n536,n479);
or (n536,n537,n542);
or (n537,n538,n541);
or (n538,n539,n540);
nor (n539,n476,n401,n409,n422,n433,n444,n455,n466);
nor (n540,n51,n400,n409,n422,n433,n444,n455,n466);
nor (n541,n476,n400,n409,n422,n433,n444,n455,n466);
nor (n542,n51,n401,n478,n422,n433,n444,n455,n466);
or (n543,n544,n549);
nor (n544,n545,n546,n548);
not (n546,n547);
and (n549,n545,n547,n548);
nor (n550,n175,n181,n178,n179);
nor (n552,n553,n555,n556,n557);
not (n553,n554);
or (n558,1'b0,n559,n561,n565,n568);
and (n559,n560,n552);
and (n561,n562,n563);
nor (n563,n554,n564,n556,n557);
not (n564,n555);
and (n565,n566,n567);
nor (n567,n553,n564,n556,n557);
and (n568,n17,n569);
and (n569,n553,n564,n556,n570);
not (n570,n557);
and (n571,n36,n572);
not (n572,n573);
wire s0n573,s1n573,notn573;
or (n573,s0n573,s1n573);
not(notn573,n586);
and (s0n573,notn573,n19);
and (s1n573,n586,n574);
or (n574,n575,n579,n582,n584);
and (n575,n22,n576);
and (n576,n577,n578);
and (n579,n27,n580);
and (n580,n581,n578);
not (n581,n577);
and (n582,n31,n583);
nor (n583,n581,n578);
and (n584,n34,n585);
nor (n585,n577,n578);
and (n586,n37,n587);
not (n587,n551);
and (n588,n589,n645);
not (n589,n590);
wire s0n590,s1n590,notn590;
or (n590,s0n590,s1n590);
not(notn590,n36);
and (s0n590,notn590,1'b0);
and (s1n590,n36,n591);
wire s0n591,s1n591,notn591;
or (n591,s0n591,s1n591);
not(notn591,n644);
and (s0n591,notn591,n592);
and (s1n591,n644,n635);
or (n592,n593,n611,n622,n633);
and (n593,n594,n23);
wire s0n594,s1n594,notn594;
or (n594,s0n594,s1n594);
not(notn594,n573);
and (s0n594,notn594,n595);
and (s1n594,n573,n596);
or (n596,n597,n602,n606,n609);
and (n597,n598,n599);
nor (n599,n600,n601);
and (n602,n603,n604);
nor (n604,n605,n601);
not (n605,n600);
and (n606,n607,n608);
and (n608,n605,n601);
and (n609,n595,n610);
and (n610,n600,n601);
and (n611,n612,n28);
wire s0n612,s1n612,notn612;
or (n612,s0n612,s1n612);
not(notn612,n573);
and (s0n612,notn612,n613);
and (s1n612,n573,n614);
or (n614,n615,n617,n619,n621);
and (n615,n616,n599);
and (n617,n618,n604);
and (n619,n620,n608);
and (n621,n613,n610);
and (n622,n623,n32);
wire s0n623,s1n623,notn623;
or (n623,s0n623,s1n623);
not(notn623,n573);
and (s0n623,notn623,n624);
and (s1n623,n573,n625);
or (n625,n626,n628,n630,n632);
and (n626,n627,n599);
and (n628,n629,n604);
and (n630,n631,n608);
and (n632,n624,n610);
and (n633,n634,n35);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n573);
and (s0n634,notn634,n635);
and (s1n634,n573,n636);
or (n636,n637,n639,n641,n643);
and (n637,n638,n599);
and (n639,n640,n604);
and (n641,n642,n608);
and (n643,n635,n610);
and (n645,n646,n694);
not (n646,n647);
wire s0n647,s1n647,notn647;
or (n647,s0n647,s1n647);
not(notn647,n36);
and (s0n647,notn647,1'b0);
and (s1n647,n36,n648);
wire s0n648,s1n648,notn648;
or (n648,s0n648,s1n648);
not(notn648,n644);
and (s0n648,notn648,n649);
and (s1n648,n644,n685);
or (n649,n650,n661,n672,n683);
and (n650,n651,n23);
wire s0n651,s1n651,notn651;
or (n651,s0n651,s1n651);
not(notn651,n573);
and (s0n651,notn651,n652);
and (s1n651,n573,n653);
or (n653,n654,n656,n658,n660);
and (n654,n655,n599);
and (n656,n657,n604);
and (n658,n659,n608);
and (n660,n652,n610);
and (n661,n662,n28);
wire s0n662,s1n662,notn662;
or (n662,s0n662,s1n662);
not(notn662,n573);
and (s0n662,notn662,n663);
and (s1n662,n573,n664);
or (n664,n665,n667,n669,n671);
and (n665,n666,n599);
and (n667,n668,n604);
and (n669,n670,n608);
and (n671,n663,n610);
and (n672,n673,n32);
wire s0n673,s1n673,notn673;
or (n673,s0n673,s1n673);
not(notn673,n573);
and (s0n673,notn673,n674);
and (s1n673,n573,n675);
or (n675,n676,n678,n680,n682);
and (n676,n677,n599);
and (n678,n679,n604);
and (n680,n681,n608);
and (n682,n674,n610);
and (n683,n684,n35);
wire s0n684,s1n684,notn684;
or (n684,s0n684,s1n684);
not(notn684,n573);
and (s0n684,notn684,n685);
and (s1n684,n573,n686);
or (n686,n687,n689,n691,n693);
and (n687,n688,n599);
and (n689,n690,n604);
and (n691,n692,n608);
and (n693,n685,n610);
not (n694,n695);
wire s0n695,s1n695,notn695;
or (n695,s0n695,s1n695);
not(notn695,n36);
and (s0n695,notn695,1'b0);
and (s1n695,n36,n696);
wire s0n696,s1n696,notn696;
or (n696,s0n696,s1n696);
not(notn696,n644);
and (s0n696,notn696,n697);
and (s1n696,n644,n733);
or (n697,n698,n709,n720,n731);
and (n698,n699,n23);
wire s0n699,s1n699,notn699;
or (n699,s0n699,s1n699);
not(notn699,n573);
and (s0n699,notn699,n700);
and (s1n699,n573,n701);
or (n701,n702,n704,n706,n708);
and (n702,n703,n599);
and (n704,n705,n604);
and (n706,n707,n608);
and (n708,n700,n610);
and (n709,n710,n28);
wire s0n710,s1n710,notn710;
or (n710,s0n710,s1n710);
not(notn710,n573);
and (s0n710,notn710,n711);
and (s1n710,n573,n712);
or (n712,n713,n715,n717,n719);
and (n713,n714,n599);
and (n715,n716,n604);
and (n717,n718,n608);
and (n719,n711,n610);
and (n720,n721,n32);
wire s0n721,s1n721,notn721;
or (n721,s0n721,s1n721);
not(notn721,n573);
and (s0n721,notn721,n722);
and (s1n721,n573,n723);
or (n723,n724,n726,n728,n730);
and (n724,n725,n599);
and (n726,n727,n604);
and (n728,n729,n608);
and (n730,n722,n610);
and (n731,n732,n35);
wire s0n732,s1n732,notn732;
or (n732,s0n732,s1n732);
not(notn732,n573);
and (s0n732,notn732,n733);
and (s1n732,n573,n734);
or (n734,n735,n737,n739,n741);
and (n735,n736,n599);
and (n737,n738,n604);
and (n739,n740,n608);
and (n741,n733,n610);
or (n742,n743,n782);
and (n743,n744,n783);
xor (n744,n745,n760);
xor (n745,n746,n758);
wire s0n746,s1n746,notn746;
or (n746,s0n746,s1n746);
not(notn746,n588);
and (s0n746,notn746,1'b0);
and (s1n746,n588,n747);
wire s0n747,s1n747,notn747;
or (n747,s0n747,s1n747);
not(notn747,n571);
and (s0n747,notn747,n748);
and (s1n747,n571,n750);
wire s0n748,s1n748,notn748;
or (n748,s0n748,s1n748);
not(notn748,n18);
and (s0n748,notn748,1'b0);
and (s1n748,n18,n749);
or (n750,1'b0,n751,n753,n755,n757);
and (n751,n752,n552);
and (n753,n754,n563);
and (n755,n756,n567);
and (n757,n749,n569);
wire s0n758,s1n758,notn758;
or (n758,s0n758,s1n758);
not(notn758,n759);
and (s0n758,notn758,1'b0);
and (s1n758,n759,n15);
xor (n759,n589,n645);
or (n760,n761,n782);
and (n761,n762,n779);
xor (n762,n763,n764);
wire s0n763,s1n763,notn763;
or (n763,s0n763,s1n763);
not(notn763,n759);
and (s0n763,notn763,1'b0);
and (s1n763,n759,n747);
xor (n764,n765,n767);
wire s0n765,s1n765,notn765;
or (n765,s0n765,s1n765);
not(notn765,n766);
and (s0n765,notn765,1'b0);
and (s1n765,n766,n15);
xor (n766,n646,n694);
wire s0n767,s1n767,notn767;
or (n767,s0n767,s1n767);
not(notn767,n588);
and (s0n767,notn767,1'b0);
and (s1n767,n588,n768);
wire s0n768,s1n768,notn768;
or (n768,s0n768,s1n768);
not(notn768,n571);
and (s0n768,notn768,n769);
and (s1n768,n571,n771);
wire s0n769,s1n769,notn769;
or (n769,s0n769,s1n769);
not(notn769,n18);
and (s0n769,notn769,1'b0);
and (s1n769,n18,n770);
or (n771,1'b0,n772,n774,n776,n778);
and (n772,n773,n552);
and (n774,n775,n563);
and (n776,n777,n567);
and (n778,n770,n569);
and (n779,n780,n781);
wire s0n780,s1n780,notn780;
or (n780,s0n780,s1n780);
not(notn780,n766);
and (s0n780,notn780,1'b0);
and (s1n780,n766,n747);
wire s0n781,s1n781,notn781;
or (n781,s0n781,s1n781);
not(notn781,n695);
and (s0n781,notn781,1'b0);
and (s1n781,n695,n15);
and (n782,n763,n764);
nand (n783,n784,n930);
or (n784,n785,n925);
nor (n785,n786,n924);
and (n786,n787,n913);
nand (n787,n788,n912);
or (n788,n789,n846);
not (n789,n790);
or (n790,n791,n824);
xor (n791,n792,n821);
xor (n792,n793,n805);
wire s0n793,s1n793,notn793;
or (n793,s0n793,s1n793);
not(notn793,n759);
and (s0n793,notn793,1'b0);
and (s1n793,n759,n794);
wire s0n794,s1n794,notn794;
or (n794,s0n794,s1n794);
not(notn794,n571);
and (s0n794,notn794,n795);
and (s1n794,n571,n797);
wire s0n795,s1n795,notn795;
or (n795,s0n795,s1n795);
not(notn795,n18);
and (s0n795,notn795,1'b0);
and (s1n795,n18,n796);
or (n797,1'b0,n798,n800,n802,n804);
and (n798,n799,n552);
and (n800,n801,n563);
and (n802,n803,n567);
and (n804,n796,n569);
xor (n805,n806,n809);
xor (n806,n807,n808);
wire s0n807,s1n807,notn807;
or (n807,s0n807,s1n807);
not(notn807,n766);
and (s0n807,notn807,1'b0);
and (s1n807,n766,n768);
wire s0n808,s1n808,notn808;
or (n808,s0n808,s1n808);
not(notn808,n695);
and (s0n808,notn808,1'b0);
and (s1n808,n695,n747);
wire s0n809,s1n809,notn809;
or (n809,s0n809,s1n809);
not(notn809,n588);
and (s0n809,notn809,1'b0);
and (s1n809,n588,n810);
wire s0n810,s1n810,notn810;
or (n810,s0n810,s1n810);
not(notn810,n571);
and (s0n810,notn810,n811);
and (s1n810,n571,n813);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n18);
and (s0n811,notn811,1'b0);
and (s1n811,n18,n812);
or (n813,1'b0,n814,n816,n818,n820);
and (n814,n815,n552);
and (n816,n817,n563);
and (n818,n819,n567);
and (n820,n812,n569);
and (n821,n822,n823);
wire s0n822,s1n822,notn822;
or (n822,s0n822,s1n822);
not(notn822,n766);
and (s0n822,notn822,1'b0);
and (s1n822,n766,n794);
wire s0n823,s1n823,notn823;
or (n823,s0n823,s1n823);
not(notn823,n695);
and (s0n823,notn823,1'b0);
and (s1n823,n695,n768);
or (n824,n825,n845);
and (n825,n826,n842);
xor (n826,n827,n828);
wire s0n827,s1n827,notn827;
or (n827,s0n827,s1n827);
not(notn827,n759);
and (s0n827,notn827,1'b0);
and (s1n827,n759,n810);
xor (n828,n829,n830);
xor (n829,n822,n823);
wire s0n830,s1n830,notn830;
or (n830,s0n830,s1n830);
not(notn830,n588);
and (s0n830,notn830,1'b0);
and (s1n830,n588,n831);
wire s0n831,s1n831,notn831;
or (n831,s0n831,s1n831);
not(notn831,n571);
and (s0n831,notn831,n832);
and (s1n831,n571,n834);
wire s0n832,s1n832,notn832;
or (n832,s0n832,s1n832);
not(notn832,n18);
and (s0n832,notn832,1'b0);
and (s1n832,n18,n833);
or (n834,1'b0,n835,n837,n839,n841);
and (n835,n836,n552);
and (n837,n838,n563);
and (n839,n840,n567);
and (n841,n833,n569);
and (n842,n843,n844);
wire s0n843,s1n843,notn843;
or (n843,s0n843,s1n843);
not(notn843,n766);
and (s0n843,notn843,1'b0);
and (s1n843,n766,n810);
wire s0n844,s1n844,notn844;
or (n844,s0n844,s1n844);
not(notn844,n695);
and (s0n844,notn844,1'b0);
and (s1n844,n695,n794);
and (n845,n827,n828);
not (n846,n847);
nand (n847,n848,n908,n911);
nand (n848,n849,n873,n905);
or (n849,n850,n851);
xor (n850,n826,n842);
or (n851,n852,n872);
and (n852,n853,n858);
xor (n853,n854,n855);
wire s0n854,s1n854,notn854;
or (n854,s0n854,s1n854);
not(notn854,n759);
and (s0n854,notn854,1'b0);
and (s1n854,n759,n831);
and (n855,n856,n857);
wire s0n856,s1n856,notn856;
or (n856,s0n856,s1n856);
not(notn856,n766);
and (s0n856,notn856,1'b0);
and (s1n856,n766,n831);
wire s0n857,s1n857,notn857;
or (n857,s0n857,s1n857);
not(notn857,n695);
and (s0n857,notn857,1'b0);
and (s1n857,n695,n810);
xor (n858,n859,n860);
xor (n859,n843,n844);
wire s0n860,s1n860,notn860;
or (n860,s0n860,s1n860);
not(notn860,n588);
and (s0n860,notn860,1'b0);
and (s1n860,n588,n861);
wire s0n861,s1n861,notn861;
or (n861,s0n861,s1n861);
not(notn861,n571);
and (s0n861,notn861,n862);
and (s1n861,n571,n864);
wire s0n862,s1n862,notn862;
or (n862,s0n862,s1n862);
not(notn862,n18);
and (s0n862,notn862,1'b0);
and (s1n862,n18,n863);
or (n864,1'b0,n865,n867,n869,n871);
and (n865,n866,n552);
and (n867,n868,n563);
and (n869,n870,n567);
and (n871,n863,n569);
and (n872,n854,n855);
or (n873,n874,n904);
and (n874,n875,n899);
xor (n875,n876,n879);
and (n876,n877,n878);
wire s0n877,s1n877,notn877;
or (n877,s0n877,s1n877);
not(notn877,n766);
and (s0n877,notn877,1'b0);
and (s1n877,n766,n861);
wire s0n878,s1n878,notn878;
or (n878,s0n878,s1n878);
not(notn878,n695);
and (s0n878,notn878,1'b0);
and (s1n878,n695,n831);
or (n879,n880,n898);
and (n880,n881,n897);
xor (n881,n882,n896);
and (n882,n883,n895);
wire s0n883,s1n883,notn883;
or (n883,s0n883,s1n883);
not(notn883,n766);
and (s0n883,notn883,1'b0);
and (s1n883,n766,n884);
wire s0n884,s1n884,notn884;
or (n884,s0n884,s1n884);
not(notn884,n571);
and (s0n884,notn884,n885);
and (s1n884,n571,n887);
wire s0n885,s1n885,notn885;
or (n885,s0n885,s1n885);
not(notn885,n18);
and (s0n885,notn885,1'b0);
and (s1n885,n18,n886);
or (n887,1'b0,n888,n890,n892,n894);
and (n888,n889,n552);
and (n890,n891,n563);
and (n892,n893,n567);
and (n894,n886,n569);
wire s0n895,s1n895,notn895;
or (n895,s0n895,s1n895);
not(notn895,n695);
and (s0n895,notn895,1'b0);
and (s1n895,n695,n861);
wire s0n896,s1n896,notn896;
or (n896,s0n896,s1n896);
not(notn896,n759);
and (s0n896,notn896,1'b0);
and (s1n896,n759,n884);
xor (n897,n877,n878);
and (n898,n882,n896);
xor (n899,n900,n903);
xor (n900,n901,n902);
wire s0n901,s1n901,notn901;
or (n901,s0n901,s1n901);
not(notn901,n588);
and (s0n901,notn901,1'b0);
and (s1n901,n588,n884);
xor (n902,n856,n857);
wire s0n903,s1n903,notn903;
or (n903,s0n903,s1n903);
not(notn903,n759);
and (s0n903,notn903,1'b0);
and (s1n903,n759,n861);
and (n904,n876,n879);
or (n905,n906,n907);
xor (n906,n853,n858);
and (n907,n900,n903);
nand (n908,n909,n849);
not (n909,n910);
nand (n910,n906,n907);
nand (n911,n850,n851);
nand (n912,n791,n824);
or (n913,n914,n921);
xor (n914,n915,n920);
xor (n915,n916,n917);
wire s0n916,s1n916,notn916;
or (n916,s0n916,s1n916);
not(notn916,n759);
and (s0n916,notn916,1'b0);
and (s1n916,n759,n768);
xor (n917,n918,n919);
xor (n918,n780,n781);
wire s0n919,s1n919,notn919;
or (n919,s0n919,s1n919);
not(notn919,n588);
and (s0n919,notn919,1'b0);
and (s1n919,n588,n794);
and (n920,n807,n808);
or (n921,n922,n923);
and (n922,n792,n821);
and (n923,n793,n805);
and (n924,n914,n921);
nor (n925,n926,n929);
or (n926,n927,n928);
and (n927,n915,n920);
and (n928,n916,n917);
xor (n929,n762,n779);
nand (n930,n926,n929);
xor (n931,n932,n980);
not (n932,n933);
wire s0n933,s1n933,notn933;
or (n933,s0n933,s1n933);
not(notn933,n36);
and (s0n933,notn933,1'b0);
and (s1n933,n36,n934);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n644);
and (s0n934,notn934,n935);
and (s1n934,n644,n971);
or (n935,n936,n947,n958,n969);
and (n936,n937,n23);
wire s0n937,s1n937,notn937;
or (n937,s0n937,s1n937);
not(notn937,n573);
and (s0n937,notn937,n938);
and (s1n937,n573,n939);
or (n939,n940,n942,n944,n946);
and (n940,n941,n599);
and (n942,n943,n604);
and (n944,n945,n608);
and (n946,n938,n610);
and (n947,n948,n28);
wire s0n948,s1n948,notn948;
or (n948,s0n948,s1n948);
not(notn948,n573);
and (s0n948,notn948,n949);
and (s1n948,n573,n950);
or (n950,n951,n953,n955,n957);
and (n951,n952,n599);
and (n953,n954,n604);
and (n955,n956,n608);
and (n957,n949,n610);
and (n958,n959,n32);
wire s0n959,s1n959,notn959;
or (n959,s0n959,s1n959);
not(notn959,n573);
and (s0n959,notn959,n960);
and (s1n959,n573,n961);
or (n961,n962,n964,n966,n968);
and (n962,n963,n599);
and (n964,n965,n604);
and (n966,n967,n608);
and (n968,n960,n610);
and (n969,n970,n35);
wire s0n970,s1n970,notn970;
or (n970,s0n970,s1n970);
not(notn970,n573);
and (s0n970,notn970,n971);
and (s1n970,n573,n972);
or (n972,n973,n975,n977,n979);
and (n973,n974,n599);
and (n975,n976,n604);
and (n977,n978,n608);
and (n979,n971,n610);
not (n980,n981);
wire s0n981,s1n981,notn981;
or (n981,s0n981,s1n981);
not(notn981,n36);
and (s0n981,notn981,1'b0);
and (s1n981,n36,n982);
wire s0n982,s1n982,notn982;
or (n982,s0n982,s1n982);
not(notn982,n644);
and (s0n982,notn982,n983);
and (s1n982,n644,n1019);
or (n983,n984,n995,n1006,n1017);
and (n984,n985,n23);
wire s0n985,s1n985,notn985;
or (n985,s0n985,s1n985);
not(notn985,n573);
and (s0n985,notn985,n986);
and (s1n985,n573,n987);
or (n987,n988,n990,n992,n994);
and (n988,n989,n599);
and (n990,n991,n604);
and (n992,n993,n608);
and (n994,n986,n610);
and (n995,n996,n28);
wire s0n996,s1n996,notn996;
or (n996,s0n996,s1n996);
not(notn996,n573);
and (s0n996,notn996,n997);
and (s1n996,n573,n998);
or (n998,n999,n1001,n1003,n1005);
and (n999,n1000,n599);
and (n1001,n1002,n604);
and (n1003,n1004,n608);
and (n1005,n997,n610);
and (n1006,n1007,n32);
wire s0n1007,s1n1007,notn1007;
or (n1007,s0n1007,s1n1007);
not(notn1007,n573);
and (s0n1007,notn1007,n1008);
and (s1n1007,n573,n1009);
or (n1009,n1010,n1012,n1014,n1016);
and (n1010,n1011,n599);
and (n1012,n1013,n604);
and (n1014,n1015,n608);
and (n1016,n1008,n610);
and (n1017,n1018,n35);
wire s0n1018,s1n1018,notn1018;
or (n1018,s0n1018,s1n1018);
not(notn1018,n573);
and (s0n1018,notn1018,n1019);
and (s1n1018,n573,n1020);
or (n1020,n1021,n1023,n1025,n1027);
and (n1021,n1022,n599);
and (n1023,n1024,n604);
and (n1025,n1026,n608);
and (n1027,n1019,n610);
and (n1028,n1029,n1224);
xor (n1029,n1030,n1078);
xor (n1030,n1031,n1056);
xor (n1031,n1032,n1044);
and (n1032,n759,n1033);
wire s0n1033,s1n1033,notn1033;
or (n1033,s0n1033,s1n1033);
not(notn1033,n571);
and (s0n1033,notn1033,n1034);
and (s1n1033,n571,n1036);
wire s0n1034,s1n1034,notn1034;
or (n1034,s0n1034,s1n1034);
not(notn1034,n18);
and (s0n1034,notn1034,1'b0);
and (s1n1034,n18,n1035);
or (n1036,1'b0,n1037,n1039,n1041,n1043);
and (n1037,n1038,n552);
and (n1039,n1040,n563);
and (n1041,n1042,n567);
and (n1043,n1035,n569);
and (n1044,n588,n1045);
wire s0n1045,s1n1045,notn1045;
or (n1045,s0n1045,s1n1045);
not(notn1045,n571);
and (s0n1045,notn1045,n1046);
and (s1n1045,n571,n1048);
wire s0n1046,s1n1046,notn1046;
or (n1046,s0n1046,s1n1046);
not(notn1046,n18);
and (s0n1046,notn1046,1'b0);
and (s1n1046,n18,n1047);
or (n1048,1'b0,n1049,n1051,n1053,n1055);
and (n1049,n1050,n552);
and (n1051,n1052,n563);
and (n1053,n1054,n567);
and (n1055,n1047,n569);
or (n1056,n1057,n1077);
and (n1057,n1058,n1074);
xor (n1058,n1059,n1073);
xor (n1059,n1060,n1061);
and (n1060,n766,n1033);
and (n1061,n588,n1062);
wire s0n1062,s1n1062,notn1062;
or (n1062,s0n1062,s1n1062);
not(notn1062,n571);
and (s0n1062,notn1062,n1063);
and (s1n1062,n571,n1065);
wire s0n1063,s1n1063,notn1063;
or (n1063,s0n1063,s1n1063);
not(notn1063,n18);
and (s0n1063,notn1063,1'b0);
and (s1n1063,n18,n1064);
or (n1065,1'b0,n1066,n1068,n1070,n1072);
and (n1066,n1067,n552);
and (n1068,n1069,n563);
and (n1070,n1071,n567);
and (n1072,n1064,n569);
and (n1073,n759,n1045);
and (n1074,n1075,n1076);
and (n1075,n766,n1045);
wire s0n1076,s1n1076,notn1076;
or (n1076,s0n1076,s1n1076);
not(notn1076,n695);
and (s0n1076,notn1076,1'b0);
and (s1n1076,n695,n1033);
and (n1077,n1059,n1073);
or (n1078,n1079,n1223);
and (n1079,n1080,n1104);
xor (n1080,n1081,n1103);
or (n1081,n1082,n1102);
and (n1082,n1083,n1099);
xor (n1083,n1084,n1098);
xor (n1084,n1085,n1086);
xor (n1085,n1075,n1076);
and (n1086,n588,n1087);
wire s0n1087,s1n1087,notn1087;
or (n1087,s0n1087,s1n1087);
not(notn1087,n571);
and (s0n1087,notn1087,n1088);
and (s1n1087,n571,n1090);
wire s0n1088,s1n1088,notn1088;
or (n1088,s0n1088,s1n1088);
not(notn1088,n18);
and (s0n1088,notn1088,1'b0);
and (s1n1088,n18,n1089);
or (n1090,1'b0,n1091,n1093,n1095,n1097);
and (n1091,n1092,n552);
and (n1093,n1094,n563);
and (n1095,n1096,n567);
and (n1097,n1089,n569);
and (n1098,n759,n1062);
and (n1099,n1100,n1101);
wire s0n1100,s1n1100,notn1100;
or (n1100,s0n1100,s1n1100);
not(notn1100,n695);
and (s0n1100,notn1100,1'b0);
and (s1n1100,n695,n1045);
and (n1101,n766,n1062);
and (n1102,n1084,n1098);
xor (n1103,n1058,n1074);
or (n1104,n1105,n1222);
and (n1105,n1106,n1130);
xor (n1106,n1107,n1129);
or (n1107,n1108,n1128);
and (n1108,n1109,n1125);
xor (n1109,n1110,n1111);
and (n1110,n759,n1087);
xor (n1111,n1112,n1113);
xor (n1112,n1100,n1101);
and (n1113,n588,n1114);
wire s0n1114,s1n1114,notn1114;
or (n1114,s0n1114,s1n1114);
not(notn1114,n571);
and (s0n1114,notn1114,n1115);
and (s1n1114,n571,n1117);
wire s0n1115,s1n1115,notn1115;
or (n1115,s0n1115,s1n1115);
not(notn1115,n18);
and (s0n1115,notn1115,1'b0);
and (s1n1115,n18,n1116);
or (n1117,1'b0,n1118,n1120,n1122,n1124);
and (n1118,n1119,n552);
and (n1120,n1121,n563);
and (n1122,n1123,n567);
and (n1124,n1116,n569);
and (n1125,n1126,n1127);
wire s0n1126,s1n1126,notn1126;
or (n1126,s0n1126,s1n1126);
not(notn1126,n695);
and (s0n1126,notn1126,1'b0);
and (s1n1126,n695,n1062);
and (n1127,n766,n1087);
and (n1128,n1110,n1111);
xor (n1129,n1083,n1099);
or (n1130,n1131,n1221);
and (n1131,n1132,n1156);
xor (n1132,n1133,n1155);
or (n1133,n1134,n1154);
and (n1134,n1135,n1151);
xor (n1135,n1136,n1137);
and (n1136,n759,n1114);
xor (n1137,n1138,n1139);
xor (n1138,n1126,n1127);
and (n1139,n588,n1140);
wire s0n1140,s1n1140,notn1140;
or (n1140,s0n1140,s1n1140);
not(notn1140,n571);
and (s0n1140,notn1140,n1141);
and (s1n1140,n571,n1143);
wire s0n1141,s1n1141,notn1141;
or (n1141,s0n1141,s1n1141);
not(notn1141,n18);
and (s0n1141,notn1141,1'b0);
and (s1n1141,n18,n1142);
or (n1143,1'b0,n1144,n1146,n1148,n1150);
and (n1144,n1145,n552);
and (n1146,n1147,n563);
and (n1148,n1149,n567);
and (n1150,n1142,n569);
and (n1151,n1152,n1153);
and (n1152,n766,n1114);
wire s0n1153,s1n1153,notn1153;
or (n1153,s0n1153,s1n1153);
not(notn1153,n695);
and (s0n1153,notn1153,1'b0);
and (s1n1153,n695,n1087);
and (n1154,n1136,n1137);
xor (n1155,n1109,n1125);
or (n1156,n1157,n1220);
and (n1157,n1158,n1182);
xor (n1158,n1159,n1181);
or (n1159,n1160,n1180);
and (n1160,n1161,n1166);
xor (n1161,n1162,n1163);
and (n1162,n759,n1140);
and (n1163,n1164,n1165);
wire s0n1164,s1n1164,notn1164;
or (n1164,s0n1164,s1n1164);
not(notn1164,n695);
and (s0n1164,notn1164,1'b0);
and (s1n1164,n695,n1114);
and (n1165,n766,n1140);
xor (n1166,n1167,n1168);
xor (n1167,n1152,n1153);
and (n1168,n588,n1169);
wire s0n1169,s1n1169,notn1169;
or (n1169,s0n1169,s1n1169);
not(notn1169,n571);
and (s0n1169,notn1169,n1170);
and (s1n1169,n571,n1172);
wire s0n1170,s1n1170,notn1170;
or (n1170,s0n1170,s1n1170);
not(notn1170,n18);
and (s0n1170,notn1170,1'b0);
and (s1n1170,n18,n1171);
or (n1172,1'b0,n1173,n1175,n1177,n1179);
and (n1173,n1174,n552);
and (n1175,n1176,n563);
and (n1177,n1178,n567);
and (n1179,n1171,n569);
and (n1180,n1162,n1163);
xor (n1181,n1135,n1151);
or (n1182,n1183,n1219);
and (n1183,n1184,n1202);
xor (n1184,n1185,n1201);
and (n1185,n1186,n1200);
xor (n1186,n1187,n1199);
and (n1187,n588,n1188);
wire s0n1188,s1n1188,notn1188;
or (n1188,s0n1188,s1n1188);
not(notn1188,n571);
and (s0n1188,notn1188,n1189);
and (s1n1188,n571,n1191);
wire s0n1189,s1n1189,notn1189;
or (n1189,s0n1189,s1n1189);
not(notn1189,n18);
and (s0n1189,notn1189,1'b0);
and (s1n1189,n18,n1190);
or (n1191,1'b0,n1192,n1194,n1196,n1198);
and (n1192,n1193,n552);
and (n1194,n1195,n563);
and (n1196,n1197,n567);
and (n1198,n1190,n569);
and (n1199,n759,n1169);
xor (n1200,n1164,n1165);
xor (n1201,n1161,n1166);
or (n1202,n1203,n1218);
and (n1203,n1204,n1217);
xor (n1204,n1205,n1208);
and (n1205,n1206,n1207);
wire s0n1206,s1n1206,notn1206;
or (n1206,s0n1206,s1n1206);
not(notn1206,n695);
and (s0n1206,notn1206,1'b0);
and (s1n1206,n695,n1140);
and (n1207,n766,n1169);
or (n1208,n1209,n1216);
and (n1209,n1210,n1215);
xor (n1210,n1211,n1214);
and (n1211,n1212,n1213);
and (n1212,n766,n1188);
wire s0n1213,s1n1213,notn1213;
or (n1213,s0n1213,s1n1213);
not(notn1213,n695);
and (s0n1213,notn1213,1'b0);
and (s1n1213,n695,n1169);
xor (n1214,n1206,n1207);
and (n1215,n759,n1188);
and (n1216,n1211,n1214);
xor (n1217,n1186,n1200);
and (n1218,n1205,n1208);
and (n1219,n1185,n1201);
and (n1220,n1159,n1181);
and (n1221,n1133,n1155);
and (n1222,n1107,n1129);
and (n1223,n1081,n1103);
wire s0n1224,s1n1224,notn1224;
or (n1224,s0n1224,s1n1224);
not(notn1224,n36);
and (s0n1224,notn1224,1'b0);
and (s1n1224,n36,n1225);
wire s0n1225,s1n1225,notn1225;
or (n1225,s0n1225,s1n1225);
not(notn1225,n644);
and (s0n1225,notn1225,n1226);
and (s1n1225,n644,n1262);
or (n1226,n1227,n1238,n1249,n1260);
and (n1227,n1228,n23);
wire s0n1228,s1n1228,notn1228;
or (n1228,s0n1228,s1n1228);
not(notn1228,n573);
and (s0n1228,notn1228,n1229);
and (s1n1228,n573,n1230);
or (n1230,n1231,n1233,n1235,n1237);
and (n1231,n1232,n599);
and (n1233,n1234,n604);
and (n1235,n1236,n608);
and (n1237,n1229,n610);
and (n1238,n1239,n28);
wire s0n1239,s1n1239,notn1239;
or (n1239,s0n1239,s1n1239);
not(notn1239,n573);
and (s0n1239,notn1239,n1240);
and (s1n1239,n573,n1241);
or (n1241,n1242,n1244,n1246,n1248);
and (n1242,n1243,n599);
and (n1244,n1245,n604);
and (n1246,n1247,n608);
and (n1248,n1240,n610);
and (n1249,n1250,n32);
wire s0n1250,s1n1250,notn1250;
or (n1250,s0n1250,s1n1250);
not(notn1250,n573);
and (s0n1250,notn1250,n1251);
and (s1n1250,n573,n1252);
or (n1252,n1253,n1255,n1257,n1259);
and (n1253,n1254,n599);
and (n1255,n1256,n604);
and (n1257,n1258,n608);
and (n1259,n1251,n610);
and (n1260,n1261,n35);
wire s0n1261,s1n1261,notn1261;
or (n1261,s0n1261,s1n1261);
not(notn1261,n573);
and (s0n1261,notn1261,n1262);
and (s1n1261,n573,n1263);
or (n1263,n1264,n1266,n1268,n1270);
and (n1264,n1265,n599);
and (n1266,n1267,n604);
and (n1268,n1269,n608);
and (n1270,n1262,n610);
and (n1271,n1272,n1273);
xor (n1272,n744,n783);
xor (n1273,n1274,n1275);
not (n1274,n1224);
and (n1275,n932,n980);
xor (n1276,n1277,n1768);
xor (n1277,n1278,n1734);
or (n1278,n1279,n1733);
and (n1279,n1280,n1602);
xor (n1280,n1281,n1589);
and (n1281,n1282,n1515);
xor (n1282,n1283,n1425);
wire s0n1283,s1n1283,notn1283;
or (n1283,s0n1283,s1n1283);
not(notn1283,n1424);
and (s0n1283,notn1283,1'b0);
and (s1n1283,n1424,n1284);
xor (n1284,n1285,n1395);
xor (n1285,n1286,n1299);
not (n1286,n1287);
nand (n1287,n590,n1288);
wire s0n1288,s1n1288,notn1288;
or (n1288,s0n1288,s1n1288);
not(notn1288,n571);
and (s0n1288,notn1288,n1289);
and (s1n1288,n571,n1291);
wire s0n1289,s1n1289,notn1289;
or (n1289,s0n1289,s1n1289);
not(notn1289,n18);
and (s0n1289,notn1289,1'b0);
and (s1n1289,n18,n1290);
or (n1291,1'b0,n1292,n1294,n1296,n1298);
and (n1292,n1293,n552);
and (n1294,n1295,n563);
and (n1296,n1297,n567);
and (n1298,n1290,n569);
xor (n1299,n1300,n1325);
xor (n1300,n1301,n1313);
wire s0n1301,s1n1301,notn1301;
or (n1301,s0n1301,s1n1301);
not(notn1301,n647);
and (s0n1301,notn1301,1'b0);
and (s1n1301,n647,n1302);
wire s0n1302,s1n1302,notn1302;
or (n1302,s0n1302,s1n1302);
not(notn1302,n571);
and (s0n1302,notn1302,n1303);
and (s1n1302,n571,n1305);
wire s0n1303,s1n1303,notn1303;
or (n1303,s0n1303,s1n1303);
not(notn1303,n18);
and (s0n1303,notn1303,1'b0);
and (s1n1303,n18,n1304);
or (n1305,1'b0,n1306,n1308,n1310,n1312);
and (n1306,n1307,n552);
and (n1308,n1309,n563);
and (n1310,n1311,n567);
and (n1312,n1304,n569);
wire s0n1313,s1n1313,notn1313;
or (n1313,s0n1313,s1n1313);
not(notn1313,n695);
and (s0n1313,notn1313,1'b0);
and (s1n1313,n695,n1314);
wire s0n1314,s1n1314,notn1314;
or (n1314,s0n1314,s1n1314);
not(notn1314,n571);
and (s0n1314,notn1314,n1315);
and (s1n1314,n571,n1317);
wire s0n1315,s1n1315,notn1315;
or (n1315,s0n1315,s1n1315);
not(notn1315,n18);
and (s0n1315,notn1315,1'b0);
and (s1n1315,n18,n1316);
or (n1317,1'b0,n1318,n1320,n1322,n1324);
and (n1318,n1319,n552);
and (n1320,n1321,n563);
and (n1322,n1323,n567);
and (n1324,n1316,n569);
or (n1325,n1326,n1329,n1394);
and (n1326,n1327,n1328);
wire s0n1327,s1n1327,notn1327;
or (n1327,s0n1327,s1n1327);
not(notn1327,n647);
and (s0n1327,notn1327,1'b0);
and (s1n1327,n647,n1288);
wire s0n1328,s1n1328,notn1328;
or (n1328,s0n1328,s1n1328);
not(notn1328,n695);
and (s0n1328,notn1328,1'b0);
and (s1n1328,n695,n1302);
and (n1329,n1328,n1330);
or (n1330,n1331,n1345,n1393);
and (n1331,n1332,n1344);
wire s0n1332,s1n1332,notn1332;
or (n1332,s0n1332,s1n1332);
not(notn1332,n647);
and (s0n1332,notn1332,1'b0);
and (s1n1332,n647,n1333);
wire s0n1333,s1n1333,notn1333;
or (n1333,s0n1333,s1n1333);
not(notn1333,n571);
and (s0n1333,notn1333,n1334);
and (s1n1333,n571,n1336);
wire s0n1334,s1n1334,notn1334;
or (n1334,s0n1334,s1n1334);
not(notn1334,n18);
and (s0n1334,notn1334,1'b0);
and (s1n1334,n18,n1335);
or (n1336,1'b0,n1337,n1339,n1341,n1343);
and (n1337,n1338,n552);
and (n1339,n1340,n563);
and (n1341,n1342,n567);
and (n1343,n1335,n569);
wire s0n1344,s1n1344,notn1344;
or (n1344,s0n1344,s1n1344);
not(notn1344,n695);
and (s0n1344,notn1344,1'b0);
and (s1n1344,n695,n1288);
and (n1345,n1344,n1346);
or (n1346,n1347,n1361,n1363);
and (n1347,n1348,n1360);
wire s0n1348,s1n1348,notn1348;
or (n1348,s0n1348,s1n1348);
not(notn1348,n647);
and (s0n1348,notn1348,1'b0);
and (s1n1348,n647,n1349);
wire s0n1349,s1n1349,notn1349;
or (n1349,s0n1349,s1n1349);
not(notn1349,n571);
and (s0n1349,notn1349,n1350);
and (s1n1349,n571,n1352);
wire s0n1350,s1n1350,notn1350;
or (n1350,s0n1350,s1n1350);
not(notn1350,n18);
and (s0n1350,notn1350,1'b0);
and (s1n1350,n18,n1351);
or (n1352,1'b0,n1353,n1355,n1357,n1359);
and (n1353,n1354,n552);
and (n1355,n1356,n563);
and (n1357,n1358,n567);
and (n1359,n1351,n569);
wire s0n1360,s1n1360,notn1360;
or (n1360,s0n1360,s1n1360);
not(notn1360,n695);
and (s0n1360,notn1360,1'b0);
and (s1n1360,n695,n1333);
and (n1361,n1360,n1362);
or (n1362,n1363,n1378,n1379);
and (n1363,n1364,n1377);
not (n1364,n1365);
nand (n1365,n647,n1366);
wire s0n1366,s1n1366,notn1366;
or (n1366,s0n1366,s1n1366);
not(notn1366,n571);
and (s0n1366,notn1366,n1367);
and (s1n1366,n571,n1369);
wire s0n1367,s1n1367,notn1367;
or (n1367,s0n1367,s1n1367);
not(notn1367,n18);
and (s0n1367,notn1367,1'b0);
and (s1n1367,n18,n1368);
or (n1369,1'b0,n1370,n1372,n1374,n1376);
and (n1370,n1371,n552);
and (n1372,n1373,n563);
and (n1374,n1375,n567);
and (n1376,n1368,n569);
wire s0n1377,s1n1377,notn1377;
or (n1377,s0n1377,s1n1377);
not(notn1377,n695);
and (s0n1377,notn1377,1'b0);
and (s1n1377,n695,n1349);
and (n1378,n1377,n1379);
and (n1379,n1380,n1392);
wire s0n1380,s1n1380,notn1380;
or (n1380,s0n1380,s1n1380);
not(notn1380,n647);
and (s0n1380,notn1380,1'b0);
and (s1n1380,n647,n1381);
wire s0n1381,s1n1381,notn1381;
or (n1381,s0n1381,s1n1381);
not(notn1381,n571);
and (s0n1381,notn1381,n1382);
and (s1n1381,n571,n1384);
wire s0n1382,s1n1382,notn1382;
or (n1382,s0n1382,s1n1382);
not(notn1382,n18);
and (s0n1382,notn1382,1'b0);
and (s1n1382,n18,n1383);
or (n1384,1'b0,n1385,n1387,n1389,n1391);
and (n1385,n1386,n552);
and (n1387,n1388,n563);
and (n1389,n1390,n567);
and (n1391,n1383,n569);
wire s0n1392,s1n1392,notn1392;
or (n1392,s0n1392,s1n1392);
not(notn1392,n695);
and (s0n1392,notn1392,1'b0);
and (s1n1392,n695,n1366);
and (n1393,n1332,n1346);
and (n1394,n1327,n1330);
or (n1395,n1396,n1401,n1423);
and (n1396,n1397,n1399);
not (n1397,n1398);
nand (n1398,n590,n1333);
xor (n1399,n1400,n1330);
xor (n1400,n1327,n1328);
and (n1401,n1399,n1402);
or (n1402,n1403,n1408,n1422);
and (n1403,n1404,n1406);
not (n1404,n1405);
nand (n1405,n590,n1349);
xor (n1406,n1407,n1346);
xor (n1407,n1332,n1344);
and (n1408,n1406,n1409);
or (n1409,n1410,n1415,n1421);
and (n1410,n1411,n1413);
not (n1411,n1412);
nand (n1412,n590,n1366);
xor (n1413,n1414,n1362);
xor (n1414,n1348,n1360);
and (n1415,n1413,n1416);
and (n1416,n1417,n1419);
not (n1417,n1418);
nand (n1418,n590,n1381);
xor (n1419,n1420,n1379);
xor (n1420,n1364,n1377);
and (n1421,n1411,n1416);
and (n1422,n1404,n1409);
and (n1423,n1397,n1402);
and (n1424,n1274,n1275);
xor (n1425,n1426,n1473);
xor (n1426,n1427,n1458);
xor (n1427,n1428,n1456);
xor (n1428,n1429,n1443);
nor (n1429,n1430,n980);
not (n1430,n1431);
wire s0n1431,s1n1431,notn1431;
or (n1431,s0n1431,s1n1431);
not(notn1431,n590);
and (s0n1431,notn1431,1'b0);
and (s1n1431,n590,n1432);
wire s0n1432,s1n1432,notn1432;
or (n1432,s0n1432,s1n1432);
not(notn1432,n571);
and (s0n1432,notn1432,n1433);
and (s1n1432,n571,n1435);
wire s0n1433,s1n1433,notn1433;
or (n1433,s0n1433,s1n1433);
not(notn1433,n18);
and (s0n1433,notn1433,1'b0);
and (s1n1433,n18,n1434);
or (n1435,1'b0,n1436,n1438,n1440,n1442);
and (n1436,n1437,n552);
and (n1438,n1439,n563);
and (n1440,n1441,n567);
and (n1442,n1434,n569);
and (n1443,n1444,n981);
and (n1444,n590,n1445);
wire s0n1445,s1n1445,notn1445;
or (n1445,s0n1445,s1n1445);
not(notn1445,n571);
and (s0n1445,notn1445,n1446);
and (s1n1445,n571,n1448);
wire s0n1446,s1n1446,notn1446;
or (n1446,s0n1446,s1n1446);
not(notn1446,n18);
and (s0n1446,notn1446,1'b0);
and (s1n1446,n18,n1447);
or (n1448,1'b0,n1449,n1451,n1453,n1455);
and (n1449,n1450,n552);
and (n1451,n1452,n563);
and (n1453,n1454,n567);
and (n1455,n1447,n569);
and (n1456,n1443,n1457);
wire s0n1457,s1n1457,notn1457;
or (n1457,s0n1457,s1n1457);
not(notn1457,n647);
and (s0n1457,notn1457,1'b0);
and (s1n1457,n647,n1314);
and (n1458,n1429,n1459);
not (n1459,n1460);
not (n1460,n1461);
wire s0n1461,s1n1461,notn1461;
or (n1461,s0n1461,s1n1461);
not(notn1461,n647);
and (s0n1461,notn1461,1'b0);
and (s1n1461,n647,n1462);
wire s0n1462,s1n1462,notn1462;
or (n1462,s0n1462,s1n1462);
not(notn1462,n571);
and (s0n1462,notn1462,n1463);
and (s1n1462,n571,n1465);
wire s0n1463,s1n1463,notn1463;
or (n1463,s0n1463,s1n1463);
not(notn1463,n18);
and (s0n1463,notn1463,1'b0);
and (s1n1463,n18,n1464);
or (n1465,1'b0,n1466,n1468,n1470,n1472);
and (n1466,n1467,n552);
and (n1468,n1469,n563);
and (n1470,n1471,n567);
and (n1472,n1464,n569);
or (n1473,n1474,n1514);
and (n1474,n1475,n1492);
xor (n1475,n1476,n1483);
nor (n1476,n1477,n980);
xnor (n1477,n1478,n1481);
not (n1478,n1479);
not (n1479,n1480);
nand (n1480,n590,n1314);
not (n1481,n1482);
wire s0n1482,s1n1482,notn1482;
or (n1482,s0n1482,s1n1482);
not(notn1482,n647);
and (s0n1482,notn1482,1'b0);
and (s1n1482,n647,n1445);
and (n1483,n1484,n981);
nand (n1484,n1485,n1491);
or (n1485,n1486,n1488);
not (n1486,n1487);
wire s0n1487,s1n1487,notn1487;
or (n1487,s0n1487,s1n1487);
not(notn1487,n647);
and (s0n1487,notn1487,1'b0);
and (s1n1487,n647,n1432);
not (n1488,n1489);
not (n1489,n1490);
wire s0n1490,s1n1490,notn1490;
or (n1490,s0n1490,s1n1490);
not(notn1490,n590);
and (s0n1490,notn1490,1'b0);
and (s1n1490,n590,n1462);
or (n1491,n1489,n1487);
and (n1492,n1493,n981);
or (n1493,n1494,n1511);
nor (n1494,n1495,n1460);
and (n1495,n1496,n1509);
not (n1496,n1497);
wire s0n1497,s1n1497,notn1497;
or (n1497,s0n1497,s1n1497);
not(notn1497,n590);
and (s0n1497,notn1497,1'b0);
and (s1n1497,n590,n1498);
wire s0n1498,s1n1498,notn1498;
or (n1498,s0n1498,s1n1498);
not(notn1498,n571);
and (s0n1498,notn1498,n1499);
and (s1n1498,n571,n1501);
wire s0n1499,s1n1499,notn1499;
or (n1499,s0n1499,s1n1499);
not(notn1499,n18);
and (s0n1499,notn1499,1'b0);
and (s1n1499,n18,n1500);
or (n1501,1'b0,n1502,n1504,n1506,n1508);
and (n1502,n1503,n552);
and (n1504,n1505,n563);
and (n1506,n1507,n567);
and (n1508,n1500,n569);
not (n1509,n1510);
wire s0n1510,s1n1510,notn1510;
or (n1510,s0n1510,s1n1510);
not(notn1510,n695);
and (s0n1510,notn1510,1'b0);
and (s1n1510,n695,n1432);
nor (n1511,n1512,n1430);
not (n1512,n1513);
wire s0n1513,s1n1513,notn1513;
or (n1513,s0n1513,s1n1513);
not(notn1513,n695);
and (s0n1513,notn1513,1'b0);
and (s1n1513,n695,n1498);
and (n1514,n1476,n1483);
and (n1515,n1516,n1273);
xor (n1516,n1517,n1534);
xor (n1517,n1518,n1527);
nor (n1518,n1519,n1524);
and (n1519,n1520,n1457);
xor (n1520,n1521,n1523);
not (n1521,n1522);
wire s0n1522,s1n1522,notn1522;
or (n1522,s0n1522,s1n1522);
not(notn1522,n695);
and (s0n1522,notn1522,1'b0);
and (s1n1522,n695,n1445);
nand (n1523,n590,n1302);
and (n1524,n1525,n1526);
not (n1525,n1520);
not (n1526,n1457);
nand (n1527,n1528,n1530,n1532);
or (n1528,n1523,n1529);
not (n1529,n1327);
or (n1530,n1287,n1531);
not (n1531,n1313);
not (n1532,n1533);
and (n1533,n1301,n1313);
nand (n1534,n1535,n1588);
or (n1535,n1536,n1549);
not (n1536,n1537);
nand (n1537,n1538,n1540);
xor (n1538,n1300,n1539);
not (n1539,n1286);
not (n1540,n1541);
nand (n1541,n1542,n1546,n1548);
or (n1542,n1543,n1544);
not (n1543,n1360);
not (n1544,n1545);
not (n1545,n1523);
or (n1546,n1539,n1547);
not (n1547,n1332);
not (n1548,n1326);
not (n1549,n1550);
or (n1550,n1551,n1587);
and (n1551,n1552,n1562);
xor (n1552,n1553,n1559);
nand (n1553,n1554,n1556,n1558);
or (n1554,n1287,n1555);
not (n1555,n1377);
or (n1556,n1398,n1557);
not (n1557,n1348);
not (n1558,n1331);
nand (n1559,n1560,n1561);
or (n1560,n1398,n1400);
nand (n1561,n1400,n1398);
or (n1562,n1563,n1586);
and (n1563,n1564,n1573);
xor (n1564,n1565,n1571);
nand (n1565,n1566,n1568,n1570);
not (n1566,n1567);
and (n1567,n1404,n1364);
or (n1568,n1398,n1569);
not (n1569,n1392);
not (n1570,n1347);
xnor (n1571,n1572,n1407);
not (n1572,n1404);
or (n1573,n1574,n1585);
and (n1574,n1575,n1581);
xor (n1575,n1576,n1577);
nor (n1576,n1418,n1555);
xnor (n1577,n1578,n1557);
nand (n1578,n1579,n1580);
or (n1579,n1411,n1543);
nand (n1580,n1411,n1543);
nand (n1581,n1582,n1584);
or (n1582,n1583,n1365);
xnor (n1583,n1555,n1418);
not (n1584,n1379);
and (n1585,n1576,n1577);
and (n1586,n1565,n1571);
and (n1587,n1553,n1559);
or (n1588,n1538,n1540);
and (n1589,n1590,n1273);
xor (n1590,n1591,n1599);
xor (n1591,n1592,n1598);
nand (n1592,n1593,n1595);
or (n1593,n1594,n1526);
and (n1594,n1521,n1523);
or (n1595,n1596,n1597);
not (n1596,n1328);
not (n1597,n1444);
not (n1598,n1477);
or (n1599,n1600,n1601);
and (n1600,n1517,n1534);
and (n1601,n1518,n1527);
wire s0n1602,s1n1602,notn1602;
or (n1602,s0n1602,s1n1602);
not(notn1602,n1224);
and (s0n1602,notn1602,1'b0);
and (s1n1602,n1224,n1603);
xor (n1603,n1604,n1695);
xor (n1604,n1490,n1605);
xor (n1605,n1487,n1606);
or (n1606,n1607,n1608,n1694);
and (n1607,n1461,n1510);
and (n1608,n1510,n1609);
or (n1609,n1610,n1613,n1693);
and (n1610,n1611,n1612);
wire s0n1611,s1n1611,notn1611;
or (n1611,s0n1611,s1n1611);
not(notn1611,n647);
and (s0n1611,notn1611,1'b0);
and (s1n1611,n647,n1498);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n695);
and (s0n1612,notn1612,1'b0);
and (s1n1612,n695,n1462);
and (n1613,n1612,n1614);
or (n1614,n1615,n1628,n1692);
and (n1615,n1616,n1513);
wire s0n1616,s1n1616,notn1616;
or (n1616,s0n1616,s1n1616);
not(notn1616,n647);
and (s0n1616,notn1616,1'b0);
and (s1n1616,n647,n1617);
wire s0n1617,s1n1617,notn1617;
or (n1617,s0n1617,s1n1617);
not(notn1617,n571);
and (s0n1617,notn1617,n1618);
and (s1n1617,n571,n1620);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n18);
and (s0n1618,notn1618,1'b0);
and (s1n1618,n18,n1619);
or (n1620,1'b0,n1621,n1623,n1625,n1627);
and (n1621,n1622,n552);
and (n1623,n1624,n563);
and (n1625,n1626,n567);
and (n1627,n1619,n569);
and (n1628,n1513,n1629);
or (n1629,n1630,n1644,n1691);
and (n1630,n1631,n1643);
wire s0n1631,s1n1631,notn1631;
or (n1631,s0n1631,s1n1631);
not(notn1631,n647);
and (s0n1631,notn1631,1'b0);
and (s1n1631,n647,n1632);
wire s0n1632,s1n1632,notn1632;
or (n1632,s0n1632,s1n1632);
not(notn1632,n571);
and (s0n1632,notn1632,n1633);
and (s1n1632,n571,n1635);
wire s0n1633,s1n1633,notn1633;
or (n1633,s0n1633,s1n1633);
not(notn1633,n18);
and (s0n1633,notn1633,1'b0);
and (s1n1633,n18,n1634);
or (n1635,1'b0,n1636,n1638,n1640,n1642);
and (n1636,n1637,n552);
and (n1638,n1639,n563);
and (n1640,n1641,n567);
and (n1642,n1634,n569);
wire s0n1643,s1n1643,notn1643;
or (n1643,s0n1643,s1n1643);
not(notn1643,n695);
and (s0n1643,notn1643,1'b0);
and (s1n1643,n695,n1617);
and (n1644,n1643,n1645);
or (n1645,n1646,n1660,n1662);
and (n1646,n1647,n1659);
wire s0n1647,s1n1647,notn1647;
or (n1647,s0n1647,s1n1647);
not(notn1647,n647);
and (s0n1647,notn1647,1'b0);
and (s1n1647,n647,n1648);
wire s0n1648,s1n1648,notn1648;
or (n1648,s0n1648,s1n1648);
not(notn1648,n571);
and (s0n1648,notn1648,n1649);
and (s1n1648,n571,n1651);
wire s0n1649,s1n1649,notn1649;
or (n1649,s0n1649,s1n1649);
not(notn1649,n18);
and (s0n1649,notn1649,1'b0);
and (s1n1649,n18,n1650);
or (n1651,1'b0,n1652,n1654,n1656,n1658);
and (n1652,n1653,n552);
and (n1654,n1655,n563);
and (n1656,n1657,n567);
and (n1658,n1650,n569);
wire s0n1659,s1n1659,notn1659;
or (n1659,s0n1659,s1n1659);
not(notn1659,n695);
and (s0n1659,notn1659,1'b0);
and (s1n1659,n695,n1632);
and (n1660,n1659,n1661);
or (n1661,n1662,n1676,n1677);
and (n1662,n1663,n1675);
wire s0n1663,s1n1663,notn1663;
or (n1663,s0n1663,s1n1663);
not(notn1663,n647);
and (s0n1663,notn1663,1'b0);
and (s1n1663,n647,n1664);
wire s0n1664,s1n1664,notn1664;
or (n1664,s0n1664,s1n1664);
not(notn1664,n571);
and (s0n1664,notn1664,n1665);
and (s1n1664,n571,n1667);
wire s0n1665,s1n1665,notn1665;
or (n1665,s0n1665,s1n1665);
not(notn1665,n18);
and (s0n1665,notn1665,1'b0);
and (s1n1665,n18,n1666);
or (n1667,1'b0,n1668,n1670,n1672,n1674);
and (n1668,n1669,n552);
and (n1670,n1671,n563);
and (n1672,n1673,n567);
and (n1674,n1666,n569);
wire s0n1675,s1n1675,notn1675;
or (n1675,s0n1675,s1n1675);
not(notn1675,n695);
and (s0n1675,notn1675,1'b0);
and (s1n1675,n695,n1648);
and (n1676,n1675,n1677);
and (n1677,n1678,n1690);
wire s0n1678,s1n1678,notn1678;
or (n1678,s0n1678,s1n1678);
not(notn1678,n647);
and (s0n1678,notn1678,1'b0);
and (s1n1678,n647,n1679);
wire s0n1679,s1n1679,notn1679;
or (n1679,s0n1679,s1n1679);
not(notn1679,n571);
and (s0n1679,notn1679,n1680);
and (s1n1679,n571,n1682);
wire s0n1680,s1n1680,notn1680;
or (n1680,s0n1680,s1n1680);
not(notn1680,n18);
and (s0n1680,notn1680,1'b0);
and (s1n1680,n18,n1681);
or (n1682,1'b0,n1683,n1685,n1687,n1689);
and (n1683,n1684,n552);
and (n1685,n1686,n563);
and (n1687,n1688,n567);
and (n1689,n1681,n569);
wire s0n1690,s1n1690,notn1690;
or (n1690,s0n1690,s1n1690);
not(notn1690,n695);
and (s0n1690,notn1690,1'b0);
and (s1n1690,n695,n1664);
and (n1691,n1631,n1645);
and (n1692,n1616,n1629);
and (n1693,n1611,n1614);
and (n1694,n1461,n1609);
or (n1695,n1696,n1699,n1732);
and (n1696,n1497,n1697);
xor (n1697,n1698,n1609);
xor (n1698,n1461,n1510);
and (n1699,n1697,n1700);
or (n1700,n1701,n1705,n1731);
and (n1701,n1702,n1703);
wire s0n1702,s1n1702,notn1702;
or (n1702,s0n1702,s1n1702);
not(notn1702,n590);
and (s0n1702,notn1702,1'b0);
and (s1n1702,n590,n1617);
xor (n1703,n1704,n1614);
xor (n1704,n1611,n1612);
and (n1705,n1703,n1706);
or (n1706,n1707,n1711,n1730);
and (n1707,n1708,n1709);
wire s0n1708,s1n1708,notn1708;
or (n1708,s0n1708,s1n1708);
not(notn1708,n590);
and (s0n1708,notn1708,1'b0);
and (s1n1708,n590,n1632);
xor (n1709,n1710,n1629);
xor (n1710,n1616,n1513);
and (n1711,n1709,n1712);
or (n1712,n1713,n1717,n1729);
and (n1713,n1714,n1715);
wire s0n1714,s1n1714,notn1714;
or (n1714,s0n1714,s1n1714);
not(notn1714,n590);
and (s0n1714,notn1714,1'b0);
and (s1n1714,n590,n1648);
xor (n1715,n1716,n1645);
xor (n1716,n1631,n1643);
and (n1717,n1715,n1718);
or (n1718,n1719,n1723,n1728);
and (n1719,n1720,n1721);
wire s0n1720,s1n1720,notn1720;
or (n1720,s0n1720,s1n1720);
not(notn1720,n590);
and (s0n1720,notn1720,1'b0);
and (s1n1720,n590,n1664);
xor (n1721,n1722,n1661);
xor (n1722,n1647,n1659);
and (n1723,n1721,n1724);
and (n1724,n1725,n1726);
wire s0n1725,s1n1725,notn1725;
or (n1725,s0n1725,s1n1725);
not(notn1725,n590);
and (s0n1725,notn1725,1'b0);
and (s1n1725,n590,n1679);
xor (n1726,n1727,n1677);
xor (n1727,n1663,n1675);
and (n1728,n1720,n1724);
and (n1729,n1714,n1718);
and (n1730,n1708,n1712);
and (n1731,n1702,n1706);
and (n1732,n1497,n1700);
and (n1733,n1281,n1589);
xor (n1734,n1735,n1765);
xor (n1735,n1736,n1764);
wire s0n1736,s1n1736,notn1736;
or (n1736,s0n1736,s1n1736);
not(notn1736,n931);
and (s0n1736,notn1736,1'b0);
and (s1n1736,n931,n1737);
or (n1737,n1738,n1747,n1763);
and (n1738,n1444,n1739);
and (n1739,n1482,n1740);
or (n1740,n1741,n1742,n1746);
and (n1741,n1457,n1522);
and (n1742,n1522,n1743);
or (n1743,n1533,n1744,n1745);
and (n1744,n1313,n1325);
and (n1745,n1301,n1325);
and (n1746,n1457,n1743);
and (n1747,n1739,n1748);
or (n1748,n1749,n1751,n1762);
and (n1749,n1479,n1750);
xor (n1750,n1482,n1740);
and (n1751,n1750,n1752);
or (n1752,n1753,n1756,n1761);
and (n1753,n1545,n1754);
xor (n1754,n1755,n1743);
xor (n1755,n1457,n1522);
and (n1756,n1754,n1757);
or (n1757,n1758,n1759,n1760);
and (n1758,n1286,n1299);
and (n1759,n1299,n1395);
and (n1760,n1286,n1395);
and (n1761,n1545,n1757);
and (n1762,n1479,n1752);
and (n1763,n1444,n1748);
and (n1764,n1590,n1424);
wire s0n1765,s1n1765,notn1765;
or (n1765,s0n1765,s1n1765);
not(notn1765,n1273);
and (s0n1765,notn1765,1'b0);
and (s1n1765,n1273,n1766);
xor (n1766,n1767,n1748);
xor (n1767,n1444,n1739);
wire s0n1768,s1n1768,notn1768;
or (n1768,s0n1768,s1n1768);
not(notn1768,n933);
and (s0n1768,notn1768,1'b0);
and (s1n1768,n933,n1769);
or (n1769,n1770,n1772,n1777);
and (n1770,n1431,n1771);
and (n1771,n1487,n1606);
and (n1772,n1771,n1773);
or (n1773,n1774,n1775,n1776);
and (n1774,n1490,n1605);
and (n1775,n1605,n1695);
and (n1776,n1490,n1695);
and (n1777,n1431,n1773);
or (n1778,n1779,n1900);
and (n1779,n1780,n1794);
xor (n1780,n1781,n1793);
or (n1781,n1782,n1792);
and (n1782,n1783,n1788);
xor (n1783,n1784,n1786);
and (n1784,n1785,n1224);
xor (n1785,n1106,n1130);
and (n1786,n1787,n933);
xor (n1787,n1080,n1104);
and (n1788,n1789,n1273);
xor (n1789,n1790,n787);
nor (n1790,n1791,n924);
not (n1791,n913);
and (n1792,n1784,n1786);
xor (n1793,n1280,n1602);
and (n1794,n1795,n1847);
xor (n1795,n1796,n1799);
and (n1796,n1797,n1424);
xnor (n1797,n847,n1798);
nand (n1798,n790,n912);
or (n1799,n1800,n1846);
and (n1800,n1801,n1826);
xor (n1801,n1802,n1805);
wire s0n1802,s1n1802,notn1802;
or (n1802,s0n1802,s1n1802);
not(notn1802,n1224);
and (s0n1802,notn1802,1'b0);
and (s1n1802,n1224,n1803);
xor (n1803,n1804,n1706);
xor (n1804,n1702,n1703);
and (n1805,n1806,n1820);
or (n1806,n1807,n1819);
and (n1807,n1808,n1818);
xor (n1808,n1809,n1817);
and (n1809,n1810,n981);
nand (n1810,n1811,n1813,n1816);
or (n1811,n1812,n1496);
not (n1812,n1659);
or (n1813,n1814,n1815);
not (n1814,n1702);
not (n1815,n1631);
not (n1816,n1615);
and (n1817,n1541,n981);
nor (n1818,n1538,n980);
and (n1819,n1809,n1817);
and (n1820,n1821,n981);
nor (n1821,n1822,n1824);
and (n1822,n1823,n1459);
xor (n1823,n1496,n1509);
and (n1824,n1825,n1460);
not (n1825,n1823);
or (n1826,n1827,n1845);
and (n1827,n1828,n1842);
xor (n1828,n1829,n1831);
and (n1829,n1830,n1273);
xor (n1830,n1552,n1562);
xor (n1831,n1832,n1841);
xor (n1832,n1833,n1834);
and (n1833,n1527,n981);
and (n1834,n1835,n981);
nand (n1835,n1836,n1840);
or (n1836,n1837,n1814);
and (n1837,n1838,n1839);
not (n1838,n1611);
not (n1839,n1612);
not (n1840,n1610);
and (n1841,n1518,n981);
wire s0n1842,s1n1842,notn1842;
or (n1842,s0n1842,s1n1842);
not(notn1842,n1224);
and (s0n1842,notn1842,1'b0);
and (s1n1842,n1224,n1843);
xor (n1843,n1844,n1712);
xor (n1844,n1708,n1709);
and (n1845,n1829,n1831);
and (n1846,n1802,n1805);
wire s0n1847,s1n1847,notn1847;
or (n1847,s0n1847,s1n1847);
not(notn1847,n931);
and (s0n1847,notn1847,1'b0);
and (s1n1847,n931,n1848);
xor (n1848,n1849,n1868);
xor (n1849,n1850,n1851);
xor (n1850,n767,n763);
xor (n1851,n765,n1852);
or (n1852,n779,n1853,n1867);
and (n1853,n781,n1854);
or (n1854,n920,n1855,n1866);
and (n1855,n808,n1856);
or (n1856,n821,n1857,n1865);
and (n1857,n823,n1858);
or (n1858,n842,n1859,n1864);
and (n1859,n844,n1860);
or (n1860,n855,n1861,n876);
and (n1861,n857,n1862);
or (n1862,n876,n1863,n882);
and (n1863,n878,n882);
and (n1864,n843,n1860);
and (n1865,n822,n1858);
and (n1866,n807,n1856);
and (n1867,n780,n1854);
or (n1868,n1869,n1872,n1899);
and (n1869,n1870,n1871);
xor (n1870,n919,n916);
xor (n1871,n918,n1854);
and (n1872,n1871,n1873);
or (n1873,n1874,n1877,n1898);
and (n1874,n1875,n1876);
xor (n1875,n809,n793);
xor (n1876,n806,n1856);
and (n1877,n1876,n1878);
or (n1878,n1879,n1882,n1897);
and (n1879,n1880,n1881);
xor (n1880,n830,n827);
xor (n1881,n829,n1858);
and (n1882,n1881,n1883);
or (n1883,n1884,n1887,n1896);
and (n1884,n1885,n1886);
xor (n1885,n860,n854);
xor (n1886,n859,n1860);
and (n1887,n1886,n1888);
or (n1888,n1889,n1892,n1895);
and (n1889,n1890,n1891);
xor (n1890,n901,n903);
xor (n1891,n902,n1862);
and (n1892,n1891,n1893);
and (n1893,n896,n1894);
xor (n1894,n897,n882);
and (n1895,n1890,n1893);
and (n1896,n1885,n1888);
and (n1897,n1880,n1883);
and (n1898,n1875,n1878);
and (n1899,n1870,n1873);
and (n1900,n1781,n1793);
xor (n1901,n1902,n1933);
xor (n1902,n1903,n1916);
xor (n1903,n1904,n1913);
xor (n1904,n1905,n1906);
wire s0n1905,s1n1905,notn1905;
or (n1905,s0n1905,s1n1905);
not(notn1905,n1424);
and (s0n1905,notn1905,1'b0);
and (s1n1905,n1424,n1848);
and (n1906,n1907,n1910);
or (n1907,n1908,n1909);
and (n1908,n1426,n1473);
and (n1909,n1427,n1458);
or (n1910,n1911,n1912);
and (n1911,n1428,n1456);
and (n1912,n1429,n1443);
wire s0n1913,s1n1913,notn1913;
or (n1913,s0n1913,s1n1913);
not(notn1913,n1224);
and (s0n1913,notn1913,1'b0);
and (s1n1913,n1224,n1914);
xor (n1914,n1915,n1773);
xor (n1915,n1431,n1771);
or (n1916,n1917,n1932);
and (n1917,n1918,n1931);
xor (n1918,n1919,n1930);
or (n1919,n1920,n1929);
and (n1920,n1921,n1928);
xor (n1921,n1922,n1923);
xor (n1922,n1282,n1515);
and (n1923,n1924,n1927);
xor (n1924,n1925,n1926);
and (n1925,n1830,n1424);
wire s0n1926,s1n1926,notn1926;
or (n1926,s0n1926,s1n1926);
not(notn1926,n1273);
and (s0n1926,notn1926,1'b0);
and (s1n1926,n1273,n1284);
and (n1927,n1516,n931);
wire s0n1928,s1n1928,notn1928;
or (n1928,s0n1928,s1n1928);
not(notn1928,n933);
and (s0n1928,notn1928,1'b0);
and (s1n1928,n933,n1603);
and (n1929,n1922,n1923);
and (n1930,n1787,n1224);
wire s0n1931,s1n1931,notn1931;
or (n1931,s0n1931,s1n1931);
not(notn1931,n1273);
and (s0n1931,notn1931,1'b0);
and (s1n1931,n1273,n1848);
and (n1932,n1919,n1930);
or (n1933,n1934,n1944);
and (n1934,n1935,n1943);
xor (n1935,n1936,n1937);
wire s0n1936,s1n1936,notn1936;
or (n1936,s0n1936,s1n1936);
not(notn1936,n981);
and (s0n1936,notn1936,1'b0);
and (s1n1936,n981,n13);
and (n1937,n1938,n981);
xnor (n1938,n1939,n1941);
not (n1939,n1940);
and (n1940,n588,n1033);
or (n1941,n1942,n1077);
and (n1942,n1030,n1078);
and (n1943,n1272,n931);
and (n1944,n1936,n1937);
or (n1945,n1946,n2119);
and (n1946,n1947,n1986);
xor (n1947,n1948,n1949);
xor (n1948,n1780,n1794);
or (n1949,n1950,n1985);
and (n1950,n1951,n1960);
xor (n1951,n1952,n1959);
or (n1952,n1953,n1958);
and (n1953,n1954,n1957);
xor (n1954,n1955,n1956);
and (n1955,n1797,n1273);
xor (n1956,n1801,n1826);
and (n1957,n1787,n981);
and (n1958,n1955,n1956);
xor (n1959,n1795,n1847);
or (n1960,n1961,n1984);
and (n1961,n1962,n1983);
xor (n1962,n1963,n1964);
and (n1963,n1785,n933);
or (n1964,n1965,n1982);
and (n1965,n1966,n1979);
xor (n1966,n1967,n1971);
xor (n1967,n1968,n1969);
xor (n1968,n1806,n1820);
and (n1969,n1970,n1424);
xor (n1970,n1564,n1573);
and (n1971,n1972,n1976);
xor (n1972,n1973,n1974);
xor (n1973,n1808,n1818);
and (n1974,n1975,n1424);
xor (n1975,n1575,n1581);
wire s0n1976,s1n1976,notn1976;
or (n1976,s0n1976,s1n1976);
not(notn1976,n1224);
and (s0n1976,notn1976,1'b0);
and (s1n1976,n1224,n1977);
xor (n1977,n1978,n1718);
xor (n1978,n1714,n1715);
wire s0n1979,s1n1979,notn1979;
or (n1979,s0n1979,s1n1979);
not(notn1979,n1424);
and (s0n1979,notn1979,1'b0);
and (s1n1979,n1424,n1980);
xor (n1980,n1981,n1888);
xor (n1981,n1885,n1886);
and (n1982,n1967,n1971);
and (n1983,n1789,n931);
and (n1984,n1963,n1964);
and (n1985,n1952,n1959);
or (n1986,n1987,n2118);
and (n1987,n1988,n2099);
xor (n1988,n1989,n2098);
or (n1989,n1990,n2097);
and (n1990,n1991,n2096);
xor (n1991,n1992,n2067);
or (n1992,n1993,n2066);
and (n1993,n1994,n2063);
xor (n1994,n1995,n2018);
xor (n1995,n1996,n2017);
xor (n1996,n1997,n1998);
wire s0n1997,s1n1997,notn1997;
or (n1997,s0n1997,s1n1997);
not(notn1997,n931);
and (s0n1997,notn1997,1'b0);
and (s1n1997,n931,n1284);
or (n1998,n1999,n2016);
and (n1999,n2000,n2015);
xor (n2000,n2001,n2013);
or (n2001,n2002,n2003);
and (n2002,n1553,n981);
and (n2003,n2004,n981);
nand (n2004,n2005,n2006);
not (n2005,n1630);
nand (n2006,n2007,n2011);
or (n2007,n2008,n2009);
not (n2008,n1815);
not (n2009,n2010);
not (n2010,n1643);
not (n2011,n2012);
not (n2012,n1714);
nor (n2013,n980,n2014);
xor (n2014,n1704,n1814);
and (n2015,n1970,n1273);
and (n2016,n2001,n2013);
wire s0n2017,s1n2017,notn2017;
or (n2017,s0n2017,s1n2017);
not(notn2017,n933);
and (s0n2017,notn2017,1'b0);
and (s1n2017,n933,n1803);
and (n2018,n2019,n2062);
xor (n2019,n2020,n2056);
or (n2020,n2021,n2055);
and (n2021,n2022,n2052);
xor (n2022,n2023,n2037);
and (n2023,n2024,n2029);
xor (n2024,n2025,n2027);
and (n2025,n2026,n981);
xnor (n2026,n2012,n1716);
and (n2027,n1424,n2028);
xor (n2028,n1380,n1392);
and (n2029,n2030,n2033);
and (n2030,n2031,n2011);
wire s0n2031,s1n2031,notn2031;
or (n2031,s0n2031,s1n2031);
not(notn2031,n981);
and (s0n2031,notn2031,1'b0);
and (s1n2031,n981,n2032);
wire s0n2032,s1n2032,notn2032;
or (n2032,s0n2032,s1n2032);
not(notn2032,n695);
and (s0n2032,notn2032,1'b0);
and (s1n2032,n695,n1679);
nor (n2033,n2034,n1572);
not (n2034,n2035);
wire s0n2035,s1n2035,notn2035;
or (n2035,s0n2035,s1n2035);
not(notn2035,n981);
and (s0n2035,notn2035,1'b0);
and (s1n2035,n981,n2036);
wire s0n2036,s1n2036,notn2036;
or (n2036,s0n2036,s1n2036);
not(notn2036,n695);
and (s0n2036,notn2036,1'b0);
and (s1n2036,n695,n1381);
or (n2037,n2038,n2051);
and (n2038,n2039,n2050);
xor (n2039,n2040,n2049);
and (n2040,n2041,n981);
not (n2041,n2042);
nor (n2042,n2043,n2044);
and (n2043,n2011,n1663);
and (n2044,n2045,n2048);
nand (n2045,n2046,n2047);
not (n2046,n1720);
not (n2047,n1647);
not (n2048,n1812);
and (n2049,n1565,n981);
and (n2050,n1571,n981);
and (n2051,n2040,n2049);
wire s0n2052,s1n2052,notn2052;
or (n2052,s0n2052,s1n2052);
not(notn2052,n1224);
and (s0n2052,notn2052,1'b0);
and (s1n2052,n1224,n2053);
xor (n2053,n2054,n1724);
xor (n2054,n1720,n1721);
and (n2055,n2023,n2037);
and (n2056,n2057,n2061);
xor (n2057,n2058,n2059);
wire s0n2058,s1n2058,notn2058;
or (n2058,s0n2058,s1n2058);
not(notn2058,n933);
and (s0n2058,notn2058,1'b0);
and (s1n2058,n933,n1977);
wire s0n2059,s1n2059,notn2059;
or (n2059,s0n2059,s1n2059);
not(notn2059,n1424);
and (s0n2059,notn2059,1'b0);
and (s1n2059,n1424,n2060);
xor (n2060,n1417,n1419);
and (n2061,n1970,n931);
xor (n2062,n1972,n1976);
wire s0n2063,s1n2063,notn2063;
or (n2063,s0n2063,s1n2063);
not(notn2063,n1273);
and (s0n2063,notn2063,1'b0);
and (s1n2063,n1273,n2064);
xor (n2064,n2065,n1883);
xor (n2065,n1880,n1881);
and (n2066,n1995,n2018);
or (n2067,n2068,n2095);
and (n2068,n2069,n2093);
xor (n2069,n2070,n2071);
xor (n2070,n1828,n1842);
or (n2071,n2072,n2092);
and (n2072,n2073,n2091);
xor (n2073,n2074,n2075);
and (n2074,n1830,n931);
or (n2075,n2076,n2090);
and (n2076,n2077,n2089);
xor (n2077,n2078,n2088);
and (n2078,n2079,n981);
not (n2079,n2080);
nor (n2080,n2081,n2087);
and (n2081,n2082,n2085);
not (n2082,n2083);
xor (n2083,n1512,n2084);
not (n2084,n1708);
not (n2085,n2086);
not (n2086,n1616);
and (n2087,n2083,n2086);
and (n2088,n1559,n981);
and (n2089,n1975,n1273);
and (n2090,n2078,n2088);
wire s0n2091,s1n2091,notn2091;
or (n2091,s0n2091,s1n2091);
not(notn2091,n933);
and (s0n2091,notn2091,1'b0);
and (s1n2091,n933,n1843);
and (n2092,n2074,n2075);
and (n2093,n2094,n1224);
xor (n2094,n1158,n1182);
and (n2095,n2070,n2071);
wire s0n2096,s1n2096,notn2096;
or (n2096,s0n2096,s1n2096);
not(notn2096,n981);
and (s0n2096,notn2096,1'b0);
and (s1n2096,n981,n1848);
and (n2097,n1992,n2067);
xor (n2098,n1783,n1788);
xor (n2099,n2100,n2117);
xor (n2100,n2101,n2102);
and (n2101,n1029,n981);
xor (n2102,n2103,n2114);
xor (n2103,n2104,n2105);
and (n2104,n1590,n931);
or (n2105,n2106,n2113);
and (n2106,n2107,n2110);
xor (n2107,n2108,n2109);
xor (n2108,n1475,n1492);
and (n2109,n1592,n981);
or (n2110,n2111,n2112);
and (n2111,n1832,n1841);
and (n2112,n1833,n1834);
and (n2113,n2108,n2109);
wire s0n2114,s1n2114,notn2114;
or (n2114,s0n2114,s1n2114);
not(notn2114,n1224);
and (s0n2114,notn2114,1'b0);
and (s1n2114,n1224,n2115);
xor (n2115,n2116,n1700);
xor (n2116,n1497,n1697);
and (n2117,n1272,n981);
and (n2118,n1989,n2098);
and (n2119,n1948,n1949);
and (n2120,n7,n1901);
xor (n2121,n2122,n2149);
xor (n2122,n2123,n2130);
xor (n2123,n2124,n2127);
xor (n2124,n2125,n2126);
and (n2125,n1904,n1913);
and (n2126,n1735,n1765);
or (n2127,n2128,n2129);
and (n2128,n10,n1271);
and (n2129,n11,n1028);
and (n2130,n2131,n2142);
xor (n2131,n2132,n2141);
or (n2132,n2133,n2140);
and (n2133,n2134,n2139);
xor (n2134,n2135,n2136);
wire s0n2135,s1n2135,notn2135;
or (n2135,s0n2135,s1n2135);
not(notn2135,n931);
and (s0n2135,notn2135,1'b0);
and (s1n2135,n931,n1766);
xor (n2136,n2137,n2138);
xor (n2137,n1907,n1910);
and (n2138,n1516,n1424);
and (n2139,n1029,n933);
and (n2140,n2135,n2136);
and (n2141,n1938,n933);
and (n2142,n2143,n2148);
xor (n2143,n2144,n2145);
and (n2144,n1789,n1424);
or (n2145,n2146,n2147);
and (n2146,n2103,n2114);
and (n2147,n2104,n2105);
wire s0n2148,s1n2148,notn2148;
or (n2148,s0n2148,s1n2148);
not(notn2148,n933);
and (s0n2148,notn2148,1'b0);
and (s1n2148,n933,n1914);
or (n2149,n2150,n2151);
and (n2150,n1902,n1933);
and (n2151,n1903,n1916);
xor (n2152,n2153,n2172);
xor (n2153,n2154,n2157);
or (n2154,n2155,n2156);
and (n2155,n8,n1778);
and (n2156,n9,n1276);
xor (n2157,n2158,n2167);
xor (n2158,n2159,n2162);
or (n2159,n2160,n2161);
and (n2160,n1277,n1768);
and (n2161,n1278,n1734);
xor (n2162,n2163,n2166);
xor (n2163,n2164,n2165);
wire s0n2164,s1n2164,notn2164;
or (n2164,s0n2164,s1n2164);
not(notn2164,n1424);
and (s0n2164,notn2164,1'b0);
and (s1n2164,n1424,n1766);
wire s0n2165,s1n2165,notn2165;
or (n2165,s0n2165,s1n2165);
not(notn2165,n1273);
and (s0n2165,notn2165,1'b0);
and (s1n2165,n1273,n1737);
and (n2166,n1272,n1424);
xor (n2167,n2168,n2171);
xor (n2168,n2169,n2170);
and (n2169,n1938,n1224);
wire s0n2170,s1n2170,notn2170;
or (n2170,s0n2170,s1n2170);
not(notn2170,n1224);
and (s0n2170,notn2170,1'b0);
and (s1n2170,n1224,n1769);
wire s0n2171,s1n2171,notn2171;
or (n2171,s0n2171,s1n2171);
not(notn2171,n1273);
and (s0n2171,notn2171,1'b0);
and (s1n2171,n1273,n13);
or (n2172,n2173,n2213);
and (n2173,n2174,n2185);
xor (n2174,n2175,n2184);
or (n2175,n2176,n2183);
and (n2176,n2177,n2182);
xor (n2177,n2178,n2181);
or (n2178,n2179,n2180);
and (n2179,n2100,n2117);
and (n2180,n2101,n2102);
xor (n2181,n2134,n2139);
xor (n2182,n1918,n1931);
and (n2183,n2178,n2181);
xor (n2184,n2131,n2142);
or (n2185,n2186,n2212);
and (n2186,n2187,n2211);
xor (n2187,n2188,n2189);
xor (n2188,n2143,n2148);
or (n2189,n2190,n2210);
and (n2190,n2191,n2202);
xor (n2191,n2192,n2193);
xor (n2192,n1921,n1928);
or (n2193,n2194,n2201);
and (n2194,n2195,n2200);
xor (n2195,n2196,n2199);
or (n2196,n2197,n2198);
and (n2197,n1996,n2017);
and (n2198,n1997,n1998);
xor (n2199,n2107,n2110);
wire s0n2200,s1n2200,notn2200;
or (n2200,s0n2200,s1n2200);
not(notn2200,n933);
and (s0n2200,notn2200,1'b0);
and (s1n2200,n933,n2115);
and (n2201,n2196,n2199);
or (n2202,n2203,n2209);
and (n2203,n2204,n2207);
xor (n2204,n2205,n2206);
wire s0n2205,s1n2205,notn2205;
or (n2205,s0n2205,s1n2205);
not(notn2205,n1424);
and (s0n2205,notn2205,1'b0);
and (s1n2205,n1424,n2064);
xor (n2206,n1924,n1927);
and (n2207,n2208,n1224);
xor (n2208,n1132,n1156);
and (n2209,n2205,n2206);
and (n2210,n2192,n2193);
xor (n2211,n1935,n1943);
and (n2212,n2188,n2189);
and (n2213,n2175,n2184);
and (n2214,n4,n2121);
nand (n2215,n2216,n2220);
not (n2216,n2217);
or (n2217,n2218,n2219);
and (n2218,n2153,n2172);
and (n2219,n2154,n2157);
nor (n2220,n2221,n2236);
not (n2221,n2222);
nor (n2222,n2223,n2233);
not (n2223,n2224);
nor (n2224,n2225,n2226);
and (n2225,n2168,n2171);
not (n2226,n2227);
nor (n2227,n2228,n2229);
and (n2228,n2163,n2166);
not (n2229,n2230);
xnor (n2230,n2231,n2232);
wire s0n2231,s1n2231,notn2231;
or (n2231,s0n2231,s1n2231);
not(notn2231,n1424);
and (s0n2231,notn2231,1'b0);
and (s1n2231,n1424,n13);
wire s0n2232,s1n2232,notn2232;
or (n2232,s0n2232,s1n2232);
not(notn2232,n1424);
and (s0n2232,notn2232,1'b0);
and (s1n2232,n1424,n1737);
or (n2233,n2234,n2235);
and (n2234,n2158,n2167);
and (n2235,n2159,n2162);
and (n2236,n2122,n2149);
or (n2237,n2238,n2770);
or (n2238,n2239,n2769);
and (n2239,n2240,n2313);
xor (n2240,n2241,n2242);
xor (n2241,n3,n2152);
or (n2242,n2243,n2312);
and (n2243,n2244,n2311);
xor (n2244,n2245,n2310);
or (n2245,n2246,n2309);
and (n2246,n2247,n2250);
xor (n2247,n2248,n2249);
xor (n2248,n2187,n2211);
xor (n2249,n2177,n2182);
or (n2250,n2251,n2308);
and (n2251,n2252,n2295);
xor (n2252,n2253,n2294);
or (n2253,n2254,n2293);
and (n2254,n2255,n2258);
xor (n2255,n2256,n2257);
xor (n2256,n2204,n2207);
xor (n2257,n2195,n2200);
or (n2258,n2259,n2292);
and (n2259,n2260,n2291);
xor (n2260,n2261,n2268);
and (n2261,n2262,n2266);
xor (n2262,n2263,n2265);
and (n2263,n2264,n1424);
xor (n2264,n875,n899);
xor (n2265,n2000,n2015);
and (n2266,n2267,n1224);
xor (n2267,n1184,n1202);
or (n2268,n2269,n2290);
and (n2269,n2270,n2289);
xor (n2270,n2271,n2272);
xor (n2271,n2073,n2091);
or (n2272,n2273,n2288);
and (n2273,n2274,n2280);
xor (n2274,n2275,n2276);
xor (n2275,n2077,n2089);
nand (n2276,n2277,n2001);
or (n2277,n2278,n2279);
not (n2278,n2003);
not (n2279,n2002);
or (n2280,n2281,n2287);
and (n2281,n2282,n2286);
xor (n2282,n2283,n2284);
wire s0n2283,s1n2283,notn2283;
or (n2283,s0n2283,s1n2283);
not(notn2283,n1273);
and (s0n2283,notn2283,1'b0);
and (s1n2283,n1273,n2060);
wire s0n2284,s1n2284,notn2284;
or (n2284,s0n2284,s1n2284);
not(notn2284,n1224);
and (s0n2284,notn2284,1'b0);
and (s1n2284,n1224,n2285);
xor (n2285,n1725,n1726);
and (n2286,n1975,n931);
and (n2287,n2283,n2284);
and (n2288,n2275,n2276);
wire s0n2289,s1n2289,notn2289;
or (n2289,s0n2289,s1n2289);
not(notn2289,n1273);
and (s0n2289,notn2289,1'b0);
and (s1n2289,n1273,n1980);
and (n2290,n2271,n2272);
and (n2291,n1785,n981);
and (n2292,n2261,n2268);
and (n2293,n2256,n2257);
xor (n2294,n2191,n2202);
or (n2295,n2296,n2307);
and (n2296,n2297,n2306);
xor (n2297,n2298,n2299);
xor (n2298,n1954,n1957);
or (n2299,n2300,n2305);
and (n2300,n2301,n2304);
xor (n2301,n2302,n2303);
and (n2302,n1797,n931);
and (n2303,n2208,n933);
and (n2304,n1789,n981);
and (n2305,n2302,n2303);
xor (n2306,n1962,n1983);
and (n2307,n2298,n2299);
and (n2308,n2253,n2294);
and (n2309,n2248,n2249);
xor (n2310,n2174,n2185);
xor (n2311,n6,n1945);
and (n2312,n2245,n2310);
or (n2313,n2314,n2768);
and (n2314,n2315,n2400);
xor (n2315,n2316,n2317);
xor (n2316,n2244,n2311);
or (n2317,n2318,n2399);
and (n2318,n2319,n2398);
xor (n2319,n2320,n2397);
or (n2320,n2321,n2396);
and (n2321,n2322,n2395);
xor (n2322,n2323,n2324);
xor (n2323,n1951,n1960);
or (n2324,n2325,n2394);
and (n2325,n2326,n2363);
xor (n2326,n2327,n2328);
xor (n2327,n1991,n2096);
or (n2328,n2329,n2362);
and (n2329,n2330,n2333);
xor (n2330,n2331,n2332);
xor (n2331,n1966,n1979);
xor (n2332,n2069,n2093);
or (n2333,n2334,n2361);
and (n2334,n2335,n2360);
xor (n2335,n2336,n2359);
and (n2336,n2337,n2358);
and (n2337,n2338,n2345);
or (n2338,n2339,n2344);
and (n2339,n2340,n2343);
xor (n2340,n2341,n2342);
and (n2341,n1273,n2028);
xor (n2342,n2030,n2033);
wire s0n2343,s1n2343,notn2343;
or (n2343,s0n2343,s1n2343);
not(notn2343,n933);
and (s0n2343,notn2343,1'b0);
and (s1n2343,n933,n2285);
and (n2344,n2341,n2342);
and (n2345,n2346,n2357);
xor (n2346,n2347,n2355);
and (n2347,n2348,n981);
nand (n2348,n2349,n2354);
or (n2349,n2047,n2350);
nand (n2350,n2351,n2353);
or (n2351,n2352,n1812);
not (n2352,n2046);
nand (n2353,n2352,n1812);
nand (n2354,n2350,n2047);
wire s0n2355,s1n2355,notn2355;
or (n2355,s0n2355,s1n2355);
not(notn2355,n1424);
and (s0n2355,notn2355,1'b0);
and (s1n2355,n1424,n2356);
wire s0n2356,s1n2356,notn2356;
or (n2356,s0n2356,s1n2356);
not(notn2356,n695);
and (s0n2356,notn2356,1'b0);
and (s1n2356,n695,n884);
and (n2357,n1577,n981);
xor (n2358,n2022,n2052);
wire s0n2359,s1n2359,notn2359;
or (n2359,s0n2359,s1n2359);
not(notn2359,n931);
and (s0n2359,notn2359,1'b0);
and (s1n2359,n931,n2064);
and (n2360,n2094,n933);
and (n2361,n2336,n2359);
and (n2362,n2331,n2332);
or (n2363,n2364,n2393);
and (n2364,n2365,n2392);
xor (n2365,n2366,n2391);
or (n2366,n2367,n2390);
and (n2367,n2368,n2389);
xor (n2368,n2369,n2388);
or (n2369,n2370,n2387);
and (n2370,n2371,n2386);
xor (n2371,n2372,n2373);
xor (n2372,n2057,n2061);
or (n2373,n2374,n2385);
and (n2374,n2375,n2384);
xor (n2375,n2376,n2377);
xor (n2376,n2039,n2050);
and (n2377,n2378,n2380);
wire s0n2378,s1n2378,notn2378;
or (n2378,s0n2378,s1n2378);
not(notn2378,n1224);
and (s0n2378,notn2378,1'b0);
and (s1n2378,n1224,n2379);
xor (n2379,n1678,n1690);
and (n2380,n2381,n2382);
wire s0n2381,s1n2381,notn2381;
or (n2381,s0n2381,s1n2381);
not(notn2381,n1224);
and (s0n2381,notn2381,1'b0);
and (s1n2381,n1224,n2032);
wire s0n2382,s1n2382,notn2382;
or (n2382,s0n2382,s1n2382);
not(notn2382,n1224);
and (s0n2382,notn2382,1'b0);
and (s1n2382,n1224,n2383);
wire s0n2383,s1n2383,notn2383;
or (n2383,s0n2383,s1n2383);
not(notn2383,n695);
and (s0n2383,notn2383,1'b0);
and (s1n2383,n695,n1188);
wire s0n2384,s1n2384,notn2384;
or (n2384,s0n2384,s1n2384);
not(notn2384,n933);
and (s0n2384,notn2384,1'b0);
and (s1n2384,n933,n2053);
and (n2385,n2376,n2377);
and (n2386,n2264,n1273);
and (n2387,n2372,n2373);
xor (n2388,n2019,n2062);
and (n2389,n1797,n981);
and (n2390,n2369,n2388);
xor (n2391,n1994,n2063);
xor (n2392,n2301,n2304);
and (n2393,n2366,n2391);
and (n2394,n2327,n2328);
xor (n2395,n1988,n2099);
and (n2396,n2323,n2324);
xor (n2397,n1947,n1986);
xor (n2398,n2247,n2250);
and (n2399,n2320,n2397);
or (n2400,n2401,n2767);
and (n2401,n2402,n2510);
xor (n2402,n2403,n2404);
xor (n2403,n2319,n2398);
or (n2404,n2405,n2509);
and (n2405,n2406,n2508);
xor (n2406,n2407,n2408);
xor (n2407,n2252,n2295);
or (n2408,n2409,n2507);
and (n2409,n2410,n2506);
xor (n2410,n2411,n2412);
xor (n2411,n2255,n2258);
or (n2412,n2413,n2505);
and (n2413,n2414,n2438);
xor (n2414,n2415,n2437);
or (n2415,n2416,n2436);
and (n2416,n2417,n2420);
xor (n2417,n2418,n2419);
and (n2418,n2208,n981);
xor (n2419,n2262,n2266);
or (n2420,n2421,n2435);
and (n2421,n2422,n2434);
xor (n2422,n2423,n2432);
or (n2423,n2424,n2431);
and (n2424,n2425,n2429);
xor (n2425,n2426,n2428);
and (n2426,n2427,n1224);
xor (n2427,n1210,n1215);
xor (n2428,n2024,n2029);
and (n2429,n2430,n1273);
xor (n2430,n881,n897);
and (n2431,n2426,n2428);
and (n2432,n2433,n1224);
xor (n2433,n1204,n1217);
wire s0n2434,s1n2434,notn2434;
or (n2434,s0n2434,s1n2434);
not(notn2434,n931);
and (s0n2434,notn2434,1'b0);
and (s1n2434,n931,n1980);
and (n2435,n2423,n2432);
and (n2436,n2418,n2419);
xor (n2437,n2260,n2291);
or (n2438,n2439,n2504);
and (n2439,n2440,n2503);
xor (n2440,n2441,n2442);
xor (n2441,n2270,n2289);
or (n2442,n2443,n2502);
and (n2443,n2444,n2501);
xor (n2444,n2445,n2446);
and (n2445,n2267,n933);
or (n2446,n2447,n2500);
and (n2447,n2448,n2473);
xor (n2448,n2449,n2450);
xor (n2449,n2282,n2286);
or (n2450,n2451,n2472);
and (n2451,n2452,n2471);
xor (n2452,n2453,n2461);
or (n2453,n2454,n2460);
and (n2454,n2455,n2458);
xor (n2455,n2456,n2457);
xor (n2456,n2381,n2382);
wire s0n2457,s1n2457,notn2457;
or (n2457,s0n2457,s1n2457);
not(notn2457,n933);
and (s0n2457,notn2457,1'b0);
and (s1n2457,n933,n2379);
and (n2458,n2459,n981);
not (n2459,n1583);
and (n2460,n2456,n2457);
or (n2461,n2462,n2470);
and (n2462,n2463,n2466);
xor (n2463,n2464,n2465);
and (n2464,n1364,n981);
and (n2465,n1663,n981);
and (n2466,n2467,n981);
xor (n2467,n2468,n2469);
not (n2468,n1675);
not (n2469,n1725);
and (n2470,n2464,n2465);
wire s0n2471,s1n2471,notn2471;
or (n2471,s0n2471,s1n2471);
not(notn2471,n931);
and (s0n2471,notn2471,1'b0);
and (s1n2471,n931,n2060);
and (n2472,n2453,n2461);
or (n2473,n2474,n2499);
and (n2474,n2475,n2497);
xor (n2475,n2476,n2494);
or (n2476,n2477,n2493);
and (n2477,n2478,n2492);
xor (n2478,n2479,n2487);
or (n2479,n2480,n2486);
and (n2480,n2481,n2484);
xor (n2481,n2482,n2483);
nor (n2482,n1569,n980);
wire s0n2483,s1n2483,notn2483;
or (n2483,s0n2483,s1n2483);
not(notn2483,n933);
and (s0n2483,notn2483,1'b0);
and (s1n2483,n933,n2032);
nor (n2484,n2485,n980);
not (n2485,n1690);
and (n2486,n2482,n2483);
and (n2487,n2488,n2490);
nor (n2488,n2489,n980);
not (n2489,n1380);
nor (n2490,n2491,n980);
not (n2491,n1678);
wire s0n2492,s1n2492,notn2492;
or (n2492,s0n2492,s1n2492);
not(notn2492,n1273);
and (s0n2492,notn2492,1'b0);
and (s1n2492,n1273,n2356);
and (n2493,n2479,n2487);
xor (n2494,n2495,n2496);
xor (n2495,n2378,n2380);
wire s0n2496,s1n2496,notn2496;
or (n2496,s0n2496,s1n2496);
not(notn2496,n1424);
and (s0n2496,notn2496,1'b0);
and (s1n2496,n1424,n2036);
and (n2497,n2498,n1224);
xor (n2498,n1212,n1213);
and (n2499,n2476,n2494);
and (n2500,n2449,n2450);
and (n2501,n2094,n981);
and (n2502,n2445,n2446);
xor (n2503,n2335,n2360);
and (n2504,n2441,n2442);
and (n2505,n2415,n2437);
xor (n2506,n2297,n2306);
and (n2507,n2411,n2412);
xor (n2508,n2322,n2395);
and (n2509,n2407,n2408);
or (n2510,n2511,n2766);
and (n2511,n2512,n2574);
xor (n2512,n2513,n2573);
or (n2513,n2514,n2572);
and (n2514,n2515,n2571);
xor (n2515,n2516,n2570);
or (n2516,n2517,n2569);
and (n2517,n2518,n2568);
xor (n2518,n2519,n2567);
or (n2519,n2520,n2566);
and (n2520,n2521,n2565);
xor (n2521,n2522,n2558);
or (n2522,n2523,n2557);
and (n2523,n2524,n2550);
xor (n2524,n2525,n2528);
xor (n2525,n2526,n2527);
xor (n2526,n2337,n2358);
and (n2527,n2430,n1424);
or (n2528,n2529,n2549);
and (n2529,n2530,n2548);
xor (n2530,n2531,n2545);
or (n2531,n2532,n2544);
and (n2532,n2533,n2543);
xor (n2533,n2534,n2536);
wire s0n2534,s1n2534,notn2534;
or (n2534,s0n2534,s1n2534);
not(notn2534,n1273);
and (s0n2534,notn2534,1'b0);
and (s1n2534,n1273,n2535);
xor (n2535,n883,n895);
or (n2536,n2537,n2542);
and (n2537,n2538,n2541);
xor (n2538,n2539,n2540);
xor (n2539,n2463,n2466);
wire s0n2540,s1n2540,notn2540;
or (n2540,s0n2540,s1n2540);
not(notn2540,n931);
and (s0n2540,notn2540,1'b0);
and (s1n2540,n931,n2028);
wire s0n2541,s1n2541,notn2541;
or (n2541,s0n2541,s1n2541);
not(notn2541,n1273);
and (s0n2541,notn2541,1'b0);
and (s1n2541,n1273,n2036);
and (n2542,n2539,n2540);
xor (n2543,n2340,n2343);
and (n2544,n2534,n2536);
xor (n2545,n2546,n2547);
xor (n2546,n2338,n2345);
wire s0n2547,s1n2547,notn2547;
or (n2547,s0n2547,s1n2547);
not(notn2547,n1424);
and (s0n2547,notn2547,1'b0);
and (s1n2547,n1424,n2535);
and (n2548,n2264,n931);
and (n2549,n2531,n2545);
or (n2550,n2551,n2556);
and (n2551,n2552,n2555);
xor (n2552,n2553,n2554);
and (n2553,n2433,n933);
xor (n2554,n2375,n2384);
wire s0n2555,s1n2555,notn2555;
or (n2555,s0n2555,s1n2555);
not(notn2555,n981);
and (s0n2555,notn2555,1'b0);
and (s1n2555,n981,n1980);
and (n2556,n2553,n2554);
and (n2557,n2525,n2528);
or (n2558,n2559,n2564);
and (n2559,n2560,n2563);
xor (n2560,n2561,n2562);
xor (n2561,n2274,n2280);
xor (n2562,n2371,n2386);
wire s0n2563,s1n2563,notn2563;
or (n2563,s0n2563,s1n2563);
not(notn2563,n981);
and (s0n2563,notn2563,1'b0);
and (s1n2563,n981,n2064);
and (n2564,n2561,n2562);
xor (n2565,n2368,n2389);
and (n2566,n2522,n2558);
xor (n2567,n2330,n2333);
xor (n2568,n2365,n2392);
and (n2569,n2519,n2567);
xor (n2570,n2326,n2363);
xor (n2571,n2410,n2506);
and (n2572,n2516,n2570);
xor (n2573,n2406,n2508);
or (n2574,n2575,n2765);
and (n2575,n2576,n2652);
xor (n2576,n2577,n2651);
or (n2577,n2578,n2650);
and (n2578,n2579,n2649);
xor (n2579,n2580,n2581);
xor (n2580,n2414,n2438);
or (n2581,n2582,n2648);
and (n2582,n2583,n2647);
xor (n2583,n2584,n2585);
xor (n2584,n2417,n2420);
or (n2585,n2586,n2646);
and (n2586,n2587,n2602);
xor (n2587,n2588,n2589);
xor (n2588,n2422,n2434);
or (n2589,n2590,n2601);
and (n2590,n2591,n2600);
xor (n2591,n2592,n2593);
xor (n2592,n2425,n2429);
or (n2593,n2594,n2599);
and (n2594,n2595,n2598);
xor (n2595,n2596,n2597);
and (n2596,n2427,n933);
xor (n2597,n2346,n2357);
and (n2598,n2430,n931);
and (n2599,n2596,n2597);
and (n2600,n2267,n981);
and (n2601,n2592,n2593);
or (n2602,n2603,n2645);
and (n2603,n2604,n2626);
xor (n2604,n2605,n2606);
xor (n2605,n2448,n2473);
or (n2606,n2607,n2625);
and (n2607,n2608,n2624);
xor (n2608,n2609,n2623);
or (n2609,n2610,n2622);
and (n2610,n2611,n2621);
xor (n2611,n2612,n2613);
xor (n2612,n2455,n2458);
or (n2613,n2614,n2620);
and (n2614,n2615,n2619);
xor (n2615,n2616,n2618);
and (n2616,n2035,n2617);
wire s0n2617,s1n2617,notn2617;
or (n2617,s0n2617,s1n2617);
not(notn2617,n981);
and (s0n2617,notn2617,1'b0);
and (s1n2617,n981,n2383);
wire s0n2618,s1n2618,notn2618;
or (n2618,s0n2618,s1n2618);
not(notn2618,n933);
and (s0n2618,notn2618,1'b0);
and (s1n2618,n933,n2383);
xor (n2619,n2488,n2490);
and (n2620,n2616,n2618);
wire s0n2621,s1n2621,notn2621;
or (n2621,s0n2621,s1n2621);
not(notn2621,n931);
and (s0n2621,notn2621,1'b0);
and (s1n2621,n931,n2535);
and (n2622,n2612,n2613);
xor (n2623,n2452,n2471);
and (n2624,n2433,n981);
and (n2625,n2609,n2623);
or (n2626,n2627,n2644);
and (n2627,n2628,n2643);
xor (n2628,n2629,n2630);
xor (n2629,n2475,n2497);
or (n2630,n2631,n2642);
and (n2631,n2632,n2641);
xor (n2632,n2633,n2634);
xor (n2633,n2538,n2541);
or (n2634,n2635,n2640);
and (n2635,n2636,n2639);
xor (n2636,n2637,n2638);
wire s0n2637,s1n2637,notn2637;
or (n2637,s0n2637,s1n2637);
not(notn2637,n931);
and (s0n2637,notn2637,1'b0);
and (s1n2637,n931,n2356);
xor (n2638,n2481,n2484);
wire s0n2639,s1n2639,notn2639;
or (n2639,s0n2639,s1n2639);
not(notn2639,n931);
and (s0n2639,notn2639,1'b0);
and (s1n2639,n931,n2036);
and (n2640,n2637,n2638);
and (n2641,n2498,n933);
and (n2642,n2633,n2634);
and (n2643,n2264,n981);
and (n2644,n2629,n2630);
and (n2645,n2605,n2606);
and (n2646,n2588,n2589);
xor (n2647,n2440,n2503);
and (n2648,n2584,n2585);
xor (n2649,n2518,n2568);
and (n2650,n2580,n2581);
xor (n2651,n2515,n2571);
nand (n2652,n2653,n2764);
or (n2653,n2654,n2669);
nor (n2654,n2655,n2656);
xor (n2655,n2579,n2649);
or (n2656,n2657,n2668);
and (n2657,n2658,n2667);
xor (n2658,n2659,n2660);
xor (n2659,n2521,n2565);
or (n2660,n2661,n2666);
and (n2661,n2662,n2665);
xor (n2662,n2663,n2664);
xor (n2663,n2444,n2501);
xor (n2664,n2560,n2563);
xor (n2665,n2524,n2550);
and (n2666,n2663,n2664);
xor (n2667,n2583,n2647);
and (n2668,n2659,n2660);
and (n2669,n2670,n2763);
nand (n2670,n2671,n2686);
or (n2671,n2672,n2673);
xor (n2672,n2658,n2667);
or (n2673,n2674,n2685);
and (n2674,n2675,n2684);
xor (n2675,n2676,n2683);
or (n2676,n2677,n2682);
and (n2677,n2678,n2681);
xor (n2678,n2679,n2680);
xor (n2679,n2552,n2555);
xor (n2680,n2530,n2548);
xor (n2681,n2591,n2600);
and (n2682,n2679,n2680);
xor (n2683,n2587,n2602);
xor (n2684,n2662,n2665);
and (n2685,n2676,n2683);
nand (n2686,n2687,n2756);
nand (n2687,n2688,n2727,n2730);
or (n2688,n2689,n2726);
or (n2689,n2690,n2725);
and (n2690,n2691,n2724);
xor (n2691,n2692,n2711);
or (n2692,n2693,n2710);
and (n2693,n2694,n2709);
xor (n2694,n2695,n2696);
xor (n2695,n2608,n2624);
or (n2696,n2697,n2708);
and (n2697,n2698,n2707);
xor (n2698,n2699,n2700);
xor (n2699,n2611,n2621);
or (n2700,n2701,n2706);
and (n2701,n2702,n2705);
xor (n2702,n2703,n2704);
xor (n2703,n2615,n2619);
wire s0n2704,s1n2704,notn2704;
or (n2704,s0n2704,s1n2704);
not(notn2704,n981);
and (s0n2704,notn2704,1'b0);
and (s1n2704,n981,n2535);
and (n2705,n2498,n981);
and (n2706,n2703,n2704);
xor (n2707,n2632,n2641);
and (n2708,n2699,n2700);
xor (n2709,n2628,n2643);
and (n2710,n2695,n2696);
or (n2711,n2712,n2723);
and (n2712,n2713,n2722);
xor (n2713,n2714,n2721);
or (n2714,n2715,n2720);
and (n2715,n2716,n2719);
xor (n2716,n2717,n2718);
and (n2717,n2427,n981);
xor (n2718,n2478,n2492);
and (n2719,n2430,n981);
and (n2720,n2717,n2718);
xor (n2721,n2533,n2543);
xor (n2722,n2595,n2598);
and (n2723,n2714,n2721);
xor (n2724,n2604,n2626);
and (n2725,n2692,n2711);
xor (n2726,n2675,n2684);
or (n2727,n2728,n2729);
xor (n2728,n2691,n2724);
xor (n2729,n2678,n2681);
nand (n2730,n2731,n2752);
or (n2731,n2732,n2735);
nor (n2732,n2733,n2734);
xor (n2733,n2694,n2709);
xor (n2734,n2713,n2722);
nand (n2735,n2736,n2739,n2742);
or (n2736,n2737,n2738);
xor (n2737,n2716,n2719);
xor (n2738,n2698,n2707);
or (n2739,n2740,n2741);
xor (n2740,n2636,n2639);
xor (n2741,n2702,n2705);
nand (n2742,n2743,n2746);
or (n2743,n2744,n2745);
not (n2744,n2740);
not (n2745,n2741);
nor (n2746,n2747,n2751);
and (n2747,n2748,n2749);
xor (n2748,n2035,n2617);
or (n2749,n2750,n2031);
wire s0n2750,s1n2750,notn2750;
or (n2750,s0n2750,s1n2750);
not(notn2750,n981);
and (s0n2750,notn2750,1'b0);
and (s1n2750,n981,n2356);
and (n2751,n2750,n2031);
nor (n2752,n2753,n2755);
and (n2753,n2754,n2737,n2738);
not (n2754,n2732);
and (n2755,n2733,n2734);
nor (n2756,n2757,n2761);
and (n2757,n2726,n2758);
nand (n2758,n2759,n2760);
not (n2759,n2689);
nand (n2760,n2728,n2729);
and (n2761,n2762,n2689);
not (n2762,n2760);
nand (n2763,n2672,n2673);
nand (n2764,n2655,n2656);
and (n2765,n2577,n2651);
and (n2766,n2513,n2573);
and (n2767,n2403,n2404);
and (n2768,n2316,n2317);
and (n2769,n2241,n2242);
not (n2770,n0);
endmodule
