module top (out,n24,n25,n26,n28,n29,n34,n35,n38,n39
        ,n47,n48,n56,n57,n65,n66,n74,n75,n83,n84
        ,n92,n93,n101,n102,n110,n111,n119,n120,n127,n128
        ,n131,n132,n198,n199,n259,n260,n314,n315,n363,n364
        ,n406,n407,n443,n444,n474,n475,n499,n500,n518,n519);
output out;
input n24;
input n25;
input n26;
input n28;
input n29;
input n34;
input n35;
input n38;
input n39;
input n47;
input n48;
input n56;
input n57;
input n65;
input n66;
input n74;
input n75;
input n83;
input n84;
input n92;
input n93;
input n101;
input n102;
input n110;
input n111;
input n119;
input n120;
input n127;
input n128;
input n131;
input n132;
input n198;
input n199;
input n259;
input n260;
input n314;
input n315;
input n363;
input n364;
input n406;
input n407;
input n443;
input n444;
input n474;
input n475;
input n499;
input n500;
input n518;
input n519;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n129;
wire n130;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
xor (out,n0,n529);
buf (n0,n1);
xor (n1,n2,n520);
xor (n2,n3,n516);
xor (n3,n4,n501);
xor (n4,n5,n497);
xor (n5,n6,n476);
xor (n6,n7,n472);
xor (n7,n8,n445);
xor (n8,n9,n441);
xor (n9,n10,n408);
xor (n10,n11,n404);
xor (n11,n12,n365);
xor (n12,n13,n361);
xor (n13,n14,n316);
xor (n14,n15,n312);
xor (n15,n16,n261);
xor (n16,n17,n257);
xor (n17,n18,n200);
xor (n18,n19,n196);
xor (n19,n20,n133);
xor (n20,n21,n129);
and (n21,n22,n30);
and (n22,n23,n27);
wire s0n23,s1n23,notn23;
or (n23,s0n23,s1n23);
not(notn23,n26);
and (s0n23,notn23,n24);
and (s1n23,n26,n25);
wire s0n27,s1n27,notn27;
or (n27,s0n27,s1n27);
not(notn27,n26);
and (s0n27,notn27,n28);
and (s1n27,n26,n29);
or (n30,n31,n40);
and (n31,n32,n36);
and (n32,n23,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n26);
and (s0n33,notn33,n34);
and (s1n33,n26,n35);
and (n36,n37,n27);
wire s0n37,s1n37,notn37;
or (n37,s0n37,s1n37);
not(notn37,n26);
and (s0n37,notn37,n38);
and (s1n37,n26,n39);
and (n40,n41,n42);
xor (n41,n32,n36);
or (n42,n43,n49);
and (n43,n44,n45);
and (n44,n37,n33);
and (n45,n46,n27);
wire s0n46,s1n46,notn46;
or (n46,s0n46,s1n46);
not(notn46,n26);
and (s0n46,notn46,n47);
and (s1n46,n26,n48);
and (n49,n50,n51);
xor (n50,n44,n45);
or (n51,n52,n58);
and (n52,n53,n54);
and (n53,n46,n33);
and (n54,n55,n27);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n26);
and (s0n55,notn55,n56);
and (s1n55,n26,n57);
and (n58,n59,n60);
xor (n59,n53,n54);
or (n60,n61,n67);
and (n61,n62,n63);
and (n62,n55,n33);
and (n63,n64,n27);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n26);
and (s0n64,notn64,n65);
and (s1n64,n26,n66);
and (n67,n68,n69);
xor (n68,n62,n63);
or (n69,n70,n76);
and (n70,n71,n72);
and (n71,n64,n33);
and (n72,n73,n27);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n26);
and (s0n73,notn73,n74);
and (s1n73,n26,n75);
and (n76,n77,n78);
xor (n77,n71,n72);
or (n78,n79,n85);
and (n79,n80,n81);
and (n80,n73,n33);
and (n81,n82,n27);
wire s0n82,s1n82,notn82;
or (n82,s0n82,s1n82);
not(notn82,n26);
and (s0n82,notn82,n83);
and (s1n82,n26,n84);
and (n85,n86,n87);
xor (n86,n80,n81);
or (n87,n88,n94);
and (n88,n89,n90);
and (n89,n82,n33);
and (n90,n91,n27);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n26);
and (s0n91,notn91,n92);
and (s1n91,n26,n93);
and (n94,n95,n96);
xor (n95,n89,n90);
or (n96,n97,n103);
and (n97,n98,n99);
and (n98,n91,n33);
and (n99,n100,n27);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n26);
and (s0n100,notn100,n101);
and (s1n100,n26,n102);
and (n103,n104,n105);
xor (n104,n98,n99);
or (n105,n106,n112);
and (n106,n107,n108);
and (n107,n100,n33);
and (n108,n109,n27);
wire s0n109,s1n109,notn109;
or (n109,s0n109,s1n109);
not(notn109,n26);
and (s0n109,notn109,n110);
and (s1n109,n26,n111);
and (n112,n113,n114);
xor (n113,n107,n108);
or (n114,n115,n121);
and (n115,n116,n117);
and (n116,n109,n33);
and (n117,n118,n27);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n26);
and (s0n118,notn118,n119);
and (s1n118,n26,n120);
and (n121,n122,n123);
xor (n122,n116,n117);
and (n123,n124,n125);
and (n124,n118,n33);
and (n125,n126,n27);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n26);
and (s0n126,notn126,n127);
and (s1n126,n26,n128);
and (n129,n23,n130);
wire s0n130,s1n130,notn130;
or (n130,s0n130,s1n130);
not(notn130,n26);
and (s0n130,notn130,n131);
and (s1n130,n26,n132);
or (n133,n134,n137);
and (n134,n135,n136);
xor (n135,n22,n30);
and (n136,n37,n130);
and (n137,n138,n139);
xor (n138,n135,n136);
or (n139,n140,n143);
and (n140,n141,n142);
xor (n141,n41,n42);
and (n142,n46,n130);
and (n143,n144,n145);
xor (n144,n141,n142);
or (n145,n146,n149);
and (n146,n147,n148);
xor (n147,n50,n51);
and (n148,n55,n130);
and (n149,n150,n151);
xor (n150,n147,n148);
or (n151,n152,n155);
and (n152,n153,n154);
xor (n153,n59,n60);
and (n154,n64,n130);
and (n155,n156,n157);
xor (n156,n153,n154);
or (n157,n158,n161);
and (n158,n159,n160);
xor (n159,n68,n69);
and (n160,n73,n130);
and (n161,n162,n163);
xor (n162,n159,n160);
or (n163,n164,n167);
and (n164,n165,n166);
xor (n165,n77,n78);
and (n166,n82,n130);
and (n167,n168,n169);
xor (n168,n165,n166);
or (n169,n170,n173);
and (n170,n171,n172);
xor (n171,n86,n87);
and (n172,n91,n130);
and (n173,n174,n175);
xor (n174,n171,n172);
or (n175,n176,n179);
and (n176,n177,n178);
xor (n177,n95,n96);
and (n178,n100,n130);
and (n179,n180,n181);
xor (n180,n177,n178);
or (n181,n182,n185);
and (n182,n183,n184);
xor (n183,n104,n105);
and (n184,n109,n130);
and (n185,n186,n187);
xor (n186,n183,n184);
or (n187,n188,n191);
and (n188,n189,n190);
xor (n189,n113,n114);
and (n190,n118,n130);
and (n191,n192,n193);
xor (n192,n189,n190);
and (n193,n194,n195);
xor (n194,n122,n123);
and (n195,n126,n130);
and (n196,n37,n197);
wire s0n197,s1n197,notn197;
or (n197,s0n197,s1n197);
not(notn197,n26);
and (s0n197,notn197,n198);
and (s1n197,n26,n199);
or (n200,n201,n204);
and (n201,n202,n203);
xor (n202,n138,n139);
and (n203,n46,n197);
and (n204,n205,n206);
xor (n205,n202,n203);
or (n206,n207,n210);
and (n207,n208,n209);
xor (n208,n144,n145);
and (n209,n55,n197);
and (n210,n211,n212);
xor (n211,n208,n209);
or (n212,n213,n216);
and (n213,n214,n215);
xor (n214,n150,n151);
and (n215,n64,n197);
and (n216,n217,n218);
xor (n217,n214,n215);
or (n218,n219,n222);
and (n219,n220,n221);
xor (n220,n156,n157);
and (n221,n73,n197);
and (n222,n223,n224);
xor (n223,n220,n221);
or (n224,n225,n228);
and (n225,n226,n227);
xor (n226,n162,n163);
and (n227,n82,n197);
and (n228,n229,n230);
xor (n229,n226,n227);
or (n230,n231,n234);
and (n231,n232,n233);
xor (n232,n168,n169);
and (n233,n91,n197);
and (n234,n235,n236);
xor (n235,n232,n233);
or (n236,n237,n240);
and (n237,n238,n239);
xor (n238,n174,n175);
and (n239,n100,n197);
and (n240,n241,n242);
xor (n241,n238,n239);
or (n242,n243,n246);
and (n243,n244,n245);
xor (n244,n180,n181);
and (n245,n109,n197);
and (n246,n247,n248);
xor (n247,n244,n245);
or (n248,n249,n252);
and (n249,n250,n251);
xor (n250,n186,n187);
and (n251,n118,n197);
and (n252,n253,n254);
xor (n253,n250,n251);
and (n254,n255,n256);
xor (n255,n192,n193);
and (n256,n126,n197);
and (n257,n46,n258);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n26);
and (s0n258,notn258,n259);
and (s1n258,n26,n260);
or (n261,n262,n265);
and (n262,n263,n264);
xor (n263,n205,n206);
and (n264,n55,n258);
and (n265,n266,n267);
xor (n266,n263,n264);
or (n267,n268,n271);
and (n268,n269,n270);
xor (n269,n211,n212);
and (n270,n64,n258);
and (n271,n272,n273);
xor (n272,n269,n270);
or (n273,n274,n277);
and (n274,n275,n276);
xor (n275,n217,n218);
and (n276,n73,n258);
and (n277,n278,n279);
xor (n278,n275,n276);
or (n279,n280,n283);
and (n280,n281,n282);
xor (n281,n223,n224);
and (n282,n82,n258);
and (n283,n284,n285);
xor (n284,n281,n282);
or (n285,n286,n289);
and (n286,n287,n288);
xor (n287,n229,n230);
and (n288,n91,n258);
and (n289,n290,n291);
xor (n290,n287,n288);
or (n291,n292,n295);
and (n292,n293,n294);
xor (n293,n235,n236);
and (n294,n100,n258);
and (n295,n296,n297);
xor (n296,n293,n294);
or (n297,n298,n301);
and (n298,n299,n300);
xor (n299,n241,n242);
and (n300,n109,n258);
and (n301,n302,n303);
xor (n302,n299,n300);
or (n303,n304,n307);
and (n304,n305,n306);
xor (n305,n247,n248);
and (n306,n118,n258);
and (n307,n308,n309);
xor (n308,n305,n306);
and (n309,n310,n311);
xor (n310,n253,n254);
and (n311,n126,n258);
and (n312,n55,n313);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n26);
and (s0n313,notn313,n314);
and (s1n313,n26,n315);
or (n316,n317,n320);
and (n317,n318,n319);
xor (n318,n266,n267);
and (n319,n64,n313);
and (n320,n321,n322);
xor (n321,n318,n319);
or (n322,n323,n326);
and (n323,n324,n325);
xor (n324,n272,n273);
and (n325,n73,n313);
and (n326,n327,n328);
xor (n327,n324,n325);
or (n328,n329,n332);
and (n329,n330,n331);
xor (n330,n278,n279);
and (n331,n82,n313);
and (n332,n333,n334);
xor (n333,n330,n331);
or (n334,n335,n338);
and (n335,n336,n337);
xor (n336,n284,n285);
and (n337,n91,n313);
and (n338,n339,n340);
xor (n339,n336,n337);
or (n340,n341,n344);
and (n341,n342,n343);
xor (n342,n290,n291);
and (n343,n100,n313);
and (n344,n345,n346);
xor (n345,n342,n343);
or (n346,n347,n350);
and (n347,n348,n349);
xor (n348,n296,n297);
and (n349,n109,n313);
and (n350,n351,n352);
xor (n351,n348,n349);
or (n352,n353,n356);
and (n353,n354,n355);
xor (n354,n302,n303);
and (n355,n118,n313);
and (n356,n357,n358);
xor (n357,n354,n355);
and (n358,n359,n360);
xor (n359,n308,n309);
and (n360,n126,n313);
and (n361,n64,n362);
wire s0n362,s1n362,notn362;
or (n362,s0n362,s1n362);
not(notn362,n26);
and (s0n362,notn362,n363);
and (s1n362,n26,n364);
or (n365,n366,n369);
and (n366,n367,n368);
xor (n367,n321,n322);
and (n368,n73,n362);
and (n369,n370,n371);
xor (n370,n367,n368);
or (n371,n372,n375);
and (n372,n373,n374);
xor (n373,n327,n328);
and (n374,n82,n362);
and (n375,n376,n377);
xor (n376,n373,n374);
or (n377,n378,n381);
and (n378,n379,n380);
xor (n379,n333,n334);
and (n380,n91,n362);
and (n381,n382,n383);
xor (n382,n379,n380);
or (n383,n384,n387);
and (n384,n385,n386);
xor (n385,n339,n340);
and (n386,n100,n362);
and (n387,n388,n389);
xor (n388,n385,n386);
or (n389,n390,n393);
and (n390,n391,n392);
xor (n391,n345,n346);
and (n392,n109,n362);
and (n393,n394,n395);
xor (n394,n391,n392);
or (n395,n396,n399);
and (n396,n397,n398);
xor (n397,n351,n352);
and (n398,n118,n362);
and (n399,n400,n401);
xor (n400,n397,n398);
and (n401,n402,n403);
xor (n402,n357,n358);
and (n403,n126,n362);
and (n404,n73,n405);
wire s0n405,s1n405,notn405;
or (n405,s0n405,s1n405);
not(notn405,n26);
and (s0n405,notn405,n406);
and (s1n405,n26,n407);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n370,n371);
and (n411,n82,n405);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n376,n377);
and (n417,n91,n405);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n382,n383);
and (n423,n100,n405);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n388,n389);
and (n429,n109,n405);
and (n430,n431,n432);
xor (n431,n428,n429);
or (n432,n433,n436);
and (n433,n434,n435);
xor (n434,n394,n395);
and (n435,n118,n405);
and (n436,n437,n438);
xor (n437,n434,n435);
and (n438,n439,n440);
xor (n439,n400,n401);
and (n440,n126,n405);
and (n441,n82,n442);
wire s0n442,s1n442,notn442;
or (n442,s0n442,s1n442);
not(notn442,n26);
and (s0n442,notn442,n443);
and (s1n442,n26,n444);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n413,n414);
and (n448,n91,n442);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n419,n420);
and (n454,n100,n442);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n425,n426);
and (n460,n109,n442);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n431,n432);
and (n466,n118,n442);
and (n467,n468,n469);
xor (n468,n465,n466);
and (n469,n470,n471);
xor (n470,n437,n438);
and (n471,n126,n442);
and (n472,n91,n473);
wire s0n473,s1n473,notn473;
or (n473,s0n473,s1n473);
not(notn473,n26);
and (s0n473,notn473,n474);
and (s1n473,n26,n475);
or (n476,n477,n480);
and (n477,n478,n479);
xor (n478,n450,n451);
and (n479,n100,n473);
and (n480,n481,n482);
xor (n481,n478,n479);
or (n482,n483,n486);
and (n483,n484,n485);
xor (n484,n456,n457);
and (n485,n109,n473);
and (n486,n487,n488);
xor (n487,n484,n485);
or (n488,n489,n492);
and (n489,n490,n491);
xor (n490,n462,n463);
and (n491,n118,n473);
and (n492,n493,n494);
xor (n493,n490,n491);
and (n494,n495,n496);
xor (n495,n468,n469);
and (n496,n126,n473);
and (n497,n100,n498);
wire s0n498,s1n498,notn498;
or (n498,s0n498,s1n498);
not(notn498,n26);
and (s0n498,notn498,n499);
and (s1n498,n26,n500);
or (n501,n502,n505);
and (n502,n503,n504);
xor (n503,n481,n482);
and (n504,n109,n498);
and (n505,n506,n507);
xor (n506,n503,n504);
or (n507,n508,n511);
and (n508,n509,n510);
xor (n509,n487,n488);
and (n510,n118,n498);
and (n511,n512,n513);
xor (n512,n509,n510);
and (n513,n514,n515);
xor (n514,n493,n494);
and (n515,n126,n498);
and (n516,n109,n517);
wire s0n517,s1n517,notn517;
or (n517,s0n517,s1n517);
not(notn517,n26);
and (s0n517,notn517,n518);
and (s1n517,n26,n519);
or (n520,n521,n524);
and (n521,n522,n523);
xor (n522,n506,n507);
and (n523,n118,n517);
and (n524,n525,n526);
xor (n525,n522,n523);
and (n526,n527,n528);
xor (n527,n512,n513);
and (n528,n126,n517);
wire s0n529,s1n529,notn529;
or (n529,s0n529,s1n529);
not(notn529,n26);
and (s0n529,notn529,n530);
and (s1n529,n26,n1010);
buf (n530,n531);
xor (n531,n532,n1001);
xor (n532,n533,n999);
xor (n533,n534,n984);
xor (n534,n535,n982);
xor (n535,n536,n961);
xor (n536,n537,n959);
xor (n537,n538,n932);
xor (n538,n539,n930);
xor (n539,n540,n897);
xor (n540,n541,n895);
xor (n541,n542,n856);
xor (n542,n543,n854);
xor (n543,n544,n809);
xor (n544,n545,n807);
xor (n545,n546,n756);
xor (n546,n547,n754);
xor (n547,n548,n697);
xor (n548,n549,n695);
xor (n549,n550,n632);
xor (n550,n551,n630);
and (n551,n552,n555);
and (n552,n553,n554);
buf (n553,n24);
buf (n554,n28);
or (n555,n556,n561);
and (n556,n557,n559);
and (n557,n553,n558);
buf (n558,n34);
and (n559,n560,n554);
buf (n560,n38);
and (n561,n562,n563);
xor (n562,n557,n559);
or (n563,n564,n568);
and (n564,n565,n566);
and (n565,n560,n558);
and (n566,n567,n554);
buf (n567,n47);
and (n568,n569,n570);
xor (n569,n565,n566);
or (n570,n571,n575);
and (n571,n572,n573);
and (n572,n567,n558);
and (n573,n574,n554);
buf (n574,n56);
and (n575,n576,n577);
xor (n576,n572,n573);
or (n577,n578,n582);
and (n578,n579,n580);
and (n579,n574,n558);
and (n580,n581,n554);
buf (n581,n65);
and (n582,n583,n584);
xor (n583,n579,n580);
or (n584,n585,n589);
and (n585,n586,n587);
and (n586,n581,n558);
and (n587,n588,n554);
buf (n588,n74);
and (n589,n590,n591);
xor (n590,n586,n587);
or (n591,n592,n596);
and (n592,n593,n594);
and (n593,n588,n558);
and (n594,n595,n554);
buf (n595,n83);
and (n596,n597,n598);
xor (n597,n593,n594);
or (n598,n599,n603);
and (n599,n600,n601);
and (n600,n595,n558);
and (n601,n602,n554);
buf (n602,n92);
and (n603,n604,n605);
xor (n604,n600,n601);
or (n605,n606,n610);
and (n606,n607,n608);
and (n607,n602,n558);
and (n608,n609,n554);
buf (n609,n101);
and (n610,n611,n612);
xor (n611,n607,n608);
or (n612,n613,n617);
and (n613,n614,n615);
and (n614,n609,n558);
and (n615,n616,n554);
buf (n616,n110);
and (n617,n618,n619);
xor (n618,n614,n615);
or (n619,n620,n624);
and (n620,n621,n622);
and (n621,n616,n558);
and (n622,n623,n554);
buf (n623,n119);
and (n624,n625,n626);
xor (n625,n621,n622);
and (n626,n627,n628);
and (n627,n623,n558);
and (n628,n629,n554);
buf (n629,n127);
and (n630,n553,n631);
buf (n631,n131);
or (n632,n633,n636);
and (n633,n634,n635);
xor (n634,n552,n555);
and (n635,n560,n631);
and (n636,n637,n638);
xor (n637,n634,n635);
or (n638,n639,n642);
and (n639,n640,n641);
xor (n640,n562,n563);
and (n641,n567,n631);
and (n642,n643,n644);
xor (n643,n640,n641);
or (n644,n645,n648);
and (n645,n646,n647);
xor (n646,n569,n570);
and (n647,n574,n631);
and (n648,n649,n650);
xor (n649,n646,n647);
or (n650,n651,n654);
and (n651,n652,n653);
xor (n652,n576,n577);
and (n653,n581,n631);
and (n654,n655,n656);
xor (n655,n652,n653);
or (n656,n657,n660);
and (n657,n658,n659);
xor (n658,n583,n584);
and (n659,n588,n631);
and (n660,n661,n662);
xor (n661,n658,n659);
or (n662,n663,n666);
and (n663,n664,n665);
xor (n664,n590,n591);
and (n665,n595,n631);
and (n666,n667,n668);
xor (n667,n664,n665);
or (n668,n669,n672);
and (n669,n670,n671);
xor (n670,n597,n598);
and (n671,n602,n631);
and (n672,n673,n674);
xor (n673,n670,n671);
or (n674,n675,n678);
and (n675,n676,n677);
xor (n676,n604,n605);
and (n677,n609,n631);
and (n678,n679,n680);
xor (n679,n676,n677);
or (n680,n681,n684);
and (n681,n682,n683);
xor (n682,n611,n612);
and (n683,n616,n631);
and (n684,n685,n686);
xor (n685,n682,n683);
or (n686,n687,n690);
and (n687,n688,n689);
xor (n688,n618,n619);
and (n689,n623,n631);
and (n690,n691,n692);
xor (n691,n688,n689);
and (n692,n693,n694);
xor (n693,n625,n626);
and (n694,n629,n631);
and (n695,n560,n696);
buf (n696,n198);
or (n697,n698,n701);
and (n698,n699,n700);
xor (n699,n637,n638);
and (n700,n567,n696);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n643,n644);
and (n706,n574,n696);
and (n707,n708,n709);
xor (n708,n705,n706);
or (n709,n710,n713);
and (n710,n711,n712);
xor (n711,n649,n650);
and (n712,n581,n696);
and (n713,n714,n715);
xor (n714,n711,n712);
or (n715,n716,n719);
and (n716,n717,n718);
xor (n717,n655,n656);
and (n718,n588,n696);
and (n719,n720,n721);
xor (n720,n717,n718);
or (n721,n722,n725);
and (n722,n723,n724);
xor (n723,n661,n662);
and (n724,n595,n696);
and (n725,n726,n727);
xor (n726,n723,n724);
or (n727,n728,n731);
and (n728,n729,n730);
xor (n729,n667,n668);
and (n730,n602,n696);
and (n731,n732,n733);
xor (n732,n729,n730);
or (n733,n734,n737);
and (n734,n735,n736);
xor (n735,n673,n674);
and (n736,n609,n696);
and (n737,n738,n739);
xor (n738,n735,n736);
or (n739,n740,n743);
and (n740,n741,n742);
xor (n741,n679,n680);
and (n742,n616,n696);
and (n743,n744,n745);
xor (n744,n741,n742);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n685,n686);
and (n748,n623,n696);
and (n749,n750,n751);
xor (n750,n747,n748);
and (n751,n752,n753);
xor (n752,n691,n692);
and (n753,n629,n696);
and (n754,n567,n755);
buf (n755,n259);
or (n756,n757,n760);
and (n757,n758,n759);
xor (n758,n702,n703);
and (n759,n574,n755);
and (n760,n761,n762);
xor (n761,n758,n759);
or (n762,n763,n766);
and (n763,n764,n765);
xor (n764,n708,n709);
and (n765,n581,n755);
and (n766,n767,n768);
xor (n767,n764,n765);
or (n768,n769,n772);
and (n769,n770,n771);
xor (n770,n714,n715);
and (n771,n588,n755);
and (n772,n773,n774);
xor (n773,n770,n771);
or (n774,n775,n778);
and (n775,n776,n777);
xor (n776,n720,n721);
and (n777,n595,n755);
and (n778,n779,n780);
xor (n779,n776,n777);
or (n780,n781,n784);
and (n781,n782,n783);
xor (n782,n726,n727);
and (n783,n602,n755);
and (n784,n785,n786);
xor (n785,n782,n783);
or (n786,n787,n790);
and (n787,n788,n789);
xor (n788,n732,n733);
and (n789,n609,n755);
and (n790,n791,n792);
xor (n791,n788,n789);
or (n792,n793,n796);
and (n793,n794,n795);
xor (n794,n738,n739);
and (n795,n616,n755);
and (n796,n797,n798);
xor (n797,n794,n795);
or (n798,n799,n802);
and (n799,n800,n801);
xor (n800,n744,n745);
and (n801,n623,n755);
and (n802,n803,n804);
xor (n803,n800,n801);
and (n804,n805,n806);
xor (n805,n750,n751);
and (n806,n629,n755);
and (n807,n574,n808);
buf (n808,n314);
or (n809,n810,n813);
and (n810,n811,n812);
xor (n811,n761,n762);
and (n812,n581,n808);
and (n813,n814,n815);
xor (n814,n811,n812);
or (n815,n816,n819);
and (n816,n817,n818);
xor (n817,n767,n768);
and (n818,n588,n808);
and (n819,n820,n821);
xor (n820,n817,n818);
or (n821,n822,n825);
and (n822,n823,n824);
xor (n823,n773,n774);
and (n824,n595,n808);
and (n825,n826,n827);
xor (n826,n823,n824);
or (n827,n828,n831);
and (n828,n829,n830);
xor (n829,n779,n780);
and (n830,n602,n808);
and (n831,n832,n833);
xor (n832,n829,n830);
or (n833,n834,n837);
and (n834,n835,n836);
xor (n835,n785,n786);
and (n836,n609,n808);
and (n837,n838,n839);
xor (n838,n835,n836);
or (n839,n840,n843);
and (n840,n841,n842);
xor (n841,n791,n792);
and (n842,n616,n808);
and (n843,n844,n845);
xor (n844,n841,n842);
or (n845,n846,n849);
and (n846,n847,n848);
xor (n847,n797,n798);
and (n848,n623,n808);
and (n849,n850,n851);
xor (n850,n847,n848);
and (n851,n852,n853);
xor (n852,n803,n804);
and (n853,n629,n808);
and (n854,n581,n855);
buf (n855,n363);
or (n856,n857,n860);
and (n857,n858,n859);
xor (n858,n814,n815);
and (n859,n588,n855);
and (n860,n861,n862);
xor (n861,n858,n859);
or (n862,n863,n866);
and (n863,n864,n865);
xor (n864,n820,n821);
and (n865,n595,n855);
and (n866,n867,n868);
xor (n867,n864,n865);
or (n868,n869,n872);
and (n869,n870,n871);
xor (n870,n826,n827);
and (n871,n602,n855);
and (n872,n873,n874);
xor (n873,n870,n871);
or (n874,n875,n878);
and (n875,n876,n877);
xor (n876,n832,n833);
and (n877,n609,n855);
and (n878,n879,n880);
xor (n879,n876,n877);
or (n880,n881,n884);
and (n881,n882,n883);
xor (n882,n838,n839);
and (n883,n616,n855);
and (n884,n885,n886);
xor (n885,n882,n883);
or (n886,n887,n890);
and (n887,n888,n889);
xor (n888,n844,n845);
and (n889,n623,n855);
and (n890,n891,n892);
xor (n891,n888,n889);
and (n892,n893,n894);
xor (n893,n850,n851);
and (n894,n629,n855);
and (n895,n588,n896);
buf (n896,n406);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n861,n862);
and (n900,n595,n896);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n867,n868);
and (n906,n602,n896);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n873,n874);
and (n912,n609,n896);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
xor (n917,n879,n880);
and (n918,n616,n896);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n925);
and (n922,n923,n924);
xor (n923,n885,n886);
and (n924,n623,n896);
and (n925,n926,n927);
xor (n926,n923,n924);
and (n927,n928,n929);
xor (n928,n891,n892);
and (n929,n629,n896);
and (n930,n595,n931);
buf (n931,n443);
or (n932,n933,n936);
and (n933,n934,n935);
xor (n934,n902,n903);
and (n935,n602,n931);
and (n936,n937,n938);
xor (n937,n934,n935);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n908,n909);
and (n941,n609,n931);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n914,n915);
and (n947,n616,n931);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n920,n921);
and (n953,n623,n931);
and (n954,n955,n956);
xor (n955,n952,n953);
and (n956,n957,n958);
xor (n957,n926,n927);
and (n958,n629,n931);
and (n959,n602,n960);
buf (n960,n474);
or (n961,n962,n965);
and (n962,n963,n964);
xor (n963,n937,n938);
and (n964,n609,n960);
and (n965,n966,n967);
xor (n966,n963,n964);
or (n967,n968,n971);
and (n968,n969,n970);
xor (n969,n943,n944);
and (n970,n616,n960);
and (n971,n972,n973);
xor (n972,n969,n970);
or (n973,n974,n977);
and (n974,n975,n976);
xor (n975,n949,n950);
and (n976,n623,n960);
and (n977,n978,n979);
xor (n978,n975,n976);
and (n979,n980,n981);
xor (n980,n955,n956);
and (n981,n629,n960);
and (n982,n609,n983);
buf (n983,n499);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n966,n967);
and (n987,n616,n983);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n972,n973);
and (n993,n623,n983);
and (n994,n995,n996);
xor (n995,n992,n993);
and (n996,n997,n998);
xor (n997,n978,n979);
and (n998,n629,n983);
and (n999,n616,n1000);
buf (n1000,n518);
or (n1001,n1002,n1005);
and (n1002,n1003,n1004);
xor (n1003,n989,n990);
and (n1004,n623,n1000);
and (n1005,n1006,n1007);
xor (n1006,n1003,n1004);
and (n1007,n1008,n1009);
xor (n1008,n995,n996);
and (n1009,n629,n1000);
buf (n1010,n1011);
xor (n1011,n1012,n1481);
xor (n1012,n1013,n1479);
xor (n1013,n1014,n1464);
xor (n1014,n1015,n1462);
xor (n1015,n1016,n1441);
xor (n1016,n1017,n1439);
xor (n1017,n1018,n1412);
xor (n1018,n1019,n1410);
xor (n1019,n1020,n1377);
xor (n1020,n1021,n1375);
xor (n1021,n1022,n1336);
xor (n1022,n1023,n1334);
xor (n1023,n1024,n1289);
xor (n1024,n1025,n1287);
xor (n1025,n1026,n1236);
xor (n1026,n1027,n1234);
xor (n1027,n1028,n1177);
xor (n1028,n1029,n1175);
xor (n1029,n1030,n1112);
xor (n1030,n1031,n1110);
and (n1031,n1032,n1035);
and (n1032,n1033,n1034);
buf (n1033,n25);
buf (n1034,n29);
or (n1035,n1036,n1041);
and (n1036,n1037,n1039);
and (n1037,n1033,n1038);
buf (n1038,n35);
and (n1039,n1040,n1034);
buf (n1040,n39);
and (n1041,n1042,n1043);
xor (n1042,n1037,n1039);
or (n1043,n1044,n1048);
and (n1044,n1045,n1046);
and (n1045,n1040,n1038);
and (n1046,n1047,n1034);
buf (n1047,n48);
and (n1048,n1049,n1050);
xor (n1049,n1045,n1046);
or (n1050,n1051,n1055);
and (n1051,n1052,n1053);
and (n1052,n1047,n1038);
and (n1053,n1054,n1034);
buf (n1054,n57);
and (n1055,n1056,n1057);
xor (n1056,n1052,n1053);
or (n1057,n1058,n1062);
and (n1058,n1059,n1060);
and (n1059,n1054,n1038);
and (n1060,n1061,n1034);
buf (n1061,n66);
and (n1062,n1063,n1064);
xor (n1063,n1059,n1060);
or (n1064,n1065,n1069);
and (n1065,n1066,n1067);
and (n1066,n1061,n1038);
and (n1067,n1068,n1034);
buf (n1068,n75);
and (n1069,n1070,n1071);
xor (n1070,n1066,n1067);
or (n1071,n1072,n1076);
and (n1072,n1073,n1074);
and (n1073,n1068,n1038);
and (n1074,n1075,n1034);
buf (n1075,n84);
and (n1076,n1077,n1078);
xor (n1077,n1073,n1074);
or (n1078,n1079,n1083);
and (n1079,n1080,n1081);
and (n1080,n1075,n1038);
and (n1081,n1082,n1034);
buf (n1082,n93);
and (n1083,n1084,n1085);
xor (n1084,n1080,n1081);
or (n1085,n1086,n1090);
and (n1086,n1087,n1088);
and (n1087,n1082,n1038);
and (n1088,n1089,n1034);
buf (n1089,n102);
and (n1090,n1091,n1092);
xor (n1091,n1087,n1088);
or (n1092,n1093,n1097);
and (n1093,n1094,n1095);
and (n1094,n1089,n1038);
and (n1095,n1096,n1034);
buf (n1096,n111);
and (n1097,n1098,n1099);
xor (n1098,n1094,n1095);
or (n1099,n1100,n1104);
and (n1100,n1101,n1102);
and (n1101,n1096,n1038);
and (n1102,n1103,n1034);
buf (n1103,n120);
and (n1104,n1105,n1106);
xor (n1105,n1101,n1102);
and (n1106,n1107,n1108);
and (n1107,n1103,n1038);
and (n1108,n1109,n1034);
buf (n1109,n128);
and (n1110,n1033,n1111);
buf (n1111,n132);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1032,n1035);
and (n1115,n1040,n1111);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1042,n1043);
and (n1121,n1047,n1111);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1049,n1050);
and (n1127,n1054,n1111);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1056,n1057);
and (n1133,n1061,n1111);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1063,n1064);
and (n1139,n1068,n1111);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1070,n1071);
and (n1145,n1075,n1111);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1077,n1078);
and (n1151,n1082,n1111);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1084,n1085);
and (n1157,n1089,n1111);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1091,n1092);
and (n1163,n1096,n1111);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1098,n1099);
and (n1169,n1103,n1111);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
and (n1172,n1173,n1174);
xor (n1173,n1105,n1106);
and (n1174,n1109,n1111);
and (n1175,n1040,n1176);
buf (n1176,n199);
or (n1177,n1178,n1181);
and (n1178,n1179,n1180);
xor (n1179,n1117,n1118);
and (n1180,n1047,n1176);
and (n1181,n1182,n1183);
xor (n1182,n1179,n1180);
or (n1183,n1184,n1187);
and (n1184,n1185,n1186);
xor (n1185,n1123,n1124);
and (n1186,n1054,n1176);
and (n1187,n1188,n1189);
xor (n1188,n1185,n1186);
or (n1189,n1190,n1193);
and (n1190,n1191,n1192);
xor (n1191,n1129,n1130);
and (n1192,n1061,n1176);
and (n1193,n1194,n1195);
xor (n1194,n1191,n1192);
or (n1195,n1196,n1199);
and (n1196,n1197,n1198);
xor (n1197,n1135,n1136);
and (n1198,n1068,n1176);
and (n1199,n1200,n1201);
xor (n1200,n1197,n1198);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1141,n1142);
and (n1204,n1075,n1176);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1147,n1148);
and (n1210,n1082,n1176);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1153,n1154);
and (n1216,n1089,n1176);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1159,n1160);
and (n1222,n1096,n1176);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1165,n1166);
and (n1228,n1103,n1176);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
and (n1231,n1232,n1233);
xor (n1232,n1171,n1172);
and (n1233,n1109,n1176);
and (n1234,n1047,n1235);
buf (n1235,n260);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1182,n1183);
and (n1239,n1054,n1235);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1246);
and (n1243,n1244,n1245);
xor (n1244,n1188,n1189);
and (n1245,n1061,n1235);
and (n1246,n1247,n1248);
xor (n1247,n1244,n1245);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1194,n1195);
and (n1251,n1068,n1235);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1200,n1201);
and (n1257,n1075,n1235);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1206,n1207);
and (n1263,n1082,n1235);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
or (n1266,n1267,n1270);
and (n1267,n1268,n1269);
xor (n1268,n1212,n1213);
and (n1269,n1089,n1235);
and (n1270,n1271,n1272);
xor (n1271,n1268,n1269);
or (n1272,n1273,n1276);
and (n1273,n1274,n1275);
xor (n1274,n1218,n1219);
and (n1275,n1096,n1235);
and (n1276,n1277,n1278);
xor (n1277,n1274,n1275);
or (n1278,n1279,n1282);
and (n1279,n1280,n1281);
xor (n1280,n1224,n1225);
and (n1281,n1103,n1235);
and (n1282,n1283,n1284);
xor (n1283,n1280,n1281);
and (n1284,n1285,n1286);
xor (n1285,n1230,n1231);
and (n1286,n1109,n1235);
and (n1287,n1054,n1288);
buf (n1288,n315);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1241,n1242);
and (n1292,n1061,n1288);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1247,n1248);
and (n1298,n1068,n1288);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1253,n1254);
and (n1304,n1075,n1288);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1259,n1260);
and (n1310,n1082,n1288);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1265,n1266);
and (n1316,n1089,n1288);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1271,n1272);
and (n1322,n1096,n1288);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
or (n1325,n1326,n1329);
and (n1326,n1327,n1328);
xor (n1327,n1277,n1278);
and (n1328,n1103,n1288);
and (n1329,n1330,n1331);
xor (n1330,n1327,n1328);
and (n1331,n1332,n1333);
xor (n1332,n1283,n1284);
and (n1333,n1109,n1288);
and (n1334,n1061,n1335);
buf (n1335,n364);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1294,n1295);
and (n1339,n1068,n1335);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1300,n1301);
and (n1345,n1075,n1335);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
or (n1348,n1349,n1352);
and (n1349,n1350,n1351);
xor (n1350,n1306,n1307);
and (n1351,n1082,n1335);
and (n1352,n1353,n1354);
xor (n1353,n1350,n1351);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1312,n1313);
and (n1357,n1089,n1335);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1318,n1319);
and (n1363,n1096,n1335);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1324,n1325);
and (n1369,n1103,n1335);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
and (n1372,n1373,n1374);
xor (n1373,n1330,n1331);
and (n1374,n1109,n1335);
and (n1375,n1068,n1376);
buf (n1376,n407);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1341,n1342);
and (n1380,n1075,n1376);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1347,n1348);
and (n1386,n1082,n1376);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1353,n1354);
and (n1392,n1089,n1376);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1359,n1360);
and (n1398,n1096,n1376);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
or (n1401,n1402,n1405);
and (n1402,n1403,n1404);
xor (n1403,n1365,n1366);
and (n1404,n1103,n1376);
and (n1405,n1406,n1407);
xor (n1406,n1403,n1404);
and (n1407,n1408,n1409);
xor (n1408,n1371,n1372);
and (n1409,n1109,n1376);
and (n1410,n1075,n1411);
buf (n1411,n444);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1382,n1383);
and (n1415,n1082,n1411);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1388,n1389);
and (n1421,n1089,n1411);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1394,n1395);
and (n1427,n1096,n1411);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1400,n1401);
and (n1433,n1103,n1411);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
and (n1436,n1437,n1438);
xor (n1437,n1406,n1407);
and (n1438,n1109,n1411);
and (n1439,n1082,n1440);
buf (n1440,n475);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1417,n1418);
and (n1444,n1089,n1440);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1423,n1424);
and (n1450,n1096,n1440);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1429,n1430);
and (n1456,n1103,n1440);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
and (n1459,n1460,n1461);
xor (n1460,n1435,n1436);
and (n1461,n1109,n1440);
and (n1462,n1089,n1463);
buf (n1463,n500);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1446,n1447);
and (n1467,n1096,n1463);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
or (n1470,n1471,n1474);
and (n1471,n1472,n1473);
xor (n1472,n1452,n1453);
and (n1473,n1103,n1463);
and (n1474,n1475,n1476);
xor (n1475,n1472,n1473);
and (n1476,n1477,n1478);
xor (n1477,n1458,n1459);
and (n1478,n1109,n1463);
and (n1479,n1096,n1480);
buf (n1480,n519);
or (n1481,n1482,n1485);
and (n1482,n1483,n1484);
xor (n1483,n1469,n1470);
and (n1484,n1103,n1480);
and (n1485,n1486,n1487);
xor (n1486,n1483,n1484);
and (n1487,n1488,n1489);
xor (n1488,n1475,n1476);
and (n1489,n1109,n1480);
endmodule
