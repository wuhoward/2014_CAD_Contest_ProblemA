module top (out,n18,n23,n24,n25,n27,n28,n39,n42,n45
        ,n48,n51,n54,n57,n60,n63,n66,n69,n72,n75
        ,n78,n81,n84,n87,n90,n92,n95,n98,n108,n118
        ,n125,n130,n165,n170,n173,n176,n179,n182,n185,n188
        ,n191,n194,n197,n200,n203,n206,n209,n212,n215,n224
        ,n492,n543,n865,n913);
output out;
input n18;
input n23;
input n24;
input n25;
input n27;
input n28;
input n39;
input n42;
input n45;
input n48;
input n51;
input n54;
input n57;
input n60;
input n63;
input n66;
input n69;
input n72;
input n75;
input n78;
input n81;
input n84;
input n87;
input n90;
input n92;
input n95;
input n98;
input n108;
input n118;
input n125;
input n130;
input n165;
input n170;
input n173;
input n176;
input n179;
input n182;
input n185;
input n188;
input n191;
input n194;
input n197;
input n200;
input n203;
input n206;
input n209;
input n212;
input n215;
input n224;
input n492;
input n543;
input n865;
input n913;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n22;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n43;
wire n44;
wire n46;
wire n47;
wire n49;
wire n50;
wire n52;
wire n53;
wire n55;
wire n56;
wire n58;
wire n59;
wire n61;
wire n62;
wire n64;
wire n65;
wire n67;
wire n68;
wire n70;
wire n71;
wire n73;
wire n74;
wire n76;
wire n77;
wire n79;
wire n80;
wire n82;
wire n83;
wire n85;
wire n86;
wire n88;
wire n89;
wire n91;
wire n93;
wire n94;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n174;
wire n175;
wire n177;
wire n178;
wire n180;
wire n181;
wire n183;
wire n184;
wire n186;
wire n187;
wire n189;
wire n190;
wire n192;
wire n193;
wire n195;
wire n196;
wire n198;
wire n199;
wire n201;
wire n202;
wire n204;
wire n205;
wire n207;
wire n208;
wire n210;
wire n211;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
xor (out,n0,n1909);
xor (n0,n1,n959);
xor (n1,n2,n830);
or (n2,n3,n829);
and (n3,n4,n744);
xor (n4,n5,n555);
xor (n5,n6,n473);
xor (n6,n7,n336);
xor (n7,n8,n230);
xor (n8,n9,n133);
nand (n9,n10,n120);
or (n10,n11,n114);
nand (n11,n12,n104);
nor (n12,n13,n102);
and (n13,n14,n96);
not (n14,n15);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n93);
and (s0n15,notn15,n16);
and (s1n15,n93,n35);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n19);
and (s0n16,notn16,1'b0);
and (s1n16,n19,n18);
or (n19,n20,n31);
or (n20,n21,n29);
nor (n21,n22,n24,n25,n26,n28);
not (n22,n23);
not (n26,n27);
nor (n29,n23,n30,n25,n26,n28);
not (n30,n24);
or (n31,n32,n34);
and (n32,n22,n24,n25,n26,n33);
not (n33,n28);
nor (n34,n22,n30,n25,n26,n28);
xor (n35,n36,n37);
not (n36,n18);
and (n37,n38,n40);
not (n38,n39);
and (n40,n41,n43);
not (n41,n42);
and (n43,n44,n46);
not (n44,n45);
and (n46,n47,n49);
not (n47,n48);
and (n49,n50,n52);
not (n50,n51);
and (n52,n53,n55);
not (n53,n54);
and (n55,n56,n58);
not (n56,n57);
and (n58,n59,n61);
not (n59,n60);
and (n61,n62,n64);
not (n62,n63);
and (n64,n65,n67);
not (n65,n66);
and (n67,n68,n70);
not (n68,n69);
and (n70,n71,n73);
not (n71,n72);
and (n73,n74,n76);
not (n74,n75);
and (n76,n77,n79);
not (n77,n78);
and (n79,n80,n82);
not (n80,n81);
and (n82,n83,n85);
not (n83,n84);
and (n85,n86,n88);
not (n86,n87);
and (n88,n89,n91);
not (n89,n90);
not (n91,n92);
and (n93,n94,n95);
or (n94,n21,n32);
wire s0n96,s1n96,notn96;
or (n96,s0n96,s1n96);
not(notn96,n93);
and (s0n96,notn96,n97);
and (s1n96,n93,n99);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n19);
and (s0n97,notn97,1'b0);
and (s1n97,n19,n98);
xor (n99,n100,n101);
not (n100,n98);
and (n101,n36,n37);
and (n102,n15,n103);
not (n103,n96);
nand (n104,n105,n112);
or (n105,n103,n106);
wire s0n106,s1n106,notn106;
or (n106,s0n106,s1n106);
not(notn106,n93);
and (s0n106,notn106,n107);
and (s1n106,n93,n109);
wire s0n107,s1n107,notn107;
or (n107,s0n107,s1n107);
not(notn107,n19);
and (s0n107,notn107,1'b0);
and (s1n107,n19,n108);
xor (n109,n110,n111);
not (n110,n108);
and (n111,n100,n101);
or (n112,n96,n113);
not (n113,n106);
nor (n114,n115,n119);
and (n115,n106,n116);
not (n116,n117);
wire s0n117,s1n117,notn117;
or (n117,s0n117,s1n117);
not(notn117,n19);
and (s0n117,notn117,1'b0);
and (s1n117,n19,n118);
and (n119,n113,n117);
or (n120,n12,n121);
nor (n121,n122,n131);
and (n122,n123,n113);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n129);
and (s0n123,notn123,n124);
and (s1n123,n129,n126);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n19);
and (s0n124,notn124,1'b0);
and (s1n124,n19,n125);
xor (n126,n127,n128);
not (n127,n125);
not (n128,n118);
and (n129,n94,n130);
and (n131,n132,n106);
not (n132,n123);
xor (n133,n134,n140);
nor (n134,n135,n113);
nor (n135,n136,n139);
and (n136,n137,n14);
not (n137,n138);
and (n138,n117,n96);
and (n139,n103,n116);
nand (n140,n141,n219);
or (n141,n142,n161);
nand (n142,n143,n154);
nor (n143,n144,n152);
and (n144,n145,n149);
not (n145,n146);
wire s0n146,s1n146,notn146;
or (n146,s0n146,s1n146);
not(notn146,n93);
and (s0n146,notn146,n147);
and (s1n146,n93,n148);
wire s0n147,s1n147,notn147;
or (n147,s0n147,s1n147);
not(notn147,n19);
and (s0n147,notn147,1'b0);
and (s1n147,n19,n90);
xor (n148,n89,n91);
wire s0n149,s1n149,notn149;
or (n149,s0n149,s1n149);
not(notn149,n93);
and (s0n149,notn149,n150);
and (s1n149,n93,n151);
wire s0n150,s1n150,notn150;
or (n150,s0n150,s1n150);
not(notn150,n19);
and (s0n150,notn150,1'b0);
and (s1n150,n19,n87);
xor (n151,n86,n88);
and (n152,n146,n153);
not (n153,n149);
nand (n154,n155,n160);
or (n155,n156,n149);
not (n156,n157);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n93);
and (s0n157,notn157,n158);
and (s1n157,n93,n159);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n19);
and (s0n158,notn158,1'b0);
and (s1n158,n19,n84);
xor (n159,n83,n85);
nand (n160,n156,n149);
nor (n161,n162,n217);
and (n162,n163,n156);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n129);
and (s0n163,notn163,n164);
and (s1n163,n129,n166);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n19);
and (s0n164,notn164,1'b0);
and (s1n164,n19,n165);
xor (n166,n167,n168);
not (n167,n165);
and (n168,n169,n171);
not (n169,n170);
and (n171,n172,n174);
not (n172,n173);
and (n174,n175,n177);
not (n175,n176);
and (n177,n178,n180);
not (n178,n179);
and (n180,n181,n183);
not (n181,n182);
and (n183,n184,n186);
not (n184,n185);
and (n186,n187,n189);
not (n187,n188);
and (n189,n190,n192);
not (n190,n191);
and (n192,n193,n195);
not (n193,n194);
and (n195,n196,n198);
not (n196,n197);
and (n198,n199,n201);
not (n199,n200);
and (n201,n202,n204);
not (n202,n203);
and (n204,n205,n207);
not (n205,n206);
and (n207,n208,n210);
not (n208,n209);
and (n210,n211,n213);
not (n211,n212);
and (n213,n214,n216);
not (n214,n215);
and (n216,n127,n128);
and (n217,n218,n157);
not (n218,n163);
or (n219,n143,n220);
nor (n220,n221,n228);
and (n221,n222,n156);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n129);
and (s0n222,notn222,n223);
and (s1n222,n129,n225);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n19);
and (s0n223,notn223,1'b0);
and (s1n223,n19,n224);
xor (n225,n226,n227);
not (n226,n224);
and (n227,n167,n168);
and (n228,n229,n157);
not (n229,n222);
or (n230,n231,n335);
and (n231,n232,n303);
xor (n232,n233,n270);
nand (n233,n234,n262);
or (n234,n235,n255);
nand (n235,n236,n247);
nor (n236,n237,n244);
and (n237,n238,n241);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n93);
and (s0n238,notn238,n239);
and (s1n238,n93,n240);
wire s0n239,s1n239,notn239;
or (n239,s0n239,s1n239);
not(notn239,n19);
and (s0n239,notn239,1'b0);
and (s1n239,n19,n69);
xor (n240,n68,n70);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n93);
and (s0n241,notn241,n242);
and (s1n241,n93,n243);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n19);
and (s0n242,notn242,1'b0);
and (s1n242,n19,n66);
xor (n243,n65,n67);
and (n244,n245,n246);
not (n245,n238);
not (n246,n241);
not (n247,n248);
nor (n248,n249,n253);
and (n249,n250,n238);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n93);
and (s0n250,notn250,n251);
and (s1n250,n93,n252);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n19);
and (s0n251,notn251,1'b0);
and (s1n251,n19,n72);
xor (n252,n71,n73);
and (n253,n254,n245);
not (n254,n250);
nor (n255,n256,n260);
and (n256,n246,n257);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n129);
and (s0n257,notn257,n258);
and (s1n257,n129,n259);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n19);
and (s0n258,notn258,1'b0);
and (s1n258,n19,n188);
xor (n259,n187,n189);
and (n260,n241,n261);
not (n261,n257);
or (n262,n263,n247);
nor (n263,n264,n268);
and (n264,n246,n265);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n129);
and (s0n265,notn265,n266);
and (s1n265,n129,n267);
wire s0n266,s1n266,notn266;
or (n266,s0n266,s1n266);
not(notn266,n19);
and (s0n266,notn266,1'b0);
and (s1n266,n19,n185);
xor (n267,n184,n186);
and (n268,n241,n269);
not (n269,n265);
nand (n270,n271,n295);
or (n271,n272,n288);
nand (n272,n273,n280);
not (n273,n274);
nand (n274,n275,n279);
or (n275,n156,n276);
wire s0n276,s1n276,notn276;
or (n276,s0n276,s1n276);
not(notn276,n93);
and (s0n276,notn276,n277);
and (s1n276,n93,n278);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n19);
and (s0n277,notn277,1'b0);
and (s1n277,n19,n81);
xor (n278,n80,n82);
nand (n279,n276,n156);
nor (n280,n281,n287);
and (n281,n282,n286);
not (n282,n283);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n93);
and (s0n283,notn283,n284);
and (s1n283,n93,n285);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n19);
and (s0n284,notn284,1'b0);
and (s1n284,n19,n78);
xor (n285,n77,n79);
not (n286,n276);
and (n287,n283,n276);
nor (n288,n289,n293);
and (n289,n290,n282);
wire s0n290,s1n290,notn290;
or (n290,s0n290,s1n290);
not(notn290,n129);
and (s0n290,notn290,n291);
and (s1n290,n129,n292);
wire s0n291,s1n291,notn291;
or (n291,s0n291,s1n291);
not(notn291,n19);
and (s0n291,notn291,1'b0);
and (s1n291,n19,n176);
xor (n292,n175,n177);
and (n293,n294,n283);
not (n294,n290);
or (n295,n273,n296);
nor (n296,n297,n301);
and (n297,n298,n282);
wire s0n298,s1n298,notn298;
or (n298,s0n298,s1n298);
not(notn298,n129);
and (s0n298,notn298,n299);
and (s1n298,n129,n300);
wire s0n299,s1n299,notn299;
or (n299,s0n299,s1n299);
not(notn299,n19);
and (s0n299,notn299,1'b0);
and (s1n299,n19,n173);
xor (n300,n172,n174);
and (n301,n302,n283);
not (n302,n298);
nand (n303,n304,n327);
or (n304,n305,n320);
nand (n305,n306,n313);
or (n306,n307,n311);
and (n307,n308,n241);
wire s0n308,s1n308,notn308;
or (n308,s0n308,s1n308);
not(notn308,n93);
and (s0n308,notn308,n309);
and (s1n308,n93,n310);
wire s0n309,s1n309,notn309;
or (n309,s0n309,s1n309);
not(notn309,n19);
and (s0n309,notn309,1'b0);
and (s1n309,n19,n63);
xor (n310,n62,n64);
and (n311,n312,n246);
not (n312,n308);
nand (n313,n314,n318);
or (n314,n312,n315);
wire s0n315,s1n315,notn315;
or (n315,s0n315,s1n315);
not(notn315,n93);
and (s0n315,notn315,n316);
and (s1n315,n93,n317);
wire s0n316,s1n316,notn316;
or (n316,s0n316,s1n316);
not(notn316,n19);
and (s0n316,notn316,1'b0);
and (s1n316,n19,n60);
xor (n317,n59,n61);
or (n318,n319,n308);
not (n319,n315);
nor (n320,n321,n325);
and (n321,n319,n322);
wire s0n322,s1n322,notn322;
or (n322,s0n322,s1n322);
not(notn322,n129);
and (s0n322,notn322,n323);
and (s1n322,n129,n324);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n19);
and (s0n323,notn323,1'b0);
and (s1n323,n19,n194);
xor (n324,n193,n195);
and (n325,n315,n326);
not (n326,n322);
or (n327,n306,n328);
nor (n328,n329,n333);
and (n329,n319,n330);
wire s0n330,s1n330,notn330;
or (n330,s0n330,s1n330);
not(notn330,n129);
and (s0n330,notn330,n331);
and (s1n330,n129,n332);
wire s0n331,s1n331,notn331;
or (n331,s0n331,s1n331);
not(notn331,n19);
and (s0n331,notn331,1'b0);
and (s1n331,n19,n191);
xor (n332,n190,n192);
and (n333,n315,n334);
not (n334,n330);
and (n335,n233,n270);
or (n336,n337,n472);
and (n337,n338,n471);
xor (n338,n339,n438);
or (n339,n340,n437);
and (n340,n341,n404);
xor (n341,n342,n366);
nand (n342,n343,n358);
or (n343,n344,n355);
nand (n344,n345,n352);
or (n345,n346,n350);
and (n346,n283,n347);
wire s0n347,s1n347,notn347;
or (n347,s0n347,s1n347);
not(notn347,n93);
and (s0n347,notn347,n348);
and (s1n347,n93,n349);
wire s0n348,s1n348,notn348;
or (n348,s0n348,s1n348);
not(notn348,n19);
and (s0n348,notn348,1'b0);
and (s1n348,n19,n75);
xor (n349,n74,n76);
and (n350,n282,n351);
not (n351,n347);
nor (n352,n353,n354);
and (n353,n250,n347);
and (n354,n254,n351);
nor (n355,n356,n357);
and (n356,n265,n254);
and (n357,n269,n250);
or (n358,n345,n359);
nor (n359,n360,n364);
and (n360,n361,n254);
wire s0n361,s1n361,notn361;
or (n361,s0n361,s1n361);
not(notn361,n129);
and (s0n361,notn361,n362);
and (s1n361,n129,n363);
wire s0n362,s1n362,notn362;
or (n362,s0n362,s1n362);
not(notn362,n19);
and (s0n362,notn362,1'b0);
and (s1n362,n19,n182);
xor (n363,n181,n183);
and (n364,n365,n250);
not (n365,n361);
nand (n366,n367,n395);
or (n367,n368,n388);
not (n368,n369);
nor (n369,n370,n380);
nand (n370,n371,n379);
or (n371,n372,n376);
not (n372,n373);
wire s0n373,s1n373,notn373;
or (n373,s0n373,s1n373);
not(notn373,n93);
and (s0n373,notn373,n374);
and (s1n373,n93,n375);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n19);
and (s0n374,notn374,1'b0);
and (s1n374,n19,n54);
xor (n375,n53,n55);
wire s0n376,s1n376,notn376;
or (n376,s0n376,s1n376);
not(notn376,n93);
and (s0n376,notn376,n377);
and (s1n376,n93,n378);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n19);
and (s0n377,notn377,1'b0);
and (s1n377,n19,n51);
xor (n378,n50,n52);
nand (n379,n372,n376);
nor (n380,n381,n386);
and (n381,n382,n376);
not (n382,n383);
wire s0n383,s1n383,notn383;
or (n383,s0n383,s1n383);
not(notn383,n93);
and (s0n383,notn383,n384);
and (s1n383,n93,n385);
wire s0n384,s1n384,notn384;
or (n384,s0n384,s1n384);
not(notn384,n19);
and (s0n384,notn384,1'b0);
and (s1n384,n19,n48);
xor (n385,n47,n49);
and (n386,n387,n383);
not (n387,n376);
nor (n388,n389,n393);
and (n389,n382,n390);
wire s0n390,s1n390,notn390;
or (n390,s0n390,s1n390);
not(notn390,n129);
and (s0n390,notn390,n391);
and (s1n390,n129,n392);
wire s0n391,s1n391,notn391;
or (n391,s0n391,s1n391);
not(notn391,n19);
and (s0n391,notn391,1'b0);
and (s1n391,n19,n209);
xor (n392,n208,n210);
and (n393,n394,n383);
not (n394,n390);
or (n395,n396,n397);
not (n396,n370);
nor (n397,n398,n402);
and (n398,n399,n382);
wire s0n399,s1n399,notn399;
or (n399,s0n399,s1n399);
not(notn399,n129);
and (s0n399,notn399,n400);
and (s1n399,n129,n401);
wire s0n400,s1n400,notn400;
or (n400,s0n400,s1n400);
not(notn400,n19);
and (s0n400,notn400,1'b0);
and (s1n400,n19,n206);
xor (n401,n205,n207);
and (n402,n403,n383);
not (n403,n399);
nand (n404,n405,n429);
or (n405,n406,n422);
not (n406,n407);
and (n407,n408,n415);
nor (n408,n409,n414);
and (n409,n383,n410);
not (n410,n411);
wire s0n411,s1n411,notn411;
or (n411,s0n411,s1n411);
not(notn411,n93);
and (s0n411,notn411,n412);
and (s1n411,n93,n413);
wire s0n412,s1n412,notn412;
or (n412,s0n412,s1n412);
not(notn412,n19);
and (s0n412,notn412,1'b0);
and (s1n412,n19,n45);
xor (n413,n44,n46);
and (n414,n382,n411);
nand (n415,n416,n420);
or (n416,n410,n417);
wire s0n417,s1n417,notn417;
or (n417,s0n417,s1n417);
not(notn417,n93);
and (s0n417,notn417,n418);
and (s1n417,n93,n419);
wire s0n418,s1n418,notn418;
or (n418,s0n418,s1n418);
not(notn418,n19);
and (s0n418,notn418,1'b0);
and (s1n418,n19,n42);
xor (n419,n41,n43);
or (n420,n421,n411);
not (n421,n417);
nor (n422,n423,n427);
and (n423,n424,n421);
wire s0n424,s1n424,notn424;
or (n424,s0n424,s1n424);
not(notn424,n129);
and (s0n424,notn424,n425);
and (s1n424,n129,n426);
wire s0n425,s1n425,notn425;
or (n425,s0n425,s1n425);
not(notn425,n19);
and (s0n425,notn425,1'b0);
and (s1n425,n19,n215);
xor (n426,n214,n216);
and (n427,n428,n417);
not (n428,n424);
or (n429,n430,n408);
nor (n430,n431,n435);
and (n431,n432,n421);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n129);
and (s0n432,notn432,n433);
and (s1n432,n129,n434);
wire s0n433,s1n433,notn433;
or (n433,s0n433,s1n433);
not(notn433,n19);
and (s0n433,notn433,1'b0);
and (s1n433,n19,n212);
xor (n434,n211,n213);
and (n435,n436,n417);
not (n436,n432);
and (n437,n342,n366);
or (n438,n439,n470);
and (n439,n440,n460);
xor (n440,n441,n454);
nand (n441,n442,n446);
or (n442,n142,n443);
nor (n443,n444,n445);
and (n444,n156,n298);
and (n445,n302,n157);
or (n446,n447,n143);
nor (n447,n448,n452);
and (n448,n449,n156);
wire s0n449,s1n449,notn449;
or (n449,s0n449,s1n449);
not(notn449,n129);
and (s0n449,notn449,n450);
and (s1n449,n129,n451);
wire s0n450,s1n450,notn450;
or (n450,s0n450,s1n450);
not(notn450,n19);
and (s0n450,notn450,1'b0);
and (s1n450,n19,n170);
xor (n451,n169,n171);
and (n452,n453,n157);
not (n453,n449);
nand (n454,n455,n459);
or (n455,n235,n456);
nor (n456,n457,n458);
and (n457,n246,n330);
and (n458,n241,n334);
or (n459,n255,n247);
nand (n460,n461,n469);
or (n461,n272,n462);
nor (n462,n463,n467);
and (n463,n464,n282);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n129);
and (s0n464,notn464,n465);
and (s1n464,n129,n466);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n19);
and (s0n465,notn465,1'b0);
and (s1n465,n19,n179);
xor (n466,n178,n180);
and (n467,n468,n283);
not (n468,n464);
or (n469,n273,n288);
and (n470,n441,n454);
xor (n471,n232,n303);
and (n472,n339,n438);
xor (n473,n474,n528);
xor (n474,n475,n505);
or (n475,n476,n504);
and (n476,n477,n498);
xor (n477,n478,n479);
nor (n478,n12,n116);
nand (n479,n480,n487);
or (n480,n481,n484);
nor (n481,n482,n483);
and (n482,n222,n145);
and (n483,n229,n146);
nand (n484,n146,n485);
not (n485,n486);
wire s0n486,s1n486,notn486;
or (n486,s0n486,s1n486);
not(notn486,n19);
and (s0n486,notn486,1'b0);
and (s1n486,n19,n92);
or (n487,n488,n485);
nor (n488,n489,n496);
and (n489,n490,n145);
wire s0n490,s1n490,notn490;
or (n490,s0n490,s1n490);
not(notn490,n129);
and (s0n490,notn490,n491);
and (s1n490,n129,n493);
wire s0n491,s1n491,notn491;
or (n491,s0n491,s1n491);
not(notn491,n19);
and (s0n491,notn491,1'b0);
and (s1n491,n19,n492);
xor (n493,n494,n495);
not (n494,n492);
and (n495,n226,n227);
and (n496,n497,n146);
not (n497,n490);
nand (n498,n499,n500);
or (n499,n344,n359);
or (n500,n345,n501);
nor (n501,n502,n503);
and (n502,n464,n254);
and (n503,n468,n250);
and (n504,n478,n479);
or (n505,n506,n527);
and (n506,n507,n524);
xor (n507,n508,n518);
nand (n508,n509,n510);
or (n509,n368,n397);
or (n510,n511,n396);
nor (n511,n512,n516);
and (n512,n382,n513);
wire s0n513,s1n513,notn513;
or (n513,s0n513,s1n513);
not(notn513,n129);
and (s0n513,notn513,n514);
and (s1n513,n129,n515);
wire s0n514,s1n514,notn514;
or (n514,s0n514,s1n514);
not(notn514,n19);
and (s0n514,notn514,1'b0);
and (s1n514,n19,n203);
xor (n515,n202,n204);
and (n516,n383,n517);
not (n517,n513);
nand (n518,n519,n520);
or (n519,n406,n430);
or (n520,n521,n408);
nor (n521,n522,n523);
and (n522,n421,n390);
and (n523,n417,n394);
nand (n524,n525,n526);
or (n525,n142,n447);
or (n526,n143,n161);
and (n527,n508,n518);
xor (n528,n529,n549);
xor (n529,n530,n536);
nand (n530,n531,n532);
or (n531,n235,n263);
or (n532,n533,n247);
nor (n533,n534,n535);
and (n534,n246,n361);
and (n535,n241,n365);
nand (n536,n537,n538);
or (n537,n488,n484);
or (n538,n539,n485);
nor (n539,n540,n547);
and (n540,n541,n145);
wire s0n541,s1n541,notn541;
or (n541,s0n541,s1n541);
not(notn541,n129);
and (s0n541,notn541,n542);
and (s1n541,n129,n544);
wire s0n542,s1n542,notn542;
or (n542,s0n542,s1n542);
not(notn542,n19);
and (s0n542,notn542,1'b0);
and (s1n542,n19,n543);
xor (n544,n545,n546);
not (n545,n543);
and (n546,n494,n495);
and (n547,n548,n146);
not (n548,n541);
nand (n549,n550,n551);
or (n550,n272,n296);
or (n551,n552,n273);
nor (n552,n553,n554);
and (n553,n449,n282);
and (n554,n453,n283);
xor (n555,n556,n694);
xor (n556,n557,n623);
or (n557,n558,n622);
and (n558,n559,n562);
xor (n559,n560,n561);
xor (n560,n477,n498);
xor (n561,n507,n524);
or (n562,n563,n621);
and (n563,n564,n600);
xor (n564,n565,n575);
nand (n565,n566,n574);
or (n566,n305,n567);
nor (n567,n568,n572);
and (n568,n319,n569);
wire s0n569,s1n569,notn569;
or (n569,s0n569,s1n569);
not(notn569,n129);
and (s0n569,notn569,n570);
and (s1n569,n129,n571);
wire s0n570,s1n570,notn570;
or (n570,s0n570,s1n570);
not(notn570,n19);
and (s0n570,notn570,1'b0);
and (s1n570,n19,n197);
xor (n571,n196,n198);
and (n572,n315,n573);
not (n573,n569);
or (n574,n306,n320);
nand (n575,n576,n591);
or (n576,n577,n588);
or (n577,n578,n585);
nor (n578,n579,n583);
and (n579,n372,n580);
wire s0n580,s1n580,notn580;
or (n580,s0n580,s1n580);
not(notn580,n93);
and (s0n580,notn580,n581);
and (s1n580,n93,n582);
wire s0n581,s1n581,notn581;
or (n581,s0n581,s1n581);
not(notn581,n19);
and (s0n581,notn581,1'b0);
and (s1n581,n19,n57);
xor (n582,n56,n58);
and (n583,n584,n373);
not (n584,n580);
nor (n585,n586,n587);
and (n586,n580,n315);
and (n587,n584,n319);
nor (n588,n589,n590);
and (n589,n372,n513);
and (n590,n373,n517);
or (n591,n592,n599);
nor (n592,n593,n597);
and (n593,n372,n594);
wire s0n594,s1n594,notn594;
or (n594,s0n594,s1n594);
not(notn594,n129);
and (s0n594,notn594,n595);
and (s1n594,n129,n596);
wire s0n595,s1n595,notn595;
or (n595,s0n595,s1n595);
not(notn595,n19);
and (s0n595,notn595,1'b0);
and (s1n595,n19,n200);
xor (n596,n199,n201);
and (n597,n373,n598);
not (n598,n594);
not (n599,n585);
nand (n600,n601,n616);
or (n601,n602,n613);
or (n602,n603,n610);
nor (n603,n604,n608);
and (n604,n605,n417);
wire s0n605,s1n605,notn605;
or (n605,s0n605,s1n605);
not(notn605,n93);
and (s0n605,notn605,n606);
and (s1n605,n93,n607);
wire s0n606,s1n606,notn606;
or (n606,s0n606,s1n606);
not(notn606,n19);
and (s0n606,notn606,1'b0);
and (s1n606,n19,n39);
xor (n607,n38,n40);
and (n608,n609,n421);
not (n609,n605);
nor (n610,n611,n612);
and (n611,n605,n14);
and (n612,n609,n15);
nor (n613,n614,n615);
and (n614,n15,n116);
and (n615,n14,n117);
or (n616,n617,n618);
not (n617,n603);
nor (n618,n619,n620);
and (n619,n123,n14);
and (n620,n132,n15);
and (n621,n565,n575);
and (n622,n560,n561);
xor (n623,n624,n671);
xor (n624,n625,n645);
xor (n625,n626,n639);
xor (n626,n627,n633);
nand (n627,n628,n629);
or (n628,n344,n501);
or (n629,n345,n630);
nor (n630,n631,n632);
and (n631,n290,n254);
and (n632,n294,n250);
nand (n633,n634,n635);
or (n634,n368,n511);
or (n635,n636,n396);
nor (n636,n637,n638);
and (n637,n382,n594);
and (n638,n383,n598);
nand (n639,n640,n641);
or (n640,n406,n521);
or (n641,n642,n408);
nor (n642,n643,n644);
and (n643,n421,n399);
and (n644,n417,n403);
xor (n645,n646,n662);
xor (n646,n647,n653);
nand (n647,n648,n649);
or (n648,n305,n328);
or (n649,n306,n650);
nor (n650,n651,n652);
and (n651,n319,n257);
and (n652,n315,n261);
nand (n653,n654,n658);
or (n654,n577,n655);
nor (n655,n656,n657);
and (n656,n372,n569);
and (n657,n373,n573);
or (n658,n599,n659);
nor (n659,n660,n661);
and (n660,n372,n322);
and (n661,n373,n326);
nand (n662,n663,n667);
or (n663,n602,n664);
nor (n664,n665,n666);
and (n665,n424,n14);
and (n666,n428,n15);
or (n667,n617,n668);
nor (n668,n669,n670);
and (n669,n432,n14);
and (n670,n436,n15);
or (n671,n672,n693);
and (n672,n673,n680);
xor (n673,n674,n677);
nand (n674,n675,n676);
or (n675,n577,n592);
or (n676,n599,n655);
nand (n677,n678,n679);
or (n678,n602,n618);
or (n679,n617,n664);
and (n680,n681,n687);
nor (n681,n682,n14);
nor (n682,n683,n686);
and (n683,n684,n421);
not (n684,n685);
and (n685,n117,n605);
and (n686,n609,n116);
nand (n687,n688,n692);
or (n688,n689,n484);
nor (n689,n690,n691);
and (n690,n163,n145);
and (n691,n218,n146);
or (n692,n481,n485);
and (n693,n674,n677);
or (n694,n695,n743);
and (n695,n696,n742);
xor (n696,n697,n698);
xor (n697,n673,n680);
or (n698,n699,n741);
and (n699,n700,n719);
xor (n700,n701,n702);
xor (n701,n681,n687);
or (n702,n703,n718);
and (n703,n704,n712);
xor (n704,n705,n706);
nor (n705,n617,n116);
nand (n706,n707,n711);
or (n707,n708,n484);
nor (n708,n709,n710);
and (n709,n449,n145);
and (n710,n453,n146);
or (n711,n689,n485);
nand (n712,n713,n714);
or (n713,n355,n345);
or (n714,n344,n715);
nor (n715,n716,n717);
and (n716,n257,n254);
and (n717,n261,n250);
and (n718,n705,n706);
or (n719,n720,n740);
and (n720,n721,n734);
xor (n721,n722,n728);
nand (n722,n723,n727);
or (n723,n368,n724);
nor (n724,n725,n726);
and (n725,n432,n382);
and (n726,n436,n383);
or (n727,n388,n396);
nand (n728,n729,n733);
or (n729,n406,n730);
nor (n730,n731,n732);
and (n731,n123,n421);
and (n732,n132,n417);
or (n733,n422,n408);
nand (n734,n735,n739);
or (n735,n142,n736);
nor (n736,n737,n738);
and (n737,n156,n290);
and (n738,n294,n157);
or (n739,n143,n443);
and (n740,n722,n728);
and (n741,n701,n702);
xor (n742,n338,n471);
and (n743,n697,n698);
or (n744,n745,n828);
and (n745,n746,n776);
xor (n746,n747,n775);
or (n747,n748,n774);
and (n748,n749,n773);
xor (n749,n750,n772);
or (n750,n751,n771);
and (n751,n752,n765);
xor (n752,n753,n759);
nand (n753,n754,n758);
or (n754,n235,n755);
nor (n755,n756,n757);
and (n756,n246,n322);
and (n757,n241,n326);
or (n758,n456,n247);
nand (n759,n760,n764);
or (n760,n272,n761);
nor (n761,n762,n763);
and (n762,n361,n282);
and (n763,n365,n283);
or (n764,n273,n462);
nand (n765,n766,n770);
or (n766,n305,n767);
nor (n767,n768,n769);
and (n768,n319,n594);
and (n769,n315,n598);
or (n770,n306,n567);
and (n771,n753,n759);
xor (n772,n440,n460);
xor (n773,n341,n404);
and (n774,n750,n772);
xor (n775,n559,n562);
or (n776,n777,n827);
and (n777,n778,n826);
xor (n778,n779,n780);
xor (n779,n564,n600);
or (n780,n781,n825);
and (n781,n782,n802);
xor (n782,n783,n789);
nand (n783,n784,n788);
or (n784,n577,n785);
nor (n785,n786,n787);
and (n786,n372,n399);
and (n787,n373,n403);
or (n788,n588,n599);
and (n789,n790,n796);
nor (n790,n791,n421);
nor (n791,n792,n795);
and (n792,n382,n793);
not (n793,n794);
and (n794,n117,n411);
and (n795,n410,n116);
nand (n796,n797,n801);
or (n797,n798,n484);
nor (n798,n799,n800);
and (n799,n298,n145);
and (n800,n302,n146);
or (n801,n708,n485);
or (n802,n803,n824);
and (n803,n804,n817);
xor (n804,n805,n811);
nand (n805,n806,n810);
or (n806,n344,n807);
nor (n807,n808,n809);
and (n808,n330,n254);
and (n809,n334,n250);
or (n810,n715,n345);
nand (n811,n812,n816);
or (n812,n368,n813);
nor (n813,n814,n815);
and (n814,n424,n382);
and (n815,n428,n383);
or (n816,n396,n724);
nand (n817,n818,n823);
or (n818,n819,n406);
not (n819,n820);
nand (n820,n821,n822);
or (n821,n421,n117);
or (n822,n417,n116);
or (n823,n730,n408);
and (n824,n805,n811);
and (n825,n783,n789);
xor (n826,n700,n719);
and (n827,n779,n780);
and (n828,n747,n775);
and (n829,n5,n555);
xor (n830,n831,n956);
xor (n831,n832,n849);
xor (n832,n833,n846);
xor (n833,n834,n843);
xor (n834,n835,n840);
xor (n835,n836,n837);
and (n836,n134,n140);
or (n837,n838,n839);
and (n838,n529,n549);
and (n839,n530,n536);
or (n840,n841,n842);
and (n841,n626,n639);
and (n842,n627,n633);
or (n843,n844,n845);
and (n844,n474,n528);
and (n845,n475,n505);
or (n846,n847,n848);
and (n847,n624,n671);
and (n848,n625,n645);
xor (n849,n850,n953);
xor (n850,n851,n903);
xor (n851,n852,n883);
xor (n852,n853,n856);
or (n853,n854,n855);
and (n854,n646,n662);
and (n855,n647,n653);
xor (n856,n857,n877);
xor (n857,n858,n871);
nand (n858,n859,n860);
or (n859,n539,n484);
or (n860,n861,n485);
nor (n861,n862,n869);
and (n862,n863,n145);
wire s0n863,s1n863,notn863;
or (n863,s0n863,s1n863);
not(notn863,n129);
and (s0n863,notn863,n864);
and (s1n863,n129,n866);
wire s0n864,s1n864,notn864;
or (n864,s0n864,s1n864);
not(notn864,n19);
and (s0n864,notn864,1'b0);
and (s1n864,n19,n865);
xor (n866,n867,n868);
not (n867,n865);
and (n868,n545,n546);
and (n869,n870,n146);
not (n870,n863);
nand (n871,n872,n873);
or (n872,n272,n552);
or (n873,n874,n273);
nor (n874,n875,n876);
and (n875,n163,n282);
and (n876,n218,n283);
nand (n877,n878,n879);
or (n878,n305,n650);
or (n879,n306,n880);
nor (n880,n881,n882);
and (n881,n319,n265);
and (n882,n315,n269);
xor (n883,n884,n897);
xor (n884,n885,n891);
nand (n885,n886,n887);
or (n886,n368,n636);
or (n887,n396,n888);
nor (n888,n889,n890);
and (n889,n382,n569);
and (n890,n383,n573);
nand (n891,n892,n893);
or (n892,n406,n642);
or (n893,n894,n408);
nor (n894,n895,n896);
and (n895,n421,n513);
and (n896,n417,n517);
nand (n897,n898,n899);
or (n898,n235,n533);
or (n899,n900,n247);
nor (n900,n901,n902);
and (n901,n246,n464);
and (n902,n241,n468);
xor (n903,n904,n950);
xor (n904,n905,n930);
xor (n905,n906,n924);
xor (n906,n907,n918);
nor (n907,n908,n116);
and (n908,n909,n917);
nand (n909,n910,n106);
not (n910,n911);
wire s0n911,s1n911,notn911;
or (n911,s0n911,s1n911);
not(notn911,n93);
and (s0n911,notn911,n912);
and (s1n911,n93,n914);
wire s0n912,s1n912,notn912;
or (n912,s0n912,s1n912);
not(notn912,n19);
and (s0n912,notn912,1'b0);
and (s1n912,n19,n913);
xor (n914,n915,n916);
not (n915,n913);
and (n916,n110,n111);
nand (n917,n911,n113);
nand (n918,n919,n920);
or (n919,n142,n220);
or (n920,n143,n921);
nor (n921,n922,n923);
and (n922,n490,n156);
and (n923,n497,n157);
nand (n924,n925,n926);
or (n925,n344,n630);
or (n926,n345,n927);
nor (n927,n928,n929);
and (n928,n298,n254);
and (n929,n302,n250);
xor (n930,n931,n944);
xor (n931,n932,n938);
nand (n932,n933,n934);
or (n933,n577,n659);
or (n934,n599,n935);
nor (n935,n936,n937);
and (n936,n372,n330);
and (n937,n373,n334);
nand (n938,n939,n940);
or (n939,n602,n668);
or (n940,n617,n941);
nor (n941,n942,n943);
and (n942,n14,n390);
and (n943,n15,n394);
nand (n944,n945,n946);
or (n945,n11,n121);
or (n946,n12,n947);
nor (n947,n948,n949);
and (n948,n424,n113);
and (n949,n428,n106);
or (n950,n951,n952);
and (n951,n8,n230);
and (n952,n9,n133);
or (n953,n954,n955);
and (n954,n6,n473);
and (n955,n7,n336);
or (n956,n957,n958);
and (n957,n556,n694);
and (n958,n557,n623);
nand (n959,n960,n1903);
or (n960,n961,n1896);
nand (n961,n962,n1885);
not (n962,n963);
nor (n963,n964,n1874);
nor (n964,n965,n1823);
nand (n965,n966,n1697);
or (n966,n967,n1696);
and (n967,n968,n1286);
xor (n968,n969,n1200);
or (n969,n970,n1199);
and (n970,n971,n1148);
xor (n971,n972,n1055);
xor (n972,n973,n1024);
xor (n973,n974,n995);
xor (n974,n975,n986);
xor (n975,n976,n977);
nor (n976,n396,n116);
nand (n977,n978,n982);
or (n978,n979,n484);
nor (n979,n980,n981);
and (n980,n145,n361);
and (n981,n365,n146);
or (n982,n983,n485);
nor (n983,n984,n985);
and (n984,n464,n145);
and (n985,n468,n146);
nand (n986,n987,n991);
or (n987,n142,n988);
nor (n988,n989,n990);
and (n989,n156,n257);
and (n990,n261,n157);
or (n991,n143,n992);
nor (n992,n993,n994);
and (n993,n265,n156);
and (n994,n269,n157);
or (n995,n996,n1023);
and (n996,n997,n1013);
xor (n997,n998,n1004);
nand (n998,n999,n1003);
or (n999,n142,n1000);
nor (n1000,n1001,n1002);
and (n1001,n156,n330);
and (n1002,n334,n157);
or (n1003,n143,n988);
nand (n1004,n1005,n1009);
or (n1005,n344,n1006);
nor (n1006,n1007,n1008);
and (n1007,n513,n254);
and (n1008,n517,n250);
or (n1009,n345,n1010);
nor (n1010,n1011,n1012);
and (n1011,n594,n254);
and (n1012,n598,n250);
nand (n1013,n1014,n1019);
or (n1014,n1015,n235);
not (n1015,n1016);
nand (n1016,n1017,n1018);
or (n1017,n241,n394);
or (n1018,n246,n390);
or (n1019,n1020,n247);
nor (n1020,n1021,n1022);
and (n1021,n246,n399);
and (n1022,n241,n403);
and (n1023,n998,n1004);
or (n1024,n1025,n1054);
and (n1025,n1026,n1045);
xor (n1026,n1027,n1036);
nand (n1027,n1028,n1032);
or (n1028,n272,n1029);
nor (n1029,n1030,n1031);
and (n1030,n569,n282);
and (n1031,n573,n283);
or (n1032,n1033,n273);
nor (n1033,n1034,n1035);
and (n1034,n322,n282);
and (n1035,n326,n283);
nand (n1036,n1037,n1041);
or (n1037,n305,n1038);
nor (n1038,n1039,n1040);
and (n1039,n424,n319);
and (n1040,n428,n315);
or (n1041,n1042,n306);
nor (n1042,n1043,n1044);
and (n1043,n432,n319);
and (n1044,n436,n315);
nand (n1045,n1046,n1050);
or (n1046,n599,n1047);
nor (n1047,n1048,n1049);
and (n1048,n123,n372);
and (n1049,n132,n373);
or (n1050,n577,n1051);
nor (n1051,n1052,n1053);
and (n1052,n373,n116);
and (n1053,n372,n117);
and (n1054,n1027,n1036);
xor (n1055,n1056,n1104);
xor (n1056,n1057,n1084);
xor (n1057,n1058,n1071);
xor (n1058,n1059,n1065);
nand (n1059,n1060,n1061);
or (n1060,n305,n1042);
or (n1061,n1062,n306);
nor (n1062,n1063,n1064);
and (n1063,n319,n390);
and (n1064,n315,n394);
nand (n1065,n1066,n1067);
or (n1066,n577,n1047);
or (n1067,n1068,n599);
nor (n1068,n1069,n1070);
and (n1069,n424,n372);
and (n1070,n428,n373);
and (n1071,n1072,n1078);
nand (n1072,n1073,n1077);
or (n1073,n1074,n484);
nor (n1074,n1075,n1076);
and (n1075,n145,n265);
and (n1076,n269,n146);
or (n1077,n979,n485);
nor (n1078,n1079,n372);
nor (n1079,n1080,n1083);
and (n1080,n319,n1081);
not (n1081,n1082);
and (n1082,n117,n580);
and (n1083,n584,n116);
xor (n1084,n1085,n1098);
xor (n1085,n1086,n1092);
nand (n1086,n1087,n1088);
or (n1087,n344,n1010);
or (n1088,n1089,n345);
nor (n1089,n1090,n1091);
and (n1090,n569,n254);
and (n1091,n573,n250);
nand (n1092,n1093,n1094);
or (n1093,n235,n1020);
or (n1094,n1095,n247);
nor (n1095,n1096,n1097);
and (n1096,n246,n513);
and (n1097,n241,n517);
nand (n1098,n1099,n1103);
or (n1099,n273,n1100);
nor (n1100,n1101,n1102);
and (n1101,n330,n282);
and (n1102,n334,n283);
or (n1103,n272,n1033);
or (n1104,n1105,n1147);
and (n1105,n1106,n1125);
xor (n1106,n1107,n1108);
xor (n1107,n1072,n1078);
or (n1108,n1109,n1124);
and (n1109,n1110,n1118);
xor (n1110,n1111,n1112);
nor (n1111,n599,n116);
nand (n1112,n1113,n1117);
or (n1113,n1114,n484);
nor (n1114,n1115,n1116);
and (n1115,n145,n257);
and (n1116,n261,n146);
or (n1117,n1074,n485);
nand (n1118,n1119,n1120);
or (n1119,n143,n1000);
or (n1120,n142,n1121);
nor (n1121,n1122,n1123);
and (n1122,n322,n156);
and (n1123,n326,n157);
and (n1124,n1111,n1112);
or (n1125,n1126,n1146);
and (n1126,n1127,n1140);
xor (n1127,n1128,n1134);
nand (n1128,n1129,n1133);
or (n1129,n344,n1130);
nor (n1130,n1131,n1132);
and (n1131,n399,n254);
and (n1132,n403,n250);
or (n1133,n1006,n345);
nand (n1134,n1135,n1136);
or (n1135,n247,n1015);
or (n1136,n235,n1137);
nor (n1137,n1138,n1139);
and (n1138,n246,n432);
and (n1139,n241,n436);
nand (n1140,n1141,n1142);
or (n1141,n306,n1038);
or (n1142,n305,n1143);
nor (n1143,n1144,n1145);
and (n1144,n123,n319);
and (n1145,n132,n315);
and (n1146,n1128,n1134);
and (n1147,n1107,n1108);
or (n1148,n1149,n1198);
and (n1149,n1150,n1153);
xor (n1150,n1151,n1152);
xor (n1151,n1026,n1045);
xor (n1152,n997,n1013);
or (n1153,n1154,n1197);
and (n1154,n1155,n1175);
xor (n1155,n1156,n1162);
nand (n1156,n1157,n1161);
or (n1157,n272,n1158);
nor (n1158,n1159,n1160);
and (n1159,n594,n282);
and (n1160,n598,n283);
or (n1161,n273,n1029);
and (n1162,n1163,n1169);
nand (n1163,n1164,n1168);
or (n1164,n1165,n484);
nor (n1165,n1166,n1167);
and (n1166,n330,n145);
and (n1167,n334,n146);
or (n1168,n1114,n485);
nor (n1169,n1170,n319);
nor (n1170,n1171,n1174);
and (n1171,n246,n1172);
not (n1172,n1173);
and (n1173,n117,n308);
and (n1174,n312,n116);
or (n1175,n1176,n1196);
and (n1176,n1177,n1190);
xor (n1177,n1178,n1184);
nand (n1178,n1179,n1183);
or (n1179,n142,n1180);
nor (n1180,n1181,n1182);
and (n1181,n569,n156);
and (n1182,n573,n157);
or (n1183,n143,n1121);
nand (n1184,n1185,n1189);
or (n1185,n344,n1186);
nor (n1186,n1187,n1188);
and (n1187,n390,n254);
and (n1188,n394,n250);
or (n1189,n1130,n345);
nand (n1190,n1191,n1195);
or (n1191,n235,n1192);
nor (n1192,n1193,n1194);
and (n1193,n424,n246);
and (n1194,n428,n241);
or (n1195,n1137,n247);
and (n1196,n1178,n1184);
and (n1197,n1156,n1162);
and (n1198,n1151,n1152);
and (n1199,n972,n1055);
xor (n1200,n1201,n1234);
xor (n1201,n1202,n1231);
xor (n1202,n1203,n1210);
xor (n1203,n1204,n1207);
or (n1204,n1205,n1206);
and (n1205,n1085,n1098);
and (n1206,n1086,n1092);
or (n1207,n1208,n1209);
and (n1208,n1058,n1071);
and (n1209,n1059,n1065);
xor (n1210,n1211,n1224);
xor (n1211,n1212,n1218);
nand (n1212,n1213,n1214);
or (n1213,n235,n1095);
or (n1214,n1215,n247);
nor (n1215,n1216,n1217);
and (n1216,n246,n594);
and (n1217,n241,n598);
nand (n1218,n1219,n1220);
or (n1219,n272,n1100);
or (n1220,n273,n1221);
nor (n1221,n1222,n1223);
and (n1222,n257,n282);
and (n1223,n261,n283);
nand (n1224,n1225,n1230);
or (n1225,n306,n1226);
not (n1226,n1227);
nand (n1227,n1228,n1229);
or (n1228,n403,n315);
or (n1229,n319,n399);
or (n1230,n305,n1062);
or (n1231,n1232,n1233);
and (n1232,n1056,n1104);
and (n1233,n1057,n1084);
xor (n1234,n1235,n1262);
xor (n1235,n1236,n1259);
xor (n1236,n1237,n1253);
xor (n1237,n1238,n1244);
nand (n1238,n1239,n1240);
or (n1239,n142,n992);
or (n1240,n143,n1241);
nor (n1241,n1242,n1243);
and (n1242,n156,n361);
and (n1243,n365,n157);
nand (n1244,n1245,n1249);
or (n1245,n368,n1246);
nor (n1246,n1247,n1248);
and (n1247,n383,n116);
and (n1248,n382,n117);
or (n1249,n1250,n396);
nor (n1250,n1251,n1252);
and (n1251,n123,n382);
and (n1252,n132,n383);
nand (n1253,n1254,n1258);
or (n1254,n1255,n345);
nor (n1255,n1256,n1257);
and (n1256,n322,n254);
and (n1257,n326,n250);
or (n1258,n344,n1089);
or (n1259,n1260,n1261);
and (n1260,n973,n1024);
and (n1261,n974,n995);
xor (n1262,n1263,n1283);
xor (n1263,n1264,n1270);
nand (n1264,n1265,n1266);
or (n1265,n577,n1068);
or (n1266,n1267,n599);
nor (n1267,n1268,n1269);
and (n1268,n432,n372);
and (n1269,n436,n373);
xor (n1270,n1271,n1277);
nand (n1271,n1272,n1273);
or (n1272,n983,n484);
or (n1273,n1274,n485);
nor (n1274,n1275,n1276);
and (n1275,n290,n145);
and (n1276,n294,n146);
nor (n1277,n1278,n382);
nor (n1278,n1279,n1282);
and (n1279,n372,n1280);
not (n1280,n1281);
and (n1281,n117,n376);
and (n1282,n387,n116);
or (n1283,n1284,n1285);
and (n1284,n975,n986);
and (n1285,n976,n977);
or (n1286,n1287,n1695);
and (n1287,n1288,n1319);
xor (n1288,n1289,n1318);
or (n1289,n1290,n1317);
and (n1290,n1291,n1316);
xor (n1291,n1292,n1315);
or (n1292,n1293,n1314);
and (n1293,n1294,n1297);
xor (n1294,n1295,n1296);
xor (n1295,n1110,n1118);
xor (n1296,n1127,n1140);
or (n1297,n1298,n1313);
and (n1298,n1299,n1312);
xor (n1299,n1300,n1306);
nand (n1300,n1301,n1305);
or (n1301,n305,n1302);
nor (n1302,n1303,n1304);
and (n1303,n315,n116);
and (n1304,n319,n117);
or (n1305,n1143,n306);
nand (n1306,n1307,n1311);
or (n1307,n272,n1308);
nor (n1308,n1309,n1310);
and (n1309,n513,n282);
and (n1310,n517,n283);
or (n1311,n1158,n273);
xor (n1312,n1163,n1169);
and (n1313,n1300,n1306);
and (n1314,n1295,n1296);
xor (n1315,n1106,n1125);
xor (n1316,n1150,n1153);
and (n1317,n1292,n1315);
xor (n1318,n971,n1148);
nand (n1319,n1320,n1692,n1694);
or (n1320,n1321,n1687);
nand (n1321,n1322,n1676);
or (n1322,n1323,n1675);
and (n1323,n1324,n1445);
xor (n1324,n1325,n1430);
or (n1325,n1326,n1429);
and (n1326,n1327,n1395);
xor (n1327,n1328,n1350);
xor (n1328,n1329,n1344);
xor (n1329,n1330,n1337);
nand (n1330,n1331,n1336);
or (n1331,n344,n1332);
not (n1332,n1333);
nor (n1333,n1334,n1335);
and (n1334,n254,n436);
and (n1335,n432,n250);
or (n1336,n1186,n345);
nand (n1337,n1338,n1343);
or (n1338,n1339,n235);
not (n1339,n1340);
nand (n1340,n1341,n1342);
or (n1341,n132,n241);
or (n1342,n123,n246);
or (n1343,n1192,n247);
nand (n1344,n1345,n1349);
or (n1345,n272,n1346);
nor (n1346,n1347,n1348);
and (n1347,n399,n282);
and (n1348,n403,n283);
or (n1349,n273,n1308);
or (n1350,n1351,n1394);
and (n1351,n1352,n1374);
xor (n1352,n1353,n1359);
nand (n1353,n1354,n1358);
or (n1354,n272,n1355);
nor (n1355,n1356,n1357);
and (n1356,n390,n282);
and (n1357,n394,n283);
or (n1358,n1346,n273);
xor (n1359,n1360,n1366);
nor (n1360,n1361,n246);
nor (n1361,n1362,n1365);
and (n1362,n1363,n254);
not (n1363,n1364);
and (n1364,n117,n238);
and (n1365,n245,n116);
nand (n1366,n1367,n1370);
or (n1367,n484,n1368);
not (n1368,n1369);
xnor (n1369,n569,n145);
or (n1370,n1371,n485);
nor (n1371,n1372,n1373);
and (n1372,n145,n322);
and (n1373,n326,n146);
or (n1374,n1375,n1393);
and (n1375,n1376,n1384);
xor (n1376,n1377,n1378);
nor (n1377,n247,n116);
nand (n1378,n1379,n1380);
or (n1379,n485,n1368);
or (n1380,n1381,n484);
nor (n1381,n1382,n1383);
and (n1382,n145,n594);
and (n1383,n598,n146);
nand (n1384,n1385,n1389);
or (n1385,n344,n1386);
nor (n1386,n1387,n1388);
and (n1387,n123,n254);
and (n1388,n132,n250);
or (n1389,n1390,n345);
nor (n1390,n1391,n1392);
and (n1391,n424,n254);
and (n1392,n428,n250);
and (n1393,n1377,n1378);
and (n1394,n1353,n1359);
xor (n1395,n1396,n1410);
xor (n1396,n1397,n1398);
and (n1397,n1360,n1366);
xor (n1398,n1399,n1404);
xor (n1399,n1400,n1401);
nor (n1400,n306,n116);
nand (n1401,n1402,n1403);
or (n1402,n1371,n484);
or (n1403,n1165,n485);
nand (n1404,n1405,n1409);
or (n1405,n142,n1406);
nor (n1406,n1407,n1408);
and (n1407,n594,n156);
and (n1408,n598,n157);
or (n1409,n143,n1180);
or (n1410,n1411,n1428);
and (n1411,n1412,n1422);
xor (n1412,n1413,n1419);
nand (n1413,n1414,n1418);
or (n1414,n142,n1415);
nor (n1415,n1416,n1417);
and (n1416,n156,n513);
and (n1417,n517,n157);
or (n1418,n1406,n143);
nand (n1419,n1420,n1421);
or (n1420,n345,n1332);
or (n1421,n1390,n344);
nand (n1422,n1423,n1424);
or (n1423,n247,n1339);
or (n1424,n235,n1425);
nor (n1425,n1426,n1427);
and (n1426,n241,n116);
and (n1427,n246,n117);
and (n1428,n1413,n1419);
and (n1429,n1328,n1350);
xor (n1430,n1431,n1436);
xor (n1431,n1432,n1433);
xor (n1432,n1177,n1190);
or (n1433,n1434,n1435);
and (n1434,n1396,n1410);
and (n1435,n1397,n1398);
xor (n1436,n1437,n1444);
xor (n1437,n1438,n1441);
or (n1438,n1439,n1440);
and (n1439,n1399,n1404);
and (n1440,n1400,n1401);
or (n1441,n1442,n1443);
and (n1442,n1329,n1344);
and (n1443,n1330,n1337);
xor (n1444,n1299,n1312);
or (n1445,n1446,n1674);
and (n1446,n1447,n1484);
xor (n1447,n1448,n1483);
or (n1448,n1449,n1482);
and (n1449,n1450,n1481);
xor (n1450,n1451,n1480);
or (n1451,n1452,n1479);
and (n1452,n1453,n1466);
xor (n1453,n1454,n1460);
nand (n1454,n1455,n1459);
or (n1455,n142,n1456);
nor (n1456,n1457,n1458);
and (n1457,n399,n156);
and (n1458,n157,n403);
or (n1459,n1415,n143);
nand (n1460,n1461,n1465);
or (n1461,n272,n1462);
nor (n1462,n1463,n1464);
and (n1463,n432,n282);
and (n1464,n436,n283);
or (n1465,n1355,n273);
and (n1466,n1467,n1473);
nor (n1467,n1468,n254);
nor (n1468,n1469,n1472);
and (n1469,n1470,n282);
not (n1470,n1471);
and (n1471,n117,n347);
and (n1472,n351,n116);
nand (n1473,n1474,n1478);
or (n1474,n1475,n484);
nor (n1475,n1476,n1477);
and (n1476,n145,n513);
and (n1477,n517,n146);
or (n1478,n1381,n485);
and (n1479,n1454,n1460);
xor (n1480,n1412,n1422);
xor (n1481,n1352,n1374);
and (n1482,n1451,n1480);
xor (n1483,n1327,n1395);
nand (n1484,n1485,n1671,n1673);
or (n1485,n1486,n1544);
nand (n1486,n1487,n1539);
not (n1487,n1488);
nor (n1488,n1489,n1515);
xor (n1489,n1490,n1514);
xor (n1490,n1491,n1513);
or (n1491,n1492,n1512);
and (n1492,n1493,n1506);
xor (n1493,n1494,n1500);
nand (n1494,n1495,n1499);
or (n1495,n344,n1496);
nor (n1496,n1497,n1498);
and (n1497,n250,n116);
and (n1498,n254,n117);
or (n1499,n1386,n345);
nand (n1500,n1501,n1505);
or (n1501,n1502,n142);
nor (n1502,n1503,n1504);
and (n1503,n157,n394);
and (n1504,n156,n390);
or (n1505,n1456,n143);
nand (n1506,n1507,n1511);
or (n1507,n272,n1508);
nor (n1508,n1509,n1510);
and (n1509,n424,n282);
and (n1510,n428,n283);
or (n1511,n1462,n273);
and (n1512,n1494,n1500);
xor (n1513,n1376,n1384);
xor (n1514,n1453,n1466);
or (n1515,n1516,n1538);
and (n1516,n1517,n1537);
xor (n1517,n1518,n1519);
xor (n1518,n1467,n1473);
or (n1519,n1520,n1536);
and (n1520,n1521,n1530);
xor (n1521,n1522,n1523);
nor (n1522,n345,n116);
nand (n1523,n1524,n1529);
or (n1524,n1525,n484);
not (n1525,n1526);
nand (n1526,n1527,n1528);
or (n1527,n146,n403);
nand (n1528,n403,n146);
or (n1529,n1475,n485);
nand (n1530,n1531,n1535);
or (n1531,n142,n1532);
nor (n1532,n1533,n1534);
and (n1533,n156,n432);
and (n1534,n157,n436);
or (n1535,n1502,n143);
and (n1536,n1522,n1523);
xor (n1537,n1493,n1506);
and (n1538,n1518,n1519);
or (n1539,n1540,n1541);
xor (n1540,n1450,n1481);
or (n1541,n1542,n1543);
and (n1542,n1490,n1514);
and (n1543,n1491,n1513);
nor (n1544,n1545,n1670);
and (n1545,n1546,n1665);
or (n1546,n1547,n1664);
and (n1547,n1548,n1589);
xor (n1548,n1549,n1582);
or (n1549,n1550,n1581);
and (n1550,n1551,n1567);
xor (n1551,n1552,n1558);
nand (n1552,n1553,n1557);
or (n1553,n142,n1554);
nor (n1554,n1555,n1556);
and (n1555,n157,n428);
and (n1556,n156,n424);
or (n1557,n1532,n143);
or (n1558,n1559,n1563);
nor (n1559,n1560,n273);
nor (n1560,n1561,n1562);
and (n1561,n282,n123);
and (n1562,n283,n132);
nor (n1563,n272,n1564);
nor (n1564,n1565,n1566);
and (n1565,n283,n116);
and (n1566,n282,n117);
xor (n1567,n1568,n1574);
nor (n1568,n1569,n282);
nor (n1569,n1570,n1573);
and (n1570,n1571,n156);
not (n1571,n1572);
and (n1572,n117,n276);
and (n1573,n286,n116);
nand (n1574,n1575,n1580);
or (n1575,n484,n1576);
not (n1576,n1577);
nand (n1577,n1578,n1579);
or (n1578,n145,n390);
nand (n1579,n390,n145);
nand (n1580,n1526,n486);
and (n1581,n1552,n1558);
xor (n1582,n1583,n1588);
xor (n1583,n1584,n1587);
nand (n1584,n1585,n1586);
or (n1585,n272,n1560);
or (n1586,n1508,n273);
and (n1587,n1568,n1574);
xor (n1588,n1521,n1530);
or (n1589,n1590,n1663);
and (n1590,n1591,n1611);
xor (n1591,n1592,n1610);
or (n1592,n1593,n1609);
and (n1593,n1594,n1603);
xor (n1594,n1595,n1596);
and (n1595,n274,n117);
nand (n1596,n1597,n1602);
or (n1597,n484,n1598);
not (n1598,n1599);
nand (n1599,n1600,n1601);
or (n1600,n146,n436);
nand (n1601,n436,n146);
nand (n1602,n1577,n486);
nand (n1603,n1604,n1608);
or (n1604,n142,n1605);
nor (n1605,n1606,n1607);
and (n1606,n156,n123);
and (n1607,n157,n132);
or (n1608,n1554,n143);
and (n1609,n1595,n1596);
xor (n1610,n1551,n1567);
or (n1611,n1612,n1662);
and (n1612,n1613,n1630);
xor (n1613,n1614,n1629);
and (n1614,n1615,n1621);
and (n1615,n1616,n157);
nand (n1616,n1617,n1620);
nand (n1617,n1618,n145);
not (n1618,n1619);
and (n1619,n117,n149);
nand (n1620,n153,n116);
nand (n1621,n1622,n1623);
or (n1622,n485,n1598);
nand (n1623,n1624,n1628);
not (n1624,n1625);
nor (n1625,n1626,n1627);
and (n1626,n428,n146);
and (n1627,n424,n145);
not (n1628,n484);
xor (n1629,n1594,n1603);
or (n1630,n1631,n1661);
and (n1631,n1632,n1640);
xor (n1632,n1633,n1639);
nand (n1633,n1634,n1638);
or (n1634,n142,n1635);
nor (n1635,n1636,n1637);
and (n1636,n157,n116);
and (n1637,n156,n117);
or (n1638,n1605,n143);
xor (n1639,n1615,n1621);
or (n1640,n1641,n1660);
and (n1641,n1642,n1650);
xor (n1642,n1643,n1644);
nor (n1643,n143,n116);
nand (n1644,n1645,n1649);
or (n1645,n1646,n484);
or (n1646,n1647,n1648);
and (n1647,n145,n132);
and (n1648,n123,n146);
or (n1649,n1625,n485);
nor (n1650,n1651,n1658);
nor (n1651,n1652,n1654);
and (n1652,n1653,n486);
not (n1653,n1646);
and (n1654,n1655,n1628);
nand (n1655,n1656,n1657);
or (n1656,n145,n117);
or (n1657,n146,n116);
or (n1658,n145,n1659);
and (n1659,n117,n486);
and (n1660,n1643,n1644);
and (n1661,n1633,n1639);
and (n1662,n1614,n1629);
and (n1663,n1592,n1610);
and (n1664,n1549,n1582);
or (n1665,n1666,n1667);
xor (n1666,n1517,n1537);
or (n1667,n1668,n1669);
and (n1668,n1583,n1588);
and (n1669,n1584,n1587);
and (n1670,n1666,n1667);
nand (n1671,n1539,n1672);
and (n1672,n1489,n1515);
nand (n1673,n1540,n1541);
and (n1674,n1448,n1483);
and (n1675,n1325,n1430);
or (n1676,n1677,n1684);
xor (n1677,n1678,n1683);
xor (n1678,n1679,n1680);
xor (n1679,n1155,n1175);
or (n1680,n1681,n1682);
and (n1681,n1437,n1444);
and (n1682,n1438,n1441);
xor (n1683,n1294,n1297);
or (n1684,n1685,n1686);
and (n1685,n1431,n1436);
and (n1686,n1432,n1433);
nor (n1687,n1688,n1689);
xor (n1688,n1291,n1316);
or (n1689,n1690,n1691);
and (n1690,n1678,n1683);
and (n1691,n1679,n1680);
or (n1692,n1687,n1693);
nand (n1693,n1677,n1684);
nand (n1694,n1688,n1689);
and (n1695,n1289,n1318);
and (n1696,n969,n1200);
nor (n1697,n1698,n1818);
nor (n1698,n1699,n1809);
xor (n1699,n1700,n1764);
xor (n1700,n1701,n1739);
xor (n1701,n1702,n1724);
xor (n1702,n1703,n1704);
xor (n1703,n804,n817);
xor (n1704,n1705,n1718);
xor (n1705,n1706,n1712);
nand (n1706,n1707,n1711);
or (n1707,n142,n1708);
nor (n1708,n1709,n1710);
and (n1709,n156,n464);
and (n1710,n468,n157);
or (n1711,n143,n736);
nand (n1712,n1713,n1717);
or (n1713,n235,n1714);
nor (n1714,n1715,n1716);
and (n1715,n246,n569);
and (n1716,n241,n573);
or (n1717,n755,n247);
nand (n1718,n1719,n1723);
or (n1719,n1720,n272);
nor (n1720,n1721,n1722);
and (n1721,n265,n282);
and (n1722,n269,n283);
or (n1723,n273,n761);
xor (n1724,n1725,n1738);
xor (n1725,n1726,n1732);
nand (n1726,n1727,n1731);
or (n1727,n305,n1728);
nor (n1728,n1729,n1730);
and (n1729,n319,n513);
and (n1730,n315,n517);
or (n1731,n767,n306);
nand (n1732,n1733,n1737);
or (n1733,n577,n1734);
nor (n1734,n1735,n1736);
and (n1735,n372,n390);
and (n1736,n394,n373);
or (n1737,n599,n785);
xor (n1738,n790,n796);
or (n1739,n1740,n1763);
and (n1740,n1741,n1748);
xor (n1741,n1742,n1745);
or (n1742,n1743,n1744);
and (n1743,n1263,n1283);
and (n1744,n1264,n1270);
or (n1745,n1746,n1747);
and (n1746,n1203,n1210);
and (n1747,n1204,n1207);
xor (n1748,n1749,n1760);
xor (n1749,n1750,n1751);
and (n1750,n1271,n1277);
xor (n1751,n1752,n1757);
xor (n1752,n1753,n1754);
nor (n1753,n408,n116);
nand (n1754,n1755,n1756);
or (n1755,n1274,n484);
or (n1756,n798,n485);
nand (n1757,n1758,n1759);
or (n1758,n142,n1241);
or (n1759,n143,n1708);
or (n1760,n1761,n1762);
and (n1761,n1237,n1253);
and (n1762,n1238,n1244);
and (n1763,n1742,n1745);
xor (n1764,n1765,n1800);
xor (n1765,n1766,n1769);
or (n1766,n1767,n1768);
and (n1767,n1749,n1760);
and (n1768,n1750,n1751);
xor (n1769,n1770,n1787);
xor (n1770,n1771,n1774);
or (n1771,n1772,n1773);
and (n1772,n1752,n1757);
and (n1773,n1753,n1754);
or (n1774,n1775,n1786);
and (n1775,n1776,n1783);
xor (n1776,n1777,n1780);
nand (n1777,n1778,n1779);
or (n1778,n272,n1221);
or (n1779,n273,n1720);
nand (n1780,n1781,n1782);
or (n1781,n1226,n305);
or (n1782,n1728,n306);
nand (n1783,n1784,n1785);
or (n1784,n577,n1267);
or (n1785,n1734,n599);
and (n1786,n1777,n1780);
or (n1787,n1788,n1799);
and (n1788,n1789,n1796);
xor (n1789,n1790,n1793);
nand (n1790,n1791,n1792);
or (n1791,n368,n1250);
or (n1792,n813,n396);
nand (n1793,n1794,n1795);
or (n1794,n344,n1255);
or (n1795,n807,n345);
nand (n1796,n1797,n1798);
or (n1797,n235,n1215);
or (n1798,n1714,n247);
and (n1799,n1790,n1793);
or (n1800,n1801,n1808);
and (n1801,n1802,n1807);
xor (n1802,n1803,n1806);
or (n1803,n1804,n1805);
and (n1804,n1211,n1224);
and (n1805,n1212,n1218);
xor (n1806,n1776,n1783);
xor (n1807,n1789,n1796);
and (n1808,n1803,n1806);
or (n1809,n1810,n1817);
and (n1810,n1811,n1816);
xor (n1811,n1812,n1813);
xor (n1812,n1802,n1807);
or (n1813,n1814,n1815);
and (n1814,n1235,n1262);
and (n1815,n1236,n1259);
xor (n1816,n1741,n1748);
and (n1817,n1812,n1813);
nor (n1818,n1819,n1820);
xor (n1819,n1811,n1816);
or (n1820,n1821,n1822);
and (n1821,n1201,n1234);
and (n1822,n1202,n1231);
or (n1823,n1824,n1869);
nor (n1824,n1825,n1860);
xor (n1825,n1826,n1845);
xor (n1826,n1827,n1828);
xor (n1827,n778,n826);
or (n1828,n1829,n1844);
and (n1829,n1830,n1837);
xor (n1830,n1831,n1834);
or (n1831,n1832,n1833);
and (n1832,n1770,n1787);
and (n1833,n1771,n1774);
or (n1834,n1835,n1836);
and (n1835,n1702,n1724);
and (n1836,n1703,n1704);
xor (n1837,n1838,n1843);
xor (n1838,n1839,n1842);
or (n1839,n1840,n1841);
and (n1840,n1705,n1718);
and (n1841,n1706,n1712);
xor (n1842,n752,n765);
xor (n1843,n704,n712);
and (n1844,n1831,n1834);
xor (n1845,n1846,n1851);
xor (n1846,n1847,n1850);
or (n1847,n1848,n1849);
and (n1848,n1838,n1843);
and (n1849,n1839,n1842);
xor (n1850,n749,n773);
or (n1851,n1852,n1859);
and (n1852,n1853,n1858);
xor (n1853,n1854,n1855);
xor (n1854,n721,n734);
or (n1855,n1856,n1857);
and (n1856,n1725,n1738);
and (n1857,n1726,n1732);
xor (n1858,n782,n802);
and (n1859,n1854,n1855);
or (n1860,n1861,n1868);
and (n1861,n1862,n1867);
xor (n1862,n1863,n1864);
xor (n1863,n1853,n1858);
or (n1864,n1865,n1866);
and (n1865,n1765,n1800);
and (n1866,n1766,n1769);
xor (n1867,n1830,n1837);
and (n1868,n1863,n1864);
nor (n1869,n1870,n1873);
or (n1870,n1871,n1872);
and (n1871,n1700,n1764);
and (n1872,n1701,n1739);
xor (n1873,n1862,n1867);
nand (n1874,n1875,n1884);
or (n1875,n1876,n1824);
nor (n1876,n1877,n1883);
and (n1877,n1878,n1882);
nand (n1878,n1879,n1881);
or (n1879,n1698,n1880);
nand (n1880,n1819,n1820);
nand (n1881,n1699,n1809);
not (n1882,n1869);
and (n1883,n1870,n1873);
nand (n1884,n1825,n1860);
or (n1885,n1886,n1893);
xor (n1886,n1887,n1892);
xor (n1887,n1888,n1889);
xor (n1888,n696,n742);
or (n1889,n1890,n1891);
and (n1890,n1846,n1851);
and (n1891,n1847,n1850);
xor (n1892,n746,n776);
or (n1893,n1894,n1895);
and (n1894,n1826,n1845);
and (n1895,n1827,n1828);
and (n1896,n1897,n1899);
not (n1897,n1898);
xor (n1898,n4,n744);
not (n1899,n1900);
or (n1900,n1901,n1902);
and (n1901,n1887,n1892);
and (n1902,n1888,n1889);
nor (n1903,n1904,n1908);
and (n1904,n1905,n1906);
not (n1905,n1896);
not (n1906,n1907);
nand (n1907,n1886,n1893);
nor (n1908,n1897,n1899);
xor (n1909,n1910,n3285);
xor (n1910,n1911,n3282);
xor (n1911,n1912,n3281);
xor (n1912,n1913,n3273);
xor (n1913,n1914,n3272);
xor (n1914,n1915,n3257);
xor (n1915,n1916,n3256);
xor (n1916,n1917,n3236);
xor (n1917,n1918,n3235);
xor (n1918,n1919,n3208);
xor (n1919,n1920,n3207);
xor (n1920,n1921,n3175);
xor (n1921,n1922,n3174);
xor (n1922,n1923,n3135);
xor (n1923,n1924,n3134);
xor (n1924,n1925,n3090);
xor (n1925,n1926,n3089);
xor (n1926,n1927,n3038);
xor (n1927,n1928,n3037);
xor (n1928,n1929,n2981);
xor (n1929,n1930,n2980);
xor (n1930,n1931,n2917);
xor (n1931,n1932,n2916);
xor (n1932,n1933,n2848);
xor (n1933,n1934,n2847);
xor (n1934,n1935,n2772);
xor (n1935,n1936,n2771);
xor (n1936,n1937,n2691);
xor (n1937,n1938,n2690);
xor (n1938,n1939,n2604);
xor (n1939,n1940,n2603);
xor (n1940,n1941,n2511);
xor (n1941,n1942,n2510);
xor (n1942,n1943,n2411);
xor (n1943,n1944,n2410);
xor (n1944,n1945,n2306);
xor (n1945,n1946,n2305);
xor (n1946,n1947,n2194);
xor (n1947,n1948,n2193);
xor (n1948,n1949,n2077);
xor (n1949,n1950,n2076);
xor (n1950,n1951,n1954);
xor (n1951,n1952,n1953);
and (n1952,n863,n486);
and (n1953,n541,n146);
or (n1954,n1955,n1958);
and (n1955,n1956,n1957);
and (n1956,n541,n486);
and (n1957,n490,n146);
and (n1958,n1959,n1960);
xor (n1959,n1956,n1957);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
and (n1962,n490,n486);
and (n1963,n222,n146);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
and (n1968,n222,n486);
and (n1969,n163,n146);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
and (n1974,n163,n486);
and (n1975,n449,n146);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
and (n1980,n449,n486);
and (n1981,n298,n146);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
and (n1986,n298,n486);
and (n1987,n290,n146);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
or (n1990,n1991,n1994);
and (n1991,n1992,n1993);
and (n1992,n290,n486);
and (n1993,n464,n146);
and (n1994,n1995,n1996);
xor (n1995,n1992,n1993);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
and (n1998,n464,n486);
and (n1999,n361,n146);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2006);
and (n2003,n2004,n2005);
and (n2004,n361,n486);
and (n2005,n265,n146);
and (n2006,n2007,n2008);
xor (n2007,n2004,n2005);
or (n2008,n2009,n2012);
and (n2009,n2010,n2011);
and (n2010,n265,n486);
and (n2011,n257,n146);
and (n2012,n2013,n2014);
xor (n2013,n2010,n2011);
or (n2014,n2015,n2018);
and (n2015,n2016,n2017);
and (n2016,n257,n486);
and (n2017,n330,n146);
and (n2018,n2019,n2020);
xor (n2019,n2016,n2017);
or (n2020,n2021,n2024);
and (n2021,n2022,n2023);
and (n2022,n330,n486);
and (n2023,n322,n146);
and (n2024,n2025,n2026);
xor (n2025,n2022,n2023);
or (n2026,n2027,n2030);
and (n2027,n2028,n2029);
and (n2028,n322,n486);
and (n2029,n569,n146);
and (n2030,n2031,n2032);
xor (n2031,n2028,n2029);
or (n2032,n2033,n2036);
and (n2033,n2034,n2035);
and (n2034,n569,n486);
and (n2035,n594,n146);
and (n2036,n2037,n2038);
xor (n2037,n2034,n2035);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
and (n2040,n594,n486);
and (n2041,n513,n146);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
or (n2044,n2045,n2048);
and (n2045,n2046,n2047);
and (n2046,n513,n486);
and (n2047,n399,n146);
and (n2048,n2049,n2050);
xor (n2049,n2046,n2047);
or (n2050,n2051,n2054);
and (n2051,n2052,n2053);
and (n2052,n399,n486);
and (n2053,n390,n146);
and (n2054,n2055,n2056);
xor (n2055,n2052,n2053);
or (n2056,n2057,n2060);
and (n2057,n2058,n2059);
and (n2058,n390,n486);
and (n2059,n432,n146);
and (n2060,n2061,n2062);
xor (n2061,n2058,n2059);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
and (n2064,n432,n486);
and (n2065,n424,n146);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2071);
and (n2069,n2070,n1648);
and (n2070,n424,n486);
and (n2071,n2072,n2073);
xor (n2072,n2070,n1648);
and (n2073,n2074,n2075);
and (n2074,n123,n486);
and (n2075,n117,n146);
and (n2076,n490,n149);
or (n2077,n2078,n2081);
and (n2078,n2079,n2080);
xor (n2079,n1959,n1960);
and (n2080,n222,n149);
and (n2081,n2082,n2083);
xor (n2082,n2079,n2080);
or (n2083,n2084,n2087);
and (n2084,n2085,n2086);
xor (n2085,n1965,n1966);
and (n2086,n163,n149);
and (n2087,n2088,n2089);
xor (n2088,n2085,n2086);
or (n2089,n2090,n2093);
and (n2090,n2091,n2092);
xor (n2091,n1971,n1972);
and (n2092,n449,n149);
and (n2093,n2094,n2095);
xor (n2094,n2091,n2092);
or (n2095,n2096,n2099);
and (n2096,n2097,n2098);
xor (n2097,n1977,n1978);
and (n2098,n298,n149);
and (n2099,n2100,n2101);
xor (n2100,n2097,n2098);
or (n2101,n2102,n2105);
and (n2102,n2103,n2104);
xor (n2103,n1983,n1984);
and (n2104,n290,n149);
and (n2105,n2106,n2107);
xor (n2106,n2103,n2104);
or (n2107,n2108,n2111);
and (n2108,n2109,n2110);
xor (n2109,n1989,n1990);
and (n2110,n464,n149);
and (n2111,n2112,n2113);
xor (n2112,n2109,n2110);
or (n2113,n2114,n2117);
and (n2114,n2115,n2116);
xor (n2115,n1995,n1996);
and (n2116,n361,n149);
and (n2117,n2118,n2119);
xor (n2118,n2115,n2116);
or (n2119,n2120,n2123);
and (n2120,n2121,n2122);
xor (n2121,n2001,n2002);
and (n2122,n265,n149);
and (n2123,n2124,n2125);
xor (n2124,n2121,n2122);
or (n2125,n2126,n2129);
and (n2126,n2127,n2128);
xor (n2127,n2007,n2008);
and (n2128,n257,n149);
and (n2129,n2130,n2131);
xor (n2130,n2127,n2128);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2013,n2014);
and (n2134,n330,n149);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2019,n2020);
and (n2140,n322,n149);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2025,n2026);
and (n2146,n569,n149);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2031,n2032);
and (n2152,n594,n149);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2037,n2038);
and (n2158,n513,n149);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2043,n2044);
and (n2164,n399,n149);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
or (n2167,n2168,n2171);
and (n2168,n2169,n2170);
xor (n2169,n2049,n2050);
and (n2170,n390,n149);
and (n2171,n2172,n2173);
xor (n2172,n2169,n2170);
or (n2173,n2174,n2177);
and (n2174,n2175,n2176);
xor (n2175,n2055,n2056);
and (n2176,n432,n149);
and (n2177,n2178,n2179);
xor (n2178,n2175,n2176);
or (n2179,n2180,n2183);
and (n2180,n2181,n2182);
xor (n2181,n2061,n2062);
and (n2182,n424,n149);
and (n2183,n2184,n2185);
xor (n2184,n2181,n2182);
or (n2185,n2186,n2189);
and (n2186,n2187,n2188);
xor (n2187,n2067,n2068);
and (n2188,n123,n149);
and (n2189,n2190,n2191);
xor (n2190,n2187,n2188);
and (n2191,n2192,n1619);
xor (n2192,n2072,n2073);
and (n2193,n222,n157);
or (n2194,n2195,n2198);
and (n2195,n2196,n2197);
xor (n2196,n2082,n2083);
and (n2197,n163,n157);
and (n2198,n2199,n2200);
xor (n2199,n2196,n2197);
or (n2200,n2201,n2204);
and (n2201,n2202,n2203);
xor (n2202,n2088,n2089);
and (n2203,n449,n157);
and (n2204,n2205,n2206);
xor (n2205,n2202,n2203);
or (n2206,n2207,n2210);
and (n2207,n2208,n2209);
xor (n2208,n2094,n2095);
and (n2209,n298,n157);
and (n2210,n2211,n2212);
xor (n2211,n2208,n2209);
or (n2212,n2213,n2216);
and (n2213,n2214,n2215);
xor (n2214,n2100,n2101);
and (n2215,n290,n157);
and (n2216,n2217,n2218);
xor (n2217,n2214,n2215);
or (n2218,n2219,n2222);
and (n2219,n2220,n2221);
xor (n2220,n2106,n2107);
and (n2221,n464,n157);
and (n2222,n2223,n2224);
xor (n2223,n2220,n2221);
or (n2224,n2225,n2228);
and (n2225,n2226,n2227);
xor (n2226,n2112,n2113);
and (n2227,n361,n157);
and (n2228,n2229,n2230);
xor (n2229,n2226,n2227);
or (n2230,n2231,n2234);
and (n2231,n2232,n2233);
xor (n2232,n2118,n2119);
and (n2233,n265,n157);
and (n2234,n2235,n2236);
xor (n2235,n2232,n2233);
or (n2236,n2237,n2240);
and (n2237,n2238,n2239);
xor (n2238,n2124,n2125);
and (n2239,n257,n157);
and (n2240,n2241,n2242);
xor (n2241,n2238,n2239);
or (n2242,n2243,n2246);
and (n2243,n2244,n2245);
xor (n2244,n2130,n2131);
and (n2245,n330,n157);
and (n2246,n2247,n2248);
xor (n2247,n2244,n2245);
or (n2248,n2249,n2252);
and (n2249,n2250,n2251);
xor (n2250,n2136,n2137);
and (n2251,n322,n157);
and (n2252,n2253,n2254);
xor (n2253,n2250,n2251);
or (n2254,n2255,n2258);
and (n2255,n2256,n2257);
xor (n2256,n2142,n2143);
and (n2257,n569,n157);
and (n2258,n2259,n2260);
xor (n2259,n2256,n2257);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2148,n2149);
and (n2263,n594,n157);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2154,n2155);
and (n2269,n513,n157);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2160,n2161);
and (n2275,n399,n157);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2282);
and (n2279,n2280,n2281);
xor (n2280,n2166,n2167);
and (n2281,n390,n157);
and (n2282,n2283,n2284);
xor (n2283,n2280,n2281);
or (n2284,n2285,n2288);
and (n2285,n2286,n2287);
xor (n2286,n2172,n2173);
and (n2287,n432,n157);
and (n2288,n2289,n2290);
xor (n2289,n2286,n2287);
or (n2290,n2291,n2294);
and (n2291,n2292,n2293);
xor (n2292,n2178,n2179);
and (n2293,n424,n157);
and (n2294,n2295,n2296);
xor (n2295,n2292,n2293);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2184,n2185);
and (n2299,n123,n157);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
and (n2302,n2303,n2304);
xor (n2303,n2190,n2191);
and (n2304,n117,n157);
and (n2305,n163,n276);
or (n2306,n2307,n2310);
and (n2307,n2308,n2309);
xor (n2308,n2199,n2200);
and (n2309,n449,n276);
and (n2310,n2311,n2312);
xor (n2311,n2308,n2309);
or (n2312,n2313,n2316);
and (n2313,n2314,n2315);
xor (n2314,n2205,n2206);
and (n2315,n298,n276);
and (n2316,n2317,n2318);
xor (n2317,n2314,n2315);
or (n2318,n2319,n2322);
and (n2319,n2320,n2321);
xor (n2320,n2211,n2212);
and (n2321,n290,n276);
and (n2322,n2323,n2324);
xor (n2323,n2320,n2321);
or (n2324,n2325,n2328);
and (n2325,n2326,n2327);
xor (n2326,n2217,n2218);
and (n2327,n464,n276);
and (n2328,n2329,n2330);
xor (n2329,n2326,n2327);
or (n2330,n2331,n2334);
and (n2331,n2332,n2333);
xor (n2332,n2223,n2224);
and (n2333,n361,n276);
and (n2334,n2335,n2336);
xor (n2335,n2332,n2333);
or (n2336,n2337,n2340);
and (n2337,n2338,n2339);
xor (n2338,n2229,n2230);
and (n2339,n265,n276);
and (n2340,n2341,n2342);
xor (n2341,n2338,n2339);
or (n2342,n2343,n2346);
and (n2343,n2344,n2345);
xor (n2344,n2235,n2236);
and (n2345,n257,n276);
and (n2346,n2347,n2348);
xor (n2347,n2344,n2345);
or (n2348,n2349,n2352);
and (n2349,n2350,n2351);
xor (n2350,n2241,n2242);
and (n2351,n330,n276);
and (n2352,n2353,n2354);
xor (n2353,n2350,n2351);
or (n2354,n2355,n2358);
and (n2355,n2356,n2357);
xor (n2356,n2247,n2248);
and (n2357,n322,n276);
and (n2358,n2359,n2360);
xor (n2359,n2356,n2357);
or (n2360,n2361,n2364);
and (n2361,n2362,n2363);
xor (n2362,n2253,n2254);
and (n2363,n569,n276);
and (n2364,n2365,n2366);
xor (n2365,n2362,n2363);
or (n2366,n2367,n2370);
and (n2367,n2368,n2369);
xor (n2368,n2259,n2260);
and (n2369,n594,n276);
and (n2370,n2371,n2372);
xor (n2371,n2368,n2369);
or (n2372,n2373,n2376);
and (n2373,n2374,n2375);
xor (n2374,n2265,n2266);
and (n2375,n513,n276);
and (n2376,n2377,n2378);
xor (n2377,n2374,n2375);
or (n2378,n2379,n2382);
and (n2379,n2380,n2381);
xor (n2380,n2271,n2272);
and (n2381,n399,n276);
and (n2382,n2383,n2384);
xor (n2383,n2380,n2381);
or (n2384,n2385,n2388);
and (n2385,n2386,n2387);
xor (n2386,n2277,n2278);
and (n2387,n390,n276);
and (n2388,n2389,n2390);
xor (n2389,n2386,n2387);
or (n2390,n2391,n2394);
and (n2391,n2392,n2393);
xor (n2392,n2283,n2284);
and (n2393,n432,n276);
and (n2394,n2395,n2396);
xor (n2395,n2392,n2393);
or (n2396,n2397,n2400);
and (n2397,n2398,n2399);
xor (n2398,n2289,n2290);
and (n2399,n424,n276);
and (n2400,n2401,n2402);
xor (n2401,n2398,n2399);
or (n2402,n2403,n2406);
and (n2403,n2404,n2405);
xor (n2404,n2295,n2296);
and (n2405,n123,n276);
and (n2406,n2407,n2408);
xor (n2407,n2404,n2405);
and (n2408,n2409,n1572);
xor (n2409,n2301,n2302);
and (n2410,n449,n283);
or (n2411,n2412,n2415);
and (n2412,n2413,n2414);
xor (n2413,n2311,n2312);
and (n2414,n298,n283);
and (n2415,n2416,n2417);
xor (n2416,n2413,n2414);
or (n2417,n2418,n2421);
and (n2418,n2419,n2420);
xor (n2419,n2317,n2318);
and (n2420,n290,n283);
and (n2421,n2422,n2423);
xor (n2422,n2419,n2420);
or (n2423,n2424,n2427);
and (n2424,n2425,n2426);
xor (n2425,n2323,n2324);
and (n2426,n464,n283);
and (n2427,n2428,n2429);
xor (n2428,n2425,n2426);
or (n2429,n2430,n2433);
and (n2430,n2431,n2432);
xor (n2431,n2329,n2330);
and (n2432,n361,n283);
and (n2433,n2434,n2435);
xor (n2434,n2431,n2432);
or (n2435,n2436,n2439);
and (n2436,n2437,n2438);
xor (n2437,n2335,n2336);
and (n2438,n265,n283);
and (n2439,n2440,n2441);
xor (n2440,n2437,n2438);
or (n2441,n2442,n2445);
and (n2442,n2443,n2444);
xor (n2443,n2341,n2342);
and (n2444,n257,n283);
and (n2445,n2446,n2447);
xor (n2446,n2443,n2444);
or (n2447,n2448,n2451);
and (n2448,n2449,n2450);
xor (n2449,n2347,n2348);
and (n2450,n330,n283);
and (n2451,n2452,n2453);
xor (n2452,n2449,n2450);
or (n2453,n2454,n2457);
and (n2454,n2455,n2456);
xor (n2455,n2353,n2354);
and (n2456,n322,n283);
and (n2457,n2458,n2459);
xor (n2458,n2455,n2456);
or (n2459,n2460,n2463);
and (n2460,n2461,n2462);
xor (n2461,n2359,n2360);
and (n2462,n569,n283);
and (n2463,n2464,n2465);
xor (n2464,n2461,n2462);
or (n2465,n2466,n2469);
and (n2466,n2467,n2468);
xor (n2467,n2365,n2366);
and (n2468,n594,n283);
and (n2469,n2470,n2471);
xor (n2470,n2467,n2468);
or (n2471,n2472,n2475);
and (n2472,n2473,n2474);
xor (n2473,n2371,n2372);
and (n2474,n513,n283);
and (n2475,n2476,n2477);
xor (n2476,n2473,n2474);
or (n2477,n2478,n2481);
and (n2478,n2479,n2480);
xor (n2479,n2377,n2378);
and (n2480,n399,n283);
and (n2481,n2482,n2483);
xor (n2482,n2479,n2480);
or (n2483,n2484,n2487);
and (n2484,n2485,n2486);
xor (n2485,n2383,n2384);
and (n2486,n390,n283);
and (n2487,n2488,n2489);
xor (n2488,n2485,n2486);
or (n2489,n2490,n2493);
and (n2490,n2491,n2492);
xor (n2491,n2389,n2390);
and (n2492,n432,n283);
and (n2493,n2494,n2495);
xor (n2494,n2491,n2492);
or (n2495,n2496,n2499);
and (n2496,n2497,n2498);
xor (n2497,n2395,n2396);
and (n2498,n424,n283);
and (n2499,n2500,n2501);
xor (n2500,n2497,n2498);
or (n2501,n2502,n2505);
and (n2502,n2503,n2504);
xor (n2503,n2401,n2402);
and (n2504,n123,n283);
and (n2505,n2506,n2507);
xor (n2506,n2503,n2504);
and (n2507,n2508,n2509);
xor (n2508,n2407,n2408);
and (n2509,n117,n283);
and (n2510,n298,n347);
or (n2511,n2512,n2515);
and (n2512,n2513,n2514);
xor (n2513,n2416,n2417);
and (n2514,n290,n347);
and (n2515,n2516,n2517);
xor (n2516,n2513,n2514);
or (n2517,n2518,n2521);
and (n2518,n2519,n2520);
xor (n2519,n2422,n2423);
and (n2520,n464,n347);
and (n2521,n2522,n2523);
xor (n2522,n2519,n2520);
or (n2523,n2524,n2527);
and (n2524,n2525,n2526);
xor (n2525,n2428,n2429);
and (n2526,n361,n347);
and (n2527,n2528,n2529);
xor (n2528,n2525,n2526);
or (n2529,n2530,n2533);
and (n2530,n2531,n2532);
xor (n2531,n2434,n2435);
and (n2532,n265,n347);
and (n2533,n2534,n2535);
xor (n2534,n2531,n2532);
or (n2535,n2536,n2539);
and (n2536,n2537,n2538);
xor (n2537,n2440,n2441);
and (n2538,n257,n347);
and (n2539,n2540,n2541);
xor (n2540,n2537,n2538);
or (n2541,n2542,n2545);
and (n2542,n2543,n2544);
xor (n2543,n2446,n2447);
and (n2544,n330,n347);
and (n2545,n2546,n2547);
xor (n2546,n2543,n2544);
or (n2547,n2548,n2551);
and (n2548,n2549,n2550);
xor (n2549,n2452,n2453);
and (n2550,n322,n347);
and (n2551,n2552,n2553);
xor (n2552,n2549,n2550);
or (n2553,n2554,n2557);
and (n2554,n2555,n2556);
xor (n2555,n2458,n2459);
and (n2556,n569,n347);
and (n2557,n2558,n2559);
xor (n2558,n2555,n2556);
or (n2559,n2560,n2563);
and (n2560,n2561,n2562);
xor (n2561,n2464,n2465);
and (n2562,n594,n347);
and (n2563,n2564,n2565);
xor (n2564,n2561,n2562);
or (n2565,n2566,n2569);
and (n2566,n2567,n2568);
xor (n2567,n2470,n2471);
and (n2568,n513,n347);
and (n2569,n2570,n2571);
xor (n2570,n2567,n2568);
or (n2571,n2572,n2575);
and (n2572,n2573,n2574);
xor (n2573,n2476,n2477);
and (n2574,n399,n347);
and (n2575,n2576,n2577);
xor (n2576,n2573,n2574);
or (n2577,n2578,n2581);
and (n2578,n2579,n2580);
xor (n2579,n2482,n2483);
and (n2580,n390,n347);
and (n2581,n2582,n2583);
xor (n2582,n2579,n2580);
or (n2583,n2584,n2587);
and (n2584,n2585,n2586);
xor (n2585,n2488,n2489);
and (n2586,n432,n347);
and (n2587,n2588,n2589);
xor (n2588,n2585,n2586);
or (n2589,n2590,n2593);
and (n2590,n2591,n2592);
xor (n2591,n2494,n2495);
and (n2592,n424,n347);
and (n2593,n2594,n2595);
xor (n2594,n2591,n2592);
or (n2595,n2596,n2599);
and (n2596,n2597,n2598);
xor (n2597,n2500,n2501);
and (n2598,n123,n347);
and (n2599,n2600,n2601);
xor (n2600,n2597,n2598);
and (n2601,n2602,n1471);
xor (n2602,n2506,n2507);
and (n2603,n290,n250);
or (n2604,n2605,n2608);
and (n2605,n2606,n2607);
xor (n2606,n2516,n2517);
and (n2607,n464,n250);
and (n2608,n2609,n2610);
xor (n2609,n2606,n2607);
or (n2610,n2611,n2614);
and (n2611,n2612,n2613);
xor (n2612,n2522,n2523);
and (n2613,n361,n250);
and (n2614,n2615,n2616);
xor (n2615,n2612,n2613);
or (n2616,n2617,n2620);
and (n2617,n2618,n2619);
xor (n2618,n2528,n2529);
and (n2619,n265,n250);
and (n2620,n2621,n2622);
xor (n2621,n2618,n2619);
or (n2622,n2623,n2626);
and (n2623,n2624,n2625);
xor (n2624,n2534,n2535);
and (n2625,n257,n250);
and (n2626,n2627,n2628);
xor (n2627,n2624,n2625);
or (n2628,n2629,n2632);
and (n2629,n2630,n2631);
xor (n2630,n2540,n2541);
and (n2631,n330,n250);
and (n2632,n2633,n2634);
xor (n2633,n2630,n2631);
or (n2634,n2635,n2638);
and (n2635,n2636,n2637);
xor (n2636,n2546,n2547);
and (n2637,n322,n250);
and (n2638,n2639,n2640);
xor (n2639,n2636,n2637);
or (n2640,n2641,n2644);
and (n2641,n2642,n2643);
xor (n2642,n2552,n2553);
and (n2643,n569,n250);
and (n2644,n2645,n2646);
xor (n2645,n2642,n2643);
or (n2646,n2647,n2650);
and (n2647,n2648,n2649);
xor (n2648,n2558,n2559);
and (n2649,n594,n250);
and (n2650,n2651,n2652);
xor (n2651,n2648,n2649);
or (n2652,n2653,n2656);
and (n2653,n2654,n2655);
xor (n2654,n2564,n2565);
and (n2655,n513,n250);
and (n2656,n2657,n2658);
xor (n2657,n2654,n2655);
or (n2658,n2659,n2662);
and (n2659,n2660,n2661);
xor (n2660,n2570,n2571);
and (n2661,n399,n250);
and (n2662,n2663,n2664);
xor (n2663,n2660,n2661);
or (n2664,n2665,n2668);
and (n2665,n2666,n2667);
xor (n2666,n2576,n2577);
and (n2667,n390,n250);
and (n2668,n2669,n2670);
xor (n2669,n2666,n2667);
or (n2670,n2671,n2673);
and (n2671,n2672,n1335);
xor (n2672,n2582,n2583);
and (n2673,n2674,n2675);
xor (n2674,n2672,n1335);
or (n2675,n2676,n2679);
and (n2676,n2677,n2678);
xor (n2677,n2588,n2589);
and (n2678,n424,n250);
and (n2679,n2680,n2681);
xor (n2680,n2677,n2678);
or (n2681,n2682,n2685);
and (n2682,n2683,n2684);
xor (n2683,n2594,n2595);
and (n2684,n123,n250);
and (n2685,n2686,n2687);
xor (n2686,n2683,n2684);
and (n2687,n2688,n2689);
xor (n2688,n2600,n2601);
and (n2689,n117,n250);
and (n2690,n464,n238);
or (n2691,n2692,n2695);
and (n2692,n2693,n2694);
xor (n2693,n2609,n2610);
and (n2694,n361,n238);
and (n2695,n2696,n2697);
xor (n2696,n2693,n2694);
or (n2697,n2698,n2701);
and (n2698,n2699,n2700);
xor (n2699,n2615,n2616);
and (n2700,n265,n238);
and (n2701,n2702,n2703);
xor (n2702,n2699,n2700);
or (n2703,n2704,n2707);
and (n2704,n2705,n2706);
xor (n2705,n2621,n2622);
and (n2706,n257,n238);
and (n2707,n2708,n2709);
xor (n2708,n2705,n2706);
or (n2709,n2710,n2713);
and (n2710,n2711,n2712);
xor (n2711,n2627,n2628);
and (n2712,n330,n238);
and (n2713,n2714,n2715);
xor (n2714,n2711,n2712);
or (n2715,n2716,n2719);
and (n2716,n2717,n2718);
xor (n2717,n2633,n2634);
and (n2718,n322,n238);
and (n2719,n2720,n2721);
xor (n2720,n2717,n2718);
or (n2721,n2722,n2725);
and (n2722,n2723,n2724);
xor (n2723,n2639,n2640);
and (n2724,n569,n238);
and (n2725,n2726,n2727);
xor (n2726,n2723,n2724);
or (n2727,n2728,n2731);
and (n2728,n2729,n2730);
xor (n2729,n2645,n2646);
and (n2730,n594,n238);
and (n2731,n2732,n2733);
xor (n2732,n2729,n2730);
or (n2733,n2734,n2737);
and (n2734,n2735,n2736);
xor (n2735,n2651,n2652);
and (n2736,n513,n238);
and (n2737,n2738,n2739);
xor (n2738,n2735,n2736);
or (n2739,n2740,n2743);
and (n2740,n2741,n2742);
xor (n2741,n2657,n2658);
and (n2742,n399,n238);
and (n2743,n2744,n2745);
xor (n2744,n2741,n2742);
or (n2745,n2746,n2749);
and (n2746,n2747,n2748);
xor (n2747,n2663,n2664);
and (n2748,n390,n238);
and (n2749,n2750,n2751);
xor (n2750,n2747,n2748);
or (n2751,n2752,n2755);
and (n2752,n2753,n2754);
xor (n2753,n2669,n2670);
and (n2754,n432,n238);
and (n2755,n2756,n2757);
xor (n2756,n2753,n2754);
or (n2757,n2758,n2761);
and (n2758,n2759,n2760);
xor (n2759,n2674,n2675);
and (n2760,n424,n238);
and (n2761,n2762,n2763);
xor (n2762,n2759,n2760);
or (n2763,n2764,n2767);
and (n2764,n2765,n2766);
xor (n2765,n2680,n2681);
and (n2766,n123,n238);
and (n2767,n2768,n2769);
xor (n2768,n2765,n2766);
and (n2769,n2770,n1364);
xor (n2770,n2686,n2687);
and (n2771,n361,n241);
or (n2772,n2773,n2776);
and (n2773,n2774,n2775);
xor (n2774,n2696,n2697);
and (n2775,n265,n241);
and (n2776,n2777,n2778);
xor (n2777,n2774,n2775);
or (n2778,n2779,n2782);
and (n2779,n2780,n2781);
xor (n2780,n2702,n2703);
and (n2781,n257,n241);
and (n2782,n2783,n2784);
xor (n2783,n2780,n2781);
or (n2784,n2785,n2788);
and (n2785,n2786,n2787);
xor (n2786,n2708,n2709);
and (n2787,n330,n241);
and (n2788,n2789,n2790);
xor (n2789,n2786,n2787);
or (n2790,n2791,n2794);
and (n2791,n2792,n2793);
xor (n2792,n2714,n2715);
and (n2793,n322,n241);
and (n2794,n2795,n2796);
xor (n2795,n2792,n2793);
or (n2796,n2797,n2800);
and (n2797,n2798,n2799);
xor (n2798,n2720,n2721);
and (n2799,n569,n241);
and (n2800,n2801,n2802);
xor (n2801,n2798,n2799);
or (n2802,n2803,n2806);
and (n2803,n2804,n2805);
xor (n2804,n2726,n2727);
and (n2805,n594,n241);
and (n2806,n2807,n2808);
xor (n2807,n2804,n2805);
or (n2808,n2809,n2812);
and (n2809,n2810,n2811);
xor (n2810,n2732,n2733);
and (n2811,n513,n241);
and (n2812,n2813,n2814);
xor (n2813,n2810,n2811);
or (n2814,n2815,n2818);
and (n2815,n2816,n2817);
xor (n2816,n2738,n2739);
and (n2817,n399,n241);
and (n2818,n2819,n2820);
xor (n2819,n2816,n2817);
or (n2820,n2821,n2824);
and (n2821,n2822,n2823);
xor (n2822,n2744,n2745);
and (n2823,n390,n241);
and (n2824,n2825,n2826);
xor (n2825,n2822,n2823);
or (n2826,n2827,n2830);
and (n2827,n2828,n2829);
xor (n2828,n2750,n2751);
and (n2829,n432,n241);
and (n2830,n2831,n2832);
xor (n2831,n2828,n2829);
or (n2832,n2833,n2836);
and (n2833,n2834,n2835);
xor (n2834,n2756,n2757);
and (n2835,n424,n241);
and (n2836,n2837,n2838);
xor (n2837,n2834,n2835);
or (n2838,n2839,n2842);
and (n2839,n2840,n2841);
xor (n2840,n2762,n2763);
and (n2841,n123,n241);
and (n2842,n2843,n2844);
xor (n2843,n2840,n2841);
and (n2844,n2845,n2846);
xor (n2845,n2768,n2769);
and (n2846,n117,n241);
and (n2847,n265,n308);
or (n2848,n2849,n2852);
and (n2849,n2850,n2851);
xor (n2850,n2777,n2778);
and (n2851,n257,n308);
and (n2852,n2853,n2854);
xor (n2853,n2850,n2851);
or (n2854,n2855,n2858);
and (n2855,n2856,n2857);
xor (n2856,n2783,n2784);
and (n2857,n330,n308);
and (n2858,n2859,n2860);
xor (n2859,n2856,n2857);
or (n2860,n2861,n2864);
and (n2861,n2862,n2863);
xor (n2862,n2789,n2790);
and (n2863,n322,n308);
and (n2864,n2865,n2866);
xor (n2865,n2862,n2863);
or (n2866,n2867,n2870);
and (n2867,n2868,n2869);
xor (n2868,n2795,n2796);
and (n2869,n569,n308);
and (n2870,n2871,n2872);
xor (n2871,n2868,n2869);
or (n2872,n2873,n2876);
and (n2873,n2874,n2875);
xor (n2874,n2801,n2802);
and (n2875,n594,n308);
and (n2876,n2877,n2878);
xor (n2877,n2874,n2875);
or (n2878,n2879,n2882);
and (n2879,n2880,n2881);
xor (n2880,n2807,n2808);
and (n2881,n513,n308);
and (n2882,n2883,n2884);
xor (n2883,n2880,n2881);
or (n2884,n2885,n2888);
and (n2885,n2886,n2887);
xor (n2886,n2813,n2814);
and (n2887,n399,n308);
and (n2888,n2889,n2890);
xor (n2889,n2886,n2887);
or (n2890,n2891,n2894);
and (n2891,n2892,n2893);
xor (n2892,n2819,n2820);
and (n2893,n390,n308);
and (n2894,n2895,n2896);
xor (n2895,n2892,n2893);
or (n2896,n2897,n2900);
and (n2897,n2898,n2899);
xor (n2898,n2825,n2826);
and (n2899,n432,n308);
and (n2900,n2901,n2902);
xor (n2901,n2898,n2899);
or (n2902,n2903,n2906);
and (n2903,n2904,n2905);
xor (n2904,n2831,n2832);
and (n2905,n424,n308);
and (n2906,n2907,n2908);
xor (n2907,n2904,n2905);
or (n2908,n2909,n2912);
and (n2909,n2910,n2911);
xor (n2910,n2837,n2838);
and (n2911,n123,n308);
and (n2912,n2913,n2914);
xor (n2913,n2910,n2911);
and (n2914,n2915,n1173);
xor (n2915,n2843,n2844);
and (n2916,n257,n315);
or (n2917,n2918,n2921);
and (n2918,n2919,n2920);
xor (n2919,n2853,n2854);
and (n2920,n330,n315);
and (n2921,n2922,n2923);
xor (n2922,n2919,n2920);
or (n2923,n2924,n2927);
and (n2924,n2925,n2926);
xor (n2925,n2859,n2860);
and (n2926,n322,n315);
and (n2927,n2928,n2929);
xor (n2928,n2925,n2926);
or (n2929,n2930,n2933);
and (n2930,n2931,n2932);
xor (n2931,n2865,n2866);
and (n2932,n569,n315);
and (n2933,n2934,n2935);
xor (n2934,n2931,n2932);
or (n2935,n2936,n2939);
and (n2936,n2937,n2938);
xor (n2937,n2871,n2872);
and (n2938,n594,n315);
and (n2939,n2940,n2941);
xor (n2940,n2937,n2938);
or (n2941,n2942,n2945);
and (n2942,n2943,n2944);
xor (n2943,n2877,n2878);
and (n2944,n513,n315);
and (n2945,n2946,n2947);
xor (n2946,n2943,n2944);
or (n2947,n2948,n2951);
and (n2948,n2949,n2950);
xor (n2949,n2883,n2884);
and (n2950,n399,n315);
and (n2951,n2952,n2953);
xor (n2952,n2949,n2950);
or (n2953,n2954,n2957);
and (n2954,n2955,n2956);
xor (n2955,n2889,n2890);
and (n2956,n390,n315);
and (n2957,n2958,n2959);
xor (n2958,n2955,n2956);
or (n2959,n2960,n2963);
and (n2960,n2961,n2962);
xor (n2961,n2895,n2896);
and (n2962,n432,n315);
and (n2963,n2964,n2965);
xor (n2964,n2961,n2962);
or (n2965,n2966,n2969);
and (n2966,n2967,n2968);
xor (n2967,n2901,n2902);
and (n2968,n424,n315);
and (n2969,n2970,n2971);
xor (n2970,n2967,n2968);
or (n2971,n2972,n2975);
and (n2972,n2973,n2974);
xor (n2973,n2907,n2908);
and (n2974,n123,n315);
and (n2975,n2976,n2977);
xor (n2976,n2973,n2974);
and (n2977,n2978,n2979);
xor (n2978,n2913,n2914);
and (n2979,n117,n315);
and (n2980,n330,n580);
or (n2981,n2982,n2985);
and (n2982,n2983,n2984);
xor (n2983,n2922,n2923);
and (n2984,n322,n580);
and (n2985,n2986,n2987);
xor (n2986,n2983,n2984);
or (n2987,n2988,n2991);
and (n2988,n2989,n2990);
xor (n2989,n2928,n2929);
and (n2990,n569,n580);
and (n2991,n2992,n2993);
xor (n2992,n2989,n2990);
or (n2993,n2994,n2997);
and (n2994,n2995,n2996);
xor (n2995,n2934,n2935);
and (n2996,n594,n580);
and (n2997,n2998,n2999);
xor (n2998,n2995,n2996);
or (n2999,n3000,n3003);
and (n3000,n3001,n3002);
xor (n3001,n2940,n2941);
and (n3002,n513,n580);
and (n3003,n3004,n3005);
xor (n3004,n3001,n3002);
or (n3005,n3006,n3009);
and (n3006,n3007,n3008);
xor (n3007,n2946,n2947);
and (n3008,n399,n580);
and (n3009,n3010,n3011);
xor (n3010,n3007,n3008);
or (n3011,n3012,n3015);
and (n3012,n3013,n3014);
xor (n3013,n2952,n2953);
and (n3014,n390,n580);
and (n3015,n3016,n3017);
xor (n3016,n3013,n3014);
or (n3017,n3018,n3021);
and (n3018,n3019,n3020);
xor (n3019,n2958,n2959);
and (n3020,n432,n580);
and (n3021,n3022,n3023);
xor (n3022,n3019,n3020);
or (n3023,n3024,n3027);
and (n3024,n3025,n3026);
xor (n3025,n2964,n2965);
and (n3026,n424,n580);
and (n3027,n3028,n3029);
xor (n3028,n3025,n3026);
or (n3029,n3030,n3033);
and (n3030,n3031,n3032);
xor (n3031,n2970,n2971);
and (n3032,n123,n580);
and (n3033,n3034,n3035);
xor (n3034,n3031,n3032);
and (n3035,n3036,n1082);
xor (n3036,n2976,n2977);
and (n3037,n322,n373);
or (n3038,n3039,n3042);
and (n3039,n3040,n3041);
xor (n3040,n2986,n2987);
and (n3041,n569,n373);
and (n3042,n3043,n3044);
xor (n3043,n3040,n3041);
or (n3044,n3045,n3048);
and (n3045,n3046,n3047);
xor (n3046,n2992,n2993);
and (n3047,n594,n373);
and (n3048,n3049,n3050);
xor (n3049,n3046,n3047);
or (n3050,n3051,n3054);
and (n3051,n3052,n3053);
xor (n3052,n2998,n2999);
and (n3053,n513,n373);
and (n3054,n3055,n3056);
xor (n3055,n3052,n3053);
or (n3056,n3057,n3060);
and (n3057,n3058,n3059);
xor (n3058,n3004,n3005);
and (n3059,n399,n373);
and (n3060,n3061,n3062);
xor (n3061,n3058,n3059);
or (n3062,n3063,n3066);
and (n3063,n3064,n3065);
xor (n3064,n3010,n3011);
and (n3065,n390,n373);
and (n3066,n3067,n3068);
xor (n3067,n3064,n3065);
or (n3068,n3069,n3072);
and (n3069,n3070,n3071);
xor (n3070,n3016,n3017);
and (n3071,n432,n373);
and (n3072,n3073,n3074);
xor (n3073,n3070,n3071);
or (n3074,n3075,n3078);
and (n3075,n3076,n3077);
xor (n3076,n3022,n3023);
and (n3077,n424,n373);
and (n3078,n3079,n3080);
xor (n3079,n3076,n3077);
or (n3080,n3081,n3084);
and (n3081,n3082,n3083);
xor (n3082,n3028,n3029);
and (n3083,n123,n373);
and (n3084,n3085,n3086);
xor (n3085,n3082,n3083);
and (n3086,n3087,n3088);
xor (n3087,n3034,n3035);
and (n3088,n117,n373);
and (n3089,n569,n376);
or (n3090,n3091,n3094);
and (n3091,n3092,n3093);
xor (n3092,n3043,n3044);
and (n3093,n594,n376);
and (n3094,n3095,n3096);
xor (n3095,n3092,n3093);
or (n3096,n3097,n3100);
and (n3097,n3098,n3099);
xor (n3098,n3049,n3050);
and (n3099,n513,n376);
and (n3100,n3101,n3102);
xor (n3101,n3098,n3099);
or (n3102,n3103,n3106);
and (n3103,n3104,n3105);
xor (n3104,n3055,n3056);
and (n3105,n399,n376);
and (n3106,n3107,n3108);
xor (n3107,n3104,n3105);
or (n3108,n3109,n3112);
and (n3109,n3110,n3111);
xor (n3110,n3061,n3062);
and (n3111,n390,n376);
and (n3112,n3113,n3114);
xor (n3113,n3110,n3111);
or (n3114,n3115,n3118);
and (n3115,n3116,n3117);
xor (n3116,n3067,n3068);
and (n3117,n432,n376);
and (n3118,n3119,n3120);
xor (n3119,n3116,n3117);
or (n3120,n3121,n3124);
and (n3121,n3122,n3123);
xor (n3122,n3073,n3074);
and (n3123,n424,n376);
and (n3124,n3125,n3126);
xor (n3125,n3122,n3123);
or (n3126,n3127,n3130);
and (n3127,n3128,n3129);
xor (n3128,n3079,n3080);
and (n3129,n123,n376);
and (n3130,n3131,n3132);
xor (n3131,n3128,n3129);
and (n3132,n3133,n1281);
xor (n3133,n3085,n3086);
and (n3134,n594,n383);
or (n3135,n3136,n3139);
and (n3136,n3137,n3138);
xor (n3137,n3095,n3096);
and (n3138,n513,n383);
and (n3139,n3140,n3141);
xor (n3140,n3137,n3138);
or (n3141,n3142,n3145);
and (n3142,n3143,n3144);
xor (n3143,n3101,n3102);
and (n3144,n399,n383);
and (n3145,n3146,n3147);
xor (n3146,n3143,n3144);
or (n3147,n3148,n3151);
and (n3148,n3149,n3150);
xor (n3149,n3107,n3108);
and (n3150,n390,n383);
and (n3151,n3152,n3153);
xor (n3152,n3149,n3150);
or (n3153,n3154,n3157);
and (n3154,n3155,n3156);
xor (n3155,n3113,n3114);
and (n3156,n432,n383);
and (n3157,n3158,n3159);
xor (n3158,n3155,n3156);
or (n3159,n3160,n3163);
and (n3160,n3161,n3162);
xor (n3161,n3119,n3120);
and (n3162,n424,n383);
and (n3163,n3164,n3165);
xor (n3164,n3161,n3162);
or (n3165,n3166,n3169);
and (n3166,n3167,n3168);
xor (n3167,n3125,n3126);
and (n3168,n123,n383);
and (n3169,n3170,n3171);
xor (n3170,n3167,n3168);
and (n3171,n3172,n3173);
xor (n3172,n3131,n3132);
and (n3173,n117,n383);
and (n3174,n513,n411);
or (n3175,n3176,n3179);
and (n3176,n3177,n3178);
xor (n3177,n3140,n3141);
and (n3178,n399,n411);
and (n3179,n3180,n3181);
xor (n3180,n3177,n3178);
or (n3181,n3182,n3185);
and (n3182,n3183,n3184);
xor (n3183,n3146,n3147);
and (n3184,n390,n411);
and (n3185,n3186,n3187);
xor (n3186,n3183,n3184);
or (n3187,n3188,n3191);
and (n3188,n3189,n3190);
xor (n3189,n3152,n3153);
and (n3190,n432,n411);
and (n3191,n3192,n3193);
xor (n3192,n3189,n3190);
or (n3193,n3194,n3197);
and (n3194,n3195,n3196);
xor (n3195,n3158,n3159);
and (n3196,n424,n411);
and (n3197,n3198,n3199);
xor (n3198,n3195,n3196);
or (n3199,n3200,n3203);
and (n3200,n3201,n3202);
xor (n3201,n3164,n3165);
and (n3202,n123,n411);
and (n3203,n3204,n3205);
xor (n3204,n3201,n3202);
and (n3205,n3206,n794);
xor (n3206,n3170,n3171);
and (n3207,n399,n417);
or (n3208,n3209,n3212);
and (n3209,n3210,n3211);
xor (n3210,n3180,n3181);
and (n3211,n390,n417);
and (n3212,n3213,n3214);
xor (n3213,n3210,n3211);
or (n3214,n3215,n3218);
and (n3215,n3216,n3217);
xor (n3216,n3186,n3187);
and (n3217,n432,n417);
and (n3218,n3219,n3220);
xor (n3219,n3216,n3217);
or (n3220,n3221,n3224);
and (n3221,n3222,n3223);
xor (n3222,n3192,n3193);
and (n3223,n424,n417);
and (n3224,n3225,n3226);
xor (n3225,n3222,n3223);
or (n3226,n3227,n3230);
and (n3227,n3228,n3229);
xor (n3228,n3198,n3199);
and (n3229,n123,n417);
and (n3230,n3231,n3232);
xor (n3231,n3228,n3229);
and (n3232,n3233,n3234);
xor (n3233,n3204,n3205);
and (n3234,n117,n417);
and (n3235,n390,n605);
or (n3236,n3237,n3240);
and (n3237,n3238,n3239);
xor (n3238,n3213,n3214);
and (n3239,n432,n605);
and (n3240,n3241,n3242);
xor (n3241,n3238,n3239);
or (n3242,n3243,n3246);
and (n3243,n3244,n3245);
xor (n3244,n3219,n3220);
and (n3245,n424,n605);
and (n3246,n3247,n3248);
xor (n3247,n3244,n3245);
or (n3248,n3249,n3252);
and (n3249,n3250,n3251);
xor (n3250,n3225,n3226);
and (n3251,n123,n605);
and (n3252,n3253,n3254);
xor (n3253,n3250,n3251);
and (n3254,n3255,n685);
xor (n3255,n3231,n3232);
and (n3256,n432,n15);
or (n3257,n3258,n3261);
and (n3258,n3259,n3260);
xor (n3259,n3241,n3242);
and (n3260,n424,n15);
and (n3261,n3262,n3263);
xor (n3262,n3259,n3260);
or (n3263,n3264,n3267);
and (n3264,n3265,n3266);
xor (n3265,n3247,n3248);
and (n3266,n123,n15);
and (n3267,n3268,n3269);
xor (n3268,n3265,n3266);
and (n3269,n3270,n3271);
xor (n3270,n3253,n3254);
and (n3271,n117,n15);
and (n3272,n424,n96);
or (n3273,n3274,n3277);
and (n3274,n3275,n3276);
xor (n3275,n3262,n3263);
and (n3276,n123,n96);
and (n3277,n3278,n3279);
xor (n3278,n3275,n3276);
and (n3279,n3280,n138);
xor (n3280,n3268,n3269);
and (n3281,n123,n106);
and (n3282,n3283,n3284);
xor (n3283,n3278,n3279);
and (n3284,n117,n106);
and (n3285,n117,n911);
endmodule
