module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n436,n501,n560,n613,n660,n722,n723,n727,n729,n736
        ,n743,n750,n757,n764,n771,n778,n785,n792,n798,n800
        ,n867,n934,n1001,n1068,n1135,n1200,n1259,n1312,n1359,n1399);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n436;
input n501;
input n560;
input n613;
input n660;
input n722;
input n723;
input n727;
input n729;
input n736;
input n743;
input n750;
input n757;
input n764;
input n771;
input n778;
input n785;
input n792;
input n798;
input n800;
input n867;
input n934;
input n1001;
input n1068;
input n1135;
input n1200;
input n1259;
input n1312;
input n1359;
input n1399;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n724;
wire n725;
wire n726;
wire n728;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n799;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
xor (out,n0,n1400);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1399);
and (s0n0,notn0,n1);
and (s1n0,n1399,n700);
xor (n1,n2,n661);
xor (n2,n3,n659);
xor (n3,n4,n614);
xor (n4,n5,n612);
xor (n5,n6,n561);
xor (n6,n7,n559);
xor (n7,n8,n502);
xor (n8,n9,n500);
xor (n9,n10,n437);
xor (n10,n11,n435);
or (n11,n12,n370);
and (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
and (n370,n371,n372);
xor (n371,n13,n368);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n304,n305);
and (n375,n30,n369);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n310,n311);
and (n381,n37,n369);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
xor (n386,n316,n317);
and (n387,n44,n369);
and (n388,n389,n390);
xor (n389,n386,n387);
or (n390,n391,n394);
and (n391,n392,n393);
xor (n392,n322,n323);
and (n393,n51,n369);
and (n394,n395,n396);
xor (n395,n392,n393);
or (n396,n397,n400);
and (n397,n398,n399);
xor (n398,n328,n329);
and (n399,n58,n369);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n334,n335);
and (n405,n65,n369);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n340,n341);
and (n411,n72,n369);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n346,n347);
and (n417,n79,n369);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n352,n353);
and (n423,n86,n369);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n358,n359);
and (n429,n93,n369);
and (n430,n431,n432);
xor (n431,n428,n429);
and (n432,n433,n434);
xor (n433,n364,n365);
and (n434,n99,n369);
and (n435,n23,n436);
or (n437,n438,n441);
and (n438,n439,n440);
xor (n439,n371,n372);
and (n440,n30,n436);
and (n441,n442,n443);
xor (n442,n439,n440);
or (n443,n444,n447);
and (n444,n445,n446);
xor (n445,n377,n378);
and (n446,n37,n436);
and (n447,n448,n449);
xor (n448,n445,n446);
or (n449,n450,n453);
and (n450,n451,n452);
xor (n451,n383,n384);
and (n452,n44,n436);
and (n453,n454,n455);
xor (n454,n451,n452);
or (n455,n456,n459);
and (n456,n457,n458);
xor (n457,n389,n390);
and (n458,n51,n436);
and (n459,n460,n461);
xor (n460,n457,n458);
or (n461,n462,n465);
and (n462,n463,n464);
xor (n463,n395,n396);
and (n464,n58,n436);
and (n465,n466,n467);
xor (n466,n463,n464);
or (n467,n468,n471);
and (n468,n469,n470);
xor (n469,n401,n402);
and (n470,n65,n436);
and (n471,n472,n473);
xor (n472,n469,n470);
or (n473,n474,n477);
and (n474,n475,n476);
xor (n475,n407,n408);
and (n476,n72,n436);
and (n477,n478,n479);
xor (n478,n475,n476);
or (n479,n480,n483);
and (n480,n481,n482);
xor (n481,n413,n414);
and (n482,n79,n436);
and (n483,n484,n485);
xor (n484,n481,n482);
or (n485,n486,n489);
and (n486,n487,n488);
xor (n487,n419,n420);
and (n488,n86,n436);
and (n489,n490,n491);
xor (n490,n487,n488);
or (n491,n492,n495);
and (n492,n493,n494);
xor (n493,n425,n426);
and (n494,n93,n436);
and (n495,n496,n497);
xor (n496,n493,n494);
and (n497,n498,n499);
xor (n498,n431,n432);
and (n499,n99,n436);
and (n500,n30,n501);
or (n502,n503,n506);
and (n503,n504,n505);
xor (n504,n442,n443);
and (n505,n37,n501);
and (n506,n507,n508);
xor (n507,n504,n505);
or (n508,n509,n512);
and (n509,n510,n511);
xor (n510,n448,n449);
and (n511,n44,n501);
and (n512,n513,n514);
xor (n513,n510,n511);
or (n514,n515,n518);
and (n515,n516,n517);
xor (n516,n454,n455);
and (n517,n51,n501);
and (n518,n519,n520);
xor (n519,n516,n517);
or (n520,n521,n524);
and (n521,n522,n523);
xor (n522,n460,n461);
and (n523,n58,n501);
and (n524,n525,n526);
xor (n525,n522,n523);
or (n526,n527,n530);
and (n527,n528,n529);
xor (n528,n466,n467);
and (n529,n65,n501);
and (n530,n531,n532);
xor (n531,n528,n529);
or (n532,n533,n536);
and (n533,n534,n535);
xor (n534,n472,n473);
and (n535,n72,n501);
and (n536,n537,n538);
xor (n537,n534,n535);
or (n538,n539,n542);
and (n539,n540,n541);
xor (n540,n478,n479);
and (n541,n79,n501);
and (n542,n543,n544);
xor (n543,n540,n541);
or (n544,n545,n548);
and (n545,n546,n547);
xor (n546,n484,n485);
and (n547,n86,n501);
and (n548,n549,n550);
xor (n549,n546,n547);
or (n550,n551,n554);
and (n551,n552,n553);
xor (n552,n490,n491);
and (n553,n93,n501);
and (n554,n555,n556);
xor (n555,n552,n553);
and (n556,n557,n558);
xor (n557,n496,n497);
and (n558,n99,n501);
and (n559,n37,n560);
or (n561,n562,n565);
and (n562,n563,n564);
xor (n563,n507,n508);
and (n564,n44,n560);
and (n565,n566,n567);
xor (n566,n563,n564);
or (n567,n568,n571);
and (n568,n569,n570);
xor (n569,n513,n514);
and (n570,n51,n560);
and (n571,n572,n573);
xor (n572,n569,n570);
or (n573,n574,n577);
and (n574,n575,n576);
xor (n575,n519,n520);
and (n576,n58,n560);
and (n577,n578,n579);
xor (n578,n575,n576);
or (n579,n580,n583);
and (n580,n581,n582);
xor (n581,n525,n526);
and (n582,n65,n560);
and (n583,n584,n585);
xor (n584,n581,n582);
or (n585,n586,n589);
and (n586,n587,n588);
xor (n587,n531,n532);
and (n588,n72,n560);
and (n589,n590,n591);
xor (n590,n587,n588);
or (n591,n592,n595);
and (n592,n593,n594);
xor (n593,n537,n538);
and (n594,n79,n560);
and (n595,n596,n597);
xor (n596,n593,n594);
or (n597,n598,n601);
and (n598,n599,n600);
xor (n599,n543,n544);
and (n600,n86,n560);
and (n601,n602,n603);
xor (n602,n599,n600);
or (n603,n604,n607);
and (n604,n605,n606);
xor (n605,n549,n550);
and (n606,n93,n560);
and (n607,n608,n609);
xor (n608,n605,n606);
and (n609,n610,n611);
xor (n610,n555,n556);
and (n611,n99,n560);
and (n612,n44,n613);
or (n614,n615,n618);
and (n615,n616,n617);
xor (n616,n566,n567);
and (n617,n51,n613);
and (n618,n619,n620);
xor (n619,n616,n617);
or (n620,n621,n624);
and (n621,n622,n623);
xor (n622,n572,n573);
and (n623,n58,n613);
and (n624,n625,n626);
xor (n625,n622,n623);
or (n626,n627,n630);
and (n627,n628,n629);
xor (n628,n578,n579);
and (n629,n65,n613);
and (n630,n631,n632);
xor (n631,n628,n629);
or (n632,n633,n636);
and (n633,n634,n635);
xor (n634,n584,n585);
and (n635,n72,n613);
and (n636,n637,n638);
xor (n637,n634,n635);
or (n638,n639,n642);
and (n639,n640,n641);
xor (n640,n590,n591);
and (n641,n79,n613);
and (n642,n643,n644);
xor (n643,n640,n641);
or (n644,n645,n648);
and (n645,n646,n647);
xor (n646,n596,n597);
and (n647,n86,n613);
and (n648,n649,n650);
xor (n649,n646,n647);
or (n650,n651,n654);
and (n651,n652,n653);
xor (n652,n602,n603);
and (n653,n93,n613);
and (n654,n655,n656);
xor (n655,n652,n653);
and (n656,n657,n658);
xor (n657,n608,n609);
and (n658,n99,n613);
and (n659,n51,n660);
or (n661,n662,n665);
and (n662,n663,n664);
xor (n663,n619,n620);
and (n664,n58,n660);
and (n665,n666,n667);
xor (n666,n663,n664);
or (n667,n668,n671);
and (n668,n669,n670);
xor (n669,n625,n626);
and (n670,n65,n660);
and (n671,n672,n673);
xor (n672,n669,n670);
or (n673,n674,n677);
and (n674,n675,n676);
xor (n675,n631,n632);
and (n676,n72,n660);
and (n677,n678,n679);
xor (n678,n675,n676);
or (n679,n680,n683);
and (n680,n681,n682);
xor (n681,n637,n638);
and (n682,n79,n660);
and (n683,n684,n685);
xor (n684,n681,n682);
or (n685,n686,n689);
and (n686,n687,n688);
xor (n687,n643,n644);
and (n688,n86,n660);
and (n689,n690,n691);
xor (n690,n687,n688);
or (n691,n692,n695);
and (n692,n693,n694);
xor (n693,n649,n650);
and (n694,n93,n660);
and (n695,n696,n697);
xor (n696,n693,n694);
and (n697,n698,n699);
xor (n698,n655,n656);
and (n699,n99,n660);
xor (n700,n701,n1360);
xor (n701,n702,n1358);
xor (n702,n703,n1313);
xor (n703,n704,n1311);
xor (n704,n705,n1260);
xor (n705,n706,n1258);
xor (n706,n707,n1201);
xor (n707,n708,n1199);
xor (n708,n709,n1136);
xor (n709,n710,n1134);
or (n710,n711,n1069);
and (n711,n712,n1067);
or (n712,n713,n1002);
and (n713,n714,n1000);
or (n714,n715,n935);
and (n715,n716,n933);
or (n716,n717,n868);
and (n717,n718,n866);
or (n718,n719,n801);
and (n719,n720,n799);
and (n720,n721,n724);
and (n721,n722,n723);
or (n724,n725,n730);
and (n725,n726,n728);
and (n726,n722,n727);
and (n728,n729,n723);
and (n730,n731,n732);
xor (n731,n726,n728);
or (n732,n733,n737);
and (n733,n734,n735);
and (n734,n729,n727);
and (n735,n736,n723);
and (n737,n738,n739);
xor (n738,n734,n735);
or (n739,n740,n744);
and (n740,n741,n742);
and (n741,n736,n727);
and (n742,n743,n723);
and (n744,n745,n746);
xor (n745,n741,n742);
or (n746,n747,n751);
and (n747,n748,n749);
and (n748,n743,n727);
and (n749,n750,n723);
and (n751,n752,n753);
xor (n752,n748,n749);
or (n753,n754,n758);
and (n754,n755,n756);
and (n755,n750,n727);
and (n756,n757,n723);
and (n758,n759,n760);
xor (n759,n755,n756);
or (n760,n761,n765);
and (n761,n762,n763);
and (n762,n757,n727);
and (n763,n764,n723);
and (n765,n766,n767);
xor (n766,n762,n763);
or (n767,n768,n772);
and (n768,n769,n770);
and (n769,n764,n727);
and (n770,n771,n723);
and (n772,n773,n774);
xor (n773,n769,n770);
or (n774,n775,n779);
and (n775,n776,n777);
and (n776,n771,n727);
and (n777,n778,n723);
and (n779,n780,n781);
xor (n780,n776,n777);
or (n781,n782,n786);
and (n782,n783,n784);
and (n783,n778,n727);
and (n784,n785,n723);
and (n786,n787,n788);
xor (n787,n783,n784);
or (n788,n789,n793);
and (n789,n790,n791);
and (n790,n785,n727);
and (n791,n792,n723);
and (n793,n794,n795);
xor (n794,n790,n791);
and (n795,n796,n797);
and (n796,n792,n727);
and (n797,n798,n723);
and (n799,n722,n800);
and (n801,n802,n803);
xor (n802,n720,n799);
or (n803,n804,n807);
and (n804,n805,n806);
xor (n805,n721,n724);
and (n806,n729,n800);
and (n807,n808,n809);
xor (n808,n805,n806);
or (n809,n810,n813);
and (n810,n811,n812);
xor (n811,n731,n732);
and (n812,n736,n800);
and (n813,n814,n815);
xor (n814,n811,n812);
or (n815,n816,n819);
and (n816,n817,n818);
xor (n817,n738,n739);
and (n818,n743,n800);
and (n819,n820,n821);
xor (n820,n817,n818);
or (n821,n822,n825);
and (n822,n823,n824);
xor (n823,n745,n746);
and (n824,n750,n800);
and (n825,n826,n827);
xor (n826,n823,n824);
or (n827,n828,n831);
and (n828,n829,n830);
xor (n829,n752,n753);
and (n830,n757,n800);
and (n831,n832,n833);
xor (n832,n829,n830);
or (n833,n834,n837);
and (n834,n835,n836);
xor (n835,n759,n760);
and (n836,n764,n800);
and (n837,n838,n839);
xor (n838,n835,n836);
or (n839,n840,n843);
and (n840,n841,n842);
xor (n841,n766,n767);
and (n842,n771,n800);
and (n843,n844,n845);
xor (n844,n841,n842);
or (n845,n846,n849);
and (n846,n847,n848);
xor (n847,n773,n774);
and (n848,n778,n800);
and (n849,n850,n851);
xor (n850,n847,n848);
or (n851,n852,n855);
and (n852,n853,n854);
xor (n853,n780,n781);
and (n854,n785,n800);
and (n855,n856,n857);
xor (n856,n853,n854);
or (n857,n858,n861);
and (n858,n859,n860);
xor (n859,n787,n788);
and (n860,n792,n800);
and (n861,n862,n863);
xor (n862,n859,n860);
and (n863,n864,n865);
xor (n864,n794,n795);
and (n865,n798,n800);
and (n866,n722,n867);
and (n868,n869,n870);
xor (n869,n718,n866);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n802,n803);
and (n873,n729,n867);
and (n874,n875,n876);
xor (n875,n872,n873);
or (n876,n877,n880);
and (n877,n878,n879);
xor (n878,n808,n809);
and (n879,n736,n867);
and (n880,n881,n882);
xor (n881,n878,n879);
or (n882,n883,n886);
and (n883,n884,n885);
xor (n884,n814,n815);
and (n885,n743,n867);
and (n886,n887,n888);
xor (n887,n884,n885);
or (n888,n889,n892);
and (n889,n890,n891);
xor (n890,n820,n821);
and (n891,n750,n867);
and (n892,n893,n894);
xor (n893,n890,n891);
or (n894,n895,n898);
and (n895,n896,n897);
xor (n896,n826,n827);
and (n897,n757,n867);
and (n898,n899,n900);
xor (n899,n896,n897);
or (n900,n901,n904);
and (n901,n902,n903);
xor (n902,n832,n833);
and (n903,n764,n867);
and (n904,n905,n906);
xor (n905,n902,n903);
or (n906,n907,n910);
and (n907,n908,n909);
xor (n908,n838,n839);
and (n909,n771,n867);
and (n910,n911,n912);
xor (n911,n908,n909);
or (n912,n913,n916);
and (n913,n914,n915);
xor (n914,n844,n845);
and (n915,n778,n867);
and (n916,n917,n918);
xor (n917,n914,n915);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n850,n851);
and (n921,n785,n867);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n856,n857);
and (n927,n792,n867);
and (n928,n929,n930);
xor (n929,n926,n927);
and (n930,n931,n932);
xor (n931,n862,n863);
and (n932,n798,n867);
and (n933,n722,n934);
and (n935,n936,n937);
xor (n936,n716,n933);
or (n937,n938,n941);
and (n938,n939,n940);
xor (n939,n869,n870);
and (n940,n729,n934);
and (n941,n942,n943);
xor (n942,n939,n940);
or (n943,n944,n947);
and (n944,n945,n946);
xor (n945,n875,n876);
and (n946,n736,n934);
and (n947,n948,n949);
xor (n948,n945,n946);
or (n949,n950,n953);
and (n950,n951,n952);
xor (n951,n881,n882);
and (n952,n743,n934);
and (n953,n954,n955);
xor (n954,n951,n952);
or (n955,n956,n959);
and (n956,n957,n958);
xor (n957,n887,n888);
and (n958,n750,n934);
and (n959,n960,n961);
xor (n960,n957,n958);
or (n961,n962,n965);
and (n962,n963,n964);
xor (n963,n893,n894);
and (n964,n757,n934);
and (n965,n966,n967);
xor (n966,n963,n964);
or (n967,n968,n971);
and (n968,n969,n970);
xor (n969,n899,n900);
and (n970,n764,n934);
and (n971,n972,n973);
xor (n972,n969,n970);
or (n973,n974,n977);
and (n974,n975,n976);
xor (n975,n905,n906);
and (n976,n771,n934);
and (n977,n978,n979);
xor (n978,n975,n976);
or (n979,n980,n983);
and (n980,n981,n982);
xor (n981,n911,n912);
and (n982,n778,n934);
and (n983,n984,n985);
xor (n984,n981,n982);
or (n985,n986,n989);
and (n986,n987,n988);
xor (n987,n917,n918);
and (n988,n785,n934);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
xor (n993,n923,n924);
and (n994,n792,n934);
and (n995,n996,n997);
xor (n996,n993,n994);
and (n997,n998,n999);
xor (n998,n929,n930);
and (n999,n798,n934);
and (n1000,n722,n1001);
and (n1002,n1003,n1004);
xor (n1003,n714,n1000);
or (n1004,n1005,n1008);
and (n1005,n1006,n1007);
xor (n1006,n936,n937);
and (n1007,n729,n1001);
and (n1008,n1009,n1010);
xor (n1009,n1006,n1007);
or (n1010,n1011,n1014);
and (n1011,n1012,n1013);
xor (n1012,n942,n943);
and (n1013,n736,n1001);
and (n1014,n1015,n1016);
xor (n1015,n1012,n1013);
or (n1016,n1017,n1020);
and (n1017,n1018,n1019);
xor (n1018,n948,n949);
and (n1019,n743,n1001);
and (n1020,n1021,n1022);
xor (n1021,n1018,n1019);
or (n1022,n1023,n1026);
and (n1023,n1024,n1025);
xor (n1024,n954,n955);
and (n1025,n750,n1001);
and (n1026,n1027,n1028);
xor (n1027,n1024,n1025);
or (n1028,n1029,n1032);
and (n1029,n1030,n1031);
xor (n1030,n960,n961);
and (n1031,n757,n1001);
and (n1032,n1033,n1034);
xor (n1033,n1030,n1031);
or (n1034,n1035,n1038);
and (n1035,n1036,n1037);
xor (n1036,n966,n967);
and (n1037,n764,n1001);
and (n1038,n1039,n1040);
xor (n1039,n1036,n1037);
or (n1040,n1041,n1044);
and (n1041,n1042,n1043);
xor (n1042,n972,n973);
and (n1043,n771,n1001);
and (n1044,n1045,n1046);
xor (n1045,n1042,n1043);
or (n1046,n1047,n1050);
and (n1047,n1048,n1049);
xor (n1048,n978,n979);
and (n1049,n778,n1001);
and (n1050,n1051,n1052);
xor (n1051,n1048,n1049);
or (n1052,n1053,n1056);
and (n1053,n1054,n1055);
xor (n1054,n984,n985);
and (n1055,n785,n1001);
and (n1056,n1057,n1058);
xor (n1057,n1054,n1055);
or (n1058,n1059,n1062);
and (n1059,n1060,n1061);
xor (n1060,n990,n991);
and (n1061,n792,n1001);
and (n1062,n1063,n1064);
xor (n1063,n1060,n1061);
and (n1064,n1065,n1066);
xor (n1065,n996,n997);
and (n1066,n798,n1001);
and (n1067,n722,n1068);
and (n1069,n1070,n1071);
xor (n1070,n712,n1067);
or (n1071,n1072,n1075);
and (n1072,n1073,n1074);
xor (n1073,n1003,n1004);
and (n1074,n729,n1068);
and (n1075,n1076,n1077);
xor (n1076,n1073,n1074);
or (n1077,n1078,n1081);
and (n1078,n1079,n1080);
xor (n1079,n1009,n1010);
and (n1080,n736,n1068);
and (n1081,n1082,n1083);
xor (n1082,n1079,n1080);
or (n1083,n1084,n1087);
and (n1084,n1085,n1086);
xor (n1085,n1015,n1016);
and (n1086,n743,n1068);
and (n1087,n1088,n1089);
xor (n1088,n1085,n1086);
or (n1089,n1090,n1093);
and (n1090,n1091,n1092);
xor (n1091,n1021,n1022);
and (n1092,n750,n1068);
and (n1093,n1094,n1095);
xor (n1094,n1091,n1092);
or (n1095,n1096,n1099);
and (n1096,n1097,n1098);
xor (n1097,n1027,n1028);
and (n1098,n757,n1068);
and (n1099,n1100,n1101);
xor (n1100,n1097,n1098);
or (n1101,n1102,n1105);
and (n1102,n1103,n1104);
xor (n1103,n1033,n1034);
and (n1104,n764,n1068);
and (n1105,n1106,n1107);
xor (n1106,n1103,n1104);
or (n1107,n1108,n1111);
and (n1108,n1109,n1110);
xor (n1109,n1039,n1040);
and (n1110,n771,n1068);
and (n1111,n1112,n1113);
xor (n1112,n1109,n1110);
or (n1113,n1114,n1117);
and (n1114,n1115,n1116);
xor (n1115,n1045,n1046);
and (n1116,n778,n1068);
and (n1117,n1118,n1119);
xor (n1118,n1115,n1116);
or (n1119,n1120,n1123);
and (n1120,n1121,n1122);
xor (n1121,n1051,n1052);
and (n1122,n785,n1068);
and (n1123,n1124,n1125);
xor (n1124,n1121,n1122);
or (n1125,n1126,n1129);
and (n1126,n1127,n1128);
xor (n1127,n1057,n1058);
and (n1128,n792,n1068);
and (n1129,n1130,n1131);
xor (n1130,n1127,n1128);
and (n1131,n1132,n1133);
xor (n1132,n1063,n1064);
and (n1133,n798,n1068);
and (n1134,n722,n1135);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1070,n1071);
and (n1139,n729,n1135);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1076,n1077);
and (n1145,n736,n1135);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1082,n1083);
and (n1151,n743,n1135);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1088,n1089);
and (n1157,n750,n1135);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1094,n1095);
and (n1163,n757,n1135);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1100,n1101);
and (n1169,n764,n1135);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
or (n1172,n1173,n1176);
and (n1173,n1174,n1175);
xor (n1174,n1106,n1107);
and (n1175,n771,n1135);
and (n1176,n1177,n1178);
xor (n1177,n1174,n1175);
or (n1178,n1179,n1182);
and (n1179,n1180,n1181);
xor (n1180,n1112,n1113);
and (n1181,n778,n1135);
and (n1182,n1183,n1184);
xor (n1183,n1180,n1181);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1118,n1119);
and (n1187,n785,n1135);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1124,n1125);
and (n1193,n792,n1135);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
and (n1196,n1197,n1198);
xor (n1197,n1130,n1131);
and (n1198,n798,n1135);
and (n1199,n729,n1200);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1141,n1142);
and (n1204,n736,n1200);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1147,n1148);
and (n1210,n743,n1200);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1153,n1154);
and (n1216,n750,n1200);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1159,n1160);
and (n1222,n757,n1200);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1165,n1166);
and (n1228,n764,n1200);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1171,n1172);
and (n1234,n771,n1200);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1177,n1178);
and (n1240,n778,n1200);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1183,n1184);
and (n1246,n785,n1200);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1189,n1190);
and (n1252,n792,n1200);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
and (n1255,n1256,n1257);
xor (n1256,n1195,n1196);
and (n1257,n798,n1200);
and (n1258,n736,n1259);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1206,n1207);
and (n1263,n743,n1259);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
or (n1266,n1267,n1270);
and (n1267,n1268,n1269);
xor (n1268,n1212,n1213);
and (n1269,n750,n1259);
and (n1270,n1271,n1272);
xor (n1271,n1268,n1269);
or (n1272,n1273,n1276);
and (n1273,n1274,n1275);
xor (n1274,n1218,n1219);
and (n1275,n757,n1259);
and (n1276,n1277,n1278);
xor (n1277,n1274,n1275);
or (n1278,n1279,n1282);
and (n1279,n1280,n1281);
xor (n1280,n1224,n1225);
and (n1281,n764,n1259);
and (n1282,n1283,n1284);
xor (n1283,n1280,n1281);
or (n1284,n1285,n1288);
and (n1285,n1286,n1287);
xor (n1286,n1230,n1231);
and (n1287,n771,n1259);
and (n1288,n1289,n1290);
xor (n1289,n1286,n1287);
or (n1290,n1291,n1294);
and (n1291,n1292,n1293);
xor (n1292,n1236,n1237);
and (n1293,n778,n1259);
and (n1294,n1295,n1296);
xor (n1295,n1292,n1293);
or (n1296,n1297,n1300);
and (n1297,n1298,n1299);
xor (n1298,n1242,n1243);
and (n1299,n785,n1259);
and (n1300,n1301,n1302);
xor (n1301,n1298,n1299);
or (n1302,n1303,n1306);
and (n1303,n1304,n1305);
xor (n1304,n1248,n1249);
and (n1305,n792,n1259);
and (n1306,n1307,n1308);
xor (n1307,n1304,n1305);
and (n1308,n1309,n1310);
xor (n1309,n1254,n1255);
and (n1310,n798,n1259);
and (n1311,n743,n1312);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1265,n1266);
and (n1316,n750,n1312);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1271,n1272);
and (n1322,n757,n1312);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
or (n1325,n1326,n1329);
and (n1326,n1327,n1328);
xor (n1327,n1277,n1278);
and (n1328,n764,n1312);
and (n1329,n1330,n1331);
xor (n1330,n1327,n1328);
or (n1331,n1332,n1335);
and (n1332,n1333,n1334);
xor (n1333,n1283,n1284);
and (n1334,n771,n1312);
and (n1335,n1336,n1337);
xor (n1336,n1333,n1334);
or (n1337,n1338,n1341);
and (n1338,n1339,n1340);
xor (n1339,n1289,n1290);
and (n1340,n778,n1312);
and (n1341,n1342,n1343);
xor (n1342,n1339,n1340);
or (n1343,n1344,n1347);
and (n1344,n1345,n1346);
xor (n1345,n1295,n1296);
and (n1346,n785,n1312);
and (n1347,n1348,n1349);
xor (n1348,n1345,n1346);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1301,n1302);
and (n1352,n792,n1312);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
and (n1355,n1356,n1357);
xor (n1356,n1307,n1308);
and (n1357,n798,n1312);
and (n1358,n750,n1359);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1318,n1319);
and (n1363,n757,n1359);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1324,n1325);
and (n1369,n764,n1359);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1330,n1331);
and (n1375,n771,n1359);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1336,n1337);
and (n1381,n778,n1359);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1342,n1343);
and (n1387,n785,n1359);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1348,n1349);
and (n1393,n792,n1359);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
and (n1396,n1397,n1398);
xor (n1397,n1354,n1355);
and (n1398,n798,n1359);
xor (n1400,n1401,n2060);
xor (n1401,n1402,n2058);
xor (n1402,n1403,n2013);
xor (n1403,n1404,n2011);
xor (n1404,n1405,n1960);
xor (n1405,n1406,n1958);
xor (n1406,n1407,n1901);
xor (n1407,n1408,n1899);
xor (n1408,n1409,n1836);
xor (n1409,n1410,n1834);
or (n1410,n1411,n1769);
and (n1411,n1412,n1767);
or (n1412,n1413,n1702);
and (n1413,n1414,n1700);
or (n1414,n1415,n1635);
and (n1415,n1416,n1633);
or (n1416,n1417,n1568);
and (n1417,n1418,n1566);
or (n1418,n1419,n1501);
and (n1419,n1420,n1499);
and (n1420,n1421,n1424);
and (n1421,n1422,n1423);
wire s0n1422,s1n1422,notn1422;
or (n1422,s0n1422,s1n1422);
not(notn1422,n1399);
and (s0n1422,notn1422,n23);
and (s1n1422,n1399,n722);
wire s0n1423,s1n1423,notn1423;
or (n1423,s0n1423,s1n1423);
not(notn1423,n1399);
and (s0n1423,notn1423,n24);
and (s1n1423,n1399,n723);
or (n1424,n1425,n1430);
and (n1425,n1426,n1428);
and (n1426,n1422,n1427);
wire s0n1427,s1n1427,notn1427;
or (n1427,s0n1427,s1n1427);
not(notn1427,n1399);
and (s0n1427,notn1427,n28);
and (s1n1427,n1399,n727);
and (n1428,n1429,n1423);
wire s0n1429,s1n1429,notn1429;
or (n1429,s0n1429,s1n1429);
not(notn1429,n1399);
and (s0n1429,notn1429,n30);
and (s1n1429,n1399,n729);
and (n1430,n1431,n1432);
xor (n1431,n1426,n1428);
or (n1432,n1433,n1437);
and (n1433,n1434,n1435);
and (n1434,n1429,n1427);
and (n1435,n1436,n1423);
wire s0n1436,s1n1436,notn1436;
or (n1436,s0n1436,s1n1436);
not(notn1436,n1399);
and (s0n1436,notn1436,n37);
and (s1n1436,n1399,n736);
and (n1437,n1438,n1439);
xor (n1438,n1434,n1435);
or (n1439,n1440,n1444);
and (n1440,n1441,n1442);
and (n1441,n1436,n1427);
and (n1442,n1443,n1423);
wire s0n1443,s1n1443,notn1443;
or (n1443,s0n1443,s1n1443);
not(notn1443,n1399);
and (s0n1443,notn1443,n44);
and (s1n1443,n1399,n743);
and (n1444,n1445,n1446);
xor (n1445,n1441,n1442);
or (n1446,n1447,n1451);
and (n1447,n1448,n1449);
and (n1448,n1443,n1427);
and (n1449,n1450,n1423);
wire s0n1450,s1n1450,notn1450;
or (n1450,s0n1450,s1n1450);
not(notn1450,n1399);
and (s0n1450,notn1450,n51);
and (s1n1450,n1399,n750);
and (n1451,n1452,n1453);
xor (n1452,n1448,n1449);
or (n1453,n1454,n1458);
and (n1454,n1455,n1456);
and (n1455,n1450,n1427);
and (n1456,n1457,n1423);
wire s0n1457,s1n1457,notn1457;
or (n1457,s0n1457,s1n1457);
not(notn1457,n1399);
and (s0n1457,notn1457,n58);
and (s1n1457,n1399,n757);
and (n1458,n1459,n1460);
xor (n1459,n1455,n1456);
or (n1460,n1461,n1465);
and (n1461,n1462,n1463);
and (n1462,n1457,n1427);
and (n1463,n1464,n1423);
wire s0n1464,s1n1464,notn1464;
or (n1464,s0n1464,s1n1464);
not(notn1464,n1399);
and (s0n1464,notn1464,n65);
and (s1n1464,n1399,n764);
and (n1465,n1466,n1467);
xor (n1466,n1462,n1463);
or (n1467,n1468,n1472);
and (n1468,n1469,n1470);
and (n1469,n1464,n1427);
and (n1470,n1471,n1423);
wire s0n1471,s1n1471,notn1471;
or (n1471,s0n1471,s1n1471);
not(notn1471,n1399);
and (s0n1471,notn1471,n72);
and (s1n1471,n1399,n771);
and (n1472,n1473,n1474);
xor (n1473,n1469,n1470);
or (n1474,n1475,n1479);
and (n1475,n1476,n1477);
and (n1476,n1471,n1427);
and (n1477,n1478,n1423);
wire s0n1478,s1n1478,notn1478;
or (n1478,s0n1478,s1n1478);
not(notn1478,n1399);
and (s0n1478,notn1478,n79);
and (s1n1478,n1399,n778);
and (n1479,n1480,n1481);
xor (n1480,n1476,n1477);
or (n1481,n1482,n1486);
and (n1482,n1483,n1484);
and (n1483,n1478,n1427);
and (n1484,n1485,n1423);
wire s0n1485,s1n1485,notn1485;
or (n1485,s0n1485,s1n1485);
not(notn1485,n1399);
and (s0n1485,notn1485,n86);
and (s1n1485,n1399,n785);
and (n1486,n1487,n1488);
xor (n1487,n1483,n1484);
or (n1488,n1489,n1493);
and (n1489,n1490,n1491);
and (n1490,n1485,n1427);
and (n1491,n1492,n1423);
wire s0n1492,s1n1492,notn1492;
or (n1492,s0n1492,s1n1492);
not(notn1492,n1399);
and (s0n1492,notn1492,n93);
and (s1n1492,n1399,n792);
and (n1493,n1494,n1495);
xor (n1494,n1490,n1491);
and (n1495,n1496,n1497);
and (n1496,n1492,n1427);
and (n1497,n1498,n1423);
wire s0n1498,s1n1498,notn1498;
or (n1498,s0n1498,s1n1498);
not(notn1498,n1399);
and (s0n1498,notn1498,n99);
and (s1n1498,n1399,n798);
and (n1499,n1422,n1500);
wire s0n1500,s1n1500,notn1500;
or (n1500,s0n1500,s1n1500);
not(notn1500,n1399);
and (s0n1500,notn1500,n101);
and (s1n1500,n1399,n800);
and (n1501,n1502,n1503);
xor (n1502,n1420,n1499);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1421,n1424);
and (n1506,n1429,n1500);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1431,n1432);
and (n1512,n1436,n1500);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1438,n1439);
and (n1518,n1443,n1500);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1445,n1446);
and (n1524,n1450,n1500);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1452,n1453);
and (n1530,n1457,n1500);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1459,n1460);
and (n1536,n1464,n1500);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1466,n1467);
and (n1542,n1471,n1500);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1473,n1474);
and (n1548,n1478,n1500);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1480,n1481);
and (n1554,n1485,n1500);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1487,n1488);
and (n1560,n1492,n1500);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
and (n1563,n1564,n1565);
xor (n1564,n1494,n1495);
and (n1565,n1498,n1500);
and (n1566,n1422,n1567);
wire s0n1567,s1n1567,notn1567;
or (n1567,s0n1567,s1n1567);
not(notn1567,n1399);
and (s0n1567,notn1567,n168);
and (s1n1567,n1399,n867);
and (n1568,n1569,n1570);
xor (n1569,n1418,n1566);
or (n1570,n1571,n1574);
and (n1571,n1572,n1573);
xor (n1572,n1502,n1503);
and (n1573,n1429,n1567);
and (n1574,n1575,n1576);
xor (n1575,n1572,n1573);
or (n1576,n1577,n1580);
and (n1577,n1578,n1579);
xor (n1578,n1508,n1509);
and (n1579,n1436,n1567);
and (n1580,n1581,n1582);
xor (n1581,n1578,n1579);
or (n1582,n1583,n1586);
and (n1583,n1584,n1585);
xor (n1584,n1514,n1515);
and (n1585,n1443,n1567);
and (n1586,n1587,n1588);
xor (n1587,n1584,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n1520,n1521);
and (n1591,n1450,n1567);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1526,n1527);
and (n1597,n1457,n1567);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1532,n1533);
and (n1603,n1464,n1567);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1538,n1539);
and (n1609,n1471,n1567);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1544,n1545);
and (n1615,n1478,n1567);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1550,n1551);
and (n1621,n1485,n1567);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1556,n1557);
and (n1627,n1492,n1567);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
and (n1630,n1631,n1632);
xor (n1631,n1562,n1563);
and (n1632,n1498,n1567);
and (n1633,n1422,n1634);
wire s0n1634,s1n1634,notn1634;
or (n1634,s0n1634,s1n1634);
not(notn1634,n1399);
and (s0n1634,notn1634,n235);
and (s1n1634,n1399,n934);
and (n1635,n1636,n1637);
xor (n1636,n1416,n1633);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1569,n1570);
and (n1640,n1429,n1634);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1575,n1576);
and (n1646,n1436,n1634);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1581,n1582);
and (n1652,n1443,n1634);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1587,n1588);
and (n1658,n1450,n1634);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1593,n1594);
and (n1664,n1457,n1634);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
or (n1667,n1668,n1671);
and (n1668,n1669,n1670);
xor (n1669,n1599,n1600);
and (n1670,n1464,n1634);
and (n1671,n1672,n1673);
xor (n1672,n1669,n1670);
or (n1673,n1674,n1677);
and (n1674,n1675,n1676);
xor (n1675,n1605,n1606);
and (n1676,n1471,n1634);
and (n1677,n1678,n1679);
xor (n1678,n1675,n1676);
or (n1679,n1680,n1683);
and (n1680,n1681,n1682);
xor (n1681,n1611,n1612);
and (n1682,n1478,n1634);
and (n1683,n1684,n1685);
xor (n1684,n1681,n1682);
or (n1685,n1686,n1689);
and (n1686,n1687,n1688);
xor (n1687,n1617,n1618);
and (n1688,n1485,n1634);
and (n1689,n1690,n1691);
xor (n1690,n1687,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
xor (n1693,n1623,n1624);
and (n1694,n1492,n1634);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
and (n1697,n1698,n1699);
xor (n1698,n1629,n1630);
and (n1699,n1498,n1634);
and (n1700,n1422,n1701);
wire s0n1701,s1n1701,notn1701;
or (n1701,s0n1701,s1n1701);
not(notn1701,n1399);
and (s0n1701,notn1701,n302);
and (s1n1701,n1399,n1001);
and (n1702,n1703,n1704);
xor (n1703,n1414,n1700);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1636,n1637);
and (n1707,n1429,n1701);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
or (n1710,n1711,n1714);
and (n1711,n1712,n1713);
xor (n1712,n1642,n1643);
and (n1713,n1436,n1701);
and (n1714,n1715,n1716);
xor (n1715,n1712,n1713);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
xor (n1718,n1648,n1649);
and (n1719,n1443,n1701);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
xor (n1724,n1654,n1655);
and (n1725,n1450,n1701);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
or (n1728,n1729,n1732);
and (n1729,n1730,n1731);
xor (n1730,n1660,n1661);
and (n1731,n1457,n1701);
and (n1732,n1733,n1734);
xor (n1733,n1730,n1731);
or (n1734,n1735,n1738);
and (n1735,n1736,n1737);
xor (n1736,n1666,n1667);
and (n1737,n1464,n1701);
and (n1738,n1739,n1740);
xor (n1739,n1736,n1737);
or (n1740,n1741,n1744);
and (n1741,n1742,n1743);
xor (n1742,n1672,n1673);
and (n1743,n1471,n1701);
and (n1744,n1745,n1746);
xor (n1745,n1742,n1743);
or (n1746,n1747,n1750);
and (n1747,n1748,n1749);
xor (n1748,n1678,n1679);
and (n1749,n1478,n1701);
and (n1750,n1751,n1752);
xor (n1751,n1748,n1749);
or (n1752,n1753,n1756);
and (n1753,n1754,n1755);
xor (n1754,n1684,n1685);
and (n1755,n1485,n1701);
and (n1756,n1757,n1758);
xor (n1757,n1754,n1755);
or (n1758,n1759,n1762);
and (n1759,n1760,n1761);
xor (n1760,n1690,n1691);
and (n1761,n1492,n1701);
and (n1762,n1763,n1764);
xor (n1763,n1760,n1761);
and (n1764,n1765,n1766);
xor (n1765,n1696,n1697);
and (n1766,n1498,n1701);
and (n1767,n1422,n1768);
wire s0n1768,s1n1768,notn1768;
or (n1768,s0n1768,s1n1768);
not(notn1768,n1399);
and (s0n1768,notn1768,n369);
and (s1n1768,n1399,n1068);
and (n1769,n1770,n1771);
xor (n1770,n1412,n1767);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1703,n1704);
and (n1774,n1429,n1768);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1709,n1710);
and (n1780,n1436,n1768);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1715,n1716);
and (n1786,n1443,n1768);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1721,n1722);
and (n1792,n1450,n1768);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1727,n1728);
and (n1798,n1457,n1768);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1733,n1734);
and (n1804,n1464,n1768);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1739,n1740);
and (n1810,n1471,n1768);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1745,n1746);
and (n1816,n1478,n1768);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1751,n1752);
and (n1822,n1485,n1768);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
xor (n1827,n1757,n1758);
and (n1828,n1492,n1768);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
and (n1831,n1832,n1833);
xor (n1832,n1763,n1764);
and (n1833,n1498,n1768);
and (n1834,n1422,n1835);
wire s0n1835,s1n1835,notn1835;
or (n1835,s0n1835,s1n1835);
not(notn1835,n1399);
and (s0n1835,notn1835,n436);
and (s1n1835,n1399,n1135);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1770,n1771);
and (n1839,n1429,n1835);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1776,n1777);
and (n1845,n1436,n1835);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1782,n1783);
and (n1851,n1443,n1835);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1788,n1789);
and (n1857,n1450,n1835);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1794,n1795);
and (n1863,n1457,n1835);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1800,n1801);
and (n1869,n1464,n1835);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1806,n1807);
and (n1875,n1471,n1835);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1812,n1813);
and (n1881,n1478,n1835);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1818,n1819);
and (n1887,n1485,n1835);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1824,n1825);
and (n1893,n1492,n1835);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
and (n1896,n1897,n1898);
xor (n1897,n1830,n1831);
and (n1898,n1498,n1835);
and (n1899,n1429,n1900);
wire s0n1900,s1n1900,notn1900;
or (n1900,s0n1900,s1n1900);
not(notn1900,n1399);
and (s0n1900,notn1900,n501);
and (s1n1900,n1399,n1200);
or (n1901,n1902,n1905);
and (n1902,n1903,n1904);
xor (n1903,n1841,n1842);
and (n1904,n1436,n1900);
and (n1905,n1906,n1907);
xor (n1906,n1903,n1904);
or (n1907,n1908,n1911);
and (n1908,n1909,n1910);
xor (n1909,n1847,n1848);
and (n1910,n1443,n1900);
and (n1911,n1912,n1913);
xor (n1912,n1909,n1910);
or (n1913,n1914,n1917);
and (n1914,n1915,n1916);
xor (n1915,n1853,n1854);
and (n1916,n1450,n1900);
and (n1917,n1918,n1919);
xor (n1918,n1915,n1916);
or (n1919,n1920,n1923);
and (n1920,n1921,n1922);
xor (n1921,n1859,n1860);
and (n1922,n1457,n1900);
and (n1923,n1924,n1925);
xor (n1924,n1921,n1922);
or (n1925,n1926,n1929);
and (n1926,n1927,n1928);
xor (n1927,n1865,n1866);
and (n1928,n1464,n1900);
and (n1929,n1930,n1931);
xor (n1930,n1927,n1928);
or (n1931,n1932,n1935);
and (n1932,n1933,n1934);
xor (n1933,n1871,n1872);
and (n1934,n1471,n1900);
and (n1935,n1936,n1937);
xor (n1936,n1933,n1934);
or (n1937,n1938,n1941);
and (n1938,n1939,n1940);
xor (n1939,n1877,n1878);
and (n1940,n1478,n1900);
and (n1941,n1942,n1943);
xor (n1942,n1939,n1940);
or (n1943,n1944,n1947);
and (n1944,n1945,n1946);
xor (n1945,n1883,n1884);
and (n1946,n1485,n1900);
and (n1947,n1948,n1949);
xor (n1948,n1945,n1946);
or (n1949,n1950,n1953);
and (n1950,n1951,n1952);
xor (n1951,n1889,n1890);
and (n1952,n1492,n1900);
and (n1953,n1954,n1955);
xor (n1954,n1951,n1952);
and (n1955,n1956,n1957);
xor (n1956,n1895,n1896);
and (n1957,n1498,n1900);
and (n1958,n1436,n1959);
wire s0n1959,s1n1959,notn1959;
or (n1959,s0n1959,s1n1959);
not(notn1959,n1399);
and (s0n1959,notn1959,n560);
and (s1n1959,n1399,n1259);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
xor (n1962,n1906,n1907);
and (n1963,n1443,n1959);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
xor (n1968,n1912,n1913);
and (n1969,n1450,n1959);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
xor (n1974,n1918,n1919);
and (n1975,n1457,n1959);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
xor (n1980,n1924,n1925);
and (n1981,n1464,n1959);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
xor (n1986,n1930,n1931);
and (n1987,n1471,n1959);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
or (n1990,n1991,n1994);
and (n1991,n1992,n1993);
xor (n1992,n1936,n1937);
and (n1993,n1478,n1959);
and (n1994,n1995,n1996);
xor (n1995,n1992,n1993);
or (n1996,n1997,n2000);
and (n1997,n1998,n1999);
xor (n1998,n1942,n1943);
and (n1999,n1485,n1959);
and (n2000,n2001,n2002);
xor (n2001,n1998,n1999);
or (n2002,n2003,n2006);
and (n2003,n2004,n2005);
xor (n2004,n1948,n1949);
and (n2005,n1492,n1959);
and (n2006,n2007,n2008);
xor (n2007,n2004,n2005);
and (n2008,n2009,n2010);
xor (n2009,n1954,n1955);
and (n2010,n1498,n1959);
and (n2011,n1443,n2012);
wire s0n2012,s1n2012,notn2012;
or (n2012,s0n2012,s1n2012);
not(notn2012,n1399);
and (s0n2012,notn2012,n613);
and (s1n2012,n1399,n1312);
or (n2013,n2014,n2017);
and (n2014,n2015,n2016);
xor (n2015,n1965,n1966);
and (n2016,n1450,n2012);
and (n2017,n2018,n2019);
xor (n2018,n2015,n2016);
or (n2019,n2020,n2023);
and (n2020,n2021,n2022);
xor (n2021,n1971,n1972);
and (n2022,n1457,n2012);
and (n2023,n2024,n2025);
xor (n2024,n2021,n2022);
or (n2025,n2026,n2029);
and (n2026,n2027,n2028);
xor (n2027,n1977,n1978);
and (n2028,n1464,n2012);
and (n2029,n2030,n2031);
xor (n2030,n2027,n2028);
or (n2031,n2032,n2035);
and (n2032,n2033,n2034);
xor (n2033,n1983,n1984);
and (n2034,n1471,n2012);
and (n2035,n2036,n2037);
xor (n2036,n2033,n2034);
or (n2037,n2038,n2041);
and (n2038,n2039,n2040);
xor (n2039,n1989,n1990);
and (n2040,n1478,n2012);
and (n2041,n2042,n2043);
xor (n2042,n2039,n2040);
or (n2043,n2044,n2047);
and (n2044,n2045,n2046);
xor (n2045,n1995,n1996);
and (n2046,n1485,n2012);
and (n2047,n2048,n2049);
xor (n2048,n2045,n2046);
or (n2049,n2050,n2053);
and (n2050,n2051,n2052);
xor (n2051,n2001,n2002);
and (n2052,n1492,n2012);
and (n2053,n2054,n2055);
xor (n2054,n2051,n2052);
and (n2055,n2056,n2057);
xor (n2056,n2007,n2008);
and (n2057,n1498,n2012);
and (n2058,n1450,n2059);
wire s0n2059,s1n2059,notn2059;
or (n2059,s0n2059,s1n2059);
not(notn2059,n1399);
and (s0n2059,notn2059,n660);
and (s1n2059,n1399,n1359);
or (n2060,n2061,n2064);
and (n2061,n2062,n2063);
xor (n2062,n2018,n2019);
and (n2063,n1457,n2059);
and (n2064,n2065,n2066);
xor (n2065,n2062,n2063);
or (n2066,n2067,n2070);
and (n2067,n2068,n2069);
xor (n2068,n2024,n2025);
and (n2069,n1464,n2059);
and (n2070,n2071,n2072);
xor (n2071,n2068,n2069);
or (n2072,n2073,n2076);
and (n2073,n2074,n2075);
xor (n2074,n2030,n2031);
and (n2075,n1471,n2059);
and (n2076,n2077,n2078);
xor (n2077,n2074,n2075);
or (n2078,n2079,n2082);
and (n2079,n2080,n2081);
xor (n2080,n2036,n2037);
and (n2081,n1478,n2059);
and (n2082,n2083,n2084);
xor (n2083,n2080,n2081);
or (n2084,n2085,n2088);
and (n2085,n2086,n2087);
xor (n2086,n2042,n2043);
and (n2087,n1485,n2059);
and (n2088,n2089,n2090);
xor (n2089,n2086,n2087);
or (n2090,n2091,n2094);
and (n2091,n2092,n2093);
xor (n2092,n2048,n2049);
and (n2093,n1492,n2059);
and (n2094,n2095,n2096);
xor (n2095,n2092,n2093);
and (n2096,n2097,n2098);
xor (n2097,n2054,n2055);
and (n2098,n1498,n2059);
endmodule
