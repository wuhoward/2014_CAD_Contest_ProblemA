module top (out,n3,n4,n5,n20,n24,n25,n33,n43,n48
        ,n50,n57,n74,n76,n81,n87,n93,n100,n102,n110
        ,n119,n126,n134,n140,n176,n181,n185,n192,n196,n207
        ,n277,n296,n350);
output out;
input n3;
input n4;
input n5;
input n20;
input n24;
input n25;
input n33;
input n43;
input n48;
input n50;
input n57;
input n74;
input n76;
input n81;
input n87;
input n93;
input n100;
input n102;
input n110;
input n119;
input n126;
input n134;
input n140;
input n176;
input n181;
input n185;
input n192;
input n196;
input n207;
input n277;
input n296;
input n350;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
xnor (out,n0,n918);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n915);
nor (n7,n8,n913);
and (n8,n9,n394);
nand (n9,n10,n393);
not (n10,n11);
nor (n11,n12,n327);
xor (n12,n13,n280);
xor (n13,n14,n166);
xor (n14,n15,n144);
xor (n15,n16,n65);
and (n16,n17,n38);
nand (n17,n18,n29);
or (n18,n19,n21);
not (n19,n20);
not (n21,n22);
nor (n22,n23,n26);
and (n23,n24,n25);
and (n26,n27,n28);
not (n27,n25);
not (n28,n24);
nand (n29,n30,n36);
not (n30,n31);
nor (n31,n32,n34);
and (n32,n28,n33);
and (n34,n24,n35);
not (n35,n33);
not (n36,n37);
nand (n37,n24,n19);
nand (n38,n39,n53);
or (n39,n40,n45);
not (n40,n41);
nand (n41,n42,n44);
or (n42,n28,n43);
nand (n44,n28,n43);
not (n45,n46);
nand (n46,n47,n51);
or (n47,n48,n49);
not (n49,n50);
or (n51,n52,n50);
not (n52,n48);
nand (n53,n54,n60);
not (n54,n55);
nor (n55,n56,n58);
and (n56,n52,n57);
and (n58,n48,n59);
not (n59,n57);
nor (n60,n41,n61);
nor (n61,n62,n63);
and (n62,n52,n43);
and (n63,n48,n64);
not (n64,n43);
or (n65,n66,n143);
and (n66,n67,n121);
xor (n67,n68,n95);
nand (n68,n69,n89);
or (n69,n70,n78);
not (n70,n71);
nor (n71,n72,n77);
and (n72,n73,n75);
not (n73,n74);
not (n75,n76);
and (n77,n76,n74);
nand (n78,n79,n83);
nand (n79,n80,n82);
or (n80,n81,n75);
nand (n82,n75,n81);
not (n83,n84);
nand (n84,n85,n88);
or (n85,n86,n81);
not (n86,n87);
nand (n88,n86,n81);
nand (n89,n90,n84);
nor (n90,n91,n94);
and (n91,n92,n75);
not (n92,n93);
and (n94,n76,n93);
nand (n95,n96,n115);
or (n96,n97,n105);
not (n97,n98);
nand (n98,n99,n103);
or (n99,n100,n101);
not (n101,n102);
or (n103,n104,n102);
not (n104,n100);
not (n105,n106);
and (n106,n107,n112);
not (n107,n108);
nand (n108,n109,n111);
or (n109,n110,n75);
nand (n111,n110,n75);
nand (n112,n113,n114);
or (n113,n110,n104);
nand (n114,n104,n110);
nand (n115,n108,n116);
nor (n116,n117,n120);
and (n117,n118,n104);
not (n118,n119);
and (n120,n100,n119);
nand (n121,n122,n137);
or (n122,n123,n132);
nand (n123,n124,n129);
nor (n124,n125,n127);
and (n125,n52,n126);
and (n127,n48,n128);
not (n128,n126);
nand (n129,n130,n131);
or (n130,n126,n86);
nand (n131,n86,n126);
nor (n132,n133,n135);
and (n133,n134,n86);
and (n135,n87,n136);
not (n136,n134);
or (n137,n138,n124);
nor (n138,n139,n141);
and (n139,n86,n140);
and (n141,n87,n142);
not (n142,n140);
and (n143,n68,n95);
xor (n144,n145,n160);
xor (n145,n146,n153);
nand (n146,n147,n149);
or (n147,n148,n78);
not (n148,n90);
nand (n149,n84,n150);
nor (n150,n151,n152);
and (n151,n136,n75);
and (n152,n76,n134);
nand (n153,n154,n156);
or (n154,n155,n105);
not (n155,n116);
nand (n156,n108,n157);
nand (n157,n158,n159);
or (n158,n100,n73);
or (n159,n104,n74);
nand (n160,n161,n162);
or (n161,n123,n138);
or (n162,n124,n163);
nor (n163,n164,n165);
and (n164,n86,n57);
and (n165,n87,n59);
or (n166,n167,n279);
and (n167,n168,n223);
xor (n168,n169,n198);
xor (n169,n170,n197);
xor (n170,n171,n195);
nand (n171,n172,n189);
or (n172,n173,n183);
nand (n173,n174,n179);
nor (n174,n175,n177);
and (n175,n104,n176);
and (n177,n100,n178);
not (n178,n176);
nand (n179,n180,n182);
or (n180,n178,n181);
nand (n182,n178,n181);
nor (n183,n184,n187);
and (n184,n185,n186);
not (n186,n181);
and (n187,n181,n188);
not (n188,n185);
or (n189,n190,n174);
nor (n190,n191,n193);
and (n191,n192,n186);
and (n193,n181,n194);
not (n194,n192);
and (n195,n181,n196);
xor (n197,n17,n38);
or (n198,n199,n222);
and (n199,n200,n208);
xor (n200,n201,n206);
nand (n201,n202,n205);
or (n202,n203,n173);
not (n203,n204);
xor (n204,n196,n181);
or (n205,n174,n183);
and (n206,n181,n207);
xor (n208,n209,n215);
nand (n209,n210,n214);
or (n210,n37,n211);
nor (n211,n212,n213);
and (n212,n28,n50);
and (n213,n24,n49);
or (n214,n31,n19);
nand (n215,n216,n221);
or (n216,n217,n218);
not (n217,n60);
nor (n218,n219,n220);
and (n219,n52,n140);
and (n220,n48,n142);
or (n221,n40,n55);
and (n222,n201,n206);
and (n223,n224,n255);
or (n224,n225,n254);
and (n225,n226,n245);
xor (n226,n227,n235);
nand (n227,n228,n233);
or (n228,n229,n217);
not (n229,n230);
nand (n230,n231,n232);
or (n231,n48,n136);
or (n232,n52,n134);
nand (n233,n234,n41);
not (n234,n218);
nand (n235,n236,n240);
or (n236,n78,n237);
nor (n237,n238,n239);
and (n238,n75,n102);
and (n239,n76,n101);
or (n240,n83,n241);
not (n241,n242);
nor (n242,n243,n244);
and (n243,n118,n75);
and (n244,n76,n119);
nand (n245,n246,n250);
or (n246,n105,n247);
nor (n247,n248,n249);
and (n248,n104,n185);
and (n249,n100,n188);
or (n250,n107,n251);
nor (n251,n252,n253);
and (n252,n104,n192);
and (n253,n100,n194);
and (n254,n227,n235);
or (n255,n256,n278);
and (n256,n257,n276);
xor (n257,n258,n267);
nand (n258,n259,n263);
or (n259,n123,n260);
nor (n260,n261,n262);
and (n261,n86,n74);
and (n262,n87,n73);
or (n263,n264,n124);
nor (n264,n265,n266);
and (n265,n93,n86);
and (n266,n87,n92);
nand (n267,n268,n269);
or (n268,n203,n174);
nand (n269,n270,n275);
not (n270,n271);
nor (n271,n272,n273);
and (n272,n207,n186);
and (n273,n274,n181);
not (n274,n207);
not (n275,n173);
and (n276,n181,n277);
and (n278,n258,n267);
and (n279,n169,n198);
xor (n280,n281,n308);
xor (n281,n282,n305);
xor (n282,n283,n290);
xor (n283,n284,n289);
nand (n284,n285,n286);
or (n285,n190,n173);
nand (n286,n287,n288);
not (n287,n174);
xor (n288,n102,n181);
and (n289,n181,n185);
xor (n290,n291,n299);
nand (n291,n292,n293);
or (n292,n37,n21);
or (n293,n294,n19);
nor (n294,n295,n297);
and (n295,n28,n296);
and (n297,n24,n298);
not (n298,n296);
nand (n299,n300,n301);
or (n300,n45,n217);
nand (n301,n41,n302);
nor (n302,n303,n304);
and (n303,n48,n33);
and (n304,n35,n52);
or (n305,n306,n307);
and (n306,n170,n197);
and (n307,n171,n195);
or (n308,n309,n326);
and (n309,n310,n325);
xor (n310,n311,n312);
and (n311,n209,n215);
or (n312,n313,n324);
and (n313,n314,n321);
xor (n314,n315,n318);
nand (n315,n316,n317);
or (n316,n241,n78);
nand (n317,n84,n71);
nand (n318,n319,n320);
or (n319,n105,n251);
nand (n320,n108,n98);
nand (n321,n322,n323);
or (n322,n123,n264);
or (n323,n124,n132);
and (n324,n315,n318);
xor (n325,n67,n121);
and (n326,n311,n312);
or (n327,n328,n392);
and (n328,n329,n332);
xor (n329,n330,n331);
xor (n330,n310,n325);
xor (n331,n168,n223);
or (n332,n333,n391);
and (n333,n334,n337);
xor (n334,n335,n336);
xor (n335,n314,n321);
xor (n336,n200,n208);
or (n337,n338,n390);
and (n338,n339,n364);
xor (n339,n340,n346);
nand (n340,n341,n345);
or (n341,n37,n342);
nor (n342,n343,n344);
and (n343,n28,n57);
and (n344,n24,n59);
or (n345,n211,n19);
or (n346,n347,n363);
and (n347,n348,n357);
xor (n348,n349,n351);
and (n349,n181,n350);
nand (n351,n352,n353);
or (n352,n40,n229);
nand (n353,n60,n354);
nand (n354,n355,n356);
or (n355,n48,n92);
or (n356,n52,n93);
nand (n357,n358,n362);
or (n358,n78,n359);
nor (n359,n360,n361);
and (n360,n75,n192);
and (n361,n76,n194);
or (n362,n237,n83);
and (n363,n349,n351);
or (n364,n365,n389);
and (n365,n366,n382);
xor (n366,n367,n376);
nand (n367,n368,n374);
or (n368,n369,n105);
not (n369,n370);
nor (n370,n371,n373);
and (n371,n372,n104);
not (n372,n196);
and (n373,n100,n196);
nand (n374,n375,n108);
not (n375,n247);
nand (n376,n377,n381);
or (n377,n378,n37);
nor (n378,n379,n380);
and (n379,n28,n140);
and (n380,n24,n142);
or (n381,n342,n19);
nand (n382,n383,n388);
or (n383,n173,n384);
nor (n384,n385,n386);
and (n385,n186,n277);
and (n386,n181,n387);
not (n387,n277);
or (n388,n174,n271);
and (n389,n367,n376);
and (n390,n340,n346);
and (n391,n335,n336);
and (n392,n330,n331);
nand (n393,n12,n327);
not (n394,n395);
nand (n395,n396,n620);
not (n396,n397);
nand (n397,n398,n613);
or (n398,n399,n591);
not (n399,n400);
nand (n400,n401,n590);
or (n401,n402,n537);
nor (n402,n403,n483);
xor (n403,n404,n449);
xor (n404,n405,n406);
xor (n405,n339,n364);
or (n406,n407,n448);
and (n407,n408,n411);
xor (n408,n409,n410);
xor (n409,n366,n382);
xor (n410,n348,n357);
or (n411,n412,n447);
and (n412,n413,n430);
xor (n413,n414,n421);
nand (n414,n415,n420);
or (n415,n173,n416);
nor (n416,n417,n418);
and (n417,n350,n186);
and (n418,n419,n181);
not (n419,n350);
or (n420,n174,n384);
nand (n421,n422,n426);
or (n422,n123,n423);
nor (n423,n424,n425);
and (n424,n86,n102);
and (n425,n87,n101);
or (n426,n124,n427);
nor (n427,n428,n429);
and (n428,n86,n119);
and (n429,n87,n118);
nand (n430,n431,n446);
or (n431,n432,n438);
not (n432,n433);
nand (n433,n434,n181);
nand (n434,n435,n436);
or (n435,n100,n176);
nand (n436,n437,n419);
or (n437,n178,n104);
not (n438,n439);
nand (n439,n440,n445);
or (n440,n441,n217);
not (n441,n442);
nand (n442,n443,n444);
or (n443,n48,n73);
or (n444,n52,n74);
nand (n445,n41,n354);
or (n446,n439,n433);
and (n447,n414,n421);
and (n448,n409,n410);
xor (n449,n450,n453);
xor (n450,n451,n452);
xor (n451,n257,n276);
xor (n452,n226,n245);
or (n453,n454,n482);
and (n454,n455,n460);
xor (n455,n456,n459);
nand (n456,n457,n458);
or (n457,n123,n427);
or (n458,n124,n260);
nor (n459,n438,n433);
or (n460,n461,n481);
and (n461,n462,n475);
xor (n462,n463,n469);
nand (n463,n464,n468);
or (n464,n78,n465);
nor (n465,n466,n467);
and (n466,n75,n185);
and (n467,n76,n188);
or (n468,n83,n359);
nand (n469,n470,n474);
or (n470,n105,n471);
nor (n471,n472,n473);
and (n472,n104,n207);
and (n473,n100,n274);
or (n474,n107,n369);
nand (n475,n476,n480);
or (n476,n477,n37);
nor (n477,n478,n479);
and (n478,n28,n134);
and (n479,n24,n136);
or (n480,n378,n19);
and (n481,n463,n469);
and (n482,n456,n459);
or (n483,n484,n536);
and (n484,n485,n535);
xor (n485,n486,n487);
xor (n486,n455,n460);
or (n487,n488,n534);
and (n488,n489,n533);
xor (n489,n490,n509);
or (n490,n491,n508);
and (n491,n492,n500);
xor (n492,n493,n494);
nor (n493,n174,n419);
nand (n494,n495,n499);
or (n495,n496,n217);
nor (n496,n497,n498);
and (n497,n118,n48);
and (n498,n119,n52);
nand (n499,n442,n41);
nand (n500,n501,n506);
or (n501,n502,n78);
not (n502,n503);
nand (n503,n504,n505);
or (n504,n76,n372);
or (n505,n75,n196);
nand (n506,n507,n84);
not (n507,n465);
and (n508,n493,n494);
or (n509,n510,n532);
and (n510,n511,n526);
xor (n511,n512,n520);
nand (n512,n513,n518);
or (n513,n514,n105);
not (n514,n515);
nand (n515,n516,n517);
or (n516,n100,n387);
or (n517,n104,n277);
nand (n518,n519,n108);
not (n519,n471);
nand (n520,n521,n525);
or (n521,n522,n37);
nor (n522,n523,n524);
and (n523,n28,n93);
and (n524,n24,n92);
or (n525,n477,n19);
nand (n526,n527,n531);
or (n527,n123,n528);
nor (n528,n529,n530);
and (n529,n86,n192);
and (n530,n87,n194);
or (n531,n124,n423);
and (n532,n512,n520);
xor (n533,n462,n475);
and (n534,n490,n509);
xor (n535,n408,n411);
and (n536,n486,n487);
nand (n537,n538,n539);
xor (n538,n485,n535);
or (n539,n540,n589);
and (n540,n541,n544);
xor (n541,n542,n543);
xor (n542,n413,n430);
xor (n543,n489,n533);
or (n544,n545,n588);
and (n545,n546,n587);
xor (n546,n547,n561);
and (n547,n548,n554);
and (n548,n549,n100);
nand (n549,n550,n551);
or (n550,n76,n110);
nand (n551,n552,n419);
or (n552,n553,n75);
not (n553,n110);
nand (n554,n555,n560);
or (n555,n556,n217);
not (n556,n557);
nand (n557,n558,n559);
or (n558,n48,n101);
or (n559,n52,n102);
or (n560,n40,n496);
or (n561,n562,n586);
and (n562,n563,n579);
xor (n563,n564,n572);
nand (n564,n565,n566);
or (n565,n83,n502);
nand (n566,n567,n571);
not (n567,n568);
nor (n568,n569,n570);
and (n569,n274,n76);
and (n570,n207,n75);
not (n571,n78);
nand (n572,n573,n578);
or (n573,n574,n105);
not (n574,n575);
nand (n575,n576,n577);
or (n576,n100,n419);
or (n577,n104,n350);
nand (n578,n515,n108);
nand (n579,n580,n585);
or (n580,n581,n37);
not (n581,n582);
nor (n582,n583,n584);
and (n583,n73,n28);
and (n584,n24,n74);
or (n585,n522,n19);
and (n586,n564,n572);
xor (n587,n492,n500);
and (n588,n547,n561);
and (n589,n542,n543);
nand (n590,n403,n483);
not (n591,n592);
nor (n592,n593,n608);
nor (n593,n594,n605);
xor (n594,n595,n602);
xor (n595,n596,n601);
nand (n596,n597,n599);
or (n597,n255,n598);
not (n598,n224);
or (n599,n224,n600);
not (n600,n255);
xor (n601,n334,n337);
or (n602,n603,n604);
and (n603,n450,n453);
and (n604,n451,n452);
or (n605,n606,n607);
and (n606,n404,n449);
and (n607,n405,n406);
nor (n608,n609,n610);
xor (n609,n329,n332);
or (n610,n611,n612);
and (n611,n595,n602);
and (n612,n596,n601);
nor (n613,n614,n619);
and (n614,n615,n616);
not (n615,n608);
nor (n616,n617,n618);
not (n617,n594);
not (n618,n605);
and (n619,n609,n610);
nand (n620,n592,n621,n910);
nand (n621,n622,n898,n909);
nand (n622,n623,n661,n760);
nand (n623,n624,n626);
not (n624,n625);
xor (n625,n541,n544);
not (n626,n627);
or (n627,n628,n660);
and (n628,n629,n659);
xor (n629,n630,n631);
xor (n630,n511,n526);
or (n631,n632,n658);
and (n632,n633,n641);
xor (n633,n634,n640);
nand (n634,n635,n639);
or (n635,n123,n636);
nor (n636,n637,n638);
and (n637,n86,n185);
and (n638,n87,n188);
or (n639,n528,n124);
xor (n640,n548,n554);
or (n641,n642,n657);
and (n642,n643,n651);
xor (n643,n644,n645);
and (n644,n108,n350);
nand (n645,n646,n647);
or (n646,n19,n581);
or (n647,n648,n37);
nor (n648,n649,n650);
and (n649,n28,n119);
and (n650,n24,n118);
nand (n651,n652,n656);
or (n652,n78,n653);
nor (n653,n654,n655);
and (n654,n75,n277);
and (n655,n76,n387);
or (n656,n83,n568);
and (n657,n644,n645);
and (n658,n634,n640);
xor (n659,n546,n587);
and (n660,n630,n631);
nor (n661,n662,n755);
not (n662,n663);
nor (n663,n664,n728);
nor (n664,n665,n700);
xor (n665,n666,n699);
xor (n666,n667,n668);
xor (n667,n563,n579);
or (n668,n669,n698);
and (n669,n670,n684);
xor (n670,n671,n678);
nand (n671,n672,n677);
or (n672,n673,n217);
not (n673,n674);
nand (n674,n675,n676);
or (n675,n48,n194);
or (n676,n52,n192);
nand (n677,n41,n557);
nand (n678,n679,n683);
or (n679,n123,n680);
nor (n680,n681,n682);
and (n681,n196,n86);
and (n682,n87,n372);
or (n683,n124,n636);
and (n684,n685,n691);
nor (n685,n686,n75);
nor (n686,n687,n689);
and (n687,n688,n419);
nand (n688,n87,n81);
and (n689,n86,n690);
not (n690,n81);
nand (n691,n692,n697);
or (n692,n37,n693);
not (n693,n694);
nor (n694,n695,n696);
and (n695,n24,n102);
and (n696,n101,n28);
or (n697,n648,n19);
and (n698,n671,n678);
xor (n699,n633,n641);
or (n700,n701,n727);
and (n701,n702,n726);
xor (n702,n703,n725);
or (n703,n704,n724);
and (n704,n705,n718);
xor (n705,n706,n712);
nand (n706,n707,n711);
or (n707,n78,n708);
nor (n708,n709,n710);
and (n709,n75,n350);
and (n710,n76,n419);
or (n711,n653,n83);
nand (n712,n713,n714);
or (n713,n673,n40);
nand (n714,n60,n715);
nand (n715,n716,n717);
or (n716,n48,n188);
or (n717,n52,n185);
nand (n718,n719,n723);
or (n719,n123,n720);
nor (n720,n721,n722);
and (n721,n86,n207);
and (n722,n87,n274);
or (n723,n124,n680);
and (n724,n706,n712);
xor (n725,n643,n651);
xor (n726,n670,n684);
and (n727,n703,n725);
nor (n728,n729,n730);
xor (n729,n702,n726);
or (n730,n731,n754);
and (n731,n732,n753);
xor (n732,n733,n734);
xor (n733,n685,n691);
or (n734,n735,n752);
and (n735,n736,n745);
xor (n736,n737,n738);
and (n737,n84,n350);
nand (n738,n739,n740);
or (n739,n19,n693);
or (n740,n741,n37);
not (n741,n742);
nand (n742,n743,n744);
or (n743,n192,n28);
nand (n744,n28,n192);
nand (n745,n746,n751);
or (n746,n747,n217);
not (n747,n748);
nor (n748,n749,n750);
and (n749,n48,n196);
and (n750,n372,n52);
nand (n751,n41,n715);
and (n752,n737,n738);
xor (n753,n705,n718);
and (n754,n733,n734);
nor (n755,n756,n757);
xor (n756,n629,n659);
or (n757,n758,n759);
and (n758,n666,n699);
and (n759,n667,n668);
or (n760,n761,n897);
and (n761,n762,n789);
xor (n762,n763,n788);
or (n763,n764,n787);
and (n764,n765,n786);
xor (n765,n766,n772);
nand (n766,n767,n771);
or (n767,n123,n768);
nor (n768,n769,n770);
and (n769,n86,n277);
and (n770,n87,n387);
or (n771,n124,n720);
nor (n772,n773,n781);
not (n773,n774);
nand (n774,n775,n780);
or (n775,n37,n776);
not (n776,n777);
nor (n777,n778,n779);
and (n778,n24,n185);
and (n779,n188,n28);
nand (n780,n742,n20);
nand (n781,n782,n87);
nand (n782,n783,n784);
or (n783,n48,n126);
nand (n784,n785,n419);
or (n785,n128,n52);
xor (n786,n736,n745);
and (n787,n766,n772);
xor (n788,n732,n753);
or (n789,n790,n896);
and (n790,n791,n815);
xor (n791,n792,n814);
or (n792,n793,n813);
and (n793,n794,n809);
xor (n794,n795,n802);
nand (n795,n796,n801);
or (n796,n797,n217);
not (n797,n798);
nand (n798,n799,n800);
or (n799,n48,n274);
or (n800,n52,n207);
nand (n801,n41,n748);
nand (n802,n803,n808);
or (n803,n804,n123);
not (n804,n805);
nand (n805,n806,n807);
or (n806,n419,n87);
or (n807,n86,n350);
or (n808,n124,n768);
nand (n809,n810,n812);
or (n810,n811,n773);
not (n811,n781);
or (n812,n774,n781);
and (n813,n795,n802);
xor (n814,n765,n786);
or (n815,n816,n895);
and (n816,n817,n838);
xor (n817,n818,n837);
or (n818,n819,n836);
and (n819,n820,n829);
xor (n820,n821,n822);
nor (n821,n124,n419);
nand (n822,n823,n828);
or (n823,n824,n217);
not (n824,n825);
nor (n825,n826,n827);
and (n826,n387,n52);
and (n827,n48,n277);
nand (n828,n41,n798);
nand (n829,n830,n835);
or (n830,n37,n831);
not (n831,n832);
nor (n832,n833,n834);
and (n833,n372,n28);
and (n834,n24,n196);
or (n835,n776,n19);
and (n836,n821,n822);
xor (n837,n794,n809);
or (n838,n839,n894);
and (n839,n840,n893);
xor (n840,n841,n854);
nor (n841,n842,n849);
not (n842,n843);
nand (n843,n844,n845);
or (n844,n19,n831);
nand (n845,n846,n36);
nor (n846,n847,n848);
and (n847,n274,n28);
and (n848,n24,n207);
nand (n849,n850,n48);
nand (n850,n851,n852);
or (n851,n43,n24);
or (n852,n853,n350);
and (n853,n24,n43);
nand (n854,n855,n892);
or (n855,n856,n880);
not (n856,n857);
nand (n857,n858,n879);
or (n858,n859,n868);
nor (n859,n860,n861);
and (n860,n41,n350);
nand (n861,n862,n864);
or (n862,n19,n863);
not (n863,n846);
nand (n864,n865,n36);
nand (n865,n866,n867);
or (n866,n387,n24);
or (n867,n28,n277);
nand (n868,n869,n872);
not (n869,n870);
nand (n870,n871,n24);
nand (n871,n350,n20);
nand (n872,n873,n875);
or (n873,n19,n874);
not (n874,n865);
nand (n875,n876,n36);
nor (n876,n877,n878);
and (n877,n419,n28);
and (n878,n24,n350);
nand (n879,n860,n861);
not (n880,n881);
nand (n881,n882,n886);
nor (n882,n883,n884);
and (n883,n849,n843);
and (n884,n885,n842);
not (n885,n849);
nor (n886,n887,n891);
and (n887,n60,n888);
nand (n888,n889,n890);
or (n889,n48,n419);
or (n890,n52,n350);
and (n891,n41,n825);
or (n892,n882,n886);
xor (n893,n820,n829);
and (n894,n841,n854);
and (n895,n818,n837);
and (n896,n792,n814);
and (n897,n763,n788);
nand (n898,n899,n623);
nand (n899,n900,n908);
or (n900,n755,n901);
nand (n901,n902,n907);
or (n902,n903,n905);
not (n903,n904);
nand (n904,n729,n730);
not (n905,n906);
nand (n906,n665,n700);
not (n907,n664);
nand (n908,n756,n757);
nand (n909,n625,n627);
nor (n910,n911,n402);
not (n911,n912);
or (n912,n539,n538);
and (n913,n914,n395);
not (n914,n9);
not (n915,n916);
nand (n916,n917,n3);
not (n917,n4);
wire s0n918,s1n918,notn918;
or (n918,s0n918,s1n918);
not(notn918,n4);
and (s0n918,notn918,n919);
and (s1n918,n4,1'b0);
wire s0n919,s1n919,notn919;
or (n919,s0n919,s1n919);
not(notn919,n3);
and (s0n919,notn919,n5);
and (s1n919,n3,n920);
xor (n920,n921,n1567);
xor (n921,n922,n1564);
xor (n922,n923,n23);
xor (n923,n924,n1555);
xor (n924,n925,n1554);
xor (n925,n926,n1539);
xor (n926,n927,n1538);
xor (n927,n928,n1517);
xor (n928,n929,n1516);
xor (n929,n930,n1489);
xor (n930,n931,n1488);
xor (n931,n932,n1455);
xor (n932,n933,n1454);
xor (n933,n934,n1415);
xor (n934,n935,n94);
xor (n935,n936,n1372);
xor (n936,n937,n1371);
xor (n937,n938,n1321);
xor (n938,n939,n120);
xor (n939,n940,n1265);
xor (n940,n941,n1264);
xor (n941,n942,n1201);
xor (n942,n943,n1200);
or (n943,n944,n1136);
and (n944,n945,n289);
or (n945,n946,n1074);
and (n946,n947,n195);
or (n947,n948,n1010);
and (n948,n949,n206);
and (n949,n276,n950);
or (n950,n951,n953);
and (n951,n349,n952);
and (n952,n176,n277);
and (n953,n954,n955);
xor (n954,n349,n952);
or (n955,n956,n959);
and (n956,n957,n958);
and (n957,n176,n350);
and (n958,n100,n277);
and (n959,n960,n961);
xor (n960,n957,n958);
or (n961,n962,n965);
and (n962,n963,n964);
and (n963,n100,n350);
and (n964,n110,n277);
and (n965,n966,n967);
xor (n966,n963,n964);
or (n967,n968,n971);
and (n968,n969,n970);
and (n969,n110,n350);
and (n970,n76,n277);
and (n971,n972,n973);
xor (n972,n969,n970);
or (n973,n974,n977);
and (n974,n975,n976);
and (n975,n76,n350);
and (n976,n81,n277);
and (n977,n978,n979);
xor (n978,n975,n976);
or (n979,n980,n983);
and (n980,n981,n982);
and (n981,n81,n350);
and (n982,n87,n277);
and (n983,n984,n985);
xor (n984,n981,n982);
or (n985,n986,n989);
and (n986,n987,n988);
and (n987,n87,n350);
and (n988,n126,n277);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n994);
and (n992,n993,n827);
and (n993,n126,n350);
and (n994,n995,n996);
xor (n995,n993,n827);
or (n996,n997,n1000);
and (n997,n998,n999);
and (n998,n48,n350);
and (n999,n43,n277);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
and (n1004,n43,n350);
and (n1005,n24,n277);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
and (n1008,n878,n1009);
and (n1009,n20,n277);
and (n1010,n1011,n1012);
xor (n1011,n949,n206);
or (n1012,n1013,n1016);
and (n1013,n1014,n1015);
xor (n1014,n276,n950);
and (n1015,n176,n207);
and (n1016,n1017,n1018);
xor (n1017,n1014,n1015);
or (n1018,n1019,n1022);
and (n1019,n1020,n1021);
xor (n1020,n954,n955);
and (n1021,n100,n207);
and (n1022,n1023,n1024);
xor (n1023,n1020,n1021);
or (n1024,n1025,n1028);
and (n1025,n1026,n1027);
xor (n1026,n960,n961);
and (n1027,n110,n207);
and (n1028,n1029,n1030);
xor (n1029,n1026,n1027);
or (n1030,n1031,n1034);
and (n1031,n1032,n1033);
xor (n1032,n966,n967);
and (n1033,n76,n207);
and (n1034,n1035,n1036);
xor (n1035,n1032,n1033);
or (n1036,n1037,n1040);
and (n1037,n1038,n1039);
xor (n1038,n972,n973);
and (n1039,n81,n207);
and (n1040,n1041,n1042);
xor (n1041,n1038,n1039);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n978,n979);
and (n1045,n87,n207);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n984,n985);
and (n1051,n126,n207);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n990,n991);
and (n1057,n48,n207);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
or (n1060,n1061,n1064);
and (n1061,n1062,n1063);
xor (n1062,n995,n996);
and (n1063,n43,n207);
and (n1064,n1065,n1066);
xor (n1065,n1062,n1063);
or (n1066,n1067,n1069);
and (n1067,n1068,n848);
xor (n1068,n1001,n1002);
and (n1069,n1070,n1071);
xor (n1070,n1068,n848);
and (n1071,n1072,n1073);
xor (n1072,n1007,n1008);
and (n1073,n20,n207);
and (n1074,n1075,n1076);
xor (n1075,n947,n195);
or (n1076,n1077,n1080);
and (n1077,n1078,n1079);
xor (n1078,n1011,n1012);
and (n1079,n176,n196);
and (n1080,n1081,n1082);
xor (n1081,n1078,n1079);
or (n1082,n1083,n1085);
and (n1083,n1084,n373);
xor (n1084,n1017,n1018);
and (n1085,n1086,n1087);
xor (n1086,n1084,n373);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
xor (n1089,n1023,n1024);
and (n1090,n110,n196);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
xor (n1095,n1029,n1030);
and (n1096,n76,n196);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
or (n1099,n1100,n1103);
and (n1100,n1101,n1102);
xor (n1101,n1035,n1036);
and (n1102,n81,n196);
and (n1103,n1104,n1105);
xor (n1104,n1101,n1102);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
xor (n1107,n1041,n1042);
and (n1108,n87,n196);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
xor (n1113,n1047,n1048);
and (n1114,n126,n196);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
or (n1117,n1118,n1120);
and (n1118,n1119,n749);
xor (n1119,n1053,n1054);
and (n1120,n1121,n1122);
xor (n1121,n1119,n749);
or (n1122,n1123,n1126);
and (n1123,n1124,n1125);
xor (n1124,n1059,n1060);
and (n1125,n43,n196);
and (n1126,n1127,n1128);
xor (n1127,n1124,n1125);
or (n1128,n1129,n1131);
and (n1129,n1130,n834);
xor (n1130,n1065,n1066);
and (n1131,n1132,n1133);
xor (n1132,n1130,n834);
and (n1133,n1134,n1135);
xor (n1134,n1070,n1071);
and (n1135,n20,n196);
and (n1136,n1137,n1138);
xor (n1137,n945,n289);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
xor (n1140,n1075,n1076);
and (n1141,n176,n185);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1081,n1082);
and (n1147,n100,n185);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1086,n1087);
and (n1153,n110,n185);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1092,n1093);
and (n1159,n76,n185);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1098,n1099);
and (n1165,n81,n185);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1104,n1105);
and (n1171,n87,n185);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1110,n1111);
and (n1177,n126,n185);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
xor (n1182,n1116,n1117);
and (n1183,n48,n185);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1121,n1122);
and (n1189,n43,n185);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1195);
and (n1193,n1194,n778);
xor (n1194,n1127,n1128);
and (n1195,n1196,n1197);
xor (n1196,n1194,n778);
and (n1197,n1198,n1199);
xor (n1198,n1132,n1133);
and (n1199,n20,n185);
and (n1200,n181,n192);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1137,n1138);
and (n1204,n176,n192);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1143,n1144);
and (n1210,n100,n192);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1149,n1150);
and (n1216,n110,n192);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1155,n1156);
and (n1222,n76,n192);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1161,n1162);
and (n1228,n81,n192);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1167,n1168);
and (n1234,n87,n192);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1173,n1174);
and (n1240,n126,n192);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1179,n1180);
and (n1246,n48,n192);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1185,n1186);
and (n1252,n43,n192);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
or (n1255,n1256,n1259);
and (n1256,n1257,n1258);
xor (n1257,n1191,n1192);
and (n1258,n24,n192);
and (n1259,n1260,n1261);
xor (n1260,n1257,n1258);
and (n1261,n1262,n1263);
xor (n1262,n1196,n1197);
and (n1263,n20,n192);
and (n1264,n176,n102);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1206,n1207);
and (n1268,n100,n102);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1212,n1213);
and (n1274,n110,n102);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1218,n1219);
and (n1280,n76,n102);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1224,n1225);
and (n1286,n81,n102);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1230,n1231);
and (n1292,n87,n102);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1236,n1237);
and (n1298,n126,n102);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1242,n1243);
and (n1304,n48,n102);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1248,n1249);
and (n1310,n43,n102);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1316);
and (n1314,n1315,n695);
xor (n1315,n1254,n1255);
and (n1316,n1317,n1318);
xor (n1317,n1315,n695);
and (n1318,n1319,n1320);
xor (n1319,n1260,n1261);
and (n1320,n20,n102);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1270,n1271);
and (n1324,n110,n119);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
or (n1327,n1328,n1330);
and (n1328,n1329,n244);
xor (n1329,n1276,n1277);
and (n1330,n1331,n1332);
xor (n1331,n1329,n244);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1282,n1283);
and (n1335,n81,n119);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1288,n1289);
and (n1341,n87,n119);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1294,n1295);
and (n1347,n126,n119);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1300,n1301);
and (n1353,n48,n119);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1306,n1307);
and (n1359,n43,n119);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1312,n1313);
and (n1365,n24,n119);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
and (n1368,n1369,n1370);
xor (n1369,n1317,n1318);
and (n1370,n20,n119);
and (n1371,n110,n74);
or (n1372,n1373,n1375);
and (n1373,n1374,n77);
xor (n1374,n1326,n1327);
and (n1375,n1376,n1377);
xor (n1376,n1374,n77);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1331,n1332);
and (n1380,n81,n74);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1337,n1338);
and (n1386,n87,n74);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1343,n1344);
and (n1392,n126,n74);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1349,n1350);
and (n1398,n48,n74);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
or (n1401,n1402,n1405);
and (n1402,n1403,n1404);
xor (n1403,n1355,n1356);
and (n1404,n43,n74);
and (n1405,n1406,n1407);
xor (n1406,n1403,n1404);
or (n1407,n1408,n1410);
and (n1408,n1409,n584);
xor (n1409,n1361,n1362);
and (n1410,n1411,n1412);
xor (n1411,n1409,n584);
and (n1412,n1413,n1414);
xor (n1413,n1367,n1368);
and (n1414,n20,n74);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1376,n1377);
and (n1418,n81,n93);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1382,n1383);
and (n1424,n87,n93);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1388,n1389);
and (n1430,n126,n93);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
or (n1433,n1434,n1437);
and (n1434,n1435,n1436);
xor (n1435,n1394,n1395);
and (n1436,n48,n93);
and (n1437,n1438,n1439);
xor (n1438,n1435,n1436);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1400,n1401);
and (n1442,n43,n93);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1406,n1407);
and (n1448,n24,n93);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
and (n1451,n1452,n1453);
xor (n1452,n1411,n1412);
and (n1453,n20,n93);
and (n1454,n81,n134);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1420,n1421);
and (n1458,n87,n134);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1426,n1427);
and (n1464,n126,n134);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1432,n1433);
and (n1470,n48,n134);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1438,n1439);
and (n1476,n43,n134);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1444,n1445);
and (n1482,n24,n134);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
and (n1485,n1486,n1487);
xor (n1486,n1450,n1451);
and (n1487,n20,n134);
and (n1488,n87,n140);
or (n1489,n1490,n1493);
and (n1490,n1491,n1492);
xor (n1491,n1460,n1461);
and (n1492,n126,n140);
and (n1493,n1494,n1495);
xor (n1494,n1491,n1492);
or (n1495,n1496,n1499);
and (n1496,n1497,n1498);
xor (n1497,n1466,n1467);
and (n1498,n48,n140);
and (n1499,n1500,n1501);
xor (n1500,n1497,n1498);
or (n1501,n1502,n1505);
and (n1502,n1503,n1504);
xor (n1503,n1472,n1473);
and (n1504,n43,n140);
and (n1505,n1506,n1507);
xor (n1506,n1503,n1504);
or (n1507,n1508,n1511);
and (n1508,n1509,n1510);
xor (n1509,n1478,n1479);
and (n1510,n24,n140);
and (n1511,n1512,n1513);
xor (n1512,n1509,n1510);
and (n1513,n1514,n1515);
xor (n1514,n1484,n1485);
and (n1515,n20,n140);
and (n1516,n126,n57);
or (n1517,n1518,n1521);
and (n1518,n1519,n1520);
xor (n1519,n1494,n1495);
and (n1520,n48,n57);
and (n1521,n1522,n1523);
xor (n1522,n1519,n1520);
or (n1523,n1524,n1527);
and (n1524,n1525,n1526);
xor (n1525,n1500,n1501);
and (n1526,n43,n57);
and (n1527,n1528,n1529);
xor (n1528,n1525,n1526);
or (n1529,n1530,n1533);
and (n1530,n1531,n1532);
xor (n1531,n1506,n1507);
and (n1532,n24,n57);
and (n1533,n1534,n1535);
xor (n1534,n1531,n1532);
and (n1535,n1536,n1537);
xor (n1536,n1512,n1513);
and (n1537,n20,n57);
and (n1538,n48,n50);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1522,n1523);
and (n1542,n43,n50);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1528,n1529);
and (n1548,n24,n50);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
and (n1551,n1552,n1553);
xor (n1552,n1534,n1535);
and (n1553,n20,n50);
and (n1554,n43,n33);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1544,n1545);
and (n1558,n24,n33);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
and (n1561,n1562,n1563);
xor (n1562,n1550,n1551);
and (n1563,n20,n33);
and (n1564,n1565,n1566);
xor (n1565,n1560,n1561);
and (n1566,n20,n25);
and (n1567,n20,n296);
endmodule
