module top (out,n4,n5,n6,n26,n28,n35,n36,n46,n54
        ,n55,n61,n62,n70,n83,n87,n90,n96,n105,n106
        ,n108,n113,n114,n118,n125,n133,n139,n148,n159,n165
        ,n174,n182,n184,n189,n195,n209,n220,n227);
output out;
input n4;
input n5;
input n6;
input n26;
input n28;
input n35;
input n36;
input n46;
input n54;
input n55;
input n61;
input n62;
input n70;
input n83;
input n87;
input n90;
input n96;
input n105;
input n106;
input n108;
input n113;
input n114;
input n118;
input n125;
input n133;
input n139;
input n148;
input n159;
input n165;
input n174;
input n182;
input n184;
input n189;
input n195;
input n209;
input n220;
input n227;
wire n0;
wire n1;
wire n2;
wire n3;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
xor (out,n0,n1019);
not (n0,n1);
nor (n1,n2,n7);
and (n2,n3,n6);
nor (n3,n4,n5);
and (n7,n8,n1016);
nand (n8,n9,n1015);
or (n9,n10,n502);
not (n10,n11);
nand (n11,n12,n501);
not (n12,n13);
nor (n13,n14,n440);
xor (n14,n15,n370);
xor (n15,n16,n229);
xor (n16,n17,n151);
xor (n17,n18,n99);
xor (n18,n19,n77);
xor (n19,n20,n48);
nand (n20,n21,n42);
or (n21,n22,n30);
not (n22,n23);
nor (n23,n24,n29);
and (n24,n25,n27);
not (n25,n26);
not (n27,n28);
and (n29,n26,n28);
not (n30,n31);
nor (n31,n32,n38);
nand (n32,n33,n37);
or (n33,n34,n36);
not (n34,n35);
nand (n37,n36,n34);
nor (n38,n39,n41);
and (n39,n40,n28);
not (n40,n36);
and (n41,n36,n27);
nand (n42,n32,n43);
nand (n43,n44,n47);
or (n44,n45,n28);
not (n45,n46);
or (n47,n27,n46);
nand (n48,n49,n65);
or (n49,n50,n57);
not (n50,n51);
nand (n51,n52,n56);
or (n52,n53,n55);
not (n53,n54);
nand (n56,n55,n53);
not (n57,n58);
nand (n58,n59,n63);
or (n59,n60,n62);
not (n60,n61);
or (n63,n64,n61);
not (n64,n62);
nand (n65,n66,n72);
not (n66,n67);
nor (n67,n68,n71);
and (n68,n62,n69);
not (n69,n70);
and (n71,n64,n70);
not (n72,n73);
nand (n73,n50,n74);
nand (n74,n75,n76);
nand (n75,n53,n62);
nand (n76,n54,n64);
nand (n77,n78,n93);
or (n78,n79,n88);
nand (n79,n80,n85);
nor (n80,n81,n84);
and (n81,n82,n62);
not (n82,n83);
and (n84,n83,n64);
xor (n85,n82,n86);
not (n86,n87);
nor (n88,n89,n91);
and (n89,n90,n86);
and (n91,n87,n92);
not (n92,n90);
or (n93,n94,n80);
nor (n94,n95,n97);
and (n95,n96,n86);
and (n97,n87,n98);
not (n98,n96);
xor (n99,n100,n127);
xor (n100,n101,n109);
and (n101,n102,n108);
nand (n102,n103,n107);
or (n103,n104,n106);
not (n104,n105);
nand (n107,n106,n104);
nand (n109,n110,n121);
or (n110,n111,n115);
nand (n111,n112,n114);
not (n112,n113);
nor (n115,n116,n119);
and (n116,n117,n118);
not (n117,n114);
and (n119,n114,n120);
not (n120,n118);
nand (n121,n122,n113);
nor (n122,n123,n126);
and (n123,n124,n117);
not (n124,n125);
and (n126,n125,n114);
nand (n127,n128,n141);
or (n128,n129,n135);
not (n129,n130);
nor (n130,n131,n134);
and (n131,n132,n34);
not (n132,n133);
and (n134,n133,n35);
not (n135,n136);
nand (n136,n137,n140);
or (n137,n138,n114);
not (n138,n139);
nand (n140,n138,n114);
or (n141,n142,n146);
nand (n142,n135,n143);
nand (n143,n144,n145);
or (n144,n35,n138);
nand (n145,n138,n35);
nor (n146,n147,n149);
and (n147,n34,n148);
and (n149,n35,n150);
not (n150,n148);
xor (n151,n152,n203);
xor (n152,n153,n176);
nand (n153,n154,n170);
or (n154,n155,n161);
not (n155,n156);
nor (n156,n157,n160);
and (n157,n158,n104);
not (n158,n159);
and (n160,n159,n105);
nand (n161,n162,n167);
not (n162,n163);
nand (n163,n164,n166);
or (n164,n86,n165);
nand (n166,n86,n165);
nand (n167,n168,n169);
or (n168,n165,n104);
nand (n169,n104,n165);
nand (n170,n163,n171);
nor (n171,n172,n175);
and (n172,n173,n104);
not (n173,n174);
and (n175,n174,n105);
nand (n176,n177,n191);
or (n177,n178,n186);
not (n178,n179);
nor (n179,n180,n185);
and (n180,n181,n183);
not (n181,n182);
not (n183,n184);
and (n185,n182,n184);
not (n186,n187);
nand (n187,n188,n190);
or (n188,n27,n189);
nand (n190,n189,n27);
nand (n191,n192,n198);
not (n192,n193);
nor (n193,n194,n196);
and (n194,n183,n195);
and (n196,n184,n197);
not (n197,n195);
not (n198,n199);
nand (n199,n200,n186);
nand (n200,n201,n202);
or (n201,n189,n183);
nand (n202,n183,n189);
nand (n203,n204,n222);
or (n204,n205,n216);
not (n205,n206);
nor (n206,n207,n213);
nor (n207,n208,n211);
and (n208,n209,n210);
not (n210,n55);
and (n211,n55,n212);
not (n212,n209);
nand (n213,n214,n215);
or (n214,n183,n209);
nand (n215,n209,n183);
not (n216,n217);
nor (n217,n218,n221);
and (n218,n219,n210);
not (n219,n220);
and (n221,n220,n55);
or (n222,n223,n224);
not (n223,n213);
nor (n224,n225,n228);
and (n225,n226,n55);
not (n226,n227);
and (n228,n227,n210);
or (n229,n230,n369);
and (n230,n231,n308);
xor (n231,n232,n271);
or (n232,n233,n270);
and (n233,n234,n253);
xor (n234,n235,n244);
nand (n235,n236,n240);
or (n236,n73,n237);
nor (n237,n238,n239);
and (n238,n64,n90);
and (n239,n62,n92);
or (n240,n50,n241);
nor (n241,n242,n243);
and (n242,n64,n96);
and (n243,n62,n98);
nand (n244,n245,n249);
or (n245,n79,n246);
nor (n246,n247,n248);
and (n247,n86,n159);
and (n248,n87,n158);
or (n249,n80,n250);
nor (n250,n251,n252);
and (n251,n86,n174);
and (n252,n87,n173);
and (n253,n254,n260);
nor (n254,n255,n86);
nor (n255,n256,n258);
and (n256,n257,n64);
nand (n257,n108,n83);
and (n258,n259,n82);
not (n259,n108);
nand (n260,n261,n266);
or (n261,n111,n262);
not (n262,n263);
nor (n263,n264,n265);
and (n264,n45,n117);
and (n265,n46,n114);
or (n266,n112,n267);
nor (n267,n268,n269);
and (n268,n117,n148);
and (n269,n114,n150);
and (n270,n235,n244);
xor (n271,n272,n290);
xor (n272,n273,n276);
nand (n273,n274,n275);
or (n274,n79,n250);
or (n275,n80,n88);
xor (n276,n277,n283);
nor (n277,n278,n104);
nor (n278,n279,n281);
and (n279,n280,n86);
nand (n280,n108,n165);
and (n281,n259,n282);
not (n282,n165);
nand (n283,n284,n289);
or (n284,n111,n285);
not (n285,n286);
nor (n286,n287,n288);
and (n287,n133,n114);
and (n288,n132,n117);
or (n289,n115,n112);
or (n290,n291,n307);
and (n291,n292,n297);
xor (n292,n293,n294);
nor (n293,n162,n259);
nand (n294,n295,n296);
or (n295,n112,n285);
or (n296,n267,n111);
nand (n297,n298,n303);
or (n298,n135,n299);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n46,n35);
and (n302,n45,n34);
or (n303,n142,n304);
nor (n304,n305,n306);
and (n305,n26,n34);
and (n306,n25,n35);
and (n307,n293,n294);
or (n308,n309,n368);
and (n309,n310,n367);
xor (n310,n311,n341);
or (n311,n312,n340);
and (n312,n313,n331);
xor (n313,n314,n321);
nand (n314,n315,n319);
or (n315,n142,n316);
nor (n316,n317,n318);
and (n317,n182,n34);
and (n318,n181,n35);
nand (n319,n320,n136);
not (n320,n304);
nand (n321,n322,n327);
or (n322,n323,n186);
not (n323,n324);
nor (n324,n325,n326);
and (n325,n220,n184);
and (n326,n219,n183);
or (n327,n199,n328);
nor (n328,n329,n330);
and (n329,n60,n184);
and (n330,n61,n183);
nand (n331,n332,n336);
or (n332,n205,n333);
nor (n333,n334,n335);
and (n334,n210,n96);
and (n335,n98,n55);
or (n336,n223,n337);
nor (n337,n338,n339);
and (n338,n210,n70);
and (n339,n55,n69);
and (n340,n314,n321);
or (n341,n342,n366);
and (n342,n343,n360);
xor (n343,n344,n354);
nand (n344,n345,n349);
or (n345,n346,n30);
nor (n346,n347,n348);
and (n347,n27,n227);
and (n348,n28,n226);
nand (n349,n350,n32);
not (n350,n351);
nor (n351,n352,n353);
and (n352,n27,n195);
and (n353,n28,n197);
nand (n354,n355,n359);
or (n355,n73,n356);
nor (n356,n357,n358);
and (n357,n64,n174);
and (n358,n62,n173);
or (n359,n50,n237);
nand (n360,n361,n365);
or (n361,n79,n362);
nor (n362,n363,n364);
and (n363,n259,n87);
and (n364,n108,n86);
or (n365,n246,n80);
and (n366,n344,n354);
xor (n367,n292,n297);
and (n368,n311,n341);
and (n369,n232,n271);
xor (n370,n371,n421);
xor (n371,n372,n375);
or (n372,n373,n374);
and (n373,n272,n290);
and (n374,n273,n276);
xor (n375,n376,n400);
xor (n376,n377,n378);
and (n377,n277,n283);
or (n378,n379,n399);
and (n379,n380,n392);
xor (n380,n381,n385);
nand (n381,n382,n383);
or (n382,n299,n142);
nand (n383,n384,n136);
not (n384,n146);
nand (n385,n386,n391);
or (n386,n387,n161);
not (n387,n388);
nand (n388,n389,n390);
or (n389,n104,n108);
or (n390,n259,n105);
nand (n391,n163,n156);
nand (n392,n393,n398);
or (n393,n199,n394);
not (n394,n395);
nor (n395,n396,n397);
and (n396,n227,n184);
and (n397,n226,n183);
or (n398,n186,n193);
and (n399,n381,n385);
or (n400,n401,n420);
and (n401,n402,n417);
xor (n402,n403,n410);
nand (n403,n404,n409);
or (n404,n405,n205);
not (n405,n406);
nor (n406,n407,n408);
and (n407,n60,n210);
and (n408,n61,n55);
nand (n409,n213,n217);
nand (n410,n411,n413);
or (n411,n22,n412);
not (n412,n32);
or (n413,n30,n414);
nor (n414,n415,n416);
and (n415,n27,n182);
and (n416,n28,n181);
nand (n417,n418,n419);
or (n418,n73,n241);
or (n419,n50,n67);
and (n420,n403,n410);
or (n421,n422,n439);
and (n422,n423,n438);
xor (n423,n424,n437);
or (n424,n425,n436);
and (n425,n426,n433);
xor (n426,n427,n430);
nand (n427,n428,n429);
or (n428,n323,n199);
nand (n429,n187,n395);
nand (n430,n431,n432);
or (n431,n205,n337);
nand (n432,n213,n406);
nand (n433,n434,n435);
or (n434,n30,n351);
or (n435,n412,n414);
and (n436,n427,n430);
xor (n437,n402,n417);
xor (n438,n380,n392);
and (n439,n424,n437);
or (n440,n441,n500);
and (n441,n442,n499);
xor (n442,n443,n444);
xor (n443,n423,n438);
or (n444,n445,n498);
and (n445,n446,n449);
xor (n446,n447,n448);
xor (n447,n426,n433);
xor (n448,n234,n253);
or (n449,n450,n497);
and (n450,n451,n472);
xor (n451,n452,n453);
xor (n452,n254,n260);
or (n453,n454,n471);
and (n454,n455,n464);
xor (n455,n456,n457);
nor (n456,n80,n259);
nand (n457,n458,n462);
or (n458,n142,n459);
nor (n459,n460,n461);
and (n460,n195,n34);
and (n461,n197,n35);
nand (n462,n463,n136);
not (n463,n316);
nand (n464,n465,n470);
or (n465,n199,n466);
not (n466,n467);
nor (n467,n468,n469);
and (n468,n69,n183);
and (n469,n70,n184);
or (n470,n186,n328);
and (n471,n456,n457);
or (n472,n473,n496);
and (n473,n474,n490);
xor (n474,n475,n483);
nand (n475,n476,n481);
or (n476,n477,n205);
not (n477,n478);
nand (n478,n479,n480);
or (n479,n55,n92);
or (n480,n90,n210);
nand (n481,n482,n213);
not (n482,n333);
nand (n483,n484,n489);
or (n484,n111,n485);
not (n485,n486);
nor (n486,n487,n488);
and (n487,n25,n117);
and (n488,n26,n114);
nand (n489,n263,n113);
nand (n490,n491,n495);
or (n491,n73,n492);
nor (n492,n493,n494);
and (n493,n64,n159);
and (n494,n62,n158);
or (n495,n50,n356);
and (n496,n475,n483);
and (n497,n452,n453);
and (n498,n447,n448);
xor (n499,n231,n308);
and (n500,n443,n444);
nand (n501,n14,n440);
not (n502,n503);
nand (n503,n504,n719);
nor (n504,n505,n718);
and (n505,n506,n570);
nand (n506,n507,n509);
not (n507,n508);
xor (n508,n442,n499);
not (n509,n510);
or (n510,n511,n569);
and (n511,n512,n515);
xor (n512,n513,n514);
xor (n513,n310,n367);
xor (n514,n446,n449);
or (n515,n516,n568);
and (n516,n517,n520);
xor (n517,n518,n519);
xor (n518,n343,n360);
xor (n519,n313,n331);
or (n520,n521,n567);
and (n521,n522,n543);
xor (n522,n523,n529);
nand (n523,n524,n528);
or (n524,n30,n525);
nor (n525,n526,n527);
and (n526,n27,n220);
and (n527,n28,n219);
or (n528,n412,n346);
and (n529,n530,n536);
nand (n530,n531,n532);
or (n531,n459,n135);
or (n532,n142,n533);
nor (n533,n534,n535);
and (n534,n227,n34);
and (n535,n226,n35);
not (n536,n537);
nand (n537,n538,n62);
nand (n538,n539,n540);
or (n539,n108,n54);
nand (n540,n541,n210);
not (n541,n542);
and (n542,n108,n54);
or (n543,n544,n566);
and (n544,n545,n560);
xor (n545,n546,n553);
nand (n546,n547,n552);
or (n547,n548,n199);
not (n548,n549);
nand (n549,n550,n551);
or (n550,n184,n98);
or (n551,n183,n96);
nand (n552,n187,n467);
nand (n553,n554,n559);
or (n554,n555,n205);
not (n555,n556);
nand (n556,n557,n558);
or (n557,n55,n173);
or (n558,n210,n174);
nand (n559,n213,n478);
nand (n560,n561,n562);
or (n561,n112,n485);
or (n562,n563,n111);
nor (n563,n564,n565);
and (n564,n117,n182);
and (n565,n114,n181);
and (n566,n546,n553);
and (n567,n523,n529);
and (n568,n518,n519);
and (n569,n513,n514);
nand (n570,n571,n717);
or (n571,n572,n709);
not (n572,n573);
nand (n573,n574,n708);
or (n574,n575,n658);
nor (n575,n576,n606);
xor (n576,n577,n605);
xor (n577,n578,n579);
xor (n578,n451,n472);
or (n579,n580,n604);
and (n580,n581,n584);
xor (n581,n582,n583);
xor (n582,n474,n490);
xor (n583,n455,n464);
or (n584,n585,n603);
and (n585,n586,n599);
xor (n586,n587,n593);
nand (n587,n588,n592);
or (n588,n73,n589);
nor (n589,n590,n591);
and (n590,n259,n62);
and (n591,n108,n64);
or (n592,n50,n492);
nand (n593,n594,n598);
or (n594,n30,n595);
nor (n595,n596,n597);
and (n596,n27,n61);
and (n597,n28,n60);
or (n598,n412,n525);
nand (n599,n600,n602);
or (n600,n536,n601);
not (n601,n530);
or (n602,n530,n537);
and (n603,n587,n593);
and (n604,n582,n583);
xor (n605,n517,n520);
or (n606,n607,n657);
and (n607,n608,n656);
xor (n608,n609,n610);
xor (n609,n522,n543);
or (n610,n611,n655);
and (n611,n612,n654);
xor (n612,n613,n631);
or (n613,n614,n630);
and (n614,n615,n624);
xor (n615,n616,n617);
nor (n616,n50,n259);
nand (n617,n618,n622);
or (n618,n619,n142);
nor (n619,n620,n621);
and (n620,n34,n220);
and (n621,n35,n219);
nand (n622,n623,n136);
not (n623,n533);
nand (n624,n625,n626);
or (n625,n548,n186);
or (n626,n199,n627);
nor (n627,n628,n629);
and (n628,n183,n90);
and (n629,n184,n92);
and (n630,n616,n617);
or (n631,n632,n653);
and (n632,n633,n647);
xor (n633,n634,n641);
nand (n634,n635,n640);
or (n635,n636,n205);
not (n636,n637);
nand (n637,n638,n639);
or (n638,n55,n158);
or (n639,n210,n159);
nand (n640,n213,n556);
nand (n641,n642,n646);
or (n642,n643,n111);
nor (n643,n644,n645);
and (n644,n117,n195);
and (n645,n114,n197);
or (n646,n563,n112);
nand (n647,n648,n652);
or (n648,n30,n649);
nor (n649,n650,n651);
and (n650,n27,n70);
and (n651,n28,n69);
or (n652,n412,n595);
and (n653,n634,n641);
xor (n654,n545,n560);
and (n655,n613,n631);
xor (n656,n581,n584);
and (n657,n609,n610);
nand (n658,n659,n707);
or (n659,n660,n706);
and (n660,n661,n664);
xor (n661,n662,n663);
xor (n662,n586,n599);
xor (n663,n612,n654);
or (n664,n665,n705);
and (n665,n666,n704);
xor (n666,n667,n680);
and (n667,n668,n674);
and (n668,n669,n55);
nand (n669,n670,n671);
or (n670,n108,n209);
nand (n671,n672,n183);
not (n672,n673);
and (n673,n108,n209);
nand (n674,n675,n679);
or (n675,n142,n676);
nor (n676,n677,n678);
and (n677,n34,n61);
and (n678,n35,n60);
or (n679,n135,n619);
or (n680,n681,n703);
and (n681,n682,n697);
xor (n682,n683,n690);
nand (n683,n684,n688);
or (n684,n685,n199);
nor (n685,n686,n687);
and (n686,n183,n174);
and (n687,n184,n173);
nand (n688,n689,n187);
not (n689,n627);
nand (n690,n691,n692);
or (n691,n636,n223);
nand (n692,n693,n206);
not (n693,n694);
nor (n694,n695,n696);
and (n695,n259,n55);
and (n696,n210,n108);
nand (n697,n698,n702);
or (n698,n111,n699);
nor (n699,n700,n701);
and (n700,n117,n227);
and (n701,n114,n226);
or (n702,n643,n112);
and (n703,n683,n690);
xor (n704,n615,n624);
and (n705,n667,n680);
and (n706,n662,n663);
xor (n707,n608,n656);
nand (n708,n576,n606);
not (n709,n710);
nand (n710,n711,n713);
not (n711,n712);
xor (n712,n512,n515);
not (n713,n714);
or (n714,n715,n716);
and (n715,n577,n605);
and (n716,n578,n579);
nand (n717,n712,n714);
nor (n718,n507,n509);
nand (n719,n720,n506,n1011);
nand (n720,n721,n1010);
or (n721,n722,n759);
not (n722,n723);
or (n723,n724,n725);
xor (n724,n661,n664);
or (n725,n726,n758);
and (n726,n727,n757);
xor (n727,n728,n729);
xor (n728,n633,n647);
or (n729,n730,n756);
and (n730,n731,n739);
xor (n731,n732,n738);
nand (n732,n733,n737);
or (n733,n30,n734);
nor (n734,n735,n736);
and (n735,n27,n96);
and (n736,n28,n98);
or (n737,n412,n649);
xor (n738,n668,n674);
or (n739,n740,n755);
and (n740,n741,n749);
xor (n741,n742,n743);
nor (n742,n223,n259);
nand (n743,n744,n748);
or (n744,n745,n111);
nor (n745,n746,n747);
and (n746,n219,n114);
and (n747,n220,n117);
or (n748,n699,n112);
nand (n749,n750,n754);
or (n750,n199,n751);
nor (n751,n752,n753);
and (n752,n183,n159);
and (n753,n184,n158);
or (n754,n186,n685);
and (n755,n742,n743);
and (n756,n732,n738);
xor (n757,n666,n704);
and (n758,n728,n729);
not (n759,n760);
or (n760,n761,n1009);
and (n761,n762,n802);
xor (n762,n763,n801);
or (n763,n764,n800);
and (n764,n765,n799);
xor (n765,n766,n767);
xor (n766,n682,n697);
or (n767,n768,n798);
and (n768,n769,n784);
xor (n769,n770,n778);
nand (n770,n771,n776);
or (n771,n772,n142);
not (n772,n773);
nand (n773,n774,n775);
or (n774,n35,n69);
or (n775,n34,n70);
nand (n776,n777,n136);
not (n777,n676);
nand (n778,n779,n783);
or (n779,n30,n780);
nor (n780,n781,n782);
and (n781,n27,n90);
and (n782,n28,n92);
or (n783,n412,n734);
and (n784,n785,n791);
nor (n785,n786,n183);
nor (n786,n787,n789);
and (n787,n259,n788);
not (n788,n189);
nor (n789,n790,n28);
and (n790,n108,n189);
nand (n791,n792,n797);
or (n792,n111,n793);
not (n793,n794);
nor (n794,n795,n796);
and (n795,n60,n117);
and (n796,n61,n114);
or (n797,n745,n112);
and (n798,n770,n778);
xor (n799,n731,n739);
and (n800,n766,n767);
xor (n801,n727,n757);
nand (n802,n803,n1006,n1008);
nand (n803,n804,n839,n999);
nand (n804,n805,n807);
not (n805,n806);
xor (n806,n765,n799);
not (n807,n808);
or (n808,n809,n838);
and (n809,n810,n837);
xor (n810,n811,n836);
or (n811,n812,n835);
and (n812,n813,n829);
xor (n813,n814,n822);
nand (n814,n815,n820);
or (n815,n816,n199);
not (n816,n817);
nand (n817,n818,n819);
or (n818,n183,n108);
or (n819,n259,n184);
nand (n820,n821,n187);
not (n821,n751);
nand (n822,n823,n828);
or (n823,n824,n142);
not (n824,n825);
nand (n825,n826,n827);
or (n826,n35,n98);
or (n827,n34,n96);
nand (n828,n136,n773);
nand (n829,n830,n834);
or (n830,n30,n831);
nor (n831,n832,n833);
and (n832,n27,n174);
and (n833,n28,n173);
or (n834,n412,n780);
and (n835,n814,n822);
xor (n836,n741,n749);
xor (n837,n769,n784);
and (n838,n811,n836);
nand (n839,n840,n998);
or (n840,n841,n891);
not (n841,n842);
nand (n842,n843,n867);
not (n843,n844);
xor (n844,n845,n866);
xor (n845,n846,n847);
xor (n846,n785,n791);
or (n847,n848,n865);
and (n848,n849,n858);
xor (n849,n850,n851);
and (n850,n187,n108);
nand (n851,n852,n857);
or (n852,n111,n853);
not (n853,n854);
nor (n854,n855,n856);
and (n855,n69,n117);
and (n856,n70,n114);
nand (n857,n794,n113);
nand (n858,n859,n864);
or (n859,n860,n142);
not (n860,n861);
nor (n861,n862,n863);
and (n862,n92,n34);
and (n863,n90,n35);
nand (n864,n136,n825);
and (n865,n850,n851);
xor (n866,n813,n829);
not (n867,n868);
or (n868,n869,n890);
and (n869,n870,n889);
xor (n870,n871,n877);
nand (n871,n872,n876);
or (n872,n30,n873);
nor (n873,n874,n875);
and (n874,n158,n28);
and (n875,n159,n27);
or (n876,n412,n831);
and (n877,n878,n883);
and (n878,n879,n28);
nand (n879,n880,n882);
or (n880,n881,n35);
and (n881,n108,n36);
or (n882,n108,n36);
nand (n883,n884,n885);
or (n884,n112,n853);
or (n885,n886,n111);
nor (n886,n887,n888);
and (n887,n117,n96);
and (n888,n114,n98);
xor (n889,n849,n858);
and (n890,n871,n877);
not (n891,n892);
nand (n892,n893,n997);
or (n893,n894,n917);
not (n894,n895);
nand (n895,n896,n898);
not (n896,n897);
xor (n897,n870,n889);
not (n898,n899);
or (n899,n900,n916);
and (n900,n901,n915);
xor (n901,n902,n909);
nand (n902,n903,n908);
or (n903,n904,n142);
not (n904,n905);
nor (n905,n906,n907);
and (n906,n173,n34);
and (n907,n174,n35);
nand (n908,n861,n136);
nand (n909,n910,n911);
or (n910,n412,n873);
nand (n911,n31,n912);
nand (n912,n913,n914);
or (n913,n108,n27);
or (n914,n259,n28);
xor (n915,n878,n883);
and (n916,n902,n909);
not (n917,n918);
or (n918,n919,n996);
and (n919,n920,n941);
xor (n920,n921,n940);
or (n921,n922,n939);
and (n922,n923,n932);
xor (n923,n924,n925);
and (n924,n32,n108);
nand (n925,n926,n931);
or (n926,n927,n142);
not (n927,n928);
nor (n928,n929,n930);
and (n929,n158,n34);
and (n930,n159,n35);
nand (n931,n905,n136);
nand (n932,n933,n938);
or (n933,n111,n934);
not (n934,n935);
nor (n935,n936,n937);
and (n936,n92,n117);
and (n937,n90,n114);
or (n938,n886,n112);
and (n939,n924,n925);
xor (n940,n901,n915);
nand (n941,n942,n995);
or (n942,n943,n959);
nor (n943,n944,n945);
xor (n944,n923,n932);
nor (n945,n946,n954);
not (n946,n947);
nand (n947,n948,n949);
or (n948,n112,n934);
nand (n949,n950,n953);
nand (n950,n951,n952);
or (n951,n174,n117);
nand (n952,n117,n174);
not (n953,n111);
nand (n954,n955,n35);
nand (n955,n956,n958);
or (n956,n957,n114);
and (n957,n108,n139);
or (n958,n108,n139);
nor (n959,n960,n994);
and (n960,n961,n973);
nand (n961,n962,n969);
not (n962,n963);
nand (n963,n964,n968);
or (n964,n142,n965);
nor (n965,n966,n967);
and (n966,n35,n259);
and (n967,n108,n34);
or (n968,n135,n927);
nor (n969,n970,n971);
and (n970,n954,n947);
and (n971,n972,n946);
not (n972,n954);
or (n973,n974,n993);
and (n974,n975,n984);
xor (n975,n976,n977);
nor (n976,n135,n259);
nand (n977,n978,n983);
or (n978,n111,n979);
not (n979,n980);
nand (n980,n981,n982);
or (n981,n158,n114);
nand (n982,n114,n158);
nand (n983,n950,n113);
nor (n984,n985,n991);
nor (n985,n986,n987);
and (n986,n980,n113);
nor (n987,n988,n111);
nor (n988,n989,n990);
and (n989,n259,n114);
and (n990,n108,n117);
or (n991,n992,n117);
and (n992,n108,n113);
and (n993,n976,n977);
nor (n994,n962,n969);
nand (n995,n944,n945);
and (n996,n921,n940);
nand (n997,n897,n899);
nand (n998,n844,n868);
nand (n999,n1000,n1004);
not (n1000,n1001);
or (n1001,n1002,n1003);
and (n1002,n845,n866);
and (n1003,n846,n847);
not (n1004,n1005);
xor (n1005,n810,n837);
nand (n1006,n804,n1007);
and (n1007,n1005,n1001);
nand (n1008,n808,n806);
and (n1009,n763,n801);
nand (n1010,n724,n725);
nor (n1011,n709,n1012);
nand (n1012,n1013,n1014);
not (n1013,n575);
or (n1014,n659,n707);
or (n1015,n503,n11);
not (n1016,n1017);
nand (n1017,n1018,n4);
not (n1018,n5);
wire s0n1019,s1n1019,notn1019;
or (n1019,s0n1019,s1n1019);
not(notn1019,n5);
and (s0n1019,notn1019,n1020);
and (s1n1019,n5,1'b0);
wire s0n1020,s1n1020,notn1020;
or (n1020,s0n1020,s1n1020);
not(notn1020,n4);
and (s0n1020,notn1020,n6);
and (s1n1020,n4,n1021);
xor (n1021,n1022,n1721);
xor (n1022,n1023,n1718);
xor (n1023,n1024,n160);
xor (n1024,n1025,n1709);
xor (n1025,n1026,n1708);
xor (n1026,n1027,n1693);
xor (n1027,n1028,n1692);
xor (n1028,n1029,n1671);
xor (n1029,n1030,n1670);
xor (n1030,n1031,n1643);
xor (n1031,n1032,n1642);
xor (n1032,n1033,n1610);
xor (n1033,n1034,n1609);
xor (n1034,n1035,n1571);
xor (n1035,n1036,n221);
xor (n1036,n1037,n1527);
xor (n1037,n1038,n1526);
xor (n1038,n1039,n1478);
xor (n1039,n1040,n1477);
xor (n1040,n1041,n1421);
xor (n1041,n1042,n1420);
xor (n1042,n1043,n1357);
xor (n1043,n1044,n29);
xor (n1044,n1045,n1289);
xor (n1045,n1046,n1288);
xor (n1046,n1047,n1217);
xor (n1047,n1048,n1216);
xor (n1048,n1049,n1136);
xor (n1049,n1050,n1135);
xor (n1050,n1051,n1054);
xor (n1051,n1052,n1053);
and (n1052,n125,n113);
and (n1053,n118,n114);
or (n1054,n1055,n1057);
and (n1055,n1056,n287);
and (n1056,n118,n113);
and (n1057,n1058,n1059);
xor (n1058,n1056,n287);
or (n1059,n1060,n1063);
and (n1060,n1061,n1062);
and (n1061,n133,n113);
and (n1062,n148,n114);
and (n1063,n1064,n1065);
xor (n1064,n1061,n1062);
or (n1065,n1066,n1068);
and (n1066,n1067,n265);
and (n1067,n148,n113);
and (n1068,n1069,n1070);
xor (n1069,n1067,n265);
or (n1070,n1071,n1073);
and (n1071,n1072,n488);
and (n1072,n46,n113);
and (n1073,n1074,n1075);
xor (n1074,n1072,n488);
or (n1075,n1076,n1079);
and (n1076,n1077,n1078);
and (n1077,n26,n113);
and (n1078,n182,n114);
and (n1079,n1080,n1081);
xor (n1080,n1077,n1078);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
and (n1083,n182,n113);
and (n1084,n195,n114);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
and (n1089,n195,n113);
and (n1090,n227,n114);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
and (n1095,n227,n113);
and (n1096,n220,n114);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
or (n1099,n1100,n1102);
and (n1100,n1101,n796);
and (n1101,n220,n113);
and (n1102,n1103,n1104);
xor (n1103,n1101,n796);
or (n1104,n1105,n1107);
and (n1105,n1106,n856);
and (n1106,n61,n113);
and (n1107,n1108,n1109);
xor (n1108,n1106,n856);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n70,n113);
and (n1112,n96,n114);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1118);
and (n1116,n1117,n937);
and (n1117,n96,n113);
and (n1118,n1119,n1120);
xor (n1119,n1117,n937);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
and (n1122,n90,n113);
and (n1123,n174,n114);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
and (n1128,n174,n113);
and (n1129,n159,n114);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
and (n1132,n1133,n1134);
and (n1133,n159,n113);
and (n1134,n108,n114);
and (n1135,n133,n139);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1058,n1059);
and (n1139,n148,n139);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1064,n1065);
and (n1145,n46,n139);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1069,n1070);
and (n1151,n26,n139);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1074,n1075);
and (n1157,n182,n139);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1080,n1081);
and (n1163,n195,n139);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1086,n1087);
and (n1169,n227,n139);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
or (n1172,n1173,n1176);
and (n1173,n1174,n1175);
xor (n1174,n1092,n1093);
and (n1175,n220,n139);
and (n1176,n1177,n1178);
xor (n1177,n1174,n1175);
or (n1178,n1179,n1182);
and (n1179,n1180,n1181);
xor (n1180,n1098,n1099);
and (n1181,n61,n139);
and (n1182,n1183,n1184);
xor (n1183,n1180,n1181);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1103,n1104);
and (n1187,n70,n139);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1108,n1109);
and (n1193,n96,n139);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
or (n1196,n1197,n1200);
and (n1197,n1198,n1199);
xor (n1198,n1114,n1115);
and (n1199,n90,n139);
and (n1200,n1201,n1202);
xor (n1201,n1198,n1199);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
xor (n1204,n1119,n1120);
and (n1205,n174,n139);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
or (n1208,n1209,n1212);
and (n1209,n1210,n1211);
xor (n1210,n1125,n1126);
and (n1211,n159,n139);
and (n1212,n1213,n1214);
xor (n1213,n1210,n1211);
and (n1214,n1215,n957);
xor (n1215,n1131,n1132);
and (n1216,n148,n35);
or (n1217,n1218,n1220);
and (n1218,n1219,n301);
xor (n1219,n1141,n1142);
and (n1220,n1221,n1222);
xor (n1221,n1219,n301);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1147,n1148);
and (n1225,n26,n35);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1153,n1154);
and (n1231,n182,n35);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1159,n1160);
and (n1237,n195,n35);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1165,n1166);
and (n1243,n227,n35);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1171,n1172);
and (n1249,n220,n35);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1177,n1178);
and (n1255,n61,n35);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1183,n1184);
and (n1261,n70,n35);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1189,n1190);
and (n1267,n96,n35);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1273);
and (n1271,n1272,n863);
xor (n1272,n1195,n1196);
and (n1273,n1274,n1275);
xor (n1274,n1272,n863);
or (n1275,n1276,n1278);
and (n1276,n1277,n907);
xor (n1277,n1201,n1202);
and (n1278,n1279,n1280);
xor (n1279,n1277,n907);
or (n1280,n1281,n1283);
and (n1281,n1282,n930);
xor (n1282,n1207,n1208);
and (n1283,n1284,n1285);
xor (n1284,n1282,n930);
and (n1285,n1286,n1287);
xor (n1286,n1213,n1214);
and (n1287,n108,n35);
and (n1288,n46,n36);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1221,n1222);
and (n1292,n26,n36);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1227,n1228);
and (n1298,n182,n36);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1233,n1234);
and (n1304,n195,n36);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1239,n1240);
and (n1310,n227,n36);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1245,n1246);
and (n1316,n220,n36);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1251,n1252);
and (n1322,n61,n36);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
or (n1325,n1326,n1329);
and (n1326,n1327,n1328);
xor (n1327,n1257,n1258);
and (n1328,n70,n36);
and (n1329,n1330,n1331);
xor (n1330,n1327,n1328);
or (n1331,n1332,n1335);
and (n1332,n1333,n1334);
xor (n1333,n1263,n1264);
and (n1334,n96,n36);
and (n1335,n1336,n1337);
xor (n1336,n1333,n1334);
or (n1337,n1338,n1341);
and (n1338,n1339,n1340);
xor (n1339,n1269,n1270);
and (n1340,n90,n36);
and (n1341,n1342,n1343);
xor (n1342,n1339,n1340);
or (n1343,n1344,n1347);
and (n1344,n1345,n1346);
xor (n1345,n1274,n1275);
and (n1346,n174,n36);
and (n1347,n1348,n1349);
xor (n1348,n1345,n1346);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1279,n1280);
and (n1352,n159,n36);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
and (n1355,n1356,n881);
xor (n1356,n1284,n1285);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1294,n1295);
and (n1360,n182,n28);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1300,n1301);
and (n1366,n195,n28);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1306,n1307);
and (n1372,n227,n28);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1312,n1313);
and (n1378,n220,n28);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1318,n1319);
and (n1384,n61,n28);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1324,n1325);
and (n1390,n70,n28);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1330,n1331);
and (n1396,n96,n28);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1336,n1337);
and (n1402,n90,n28);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1342,n1343);
and (n1408,n174,n28);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1348,n1349);
and (n1414,n159,n28);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
and (n1417,n1418,n1419);
xor (n1418,n1354,n1355);
and (n1419,n108,n28);
and (n1420,n182,n189);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1362,n1363);
and (n1424,n195,n189);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1368,n1369);
and (n1430,n227,n189);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
or (n1433,n1434,n1437);
and (n1434,n1435,n1436);
xor (n1435,n1374,n1375);
and (n1436,n220,n189);
and (n1437,n1438,n1439);
xor (n1438,n1435,n1436);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1380,n1381);
and (n1442,n61,n189);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1386,n1387);
and (n1448,n70,n189);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1392,n1393);
and (n1454,n96,n189);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
or (n1457,n1458,n1461);
and (n1458,n1459,n1460);
xor (n1459,n1398,n1399);
and (n1460,n90,n189);
and (n1461,n1462,n1463);
xor (n1462,n1459,n1460);
or (n1463,n1464,n1467);
and (n1464,n1465,n1466);
xor (n1465,n1404,n1405);
and (n1466,n174,n189);
and (n1467,n1468,n1469);
xor (n1468,n1465,n1466);
or (n1469,n1470,n1473);
and (n1470,n1471,n1472);
xor (n1471,n1410,n1411);
and (n1472,n159,n189);
and (n1473,n1474,n1475);
xor (n1474,n1471,n1472);
and (n1475,n1476,n790);
xor (n1476,n1416,n1417);
and (n1477,n195,n184);
or (n1478,n1479,n1481);
and (n1479,n1480,n396);
xor (n1480,n1426,n1427);
and (n1481,n1482,n1483);
xor (n1482,n1480,n396);
or (n1483,n1484,n1486);
and (n1484,n1485,n325);
xor (n1485,n1432,n1433);
and (n1486,n1487,n1488);
xor (n1487,n1485,n325);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1438,n1439);
and (n1491,n61,n184);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1497);
and (n1495,n1496,n469);
xor (n1496,n1444,n1445);
and (n1497,n1498,n1499);
xor (n1498,n1496,n469);
or (n1499,n1500,n1503);
and (n1500,n1501,n1502);
xor (n1501,n1450,n1451);
and (n1502,n96,n184);
and (n1503,n1504,n1505);
xor (n1504,n1501,n1502);
or (n1505,n1506,n1509);
and (n1506,n1507,n1508);
xor (n1507,n1456,n1457);
and (n1508,n90,n184);
and (n1509,n1510,n1511);
xor (n1510,n1507,n1508);
or (n1511,n1512,n1515);
and (n1512,n1513,n1514);
xor (n1513,n1462,n1463);
and (n1514,n174,n184);
and (n1515,n1516,n1517);
xor (n1516,n1513,n1514);
or (n1517,n1518,n1521);
and (n1518,n1519,n1520);
xor (n1519,n1468,n1469);
and (n1520,n159,n184);
and (n1521,n1522,n1523);
xor (n1522,n1519,n1520);
and (n1523,n1524,n1525);
xor (n1524,n1474,n1475);
and (n1525,n108,n184);
and (n1526,n227,n209);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1482,n1483);
and (n1530,n220,n209);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1487,n1488);
and (n1536,n61,n209);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1493,n1494);
and (n1542,n70,n209);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1498,n1499);
and (n1548,n96,n209);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1504,n1505);
and (n1554,n90,n209);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1510,n1511);
and (n1560,n174,n209);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1516,n1517);
and (n1566,n159,n209);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
and (n1569,n1570,n673);
xor (n1570,n1522,n1523);
or (n1571,n1572,n1574);
and (n1572,n1573,n408);
xor (n1573,n1532,n1533);
and (n1574,n1575,n1576);
xor (n1575,n1573,n408);
or (n1576,n1577,n1580);
and (n1577,n1578,n1579);
xor (n1578,n1538,n1539);
and (n1579,n70,n55);
and (n1580,n1581,n1582);
xor (n1581,n1578,n1579);
or (n1582,n1583,n1586);
and (n1583,n1584,n1585);
xor (n1584,n1544,n1545);
and (n1585,n96,n55);
and (n1586,n1587,n1588);
xor (n1587,n1584,n1585);
or (n1588,n1589,n1592);
and (n1589,n1590,n1591);
xor (n1590,n1550,n1551);
and (n1591,n90,n55);
and (n1592,n1593,n1594);
xor (n1593,n1590,n1591);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1556,n1557);
and (n1597,n174,n55);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1562,n1563);
and (n1603,n159,n55);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
and (n1606,n1607,n1608);
xor (n1607,n1568,n1569);
and (n1608,n108,n55);
and (n1609,n61,n54);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1575,n1576);
and (n1613,n70,n54);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
xor (n1618,n1581,n1582);
and (n1619,n96,n54);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
xor (n1624,n1587,n1588);
and (n1625,n90,n54);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1593,n1594);
and (n1631,n174,n54);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1599,n1600);
and (n1637,n159,n54);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
and (n1640,n1641,n542);
xor (n1641,n1605,n1606);
and (n1642,n70,n62);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1615,n1616);
and (n1646,n96,n62);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1621,n1622);
and (n1652,n90,n62);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1627,n1628);
and (n1658,n174,n62);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1633,n1634);
and (n1664,n159,n62);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
and (n1667,n1668,n1669);
xor (n1668,n1639,n1640);
and (n1669,n108,n62);
and (n1670,n96,n83);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1648,n1649);
and (n1674,n90,n83);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1654,n1655);
and (n1680,n174,n83);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1660,n1661);
and (n1686,n159,n83);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
and (n1689,n1690,n1691);
xor (n1690,n1666,n1667);
not (n1691,n257);
and (n1692,n90,n87);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1676,n1677);
and (n1696,n174,n87);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1682,n1683);
and (n1702,n159,n87);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
and (n1705,n1706,n1707);
xor (n1706,n1688,n1689);
and (n1707,n108,n87);
and (n1708,n174,n165);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1698,n1699);
and (n1712,n159,n165);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
and (n1715,n1716,n1717);
xor (n1716,n1704,n1705);
not (n1717,n280);
and (n1718,n1719,n1720);
xor (n1719,n1714,n1715);
and (n1720,n108,n105);
and (n1721,n108,n106);
endmodule
