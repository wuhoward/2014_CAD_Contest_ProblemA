module top (out,n14,n19,n21,n22,n24,n28,n31,n37,n55
        ,n69,n70,n71,n72,n73,n74,n75,n76,n80,n81
        ,n82,n86,n88,n90,n127,n129,n130,n131,n142,n143
        ,n144,n145,n157,n158,n159,n160,n173,n174,n175,n176
        ,n182,n184,n185,n188,n190,n193,n195,n196,n197,n277
        ,n383,n386,n388,n542,n544,n545,n548,n551,n552,n553
        ,n554,n557,n559,n563,n574,n575,n592,n595,n597,n598
        ,n600,n604,n610,n613,n615,n617,n621,n624,n626,n628
        ,n632,n635,n637,n639,n641,n649,n652,n654,n656,n660
        ,n663,n665,n667,n671,n674,n676,n678,n682,n685,n687
        ,n689,n697,n700,n702,n704,n708,n711,n713,n715,n719
        ,n722,n724,n726,n730,n733,n735,n737,n746,n749,n751
        ,n753,n767,n770,n772,n774,n793,n796,n798,n800,n809
        ,n812,n814,n816,n830,n833,n835,n837,n860,n863,n865
        ,n867,n883,n886,n888,n890,n935,n938,n940,n942,n946
        ,n949,n951,n953,n957,n960,n962,n964,n968,n971,n973
        ,n975,n984,n987,n989,n991,n995,n998,n1000,n1002,n1006
        ,n1009,n1011,n1013,n1017,n1020,n1022,n1024,n1032,n1035,n1037
        ,n1039,n1043,n1046,n1048,n1050,n1054,n1057,n1059,n1061,n1065
        ,n1068,n1070,n1072,n1297,n1300,n1302,n1304,n1313,n1316,n1318
        ,n1320,n1329,n1332,n1334,n1336,n1345,n1348,n1350,n1352,n1361
        ,n1364,n1366,n1368,n1377,n1380,n1382,n1384,n1394,n1397,n1399
        ,n1401,n1409,n1412,n1414,n1416,n1824,n1827,n1829,n1831,n1841
        ,n1844,n1846,n1848,n1858,n1861,n1863,n1865,n1883,n1886,n1888
        ,n1890,n1910,n1913,n1915,n1917,n1936,n1939,n1941,n1943,n1965
        ,n1968,n1970,n1972,n1984,n1987,n1989,n1991,n2161,n2164,n2166
        ,n2168,n2177,n2180,n2182,n2184,n2193,n2196,n2198,n2200,n2209
        ,n2212,n2214,n2216,n2225,n2228,n2230,n2232,n2241,n2244,n2246
        ,n2248,n2257,n2260,n2262,n2264,n2272,n2275,n2277,n2279,n2703
        ,n2705,n2707,n2709,n2715,n2717,n2719,n2721,n2727,n2729,n2731
        ,n2733,n2739,n2741,n2882,n2893,n2920,n2946,n2954,n2963,n2974
        ,n2977,n2980,n2983,n2988,n2991,n2994,n2997,n3002,n3005,n3008
        ,n3011,n3017,n3018,n3032,n3033,n3051,n3052,n3055,n3056,n3059
        ,n3060,n3063,n3064,n3069,n3070,n3073,n3074,n3077,n3078,n3081
        ,n3082,n3087,n3088,n3091,n3092,n3095,n3096,n3099,n3100,n3105
        ,n3106,n3109,n3110,n3113,n3116,n3122,n3123,n3137,n3138,n3156
        ,n3157,n3160,n3161,n3164,n3165,n3168,n3169,n3174,n3175,n3178
        ,n3179,n3182,n3183,n3186,n3187,n3192,n3193,n3196,n3197,n3200
        ,n3201,n3204,n3205,n3210,n3211,n3214,n3215,n3218,n3221,n3227
        ,n3228,n3242,n3243,n3261,n3262,n3265,n3266,n3269,n3270,n3273
        ,n3274,n3279,n3280,n3283,n3284,n3287,n3288,n3291,n3292,n3297
        ,n3298,n3301,n3302,n3305,n3306,n3309,n3310,n3315,n3316,n3319
        ,n3320,n3323,n3326,n3332,n3333,n3347,n3348,n3366,n3367,n3370
        ,n3371,n3374,n3375,n3378,n3379,n3384,n3385,n3388,n3389,n3392
        ,n3393,n3396,n3397,n3402,n3403,n3406,n3407,n3410,n3411,n3414
        ,n3415,n3420,n3421,n3424,n3425,n3428,n3431,n3437,n3438,n3452
        ,n3453,n3471,n3472,n3475,n3476,n3479,n3480,n3483,n3484,n3489
        ,n3490,n3493,n3494,n3497,n3498,n3501,n3502,n3507,n3508,n3511
        ,n3512,n3515,n3516,n3519,n3520,n3525,n3526,n3529,n3530,n3533
        ,n3536,n3542,n3543,n3557,n3558,n3576,n3577,n3580,n3581,n3584
        ,n3585,n3588,n3589,n3594,n3595,n3598,n3599,n3602,n3603,n3606
        ,n3607,n3612,n3613,n3616,n3617,n3620,n3621,n3624,n3625,n3630
        ,n3631,n3634,n3635,n3638,n3641,n3647,n3648,n3662,n3663,n3680
        ,n3681,n3684,n3685,n3688,n3689,n3692,n3693,n3698,n3699,n3702
        ,n3703,n3706,n3707,n3710,n3711,n3716,n3717,n3720,n3721,n3724
        ,n3725,n3728,n3729,n3734,n3735,n3738,n3739,n3742,n3745,n3751
        ,n3752,n3766,n3767,n3808,n3809,n3823,n3829,n3830,n3844,n3845
        ,n3872,n3873,n3887,n3893,n3894,n3908,n3909,n3936,n3937,n3951
        ,n3957,n3958,n3972,n3973,n4000,n4001,n4015,n4021,n4022,n4036
        ,n4037,n4065,n4066,n4080,n4086,n4087,n4102,n4103,n4132,n4133
        ,n4148,n4154,n4155,n4169,n4170,n4197,n4198,n4212,n4218,n4219
        ,n4233,n4234,n4261,n4262,n4277,n4283,n4284,n4299,n4300,n4418
        ,n4419,n4429,n4435,n4436,n4446,n4447,n4465,n4466,n4476,n4482
        ,n4483,n4493,n4494,n4512,n4513,n4523,n4529,n4530,n4540,n4541
        ,n4559,n4560,n4570,n4576,n4577,n4587,n4588,n4606,n4607,n4617
        ,n4623,n4624,n4633,n4634,n4651,n4652,n4662,n4668,n4669,n4679
        ,n4680,n4698,n4699,n4709,n4715,n4716,n4726,n4727,n4744,n4745
        ,n4755,n4761,n4762,n4772,n4773,n5020,n5030,n5034,n5036,n5041
        ,n5043,n5048,n5050,n5055,n5057,n5067,n5068,n5082,n5087,n5092
        ,n5099,n5102,n5105,n5108,n5113,n5114,n5117,n5120,n5123,n5128
        ,n5131,n5136,n5143,n5144,n5147,n5150,n5153,n5158,n5161,n5164
        ,n5167,n5172,n5173,n5176,n5179,n5182,n5187,n5190,n5193,n5196
        ,n5197,n5207,n5208,n5211,n5214,n5217,n5222,n5225,n5228,n5231
        ,n5236,n5237,n5240,n5243,n5246,n5251,n5254,n5259,n5266,n5267
        ,n5270,n5273,n5276,n5281,n5284,n5287,n5290,n5295,n5296,n5299
        ,n5302,n5305,n5310,n5313,n5316,n5319,n5320,n5330,n5331,n5334
        ,n5337,n5340,n5345,n5348,n5351,n5354,n5359,n5360,n5363,n5366
        ,n5369,n5374,n5377,n5382,n5389,n5390,n5393,n5396,n5399,n5404
        ,n5407,n5410,n5413,n5418,n5419,n5422,n5425,n5428,n5433,n5436
        ,n5439,n5442,n5443,n5453,n5454,n5457,n5460,n5463,n5468,n5471
        ,n5474,n5477,n5482,n5483,n5486,n5489,n5492,n5497,n5500,n5505
        ,n5512,n5513,n5516,n5519,n5522,n5527,n5530,n5533,n5536,n5541
        ,n5542,n5545,n5548,n5551,n5556,n5559,n5562,n5565,n5566,n5576
        ,n5577,n5580,n5583,n5586,n5591,n5594,n5597,n5600,n5605,n5606
        ,n5609,n5612,n5615,n5620,n5623,n5628,n5635,n5636,n5639,n5642
        ,n5645,n5650,n5653,n5656,n5659,n5664,n5665,n5668,n5671,n5674
        ,n5679,n5682,n5685,n5688,n5689,n5699,n5700,n5703,n5706,n5709
        ,n5714,n5717,n5720,n5723,n5728,n5729,n5732,n5735,n5738,n5743
        ,n5746,n5751,n5758,n5759,n5762,n5765,n5768,n5773,n5776,n5779
        ,n5782,n5787,n5788,n5791,n5794,n5797,n5802,n5805,n5808,n5811
        ,n5812,n5822,n5823,n5826,n5829,n5832,n5837,n5840,n5843,n5846
        ,n5851,n5852,n5855,n5858,n5861,n5866,n5869,n5874,n5881,n5882
        ,n5885,n5888,n5891,n5896,n5899,n5902,n5905,n5910,n5911,n5914
        ,n5917,n5920,n5925,n5928,n5931,n5934,n5935,n5944,n5945,n5948
        ,n5951,n5954,n5959,n5962,n5965,n5968,n5973,n5974,n5977,n5980
        ,n5983,n5988,n5991,n5996,n6003,n6004,n6007,n6010,n6013,n6018
        ,n6021,n6024,n6027,n6032,n6033,n6036,n6039,n6042,n6047,n6050
        ,n6053,n6056,n6057,n6075,n6077,n6081,n6083,n6088,n6090,n6136
        ,n6179,n6225,n6268,n6314,n6357,n6403,n6446,n6492,n6535,n6581
        ,n6624,n6670,n6713,n6758,n6801,n6820,n6822,n6825,n6827,n6831
        ,n6833,n6836,n6838,n6850,n6851,n6854,n6857,n6860,n6865,n6868
        ,n6873,n6880,n6881,n6884,n6887,n6890,n6895,n6898,n6901,n6904
        ,n6907,n6919,n6920,n6923,n6926,n6929,n6934,n6937,n6942,n6949
        ,n6950,n6953,n6956,n6959,n6964,n6967,n6970,n6973,n6976,n6988
        ,n6989,n6992,n6995,n6998,n7003,n7006,n7011,n7018,n7019,n7022
        ,n7025,n7028,n7033,n7036,n7039,n7042,n7045,n7057,n7058,n7061
        ,n7064,n7067,n7072,n7075,n7080,n7087,n7088,n7091,n7094,n7097
        ,n7102,n7105,n7108,n7111,n7114,n7126,n7127,n7130,n7133,n7136
        ,n7141,n7144,n7149,n7156,n7157,n7160,n7163,n7166,n7171,n7174
        ,n7177,n7180,n7183,n7195,n7196,n7199,n7202,n7205,n7210,n7213
        ,n7218,n7225,n7226,n7229,n7232,n7235,n7240,n7243,n7246,n7249
        ,n7252,n7264,n7265,n7268,n7271,n7274,n7279,n7282,n7287,n7294
        ,n7295,n7298,n7301,n7304,n7309,n7312,n7315,n7318,n7321,n7332
        ,n7333,n7336,n7339,n7342,n7347,n7350,n7355,n7362,n7363,n7366
        ,n7369,n7372,n7377,n7380,n7383,n7386,n7389,n7415,n7417,n7786
        ,n7788,n7795,n7797,n7811,n7813,n7820,n7822,n7827,n7829,n7834
        ,n7836,n7856,n7858,n7861,n7863,n8056,n8059,n8168,n8171,n8280
        ,n8283,n8392,n8395,n8500,n8503,n8608,n8611,n8715,n8718);
output out;
input n14;
input n19;
input n21;
input n22;
input n24;
input n28;
input n31;
input n37;
input n55;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n80;
input n81;
input n82;
input n86;
input n88;
input n90;
input n127;
input n129;
input n130;
input n131;
input n142;
input n143;
input n144;
input n145;
input n157;
input n158;
input n159;
input n160;
input n173;
input n174;
input n175;
input n176;
input n182;
input n184;
input n185;
input n188;
input n190;
input n193;
input n195;
input n196;
input n197;
input n277;
input n383;
input n386;
input n388;
input n542;
input n544;
input n545;
input n548;
input n551;
input n552;
input n553;
input n554;
input n557;
input n559;
input n563;
input n574;
input n575;
input n592;
input n595;
input n597;
input n598;
input n600;
input n604;
input n610;
input n613;
input n615;
input n617;
input n621;
input n624;
input n626;
input n628;
input n632;
input n635;
input n637;
input n639;
input n641;
input n649;
input n652;
input n654;
input n656;
input n660;
input n663;
input n665;
input n667;
input n671;
input n674;
input n676;
input n678;
input n682;
input n685;
input n687;
input n689;
input n697;
input n700;
input n702;
input n704;
input n708;
input n711;
input n713;
input n715;
input n719;
input n722;
input n724;
input n726;
input n730;
input n733;
input n735;
input n737;
input n746;
input n749;
input n751;
input n753;
input n767;
input n770;
input n772;
input n774;
input n793;
input n796;
input n798;
input n800;
input n809;
input n812;
input n814;
input n816;
input n830;
input n833;
input n835;
input n837;
input n860;
input n863;
input n865;
input n867;
input n883;
input n886;
input n888;
input n890;
input n935;
input n938;
input n940;
input n942;
input n946;
input n949;
input n951;
input n953;
input n957;
input n960;
input n962;
input n964;
input n968;
input n971;
input n973;
input n975;
input n984;
input n987;
input n989;
input n991;
input n995;
input n998;
input n1000;
input n1002;
input n1006;
input n1009;
input n1011;
input n1013;
input n1017;
input n1020;
input n1022;
input n1024;
input n1032;
input n1035;
input n1037;
input n1039;
input n1043;
input n1046;
input n1048;
input n1050;
input n1054;
input n1057;
input n1059;
input n1061;
input n1065;
input n1068;
input n1070;
input n1072;
input n1297;
input n1300;
input n1302;
input n1304;
input n1313;
input n1316;
input n1318;
input n1320;
input n1329;
input n1332;
input n1334;
input n1336;
input n1345;
input n1348;
input n1350;
input n1352;
input n1361;
input n1364;
input n1366;
input n1368;
input n1377;
input n1380;
input n1382;
input n1384;
input n1394;
input n1397;
input n1399;
input n1401;
input n1409;
input n1412;
input n1414;
input n1416;
input n1824;
input n1827;
input n1829;
input n1831;
input n1841;
input n1844;
input n1846;
input n1848;
input n1858;
input n1861;
input n1863;
input n1865;
input n1883;
input n1886;
input n1888;
input n1890;
input n1910;
input n1913;
input n1915;
input n1917;
input n1936;
input n1939;
input n1941;
input n1943;
input n1965;
input n1968;
input n1970;
input n1972;
input n1984;
input n1987;
input n1989;
input n1991;
input n2161;
input n2164;
input n2166;
input n2168;
input n2177;
input n2180;
input n2182;
input n2184;
input n2193;
input n2196;
input n2198;
input n2200;
input n2209;
input n2212;
input n2214;
input n2216;
input n2225;
input n2228;
input n2230;
input n2232;
input n2241;
input n2244;
input n2246;
input n2248;
input n2257;
input n2260;
input n2262;
input n2264;
input n2272;
input n2275;
input n2277;
input n2279;
input n2703;
input n2705;
input n2707;
input n2709;
input n2715;
input n2717;
input n2719;
input n2721;
input n2727;
input n2729;
input n2731;
input n2733;
input n2739;
input n2741;
input n2882;
input n2893;
input n2920;
input n2946;
input n2954;
input n2963;
input n2974;
input n2977;
input n2980;
input n2983;
input n2988;
input n2991;
input n2994;
input n2997;
input n3002;
input n3005;
input n3008;
input n3011;
input n3017;
input n3018;
input n3032;
input n3033;
input n3051;
input n3052;
input n3055;
input n3056;
input n3059;
input n3060;
input n3063;
input n3064;
input n3069;
input n3070;
input n3073;
input n3074;
input n3077;
input n3078;
input n3081;
input n3082;
input n3087;
input n3088;
input n3091;
input n3092;
input n3095;
input n3096;
input n3099;
input n3100;
input n3105;
input n3106;
input n3109;
input n3110;
input n3113;
input n3116;
input n3122;
input n3123;
input n3137;
input n3138;
input n3156;
input n3157;
input n3160;
input n3161;
input n3164;
input n3165;
input n3168;
input n3169;
input n3174;
input n3175;
input n3178;
input n3179;
input n3182;
input n3183;
input n3186;
input n3187;
input n3192;
input n3193;
input n3196;
input n3197;
input n3200;
input n3201;
input n3204;
input n3205;
input n3210;
input n3211;
input n3214;
input n3215;
input n3218;
input n3221;
input n3227;
input n3228;
input n3242;
input n3243;
input n3261;
input n3262;
input n3265;
input n3266;
input n3269;
input n3270;
input n3273;
input n3274;
input n3279;
input n3280;
input n3283;
input n3284;
input n3287;
input n3288;
input n3291;
input n3292;
input n3297;
input n3298;
input n3301;
input n3302;
input n3305;
input n3306;
input n3309;
input n3310;
input n3315;
input n3316;
input n3319;
input n3320;
input n3323;
input n3326;
input n3332;
input n3333;
input n3347;
input n3348;
input n3366;
input n3367;
input n3370;
input n3371;
input n3374;
input n3375;
input n3378;
input n3379;
input n3384;
input n3385;
input n3388;
input n3389;
input n3392;
input n3393;
input n3396;
input n3397;
input n3402;
input n3403;
input n3406;
input n3407;
input n3410;
input n3411;
input n3414;
input n3415;
input n3420;
input n3421;
input n3424;
input n3425;
input n3428;
input n3431;
input n3437;
input n3438;
input n3452;
input n3453;
input n3471;
input n3472;
input n3475;
input n3476;
input n3479;
input n3480;
input n3483;
input n3484;
input n3489;
input n3490;
input n3493;
input n3494;
input n3497;
input n3498;
input n3501;
input n3502;
input n3507;
input n3508;
input n3511;
input n3512;
input n3515;
input n3516;
input n3519;
input n3520;
input n3525;
input n3526;
input n3529;
input n3530;
input n3533;
input n3536;
input n3542;
input n3543;
input n3557;
input n3558;
input n3576;
input n3577;
input n3580;
input n3581;
input n3584;
input n3585;
input n3588;
input n3589;
input n3594;
input n3595;
input n3598;
input n3599;
input n3602;
input n3603;
input n3606;
input n3607;
input n3612;
input n3613;
input n3616;
input n3617;
input n3620;
input n3621;
input n3624;
input n3625;
input n3630;
input n3631;
input n3634;
input n3635;
input n3638;
input n3641;
input n3647;
input n3648;
input n3662;
input n3663;
input n3680;
input n3681;
input n3684;
input n3685;
input n3688;
input n3689;
input n3692;
input n3693;
input n3698;
input n3699;
input n3702;
input n3703;
input n3706;
input n3707;
input n3710;
input n3711;
input n3716;
input n3717;
input n3720;
input n3721;
input n3724;
input n3725;
input n3728;
input n3729;
input n3734;
input n3735;
input n3738;
input n3739;
input n3742;
input n3745;
input n3751;
input n3752;
input n3766;
input n3767;
input n3808;
input n3809;
input n3823;
input n3829;
input n3830;
input n3844;
input n3845;
input n3872;
input n3873;
input n3887;
input n3893;
input n3894;
input n3908;
input n3909;
input n3936;
input n3937;
input n3951;
input n3957;
input n3958;
input n3972;
input n3973;
input n4000;
input n4001;
input n4015;
input n4021;
input n4022;
input n4036;
input n4037;
input n4065;
input n4066;
input n4080;
input n4086;
input n4087;
input n4102;
input n4103;
input n4132;
input n4133;
input n4148;
input n4154;
input n4155;
input n4169;
input n4170;
input n4197;
input n4198;
input n4212;
input n4218;
input n4219;
input n4233;
input n4234;
input n4261;
input n4262;
input n4277;
input n4283;
input n4284;
input n4299;
input n4300;
input n4418;
input n4419;
input n4429;
input n4435;
input n4436;
input n4446;
input n4447;
input n4465;
input n4466;
input n4476;
input n4482;
input n4483;
input n4493;
input n4494;
input n4512;
input n4513;
input n4523;
input n4529;
input n4530;
input n4540;
input n4541;
input n4559;
input n4560;
input n4570;
input n4576;
input n4577;
input n4587;
input n4588;
input n4606;
input n4607;
input n4617;
input n4623;
input n4624;
input n4633;
input n4634;
input n4651;
input n4652;
input n4662;
input n4668;
input n4669;
input n4679;
input n4680;
input n4698;
input n4699;
input n4709;
input n4715;
input n4716;
input n4726;
input n4727;
input n4744;
input n4745;
input n4755;
input n4761;
input n4762;
input n4772;
input n4773;
input n5020;
input n5030;
input n5034;
input n5036;
input n5041;
input n5043;
input n5048;
input n5050;
input n5055;
input n5057;
input n5067;
input n5068;
input n5082;
input n5087;
input n5092;
input n5099;
input n5102;
input n5105;
input n5108;
input n5113;
input n5114;
input n5117;
input n5120;
input n5123;
input n5128;
input n5131;
input n5136;
input n5143;
input n5144;
input n5147;
input n5150;
input n5153;
input n5158;
input n5161;
input n5164;
input n5167;
input n5172;
input n5173;
input n5176;
input n5179;
input n5182;
input n5187;
input n5190;
input n5193;
input n5196;
input n5197;
input n5207;
input n5208;
input n5211;
input n5214;
input n5217;
input n5222;
input n5225;
input n5228;
input n5231;
input n5236;
input n5237;
input n5240;
input n5243;
input n5246;
input n5251;
input n5254;
input n5259;
input n5266;
input n5267;
input n5270;
input n5273;
input n5276;
input n5281;
input n5284;
input n5287;
input n5290;
input n5295;
input n5296;
input n5299;
input n5302;
input n5305;
input n5310;
input n5313;
input n5316;
input n5319;
input n5320;
input n5330;
input n5331;
input n5334;
input n5337;
input n5340;
input n5345;
input n5348;
input n5351;
input n5354;
input n5359;
input n5360;
input n5363;
input n5366;
input n5369;
input n5374;
input n5377;
input n5382;
input n5389;
input n5390;
input n5393;
input n5396;
input n5399;
input n5404;
input n5407;
input n5410;
input n5413;
input n5418;
input n5419;
input n5422;
input n5425;
input n5428;
input n5433;
input n5436;
input n5439;
input n5442;
input n5443;
input n5453;
input n5454;
input n5457;
input n5460;
input n5463;
input n5468;
input n5471;
input n5474;
input n5477;
input n5482;
input n5483;
input n5486;
input n5489;
input n5492;
input n5497;
input n5500;
input n5505;
input n5512;
input n5513;
input n5516;
input n5519;
input n5522;
input n5527;
input n5530;
input n5533;
input n5536;
input n5541;
input n5542;
input n5545;
input n5548;
input n5551;
input n5556;
input n5559;
input n5562;
input n5565;
input n5566;
input n5576;
input n5577;
input n5580;
input n5583;
input n5586;
input n5591;
input n5594;
input n5597;
input n5600;
input n5605;
input n5606;
input n5609;
input n5612;
input n5615;
input n5620;
input n5623;
input n5628;
input n5635;
input n5636;
input n5639;
input n5642;
input n5645;
input n5650;
input n5653;
input n5656;
input n5659;
input n5664;
input n5665;
input n5668;
input n5671;
input n5674;
input n5679;
input n5682;
input n5685;
input n5688;
input n5689;
input n5699;
input n5700;
input n5703;
input n5706;
input n5709;
input n5714;
input n5717;
input n5720;
input n5723;
input n5728;
input n5729;
input n5732;
input n5735;
input n5738;
input n5743;
input n5746;
input n5751;
input n5758;
input n5759;
input n5762;
input n5765;
input n5768;
input n5773;
input n5776;
input n5779;
input n5782;
input n5787;
input n5788;
input n5791;
input n5794;
input n5797;
input n5802;
input n5805;
input n5808;
input n5811;
input n5812;
input n5822;
input n5823;
input n5826;
input n5829;
input n5832;
input n5837;
input n5840;
input n5843;
input n5846;
input n5851;
input n5852;
input n5855;
input n5858;
input n5861;
input n5866;
input n5869;
input n5874;
input n5881;
input n5882;
input n5885;
input n5888;
input n5891;
input n5896;
input n5899;
input n5902;
input n5905;
input n5910;
input n5911;
input n5914;
input n5917;
input n5920;
input n5925;
input n5928;
input n5931;
input n5934;
input n5935;
input n5944;
input n5945;
input n5948;
input n5951;
input n5954;
input n5959;
input n5962;
input n5965;
input n5968;
input n5973;
input n5974;
input n5977;
input n5980;
input n5983;
input n5988;
input n5991;
input n5996;
input n6003;
input n6004;
input n6007;
input n6010;
input n6013;
input n6018;
input n6021;
input n6024;
input n6027;
input n6032;
input n6033;
input n6036;
input n6039;
input n6042;
input n6047;
input n6050;
input n6053;
input n6056;
input n6057;
input n6075;
input n6077;
input n6081;
input n6083;
input n6088;
input n6090;
input n6136;
input n6179;
input n6225;
input n6268;
input n6314;
input n6357;
input n6403;
input n6446;
input n6492;
input n6535;
input n6581;
input n6624;
input n6670;
input n6713;
input n6758;
input n6801;
input n6820;
input n6822;
input n6825;
input n6827;
input n6831;
input n6833;
input n6836;
input n6838;
input n6850;
input n6851;
input n6854;
input n6857;
input n6860;
input n6865;
input n6868;
input n6873;
input n6880;
input n6881;
input n6884;
input n6887;
input n6890;
input n6895;
input n6898;
input n6901;
input n6904;
input n6907;
input n6919;
input n6920;
input n6923;
input n6926;
input n6929;
input n6934;
input n6937;
input n6942;
input n6949;
input n6950;
input n6953;
input n6956;
input n6959;
input n6964;
input n6967;
input n6970;
input n6973;
input n6976;
input n6988;
input n6989;
input n6992;
input n6995;
input n6998;
input n7003;
input n7006;
input n7011;
input n7018;
input n7019;
input n7022;
input n7025;
input n7028;
input n7033;
input n7036;
input n7039;
input n7042;
input n7045;
input n7057;
input n7058;
input n7061;
input n7064;
input n7067;
input n7072;
input n7075;
input n7080;
input n7087;
input n7088;
input n7091;
input n7094;
input n7097;
input n7102;
input n7105;
input n7108;
input n7111;
input n7114;
input n7126;
input n7127;
input n7130;
input n7133;
input n7136;
input n7141;
input n7144;
input n7149;
input n7156;
input n7157;
input n7160;
input n7163;
input n7166;
input n7171;
input n7174;
input n7177;
input n7180;
input n7183;
input n7195;
input n7196;
input n7199;
input n7202;
input n7205;
input n7210;
input n7213;
input n7218;
input n7225;
input n7226;
input n7229;
input n7232;
input n7235;
input n7240;
input n7243;
input n7246;
input n7249;
input n7252;
input n7264;
input n7265;
input n7268;
input n7271;
input n7274;
input n7279;
input n7282;
input n7287;
input n7294;
input n7295;
input n7298;
input n7301;
input n7304;
input n7309;
input n7312;
input n7315;
input n7318;
input n7321;
input n7332;
input n7333;
input n7336;
input n7339;
input n7342;
input n7347;
input n7350;
input n7355;
input n7362;
input n7363;
input n7366;
input n7369;
input n7372;
input n7377;
input n7380;
input n7383;
input n7386;
input n7389;
input n7415;
input n7417;
input n7786;
input n7788;
input n7795;
input n7797;
input n7811;
input n7813;
input n7820;
input n7822;
input n7827;
input n7829;
input n7834;
input n7836;
input n7856;
input n7858;
input n7861;
input n7863;
input n8056;
input n8059;
input n8168;
input n8171;
input n8280;
input n8283;
input n8392;
input n8395;
input n8500;
input n8503;
input n8608;
input n8611;
input n8715;
input n8718;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n16;
wire n17;
wire n18;
wire n20;
wire n23;
wire n25;
wire n26;
wire n27;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n77;
wire n78;
wire n79;
wire n83;
wire n84;
wire n85;
wire n87;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n186;
wire n187;
wire n189;
wire n191;
wire n192;
wire n194;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n384;
wire n385;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n543;
wire n546;
wire n547;
wire n549;
wire n550;
wire n555;
wire n556;
wire n558;
wire n560;
wire n561;
wire n562;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n593;
wire n594;
wire n596;
wire n599;
wire n601;
wire n602;
wire n603;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n611;
wire n612;
wire n614;
wire n616;
wire n618;
wire n619;
wire n620;
wire n622;
wire n623;
wire n625;
wire n627;
wire n629;
wire n630;
wire n631;
wire n633;
wire n634;
wire n636;
wire n638;
wire n640;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n650;
wire n651;
wire n653;
wire n655;
wire n657;
wire n658;
wire n659;
wire n661;
wire n662;
wire n664;
wire n666;
wire n668;
wire n669;
wire n670;
wire n672;
wire n673;
wire n675;
wire n677;
wire n679;
wire n680;
wire n681;
wire n683;
wire n684;
wire n686;
wire n688;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n698;
wire n699;
wire n701;
wire n703;
wire n705;
wire n706;
wire n707;
wire n709;
wire n710;
wire n712;
wire n714;
wire n716;
wire n717;
wire n718;
wire n720;
wire n721;
wire n723;
wire n725;
wire n727;
wire n728;
wire n729;
wire n731;
wire n732;
wire n734;
wire n736;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n747;
wire n748;
wire n750;
wire n752;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n768;
wire n769;
wire n771;
wire n773;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n794;
wire n795;
wire n797;
wire n799;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n810;
wire n811;
wire n813;
wire n815;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n831;
wire n832;
wire n834;
wire n836;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n861;
wire n862;
wire n864;
wire n866;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n884;
wire n885;
wire n887;
wire n889;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n937;
wire n939;
wire n941;
wire n943;
wire n944;
wire n945;
wire n947;
wire n948;
wire n950;
wire n952;
wire n954;
wire n955;
wire n956;
wire n958;
wire n959;
wire n961;
wire n963;
wire n965;
wire n966;
wire n967;
wire n969;
wire n970;
wire n972;
wire n974;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n985;
wire n986;
wire n988;
wire n990;
wire n992;
wire n993;
wire n994;
wire n996;
wire n997;
wire n999;
wire n1001;
wire n1003;
wire n1004;
wire n1005;
wire n1007;
wire n1008;
wire n1010;
wire n1012;
wire n1014;
wire n1015;
wire n1016;
wire n1018;
wire n1019;
wire n1021;
wire n1023;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1033;
wire n1034;
wire n1036;
wire n1038;
wire n1040;
wire n1041;
wire n1042;
wire n1044;
wire n1045;
wire n1047;
wire n1049;
wire n1051;
wire n1052;
wire n1053;
wire n1055;
wire n1056;
wire n1058;
wire n1060;
wire n1062;
wire n1063;
wire n1064;
wire n1066;
wire n1067;
wire n1069;
wire n1071;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1298;
wire n1299;
wire n1301;
wire n1303;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1314;
wire n1315;
wire n1317;
wire n1319;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1330;
wire n1331;
wire n1333;
wire n1335;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1346;
wire n1347;
wire n1349;
wire n1351;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1362;
wire n1363;
wire n1365;
wire n1367;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1378;
wire n1379;
wire n1381;
wire n1383;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1395;
wire n1396;
wire n1398;
wire n1400;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1410;
wire n1411;
wire n1413;
wire n1415;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1825;
wire n1826;
wire n1828;
wire n1830;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1842;
wire n1843;
wire n1845;
wire n1847;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1859;
wire n1860;
wire n1862;
wire n1864;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1884;
wire n1885;
wire n1887;
wire n1889;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1911;
wire n1912;
wire n1914;
wire n1916;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1937;
wire n1938;
wire n1940;
wire n1942;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1966;
wire n1967;
wire n1969;
wire n1971;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1985;
wire n1986;
wire n1988;
wire n1990;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2162;
wire n2163;
wire n2165;
wire n2167;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2178;
wire n2179;
wire n2181;
wire n2183;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2194;
wire n2195;
wire n2197;
wire n2199;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2210;
wire n2211;
wire n2213;
wire n2215;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2226;
wire n2227;
wire n2229;
wire n2231;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2242;
wire n2243;
wire n2245;
wire n2247;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2258;
wire n2259;
wire n2261;
wire n2263;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2273;
wire n2274;
wire n2276;
wire n2278;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2704;
wire n2706;
wire n2708;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2716;
wire n2718;
wire n2720;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2728;
wire n2730;
wire n2732;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2740;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2975;
wire n2976;
wire n2978;
wire n2979;
wire n2981;
wire n2982;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2989;
wire n2990;
wire n2992;
wire n2993;
wire n2995;
wire n2996;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3003;
wire n3004;
wire n3006;
wire n3007;
wire n3009;
wire n3010;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3053;
wire n3054;
wire n3057;
wire n3058;
wire n3061;
wire n3062;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3071;
wire n3072;
wire n3075;
wire n3076;
wire n3079;
wire n3080;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3089;
wire n3090;
wire n3093;
wire n3094;
wire n3097;
wire n3098;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3107;
wire n3108;
wire n3111;
wire n3112;
wire n3114;
wire n3115;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3158;
wire n3159;
wire n3162;
wire n3163;
wire n3166;
wire n3167;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3176;
wire n3177;
wire n3180;
wire n3181;
wire n3184;
wire n3185;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3194;
wire n3195;
wire n3198;
wire n3199;
wire n3202;
wire n3203;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3212;
wire n3213;
wire n3216;
wire n3217;
wire n3219;
wire n3220;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3263;
wire n3264;
wire n3267;
wire n3268;
wire n3271;
wire n3272;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3281;
wire n3282;
wire n3285;
wire n3286;
wire n3289;
wire n3290;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3299;
wire n3300;
wire n3303;
wire n3304;
wire n3307;
wire n3308;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3317;
wire n3318;
wire n3321;
wire n3322;
wire n3324;
wire n3325;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3368;
wire n3369;
wire n3372;
wire n3373;
wire n3376;
wire n3377;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3386;
wire n3387;
wire n3390;
wire n3391;
wire n3394;
wire n3395;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3404;
wire n3405;
wire n3408;
wire n3409;
wire n3412;
wire n3413;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3422;
wire n3423;
wire n3426;
wire n3427;
wire n3429;
wire n3430;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3473;
wire n3474;
wire n3477;
wire n3478;
wire n3481;
wire n3482;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3491;
wire n3492;
wire n3495;
wire n3496;
wire n3499;
wire n3500;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3509;
wire n3510;
wire n3513;
wire n3514;
wire n3517;
wire n3518;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3527;
wire n3528;
wire n3531;
wire n3532;
wire n3534;
wire n3535;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3578;
wire n3579;
wire n3582;
wire n3583;
wire n3586;
wire n3587;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3596;
wire n3597;
wire n3600;
wire n3601;
wire n3604;
wire n3605;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3614;
wire n3615;
wire n3618;
wire n3619;
wire n3622;
wire n3623;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3632;
wire n3633;
wire n3636;
wire n3637;
wire n3639;
wire n3640;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3682;
wire n3683;
wire n3686;
wire n3687;
wire n3690;
wire n3691;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3700;
wire n3701;
wire n3704;
wire n3705;
wire n3708;
wire n3709;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3718;
wire n3719;
wire n3722;
wire n3723;
wire n3726;
wire n3727;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3736;
wire n3737;
wire n3740;
wire n3741;
wire n3743;
wire n3744;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5031;
wire n5032;
wire n5033;
wire n5035;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5042;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5049;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5056;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5100;
wire n5101;
wire n5103;
wire n5104;
wire n5106;
wire n5107;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5115;
wire n5116;
wire n5118;
wire n5119;
wire n5121;
wire n5122;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5129;
wire n5130;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5145;
wire n5146;
wire n5148;
wire n5149;
wire n5151;
wire n5152;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5159;
wire n5160;
wire n5162;
wire n5163;
wire n5165;
wire n5166;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5174;
wire n5175;
wire n5177;
wire n5178;
wire n5180;
wire n5181;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5188;
wire n5189;
wire n5191;
wire n5192;
wire n5194;
wire n5195;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5209;
wire n5210;
wire n5212;
wire n5213;
wire n5215;
wire n5216;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5223;
wire n5224;
wire n5226;
wire n5227;
wire n5229;
wire n5230;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5238;
wire n5239;
wire n5241;
wire n5242;
wire n5244;
wire n5245;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5252;
wire n5253;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5268;
wire n5269;
wire n5271;
wire n5272;
wire n5274;
wire n5275;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5282;
wire n5283;
wire n5285;
wire n5286;
wire n5288;
wire n5289;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5297;
wire n5298;
wire n5300;
wire n5301;
wire n5303;
wire n5304;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5311;
wire n5312;
wire n5314;
wire n5315;
wire n5317;
wire n5318;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5332;
wire n5333;
wire n5335;
wire n5336;
wire n5338;
wire n5339;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5346;
wire n5347;
wire n5349;
wire n5350;
wire n5352;
wire n5353;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5361;
wire n5362;
wire n5364;
wire n5365;
wire n5367;
wire n5368;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5375;
wire n5376;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5391;
wire n5392;
wire n5394;
wire n5395;
wire n5397;
wire n5398;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5405;
wire n5406;
wire n5408;
wire n5409;
wire n5411;
wire n5412;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5420;
wire n5421;
wire n5423;
wire n5424;
wire n5426;
wire n5427;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5434;
wire n5435;
wire n5437;
wire n5438;
wire n5440;
wire n5441;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5455;
wire n5456;
wire n5458;
wire n5459;
wire n5461;
wire n5462;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5469;
wire n5470;
wire n5472;
wire n5473;
wire n5475;
wire n5476;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5484;
wire n5485;
wire n5487;
wire n5488;
wire n5490;
wire n5491;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5498;
wire n5499;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5514;
wire n5515;
wire n5517;
wire n5518;
wire n5520;
wire n5521;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5528;
wire n5529;
wire n5531;
wire n5532;
wire n5534;
wire n5535;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5543;
wire n5544;
wire n5546;
wire n5547;
wire n5549;
wire n5550;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5557;
wire n5558;
wire n5560;
wire n5561;
wire n5563;
wire n5564;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5578;
wire n5579;
wire n5581;
wire n5582;
wire n5584;
wire n5585;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5592;
wire n5593;
wire n5595;
wire n5596;
wire n5598;
wire n5599;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5607;
wire n5608;
wire n5610;
wire n5611;
wire n5613;
wire n5614;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5621;
wire n5622;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5637;
wire n5638;
wire n5640;
wire n5641;
wire n5643;
wire n5644;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5651;
wire n5652;
wire n5654;
wire n5655;
wire n5657;
wire n5658;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5666;
wire n5667;
wire n5669;
wire n5670;
wire n5672;
wire n5673;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5680;
wire n5681;
wire n5683;
wire n5684;
wire n5686;
wire n5687;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5701;
wire n5702;
wire n5704;
wire n5705;
wire n5707;
wire n5708;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5715;
wire n5716;
wire n5718;
wire n5719;
wire n5721;
wire n5722;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5730;
wire n5731;
wire n5733;
wire n5734;
wire n5736;
wire n5737;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5744;
wire n5745;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5760;
wire n5761;
wire n5763;
wire n5764;
wire n5766;
wire n5767;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5774;
wire n5775;
wire n5777;
wire n5778;
wire n5780;
wire n5781;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5789;
wire n5790;
wire n5792;
wire n5793;
wire n5795;
wire n5796;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5803;
wire n5804;
wire n5806;
wire n5807;
wire n5809;
wire n5810;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5824;
wire n5825;
wire n5827;
wire n5828;
wire n5830;
wire n5831;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5838;
wire n5839;
wire n5841;
wire n5842;
wire n5844;
wire n5845;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5853;
wire n5854;
wire n5856;
wire n5857;
wire n5859;
wire n5860;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5867;
wire n5868;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5883;
wire n5884;
wire n5886;
wire n5887;
wire n5889;
wire n5890;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5897;
wire n5898;
wire n5900;
wire n5901;
wire n5903;
wire n5904;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5912;
wire n5913;
wire n5915;
wire n5916;
wire n5918;
wire n5919;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5926;
wire n5927;
wire n5929;
wire n5930;
wire n5932;
wire n5933;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5946;
wire n5947;
wire n5949;
wire n5950;
wire n5952;
wire n5953;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5960;
wire n5961;
wire n5963;
wire n5964;
wire n5966;
wire n5967;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5975;
wire n5976;
wire n5978;
wire n5979;
wire n5981;
wire n5982;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5989;
wire n5990;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6005;
wire n6006;
wire n6008;
wire n6009;
wire n6011;
wire n6012;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6019;
wire n6020;
wire n6022;
wire n6023;
wire n6025;
wire n6026;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6034;
wire n6035;
wire n6037;
wire n6038;
wire n6040;
wire n6041;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6048;
wire n6049;
wire n6051;
wire n6052;
wire n6054;
wire n6055;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6076;
wire n6078;
wire n6079;
wire n6080;
wire n6082;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6089;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6821;
wire n6823;
wire n6824;
wire n6826;
wire n6828;
wire n6829;
wire n6830;
wire n6832;
wire n6834;
wire n6835;
wire n6837;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6852;
wire n6853;
wire n6855;
wire n6856;
wire n6858;
wire n6859;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6866;
wire n6867;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6882;
wire n6883;
wire n6885;
wire n6886;
wire n6888;
wire n6889;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6896;
wire n6897;
wire n6899;
wire n6900;
wire n6902;
wire n6903;
wire n6905;
wire n6906;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6921;
wire n6922;
wire n6924;
wire n6925;
wire n6927;
wire n6928;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6935;
wire n6936;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6951;
wire n6952;
wire n6954;
wire n6955;
wire n6957;
wire n6958;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6965;
wire n6966;
wire n6968;
wire n6969;
wire n6971;
wire n6972;
wire n6974;
wire n6975;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6990;
wire n6991;
wire n6993;
wire n6994;
wire n6996;
wire n6997;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7004;
wire n7005;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7020;
wire n7021;
wire n7023;
wire n7024;
wire n7026;
wire n7027;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7034;
wire n7035;
wire n7037;
wire n7038;
wire n7040;
wire n7041;
wire n7043;
wire n7044;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7059;
wire n7060;
wire n7062;
wire n7063;
wire n7065;
wire n7066;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7073;
wire n7074;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7089;
wire n7090;
wire n7092;
wire n7093;
wire n7095;
wire n7096;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7103;
wire n7104;
wire n7106;
wire n7107;
wire n7109;
wire n7110;
wire n7112;
wire n7113;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7128;
wire n7129;
wire n7131;
wire n7132;
wire n7134;
wire n7135;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7142;
wire n7143;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7158;
wire n7159;
wire n7161;
wire n7162;
wire n7164;
wire n7165;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7172;
wire n7173;
wire n7175;
wire n7176;
wire n7178;
wire n7179;
wire n7181;
wire n7182;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7197;
wire n7198;
wire n7200;
wire n7201;
wire n7203;
wire n7204;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7211;
wire n7212;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7227;
wire n7228;
wire n7230;
wire n7231;
wire n7233;
wire n7234;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7241;
wire n7242;
wire n7244;
wire n7245;
wire n7247;
wire n7248;
wire n7250;
wire n7251;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7266;
wire n7267;
wire n7269;
wire n7270;
wire n7272;
wire n7273;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7280;
wire n7281;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7296;
wire n7297;
wire n7299;
wire n7300;
wire n7302;
wire n7303;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7310;
wire n7311;
wire n7313;
wire n7314;
wire n7316;
wire n7317;
wire n7319;
wire n7320;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7334;
wire n7335;
wire n7337;
wire n7338;
wire n7340;
wire n7341;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7348;
wire n7349;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7364;
wire n7365;
wire n7367;
wire n7368;
wire n7370;
wire n7371;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7378;
wire n7379;
wire n7381;
wire n7382;
wire n7384;
wire n7385;
wire n7387;
wire n7388;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7416;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7787;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7796;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7812;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7821;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7828;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7835;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7857;
wire n7859;
wire n7860;
wire n7862;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8057;
wire n8058;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8169;
wire n8170;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8281;
wire n8282;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8393;
wire n8394;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8501;
wire n8502;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8609;
wire n8610;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8716;
wire n8717;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
xor (out,n0,n8861);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n8860);
and (s0n0,notn0,n1);
and (s1n0,n8860,n2870);
wire s0n1,s1n1,notn1;
or (n1,s0n1,s1n1);
not(notn1,n2697);
and (s0n1,notn1,n2);
and (s1n1,n2697,n2692);
xor (n2,n3,n2669);
xor (n3,n4,n2570);
xor (n4,n5,n1814);
xor (n5,n6,n1719);
xor (n6,n7,n1290);
xor (n7,n8,n1074);
wire s0n8,s1n8,notn8;
or (n8,s0n8,s1n8);
not(notn8,n928);
and (s0n8,notn8,1'b0);
and (s1n8,n928,n10);
xor (n10,n11,n739);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n585);
and (s0n11,notn11,1'b0);
and (s1n11,n585,n12);
wire s0n12,s1n12,notn12;
or (n12,s0n12,s1n12);
not(notn12,n568);
and (s0n12,notn12,n13);
and (s1n12,n568,n555);
wire s0n13,s1n13,notn13;
or (n13,s0n13,s1n13);
not(notn13,n15);
and (s0n13,notn13,1'b0);
and (s1n13,n15,n14);
and (n15,n16,n549);
and (n16,n17,n33);
or (n17,n18,n23,n27,n30);
and (n18,n19,n20);
and (n20,n21,n22);
and (n23,n24,n25);
and (n25,n26,n22);
not (n26,n21);
and (n27,n28,n29);
nor (n29,n26,n22);
and (n30,n31,n32);
nor (n32,n21,n22);
and (n33,n34,n548);
not (n34,n35);
wire s0n35,s1n35,notn35;
or (n35,s0n35,s1n35);
not(notn35,n547);
and (s0n35,notn35,n36);
and (s1n35,n547,1'b0);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n177);
and (s0n36,notn36,n37);
and (s1n36,n177,n38);
wire s0n38,s1n38,notn38;
or (n38,s0n38,s1n38);
not(notn38,n540);
and (s0n38,notn38,n39);
and (s1n38,n540,n514);
or (n39,n40,n482,n513,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n40,n41,n481);
or (n41,n42,n480);
or (n42,n43,n479);
or (n43,n44,n477);
or (n44,n45,n476);
or (n45,n46,n474);
or (n46,n47,n472);
nor (n47,n48,n397,n406,n418,n430,n441,n452,n463);
or (n48,1'b0,n49,n391,n395);
and (n49,n50,n390);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n381);
and (s0n50,notn50,n51);
and (s1n50,n381,n289);
wire s0n51,s1n51,notn51;
or (n51,s0n51,s1n51);
not(notn51,n248);
and (s0n51,notn51,1'b0);
and (s1n51,n248,n52);
or (n52,n53,n229,n233,n237,n240,n243,n245,1'b0);
and (n53,n54,n56);
not (n54,n55);
and (n56,n57,n202,n213,n223);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n91);
and (s0n57,notn57,n58);
and (s1n57,n91,1'b0);
wire s0n58,s1n58,notn58;
or (n58,s0n58,s1n58);
not(notn58,n89);
and (s0n58,notn58,n59);
and (s1n58,n89,n87);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n83);
and (s0n59,notn59,n60);
and (s1n59,n83,n77);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n76);
and (s0n60,notn60,n61);
and (s1n60,n76,1'b0);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n75);
and (s0n61,notn61,n62);
and (s1n61,n75,1'b1);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n74);
and (s0n62,notn62,n63);
and (s1n62,n74,1'b0);
wire s0n63,s1n63,notn63;
or (n63,s0n63,s1n63);
not(notn63,n73);
and (s0n63,notn63,n64);
and (s1n63,n73,1'b1);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n72);
and (s0n64,notn64,n65);
and (s1n64,n72,1'b0);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n71);
and (s0n65,notn65,n66);
and (s1n65,n71,1'b1);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n70);
and (s0n66,notn66,n67);
and (s1n66,n70,1'b0);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n69);
and (s0n67,notn67,n54);
and (s1n67,n69,1'b1);
wire s0n77,s1n77,notn77;
or (n77,s0n77,s1n77);
not(notn77,n82);
and (s0n77,notn77,n78);
and (s1n77,n82,1'b0);
wire s0n78,s1n78,notn78;
or (n78,s0n78,s1n78);
not(notn78,n81);
and (s0n78,notn78,n79);
and (s1n78,n81,1'b1);
not (n79,n80);
or (n83,n84,n86);
or (n84,n85,n80);
or (n85,n82,n81);
not (n87,n88);
or (n89,n88,n90);
not (n91,n92);
or (n92,n93,n200);
or (n93,n94,n198);
or (n94,n95,n192);
or (n95,n96,n191);
or (n96,n97,n187);
or (n97,n98,n186);
or (n98,n99,n181);
or (n99,n100,n180);
or (n100,n101,n179);
or (n101,n102,n177);
or (n102,n103,n171);
or (n103,n104,n170);
or (n104,n105,n169);
or (n105,n106,n168);
or (n106,n107,n167);
or (n107,n108,n166);
or (n108,n109,n165);
or (n109,n110,n164);
or (n110,n111,n161);
or (n111,n112,n155);
or (n112,n113,n154);
or (n113,n114,n153);
or (n114,n115,n152);
or (n115,n116,n151);
or (n116,n117,n150);
or (n117,n118,n148);
or (n118,n119,n146);
or (n119,n120,n140);
or (n120,n121,n139);
or (n121,n122,n138);
or (n122,n123,n137);
or (n123,n124,n136);
or (n124,n125,n134);
or (n125,n126,n132);
nor (n126,n127,n128,n130,n131);
not (n128,n129);
nor (n132,n127,n128,n133,n131);
not (n133,n130);
and (n134,n127,n129,n130,n135);
not (n135,n131);
and (n136,n127,n128,n130,n135);
nor (n137,n127,n129,n133,n131);
and (n138,n127,n128,n130,n131);
and (n139,n127,n129,n130,n131);
nor (n140,n141,n143,n144,n145);
not (n141,n142);
nor (n146,n141,n147,n144,n145);
not (n147,n143);
and (n148,n141,n143,n144,n149);
not (n149,n145);
and (n150,n142,n143,n144,n149);
and (n151,n142,n147,n144,n149);
and (n152,n141,n147,n144,n145);
and (n153,n142,n147,n144,n145);
and (n154,n142,n143,n144,n145);
nor (n155,n156,n158,n159,n160);
not (n156,n157);
and (n161,n157,n158,n162,n163);
not (n162,n159);
not (n163,n160);
and (n164,n156,n158,n162,n163);
and (n165,n157,n158,n159,n163);
nor (n166,n157,n158,n162,n163);
and (n167,n156,n158,n159,n160);
and (n168,n156,n158,n162,n160);
and (n169,n157,n158,n162,n160);
nor (n170,n156,n158,n159,n163);
nor (n171,n172,n174,n175,n176);
not (n172,n173);
nor (n177,n173,n178,n175,n176);
not (n178,n174);
and (n179,n172,n178,n175,n176);
and (n180,n173,n178,n175,n176);
nor (n181,n182,n183,n185);
not (n183,n184);
and (n186,n182,n184,n185);
and (n187,n188,n189);
not (n189,n190);
nor (n191,n188,n189);
nor (n192,n193,n194,n196,n197);
not (n194,n195);
and (n198,n193,n195,n196,n199);
not (n199,n197);
and (n200,n201,n194,n196,n199);
not (n201,n193);
wire s0n202,s1n202,notn202;
or (n202,s0n202,s1n202);
not(notn202,n91);
and (s0n202,notn202,n203);
and (s1n202,n91,1'b0);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n89);
and (s0n203,notn203,n204);
and (s1n203,n89,1'b0);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n83);
and (s0n204,notn204,n205);
and (s1n204,n83,n85);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n76);
and (s0n205,notn205,n206);
and (s1n205,n76,1'b1);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n75);
and (s0n206,notn206,n207);
and (s1n206,n75,1'b1);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n74);
and (s0n207,notn207,n208);
and (s1n207,n74,1'b0);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n73);
and (s0n208,notn208,n209);
and (s1n208,n73,1'b0);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n72);
and (s0n209,notn209,n210);
and (s1n209,n72,1'b1);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n71);
and (s0n210,notn210,n211);
and (s1n210,n71,1'b1);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n70);
and (s0n211,notn211,n212);
and (s1n211,n70,1'b0);
not (n212,n69);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n91);
and (s0n213,notn213,n214);
and (s1n213,n91,1'b0);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n89);
and (s0n214,notn214,n215);
and (s1n214,n89,1'b0);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n83);
and (s0n215,notn215,n216);
and (s1n215,n83,n222);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n76);
and (s0n216,notn216,n217);
and (s1n216,n76,1'b1);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n75);
and (s0n217,notn217,n218);
and (s1n217,n75,1'b1);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n74);
and (s0n218,notn218,n219);
and (s1n218,n74,1'b0);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n73);
and (s0n219,notn219,n220);
and (s1n219,n73,1'b0);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n72);
and (s0n220,notn220,n221);
and (s1n220,n72,1'b0);
not (n221,n71);
not (n222,n85);
not (n223,n224);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n91);
and (s0n224,notn224,n225);
and (s1n224,n91,1'b0);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n89);
and (s0n225,notn225,n226);
and (s1n225,n89,1'b0);
wire s0n226,s1n226,notn226;
or (n226,s0n226,s1n226);
not(notn226,n83);
and (s0n226,notn226,n227);
and (s1n226,n83,1'b0);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n76);
and (s0n227,notn227,n228);
and (s1n227,n76,1'b0);
not (n228,n75);
and (n229,n230,n231);
not (n230,n70);
and (n231,n232,n202,n213,n223);
not (n232,n57);
and (n233,n234,n235);
not (n234,n72);
and (n235,n57,n236,n213,n223);
not (n236,n202);
and (n237,n238,n239);
not (n238,n74);
and (n239,n232,n236,n213,n223);
and (n240,n241,n242);
not (n241,n76);
nor (n242,n232,n236,n213,n224);
and (n243,n79,n244);
nor (n244,n57,n236,n213,n224);
and (n245,n246,n247);
not (n246,n82);
nor (n247,n232,n202,n213,n224);
or (n248,n249,n278);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n276);
and (s0n249,notn249,n250);
and (s1n249,n276,1'b0);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n275);
and (s0n250,notn250,n251);
and (s1n250,n275,n270);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n269);
and (s0n251,notn251,n252);
and (s1n251,n269,n258);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n257);
and (s0n252,notn252,n253);
and (s1n252,n257,n120);
or (n253,n254,n151);
or (n254,n255,n150);
or (n255,n256,n148);
or (n256,n140,n146);
or (n257,n127,n129,n130,n131);
or (n258,1'b0,1'b0,n259,n265,n267);
and (n259,n260,n263);
or (n260,1'b0,1'b0,n261,n181);
and (n261,n262,n184,n185);
not (n262,n182);
and (n263,n172,n178,n175,n264);
not (n264,n176);
and (n265,n188,n266);
and (n266,n173,n178,n175,n264);
or (n267,n268,n179);
or (n268,n171,n177);
or (n269,n173,n174,n175,n176);
or (n270,n271,n170);
or (n271,n272,n168);
or (n272,n273,n165);
or (n273,n274,n164);
or (n274,n155,n161);
or (n275,n157,n158,n159,n160);
not (n276,n277);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n276);
and (s0n278,notn278,n279);
and (s1n278,n276,1'b0);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n275);
and (s0n279,notn279,n280);
and (s1n279,n275,n288);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n269);
and (s0n280,notn280,n281);
and (s1n280,n269,n284);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n257);
and (s0n281,notn281,n282);
and (s1n281,n257,1'b0);
or (n282,n283,n154);
or (n283,n152,n153);
or (n284,1'b0,n180,n285,n287,1'b0);
and (n285,n286,n263);
or (n286,1'b0,n186,n261,1'b0);
and (n287,n190,n266);
or (n288,n167,n169);
not (n289,n290);
nor (n290,n51,n291,n307,n327,n344,n358,n369,n377);
wire s0n291,s1n291,notn291;
or (n291,s0n291,s1n291);
not(notn291,n248);
and (s0n291,notn291,1'b0);
and (s1n291,n248,n292);
or (n292,n293,n295,n297,n299,n301,n303,n305,1'b0);
and (n293,n294,n56);
xnor (n294,n69,n55);
and (n295,n296,n231);
xnor (n296,n71,n70);
and (n297,n298,n235);
xnor (n298,n73,n72);
and (n299,n300,n239);
xnor (n300,n75,n74);
and (n301,n302,n242);
xnor (n302,n86,n76);
and (n303,n304,n244);
xnor (n304,n81,n80);
and (n305,n306,n247);
xnor (n306,n90,n82);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n248);
and (s0n307,notn307,1'b0);
and (s1n307,n248,n308);
or (n308,n309,n312,n315,n318,n321,n324,1'b0,1'b0);
and (n309,n310,n56);
xnor (n310,n70,n311);
or (n311,n69,n55);
and (n312,n313,n231);
xnor (n313,n72,n314);
or (n314,n71,n70);
and (n315,n316,n235);
xnor (n316,n74,n317);
or (n317,n73,n72);
and (n318,n319,n239);
xnor (n319,n76,n320);
or (n320,n75,n74);
and (n321,n322,n242);
xnor (n322,n80,n323);
or (n323,n86,n76);
and (n324,n325,n244);
xnor (n325,n82,n326);
or (n326,n81,n80);
wire s0n327,s1n327,notn327;
or (n327,s0n327,s1n327);
not(notn327,n248);
and (s0n327,notn327,1'b0);
and (s1n327,n248,n328);
or (n328,n329,n332,n335,n338,n341,1'b0,1'b0,1'b0);
and (n329,n330,n56);
xnor (n330,n71,n331);
or (n331,n70,n311);
and (n332,n333,n231);
xnor (n333,n73,n334);
or (n334,n72,n314);
and (n335,n336,n235);
xnor (n336,n75,n337);
or (n337,n74,n317);
and (n338,n339,n239);
xnor (n339,n86,n340);
or (n340,n76,n320);
and (n341,n342,n242);
xnor (n342,n81,n343);
or (n343,n80,n323);
wire s0n344,s1n344,notn344;
or (n344,s0n344,s1n344);
not(notn344,n248);
and (s0n344,notn344,1'b0);
and (s1n344,n248,n345);
or (n345,n346,n349,n352,n355,1'b0,1'b0,1'b0,1'b0);
and (n346,n347,n56);
xnor (n347,n72,n348);
or (n348,n71,n331);
and (n349,n350,n231);
xnor (n350,n74,n351);
or (n351,n73,n334);
and (n352,n353,n235);
xnor (n353,n76,n354);
or (n354,n75,n337);
and (n355,n356,n239);
xnor (n356,n80,n357);
or (n357,n86,n340);
wire s0n358,s1n358,notn358;
or (n358,s0n358,s1n358);
not(notn358,n248);
and (s0n358,notn358,1'b0);
and (s1n358,n248,n359);
or (n359,n360,n363,n366,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n360,n361,n56);
xnor (n361,n73,n362);
or (n362,n72,n348);
and (n363,n364,n231);
xnor (n364,n75,n365);
or (n365,n74,n351);
and (n366,n367,n235);
xnor (n367,n86,n368);
or (n368,n76,n354);
wire s0n369,s1n369,notn369;
or (n369,s0n369,s1n369);
not(notn369,n248);
and (s0n369,notn369,1'b0);
and (s1n369,n248,n370);
or (n370,n371,n374,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n371,n372,n56);
xnor (n372,n74,n373);
or (n373,n73,n362);
and (n374,n375,n231);
xnor (n375,n76,n376);
or (n376,n75,n365);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n248);
and (s0n377,notn377,1'b0);
and (s1n377,n248,n378);
and (n378,n379,n56);
xnor (n379,n75,n380);
or (n380,n74,n373);
nor (n381,n382,n384,n387);
not (n382,n383);
not (n384,n385);
xor (n385,n386,n383);
xor (n387,n388,n389);
and (n389,n386,n383);
and (n390,n249,n278);
and (n391,n392,n393);
xor (n392,n291,n51);
nor (n393,n249,n394);
not (n394,n278);
and (n395,n51,n396);
and (n396,n249,n394);
not (n397,n398);
or (n398,1'b0,n399,n401,n405);
and (n399,n400,n390);
wire s0n400,s1n400,notn400;
or (n400,s0n400,s1n400);
not(notn400,n381);
and (s0n400,notn400,n291);
and (s1n400,n381,1'b0);
and (n401,n402,n393);
xor (n402,n403,n404);
not (n403,n307);
not (n404,n291);
and (n405,n291,n396);
or (n406,1'b0,n407,n409,n417);
and (n407,n408,n390);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n381);
and (s0n408,notn408,n307);
and (s1n408,n381,1'b0);
and (n409,n410,n393);
wire s0n410,s1n410,notn410;
or (n410,s0n410,s1n410);
not(notn410,n51);
and (s0n410,notn410,n411);
and (s1n410,n51,n414);
xor (n411,n412,n413);
not (n412,n327);
and (n413,n403,n404);
xor (n414,n327,n415);
and (n415,n307,n416);
and (n416,n291,n51);
and (n417,n307,n396);
not (n418,n419);
or (n419,1'b0,n420,n422,n429);
and (n420,n421,n390);
wire s0n421,s1n421,notn421;
or (n421,s0n421,s1n421);
not(notn421,n381);
and (s0n421,notn421,n327);
and (s1n421,n381,1'b0);
and (n422,n423,n393);
wire s0n423,s1n423,notn423;
or (n423,s0n423,s1n423);
not(notn423,n51);
and (s0n423,notn423,n424);
and (s1n423,n51,n427);
xor (n424,n425,n426);
not (n425,n344);
and (n426,n412,n413);
xor (n427,n344,n428);
and (n428,n327,n415);
and (n429,n327,n396);
or (n430,1'b0,n431,n433,n440);
and (n431,n432,n390);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n381);
and (s0n432,notn432,n344);
and (s1n432,n381,1'b0);
and (n433,n434,n393);
wire s0n434,s1n434,notn434;
or (n434,s0n434,s1n434);
not(notn434,n51);
and (s0n434,notn434,n435);
and (s1n434,n51,n438);
xor (n435,n436,n437);
not (n436,n358);
and (n437,n425,n426);
xor (n438,n358,n439);
and (n439,n344,n428);
and (n440,n344,n396);
or (n441,1'b0,n442,n444,n451);
and (n442,n443,n390);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n381);
and (s0n443,notn443,n358);
and (s1n443,n381,1'b0);
and (n444,n445,n393);
wire s0n445,s1n445,notn445;
or (n445,s0n445,s1n445);
not(notn445,n51);
and (s0n445,notn445,n446);
and (s1n445,n51,n449);
xor (n446,n447,n448);
not (n447,n369);
and (n448,n436,n437);
xor (n449,n369,n450);
and (n450,n358,n439);
and (n451,n358,n396);
or (n452,1'b0,n453,n455,n462);
and (n453,n454,n390);
wire s0n454,s1n454,notn454;
or (n454,s0n454,s1n454);
not(notn454,n381);
and (s0n454,notn454,n369);
and (s1n454,n381,1'b0);
and (n455,n456,n393);
wire s0n456,s1n456,notn456;
or (n456,s0n456,s1n456);
not(notn456,n51);
and (s0n456,notn456,n457);
and (s1n456,n51,n460);
xor (n457,n458,n459);
not (n458,n377);
and (n459,n447,n448);
xor (n460,n377,n461);
and (n461,n369,n450);
and (n462,n369,n396);
or (n463,1'b0,n464,n466,n471);
and (n464,n465,n390);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n381);
and (s0n465,notn465,n377);
and (s1n465,n381,1'b0);
and (n466,n467,n393);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n51);
and (s0n467,notn467,n468);
and (s1n467,n51,n470);
not (n468,n469);
and (n469,n458,n459);
and (n470,n377,n461);
and (n471,n377,n396);
nor (n472,n473,n397,n406,n418,n430,n441,n452,n463);
not (n473,n48);
nor (n474,n48,n398,n475,n418,n430,n441,n452,n463);
not (n475,n406);
nor (n476,n473,n398,n475,n418,n430,n441,n452,n463);
nor (n477,n48,n397,n475,n419,n478,n441,n452,n463);
not (n478,n430);
nor (n479,n473,n397,n475,n419,n478,n441,n452,n463);
nor (n480,n48,n398,n406,n418,n478,n441,n452,n463);
nor (n481,n473,n398,n406,n418,n478,n441,n452,n463);
or (n482,n483,n498);
or (n483,n484,n497);
or (n484,n485,n496);
or (n485,n486,n495);
or (n486,n487,n494);
or (n487,n488,n493);
or (n488,n489,n492);
or (n489,n490,n491);
nor (n490,n48,n397,n475,n419,n430,n441,n452,n463);
nor (n491,n473,n397,n475,n419,n430,n441,n452,n463);
nor (n492,n48,n398,n406,n418,n430,n441,n452,n463);
nor (n493,n473,n398,n406,n418,n430,n441,n452,n463);
nor (n494,n48,n397,n406,n419,n478,n441,n452,n463);
nor (n495,n473,n397,n406,n419,n478,n441,n452,n463);
nor (n496,n48,n398,n475,n419,n478,n441,n452,n463);
nor (n497,n473,n398,n475,n419,n478,n441,n452,n463);
or (n498,n499,n512);
or (n499,n500,n511);
or (n500,n501,n510);
or (n501,n502,n509);
or (n502,n503,n508);
or (n503,n504,n507);
or (n504,n505,n506);
nor (n505,n48,n397,n475,n418,n430,n441,n452,n463);
nor (n506,n473,n397,n475,n418,n430,n441,n452,n463);
nor (n507,n48,n398,n406,n419,n478,n441,n452,n463);
nor (n508,n473,n398,n406,n419,n478,n441,n452,n463);
nor (n509,n48,n397,n406,n418,n478,n441,n452,n463);
nor (n510,n473,n397,n406,n418,n478,n441,n452,n463);
nor (n511,n48,n398,n475,n418,n478,n441,n452,n463);
nor (n512,n473,n398,n475,n418,n478,n441,n452,n463);
nor (n513,n473,n398,n475,n419,n430,n441,n452,n463);
or (n514,1'b0,n515,n522,n529,n290);
or (n515,n516,n480);
or (n516,n517,n479);
or (n517,n518,n477);
or (n518,n519,n497);
or (n519,n520,n474);
or (n520,n521,n472);
or (n521,n493,n47);
or (n522,n523,n496);
or (n523,n524,n495);
or (n524,n525,n494);
or (n525,n526,n508);
or (n526,n527,n492);
or (n527,n528,n491);
or (n528,n513,n490);
or (n529,n530,n507);
or (n530,n531,n506);
or (n531,n532,n505);
or (n532,n533,n476);
or (n533,n534,n539);
or (n534,n535,n538);
or (n535,n536,n537);
nor (n536,n473,n398,n406,n419,n430,n441,n452,n463);
nor (n537,n48,n397,n406,n419,n430,n441,n452,n463);
nor (n538,n473,n397,n406,n419,n430,n441,n452,n463);
nor (n539,n48,n398,n475,n419,n430,n441,n452,n463);
or (n540,n541,n546);
nor (n541,n542,n543,n545);
not (n543,n544);
and (n546,n542,n544,n545);
nor (n547,n172,n178,n175,n176);
nor (n549,n550,n552,n553,n554);
not (n550,n551);
or (n555,1'b0,n556,n558,n562,n565);
and (n556,n557,n549);
and (n558,n559,n560);
nor (n560,n551,n561,n553,n554);
not (n561,n552);
and (n562,n563,n564);
nor (n564,n550,n561,n553,n554);
and (n565,n14,n566);
and (n566,n550,n561,n553,n567);
not (n567,n554);
and (n568,n33,n569);
not (n569,n570);
wire s0n570,s1n570,notn570;
or (n570,s0n570,s1n570);
not(notn570,n583);
and (s0n570,notn570,n16);
and (s1n570,n583,n571);
or (n571,n572,n576,n579,n581);
and (n572,n19,n573);
and (n573,n574,n575);
and (n576,n24,n577);
and (n577,n578,n575);
not (n578,n574);
and (n579,n28,n580);
nor (n580,n578,n575);
and (n581,n31,n582);
nor (n582,n574,n575);
and (n583,n34,n584);
not (n584,n548);
and (n585,n586,n642);
not (n586,n587);
wire s0n587,s1n587,notn587;
or (n587,s0n587,s1n587);
not(notn587,n33);
and (s0n587,notn587,1'b0);
and (s1n587,n33,n588);
wire s0n588,s1n588,notn588;
or (n588,s0n588,s1n588);
not(notn588,n641);
and (s0n588,notn588,n589);
and (s1n588,n641,n632);
or (n589,n590,n608,n619,n630);
and (n590,n591,n20);
wire s0n591,s1n591,notn591;
or (n591,s0n591,s1n591);
not(notn591,n570);
and (s0n591,notn591,n592);
and (s1n591,n570,n593);
or (n593,n594,n599,n603,n606);
and (n594,n595,n596);
nor (n596,n597,n598);
and (n599,n600,n601);
nor (n601,n602,n598);
not (n602,n597);
and (n603,n604,n605);
and (n605,n602,n598);
and (n606,n592,n607);
and (n607,n597,n598);
and (n608,n609,n25);
wire s0n609,s1n609,notn609;
or (n609,s0n609,s1n609);
not(notn609,n570);
and (s0n609,notn609,n610);
and (s1n609,n570,n611);
or (n611,n612,n614,n616,n618);
and (n612,n613,n596);
and (n614,n615,n601);
and (n616,n617,n605);
and (n618,n610,n607);
and (n619,n620,n29);
wire s0n620,s1n620,notn620;
or (n620,s0n620,s1n620);
not(notn620,n570);
and (s0n620,notn620,n621);
and (s1n620,n570,n622);
or (n622,n623,n625,n627,n629);
and (n623,n624,n596);
and (n625,n626,n601);
and (n627,n628,n605);
and (n629,n621,n607);
and (n630,n631,n32);
wire s0n631,s1n631,notn631;
or (n631,s0n631,s1n631);
not(notn631,n570);
and (s0n631,notn631,n632);
and (s1n631,n570,n633);
or (n633,n634,n636,n638,n640);
and (n634,n635,n596);
and (n636,n637,n601);
and (n638,n639,n605);
and (n640,n632,n607);
and (n642,n643,n691);
not (n643,n644);
wire s0n644,s1n644,notn644;
or (n644,s0n644,s1n644);
not(notn644,n33);
and (s0n644,notn644,1'b0);
and (s1n644,n33,n645);
wire s0n645,s1n645,notn645;
or (n645,s0n645,s1n645);
not(notn645,n641);
and (s0n645,notn645,n646);
and (s1n645,n641,n682);
or (n646,n647,n658,n669,n680);
and (n647,n648,n20);
wire s0n648,s1n648,notn648;
or (n648,s0n648,s1n648);
not(notn648,n570);
and (s0n648,notn648,n649);
and (s1n648,n570,n650);
or (n650,n651,n653,n655,n657);
and (n651,n652,n596);
and (n653,n654,n601);
and (n655,n656,n605);
and (n657,n649,n607);
and (n658,n659,n25);
wire s0n659,s1n659,notn659;
or (n659,s0n659,s1n659);
not(notn659,n570);
and (s0n659,notn659,n660);
and (s1n659,n570,n661);
or (n661,n662,n664,n666,n668);
and (n662,n663,n596);
and (n664,n665,n601);
and (n666,n667,n605);
and (n668,n660,n607);
and (n669,n670,n29);
wire s0n670,s1n670,notn670;
or (n670,s0n670,s1n670);
not(notn670,n570);
and (s0n670,notn670,n671);
and (s1n670,n570,n672);
or (n672,n673,n675,n677,n679);
and (n673,n674,n596);
and (n675,n676,n601);
and (n677,n678,n605);
and (n679,n671,n607);
and (n680,n681,n32);
wire s0n681,s1n681,notn681;
or (n681,s0n681,s1n681);
not(notn681,n570);
and (s0n681,notn681,n682);
and (s1n681,n570,n683);
or (n683,n684,n686,n688,n690);
and (n684,n685,n596);
and (n686,n687,n601);
and (n688,n689,n605);
and (n690,n682,n607);
not (n691,n692);
wire s0n692,s1n692,notn692;
or (n692,s0n692,s1n692);
not(notn692,n33);
and (s0n692,notn692,1'b0);
and (s1n692,n33,n693);
wire s0n693,s1n693,notn693;
or (n693,s0n693,s1n693);
not(notn693,n641);
and (s0n693,notn693,n694);
and (s1n693,n641,n730);
or (n694,n695,n706,n717,n728);
and (n695,n696,n20);
wire s0n696,s1n696,notn696;
or (n696,s0n696,s1n696);
not(notn696,n570);
and (s0n696,notn696,n697);
and (s1n696,n570,n698);
or (n698,n699,n701,n703,n705);
and (n699,n700,n596);
and (n701,n702,n601);
and (n703,n704,n605);
and (n705,n697,n607);
and (n706,n707,n25);
wire s0n707,s1n707,notn707;
or (n707,s0n707,s1n707);
not(notn707,n570);
and (s0n707,notn707,n708);
and (s1n707,n570,n709);
or (n709,n710,n712,n714,n716);
and (n710,n711,n596);
and (n712,n713,n601);
and (n714,n715,n605);
and (n716,n708,n607);
and (n717,n718,n29);
wire s0n718,s1n718,notn718;
or (n718,s0n718,s1n718);
not(notn718,n570);
and (s0n718,notn718,n719);
and (s1n718,n570,n720);
or (n720,n721,n723,n725,n727);
and (n721,n722,n596);
and (n723,n724,n601);
and (n725,n726,n605);
and (n727,n719,n607);
and (n728,n729,n32);
wire s0n729,s1n729,notn729;
or (n729,s0n729,s1n729);
not(notn729,n570);
and (s0n729,notn729,n730);
and (s1n729,n570,n731);
or (n731,n732,n734,n736,n738);
and (n732,n733,n596);
and (n734,n735,n601);
and (n736,n737,n605);
and (n738,n730,n607);
or (n739,n740,n779);
and (n740,n741,n780);
xor (n741,n742,n757);
xor (n742,n743,n755);
wire s0n743,s1n743,notn743;
or (n743,s0n743,s1n743);
not(notn743,n585);
and (s0n743,notn743,1'b0);
and (s1n743,n585,n744);
wire s0n744,s1n744,notn744;
or (n744,s0n744,s1n744);
not(notn744,n568);
and (s0n744,notn744,n745);
and (s1n744,n568,n747);
wire s0n745,s1n745,notn745;
or (n745,s0n745,s1n745);
not(notn745,n15);
and (s0n745,notn745,1'b0);
and (s1n745,n15,n746);
or (n747,1'b0,n748,n750,n752,n754);
and (n748,n749,n549);
and (n750,n751,n560);
and (n752,n753,n564);
and (n754,n746,n566);
wire s0n755,s1n755,notn755;
or (n755,s0n755,s1n755);
not(notn755,n756);
and (s0n755,notn755,1'b0);
and (s1n755,n756,n12);
xor (n756,n586,n642);
or (n757,n758,n779);
and (n758,n759,n776);
xor (n759,n760,n761);
wire s0n760,s1n760,notn760;
or (n760,s0n760,s1n760);
not(notn760,n756);
and (s0n760,notn760,1'b0);
and (s1n760,n756,n744);
xor (n761,n762,n764);
wire s0n762,s1n762,notn762;
or (n762,s0n762,s1n762);
not(notn762,n763);
and (s0n762,notn762,1'b0);
and (s1n762,n763,n12);
xor (n763,n643,n691);
wire s0n764,s1n764,notn764;
or (n764,s0n764,s1n764);
not(notn764,n585);
and (s0n764,notn764,1'b0);
and (s1n764,n585,n765);
wire s0n765,s1n765,notn765;
or (n765,s0n765,s1n765);
not(notn765,n568);
and (s0n765,notn765,n766);
and (s1n765,n568,n768);
wire s0n766,s1n766,notn766;
or (n766,s0n766,s1n766);
not(notn766,n15);
and (s0n766,notn766,1'b0);
and (s1n766,n15,n767);
or (n768,1'b0,n769,n771,n773,n775);
and (n769,n770,n549);
and (n771,n772,n560);
and (n773,n774,n564);
and (n775,n767,n566);
and (n776,n777,n778);
wire s0n777,s1n777,notn777;
or (n777,s0n777,s1n777);
not(notn777,n763);
and (s0n777,notn777,1'b0);
and (s1n777,n763,n744);
wire s0n778,s1n778,notn778;
or (n778,s0n778,s1n778);
not(notn778,n692);
and (s0n778,notn778,1'b0);
and (s1n778,n692,n12);
and (n779,n760,n761);
nand (n780,n781,n927);
or (n781,n782,n922);
nor (n782,n783,n921);
and (n783,n784,n910);
nand (n784,n785,n909);
or (n785,n786,n843);
not (n786,n787);
or (n787,n788,n821);
xor (n788,n789,n818);
xor (n789,n790,n802);
wire s0n790,s1n790,notn790;
or (n790,s0n790,s1n790);
not(notn790,n756);
and (s0n790,notn790,1'b0);
and (s1n790,n756,n791);
wire s0n791,s1n791,notn791;
or (n791,s0n791,s1n791);
not(notn791,n568);
and (s0n791,notn791,n792);
and (s1n791,n568,n794);
wire s0n792,s1n792,notn792;
or (n792,s0n792,s1n792);
not(notn792,n15);
and (s0n792,notn792,1'b0);
and (s1n792,n15,n793);
or (n794,1'b0,n795,n797,n799,n801);
and (n795,n796,n549);
and (n797,n798,n560);
and (n799,n800,n564);
and (n801,n793,n566);
xor (n802,n803,n806);
xor (n803,n804,n805);
wire s0n804,s1n804,notn804;
or (n804,s0n804,s1n804);
not(notn804,n763);
and (s0n804,notn804,1'b0);
and (s1n804,n763,n765);
wire s0n805,s1n805,notn805;
or (n805,s0n805,s1n805);
not(notn805,n692);
and (s0n805,notn805,1'b0);
and (s1n805,n692,n744);
wire s0n806,s1n806,notn806;
or (n806,s0n806,s1n806);
not(notn806,n585);
and (s0n806,notn806,1'b0);
and (s1n806,n585,n807);
wire s0n807,s1n807,notn807;
or (n807,s0n807,s1n807);
not(notn807,n568);
and (s0n807,notn807,n808);
and (s1n807,n568,n810);
wire s0n808,s1n808,notn808;
or (n808,s0n808,s1n808);
not(notn808,n15);
and (s0n808,notn808,1'b0);
and (s1n808,n15,n809);
or (n810,1'b0,n811,n813,n815,n817);
and (n811,n812,n549);
and (n813,n814,n560);
and (n815,n816,n564);
and (n817,n809,n566);
and (n818,n819,n820);
wire s0n819,s1n819,notn819;
or (n819,s0n819,s1n819);
not(notn819,n763);
and (s0n819,notn819,1'b0);
and (s1n819,n763,n791);
wire s0n820,s1n820,notn820;
or (n820,s0n820,s1n820);
not(notn820,n692);
and (s0n820,notn820,1'b0);
and (s1n820,n692,n765);
or (n821,n822,n842);
and (n822,n823,n839);
xor (n823,n824,n825);
wire s0n824,s1n824,notn824;
or (n824,s0n824,s1n824);
not(notn824,n756);
and (s0n824,notn824,1'b0);
and (s1n824,n756,n807);
xor (n825,n826,n827);
xor (n826,n819,n820);
wire s0n827,s1n827,notn827;
or (n827,s0n827,s1n827);
not(notn827,n585);
and (s0n827,notn827,1'b0);
and (s1n827,n585,n828);
wire s0n828,s1n828,notn828;
or (n828,s0n828,s1n828);
not(notn828,n568);
and (s0n828,notn828,n829);
and (s1n828,n568,n831);
wire s0n829,s1n829,notn829;
or (n829,s0n829,s1n829);
not(notn829,n15);
and (s0n829,notn829,1'b0);
and (s1n829,n15,n830);
or (n831,1'b0,n832,n834,n836,n838);
and (n832,n833,n549);
and (n834,n835,n560);
and (n836,n837,n564);
and (n838,n830,n566);
and (n839,n840,n841);
wire s0n840,s1n840,notn840;
or (n840,s0n840,s1n840);
not(notn840,n763);
and (s0n840,notn840,1'b0);
and (s1n840,n763,n807);
wire s0n841,s1n841,notn841;
or (n841,s0n841,s1n841);
not(notn841,n692);
and (s0n841,notn841,1'b0);
and (s1n841,n692,n791);
and (n842,n824,n825);
not (n843,n844);
nand (n844,n845,n905,n908);
nand (n845,n846,n870,n902);
or (n846,n847,n848);
xor (n847,n823,n839);
or (n848,n849,n869);
and (n849,n850,n855);
xor (n850,n851,n852);
wire s0n851,s1n851,notn851;
or (n851,s0n851,s1n851);
not(notn851,n756);
and (s0n851,notn851,1'b0);
and (s1n851,n756,n828);
and (n852,n853,n854);
wire s0n853,s1n853,notn853;
or (n853,s0n853,s1n853);
not(notn853,n763);
and (s0n853,notn853,1'b0);
and (s1n853,n763,n828);
wire s0n854,s1n854,notn854;
or (n854,s0n854,s1n854);
not(notn854,n692);
and (s0n854,notn854,1'b0);
and (s1n854,n692,n807);
xor (n855,n856,n857);
xor (n856,n840,n841);
wire s0n857,s1n857,notn857;
or (n857,s0n857,s1n857);
not(notn857,n585);
and (s0n857,notn857,1'b0);
and (s1n857,n585,n858);
wire s0n858,s1n858,notn858;
or (n858,s0n858,s1n858);
not(notn858,n568);
and (s0n858,notn858,n859);
and (s1n858,n568,n861);
wire s0n859,s1n859,notn859;
or (n859,s0n859,s1n859);
not(notn859,n15);
and (s0n859,notn859,1'b0);
and (s1n859,n15,n860);
or (n861,1'b0,n862,n864,n866,n868);
and (n862,n863,n549);
and (n864,n865,n560);
and (n866,n867,n564);
and (n868,n860,n566);
and (n869,n851,n852);
or (n870,n871,n901);
and (n871,n872,n896);
xor (n872,n873,n876);
and (n873,n874,n875);
wire s0n874,s1n874,notn874;
or (n874,s0n874,s1n874);
not(notn874,n763);
and (s0n874,notn874,1'b0);
and (s1n874,n763,n858);
wire s0n875,s1n875,notn875;
or (n875,s0n875,s1n875);
not(notn875,n692);
and (s0n875,notn875,1'b0);
and (s1n875,n692,n828);
or (n876,n877,n895);
and (n877,n878,n894);
xor (n878,n879,n893);
and (n879,n880,n892);
wire s0n880,s1n880,notn880;
or (n880,s0n880,s1n880);
not(notn880,n763);
and (s0n880,notn880,1'b0);
and (s1n880,n763,n881);
wire s0n881,s1n881,notn881;
or (n881,s0n881,s1n881);
not(notn881,n568);
and (s0n881,notn881,n882);
and (s1n881,n568,n884);
wire s0n882,s1n882,notn882;
or (n882,s0n882,s1n882);
not(notn882,n15);
and (s0n882,notn882,1'b0);
and (s1n882,n15,n883);
or (n884,1'b0,n885,n887,n889,n891);
and (n885,n886,n549);
and (n887,n888,n560);
and (n889,n890,n564);
and (n891,n883,n566);
wire s0n892,s1n892,notn892;
or (n892,s0n892,s1n892);
not(notn892,n692);
and (s0n892,notn892,1'b0);
and (s1n892,n692,n858);
wire s0n893,s1n893,notn893;
or (n893,s0n893,s1n893);
not(notn893,n756);
and (s0n893,notn893,1'b0);
and (s1n893,n756,n881);
xor (n894,n874,n875);
and (n895,n879,n893);
xor (n896,n897,n900);
xor (n897,n898,n899);
wire s0n898,s1n898,notn898;
or (n898,s0n898,s1n898);
not(notn898,n585);
and (s0n898,notn898,1'b0);
and (s1n898,n585,n881);
xor (n899,n853,n854);
wire s0n900,s1n900,notn900;
or (n900,s0n900,s1n900);
not(notn900,n756);
and (s0n900,notn900,1'b0);
and (s1n900,n756,n858);
and (n901,n873,n876);
or (n902,n903,n904);
xor (n903,n850,n855);
and (n904,n897,n900);
nand (n905,n906,n846);
not (n906,n907);
nand (n907,n903,n904);
nand (n908,n847,n848);
nand (n909,n788,n821);
or (n910,n911,n918);
xor (n911,n912,n917);
xor (n912,n913,n914);
wire s0n913,s1n913,notn913;
or (n913,s0n913,s1n913);
not(notn913,n756);
and (s0n913,notn913,1'b0);
and (s1n913,n756,n765);
xor (n914,n915,n916);
xor (n915,n777,n778);
wire s0n916,s1n916,notn916;
or (n916,s0n916,s1n916);
not(notn916,n585);
and (s0n916,notn916,1'b0);
and (s1n916,n585,n791);
and (n917,n804,n805);
or (n918,n919,n920);
and (n919,n789,n818);
and (n920,n790,n802);
and (n921,n911,n918);
nor (n922,n923,n926);
or (n923,n924,n925);
and (n924,n912,n917);
and (n925,n913,n914);
xor (n926,n759,n776);
nand (n927,n923,n926);
and (n928,n929,n977);
not (n929,n930);
wire s0n930,s1n930,notn930;
or (n930,s0n930,s1n930);
not(notn930,n33);
and (s0n930,notn930,1'b0);
and (s1n930,n33,n931);
wire s0n931,s1n931,notn931;
or (n931,s0n931,s1n931);
not(notn931,n641);
and (s0n931,notn931,n932);
and (s1n931,n641,n968);
or (n932,n933,n944,n955,n966);
and (n933,n934,n20);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n570);
and (s0n934,notn934,n935);
and (s1n934,n570,n936);
or (n936,n937,n939,n941,n943);
and (n937,n938,n596);
and (n939,n940,n601);
and (n941,n942,n605);
and (n943,n935,n607);
and (n944,n945,n25);
wire s0n945,s1n945,notn945;
or (n945,s0n945,s1n945);
not(notn945,n570);
and (s0n945,notn945,n946);
and (s1n945,n570,n947);
or (n947,n948,n950,n952,n954);
and (n948,n949,n596);
and (n950,n951,n601);
and (n952,n953,n605);
and (n954,n946,n607);
and (n955,n956,n29);
wire s0n956,s1n956,notn956;
or (n956,s0n956,s1n956);
not(notn956,n570);
and (s0n956,notn956,n957);
and (s1n956,n570,n958);
or (n958,n959,n961,n963,n965);
and (n959,n960,n596);
and (n961,n962,n601);
and (n963,n964,n605);
and (n965,n957,n607);
and (n966,n967,n32);
wire s0n967,s1n967,notn967;
or (n967,s0n967,s1n967);
not(notn967,n570);
and (s0n967,notn967,n968);
and (s1n967,n570,n969);
or (n969,n970,n972,n974,n976);
and (n970,n971,n596);
and (n972,n973,n601);
and (n974,n975,n605);
and (n976,n968,n607);
and (n977,n978,n1026);
not (n978,n979);
wire s0n979,s1n979,notn979;
or (n979,s0n979,s1n979);
not(notn979,n33);
and (s0n979,notn979,1'b0);
and (s1n979,n33,n980);
wire s0n980,s1n980,notn980;
or (n980,s0n980,s1n980);
not(notn980,n641);
and (s0n980,notn980,n981);
and (s1n980,n641,n1017);
or (n981,n982,n993,n1004,n1015);
and (n982,n983,n20);
wire s0n983,s1n983,notn983;
or (n983,s0n983,s1n983);
not(notn983,n570);
and (s0n983,notn983,n984);
and (s1n983,n570,n985);
or (n985,n986,n988,n990,n992);
and (n986,n987,n596);
and (n988,n989,n601);
and (n990,n991,n605);
and (n992,n984,n607);
and (n993,n994,n25);
wire s0n994,s1n994,notn994;
or (n994,s0n994,s1n994);
not(notn994,n570);
and (s0n994,notn994,n995);
and (s1n994,n570,n996);
or (n996,n997,n999,n1001,n1003);
and (n997,n998,n596);
and (n999,n1000,n601);
and (n1001,n1002,n605);
and (n1003,n995,n607);
and (n1004,n1005,n29);
wire s0n1005,s1n1005,notn1005;
or (n1005,s0n1005,s1n1005);
not(notn1005,n570);
and (s0n1005,notn1005,n1006);
and (s1n1005,n570,n1007);
or (n1007,n1008,n1010,n1012,n1014);
and (n1008,n1009,n596);
and (n1010,n1011,n601);
and (n1012,n1013,n605);
and (n1014,n1006,n607);
and (n1015,n1016,n32);
wire s0n1016,s1n1016,notn1016;
or (n1016,s0n1016,s1n1016);
not(notn1016,n570);
and (s0n1016,notn1016,n1017);
and (s1n1016,n570,n1018);
or (n1018,n1019,n1021,n1023,n1025);
and (n1019,n1020,n596);
and (n1021,n1022,n601);
and (n1023,n1024,n605);
and (n1025,n1017,n607);
not (n1026,n1027);
wire s0n1027,s1n1027,notn1027;
or (n1027,s0n1027,s1n1027);
not(notn1027,n33);
and (s0n1027,notn1027,1'b0);
and (s1n1027,n33,n1028);
wire s0n1028,s1n1028,notn1028;
or (n1028,s0n1028,s1n1028);
not(notn1028,n641);
and (s0n1028,notn1028,n1029);
and (s1n1028,n641,n1065);
or (n1029,n1030,n1041,n1052,n1063);
and (n1030,n1031,n20);
wire s0n1031,s1n1031,notn1031;
or (n1031,s0n1031,s1n1031);
not(notn1031,n570);
and (s0n1031,notn1031,n1032);
and (s1n1031,n570,n1033);
or (n1033,n1034,n1036,n1038,n1040);
and (n1034,n1035,n596);
and (n1036,n1037,n601);
and (n1038,n1039,n605);
and (n1040,n1032,n607);
and (n1041,n1042,n25);
wire s0n1042,s1n1042,notn1042;
or (n1042,s0n1042,s1n1042);
not(notn1042,n570);
and (s0n1042,notn1042,n1043);
and (s1n1042,n570,n1044);
or (n1044,n1045,n1047,n1049,n1051);
and (n1045,n1046,n596);
and (n1047,n1048,n601);
and (n1049,n1050,n605);
and (n1051,n1043,n607);
and (n1052,n1053,n29);
wire s0n1053,s1n1053,notn1053;
or (n1053,s0n1053,s1n1053);
not(notn1053,n570);
and (s0n1053,notn1053,n1054);
and (s1n1053,n570,n1055);
or (n1055,n1056,n1058,n1060,n1062);
and (n1056,n1057,n596);
and (n1058,n1059,n601);
and (n1060,n1061,n605);
and (n1062,n1054,n607);
and (n1063,n1064,n32);
wire s0n1064,s1n1064,notn1064;
or (n1064,s0n1064,s1n1064);
not(notn1064,n570);
and (s0n1064,notn1064,n1065);
and (s1n1064,n570,n1066);
or (n1066,n1067,n1069,n1071,n1073);
and (n1067,n1068,n596);
and (n1069,n1070,n601);
and (n1071,n1072,n605);
and (n1073,n1065,n607);
or (n1074,n1075,n1204,n1289);
and (n1075,n1076,n1081);
xor (n1076,n1077,n1079);
and (n1077,n1078,n928);
xor (n1078,n741,n780);
wire s0n1079,s1n1079,notn1079;
or (n1079,s0n1079,s1n1079);
not(notn1079,n1080);
and (s0n1079,notn1079,1'b0);
and (s1n1079,n1080,n10);
xor (n1080,n929,n977);
and (n1081,n1082,n1084);
wire s0n1082,s1n1082,notn1082;
or (n1082,s0n1082,s1n1082);
not(notn1082,n1083);
and (s0n1082,notn1082,1'b0);
and (s1n1082,n1083,n10);
xor (n1083,n978,n1026);
or (n1084,n1085,n1088,n1203);
and (n1085,n1086,n1087);
and (n1086,n1078,n1083);
wire s0n1087,s1n1087,notn1087;
or (n1087,s0n1087,s1n1087);
not(notn1087,n1027);
and (s0n1087,notn1087,1'b0);
and (s1n1087,n1027,n10);
and (n1088,n1087,n1089);
or (n1089,n1090,n1145,n1202);
and (n1090,n1091,n1144);
wire s0n1091,s1n1091,notn1091;
or (n1091,s0n1091,s1n1091);
not(notn1091,n1083);
and (s0n1091,notn1091,1'b0);
and (s1n1091,n1083,n1092);
xor (n1092,n1093,n1112);
xor (n1093,n1094,n1095);
xor (n1094,n764,n760);
xor (n1095,n762,n1096);
or (n1096,n776,n1097,n1111);
and (n1097,n778,n1098);
or (n1098,n917,n1099,n1110);
and (n1099,n805,n1100);
or (n1100,n818,n1101,n1109);
and (n1101,n820,n1102);
or (n1102,n839,n1103,n1108);
and (n1103,n841,n1104);
or (n1104,n852,n1105,n873);
and (n1105,n854,n1106);
or (n1106,n873,n1107,n879);
and (n1107,n875,n879);
and (n1108,n840,n1104);
and (n1109,n819,n1102);
and (n1110,n804,n1100);
and (n1111,n777,n1098);
or (n1112,n1113,n1116,n1143);
and (n1113,n1114,n1115);
xor (n1114,n916,n913);
xor (n1115,n915,n1098);
and (n1116,n1115,n1117);
or (n1117,n1118,n1121,n1142);
and (n1118,n1119,n1120);
xor (n1119,n806,n790);
xor (n1120,n803,n1100);
and (n1121,n1120,n1122);
or (n1122,n1123,n1126,n1141);
and (n1123,n1124,n1125);
xor (n1124,n827,n824);
xor (n1125,n826,n1102);
and (n1126,n1125,n1127);
or (n1127,n1128,n1131,n1140);
and (n1128,n1129,n1130);
xor (n1129,n857,n851);
xor (n1130,n856,n1104);
and (n1131,n1130,n1132);
or (n1132,n1133,n1136,n1139);
and (n1133,n1134,n1135);
xor (n1134,n898,n900);
xor (n1135,n899,n1106);
and (n1136,n1135,n1137);
and (n1137,n893,n1138);
xor (n1138,n894,n879);
and (n1139,n1134,n1137);
and (n1140,n1129,n1132);
and (n1141,n1124,n1127);
and (n1142,n1119,n1122);
and (n1143,n1114,n1117);
and (n1144,n1078,n1027);
and (n1145,n1144,n1146);
or (n1146,n1147,n1153,n1201);
and (n1147,n1148,n1152);
and (n1148,n1149,n1083);
xor (n1149,n1150,n784);
nor (n1150,n1151,n921);
not (n1151,n910);
wire s0n1152,s1n1152,notn1152;
or (n1152,s0n1152,s1n1152);
not(notn1152,n1027);
and (s0n1152,notn1152,1'b0);
and (s1n1152,n1027,n1092);
and (n1153,n1152,n1154);
or (n1154,n1155,n1160,n1200);
and (n1155,n1156,n1159);
and (n1156,n1157,n1083);
xnor (n1157,n844,n1158);
nand (n1158,n787,n909);
and (n1159,n1149,n1027);
and (n1160,n1159,n1161);
or (n1161,n1162,n1167,n1199);
and (n1162,n1163,n1166);
wire s0n1163,s1n1163,notn1163;
or (n1163,s0n1163,s1n1163);
not(notn1163,n1083);
and (s0n1163,notn1163,1'b0);
and (s1n1163,n1083,n1164);
xor (n1164,n1165,n1127);
xor (n1165,n1124,n1125);
and (n1166,n1157,n1027);
and (n1167,n1166,n1168);
or (n1168,n1169,n1174,n1198);
and (n1169,n1170,n1173);
wire s0n1170,s1n1170,notn1170;
or (n1170,s0n1170,s1n1170);
not(notn1170,n1083);
and (s0n1170,notn1170,1'b0);
and (s1n1170,n1083,n1171);
xor (n1171,n1172,n1132);
xor (n1172,n1129,n1130);
wire s0n1173,s1n1173,notn1173;
or (n1173,s0n1173,s1n1173);
not(notn1173,n1027);
and (s0n1173,notn1173,1'b0);
and (s1n1173,n1027,n1164);
and (n1174,n1173,n1175);
or (n1175,n1176,n1180,n1197);
and (n1176,n1177,n1179);
and (n1177,n1178,n1083);
xor (n1178,n872,n896);
wire s0n1179,s1n1179,notn1179;
or (n1179,s0n1179,s1n1179);
not(notn1179,n1027);
and (s0n1179,notn1179,1'b0);
and (s1n1179,n1027,n1171);
and (n1180,n1179,n1181);
or (n1181,n1182,n1186,n1188);
and (n1182,n1183,n1185);
and (n1183,n1184,n1083);
xor (n1184,n878,n894);
and (n1185,n1178,n1027);
and (n1186,n1185,n1187);
or (n1187,n1188,n1192,n1193);
and (n1188,n1189,n1191);
wire s0n1189,s1n1189,notn1189;
or (n1189,s0n1189,s1n1189);
not(notn1189,n1083);
and (s0n1189,notn1189,1'b0);
and (s1n1189,n1083,n1190);
xor (n1190,n880,n892);
and (n1191,n1184,n1027);
and (n1192,n1191,n1193);
and (n1193,n1194,n1196);
wire s0n1194,s1n1194,notn1194;
or (n1194,s0n1194,s1n1194);
not(notn1194,n1083);
and (s0n1194,notn1194,1'b0);
and (s1n1194,n1083,n1195);
wire s0n1195,s1n1195,notn1195;
or (n1195,s0n1195,s1n1195);
not(notn1195,n692);
and (s0n1195,notn1195,1'b0);
and (s1n1195,n692,n881);
wire s0n1196,s1n1196,notn1196;
or (n1196,s0n1196,s1n1196);
not(notn1196,n1027);
and (s0n1196,notn1196,1'b0);
and (s1n1196,n1027,n1190);
and (n1197,n1177,n1181);
and (n1198,n1170,n1175);
and (n1199,n1163,n1168);
and (n1200,n1156,n1161);
and (n1201,n1148,n1154);
and (n1202,n1091,n1146);
and (n1203,n1086,n1089);
and (n1204,n1081,n1205);
or (n1205,n1206,n1211,n1288);
and (n1206,n1207,n1210);
xor (n1207,n1208,n1209);
wire s0n1208,s1n1208,notn1208;
or (n1208,s0n1208,s1n1208);
not(notn1208,n928);
and (s0n1208,notn1208,1'b0);
and (s1n1208,n928,n1092);
and (n1209,n1078,n1080);
xor (n1210,n1082,n1084);
and (n1211,n1210,n1212);
or (n1212,n1213,n1219,n1287);
and (n1213,n1214,n1217);
xor (n1214,n1215,n1216);
and (n1215,n1149,n928);
wire s0n1216,s1n1216,notn1216;
or (n1216,s0n1216,s1n1216);
not(notn1216,n1080);
and (s0n1216,notn1216,1'b0);
and (s1n1216,n1080,n1092);
xor (n1217,n1218,n1089);
xor (n1218,n1086,n1087);
and (n1219,n1217,n1220);
or (n1220,n1221,n1227,n1286);
and (n1221,n1222,n1225);
xor (n1222,n1223,n1224);
and (n1223,n1157,n928);
and (n1224,n1149,n1080);
xor (n1225,n1226,n1146);
xor (n1226,n1091,n1144);
and (n1227,n1225,n1228);
or (n1228,n1229,n1235,n1285);
and (n1229,n1230,n1233);
xor (n1230,n1231,n1232);
wire s0n1231,s1n1231,notn1231;
or (n1231,s0n1231,s1n1231);
not(notn1231,n928);
and (s0n1231,notn1231,1'b0);
and (s1n1231,n928,n1164);
and (n1232,n1157,n1080);
xor (n1233,n1234,n1154);
xor (n1234,n1148,n1152);
and (n1235,n1233,n1236);
or (n1236,n1237,n1243,n1284);
and (n1237,n1238,n1241);
xor (n1238,n1239,n1240);
wire s0n1239,s1n1239,notn1239;
or (n1239,s0n1239,s1n1239);
not(notn1239,n928);
and (s0n1239,notn1239,1'b0);
and (s1n1239,n928,n1171);
wire s0n1240,s1n1240,notn1240;
or (n1240,s0n1240,s1n1240);
not(notn1240,n1080);
and (s0n1240,notn1240,1'b0);
and (s1n1240,n1080,n1164);
xor (n1241,n1242,n1161);
xor (n1242,n1156,n1159);
and (n1243,n1241,n1244);
or (n1244,n1245,n1251,n1283);
and (n1245,n1246,n1249);
xor (n1246,n1247,n1248);
and (n1247,n1178,n928);
wire s0n1248,s1n1248,notn1248;
or (n1248,s0n1248,s1n1248);
not(notn1248,n1080);
and (s0n1248,notn1248,1'b0);
and (s1n1248,n1080,n1171);
xor (n1249,n1250,n1168);
xor (n1250,n1163,n1166);
and (n1251,n1249,n1252);
or (n1252,n1253,n1259,n1282);
and (n1253,n1254,n1257);
xor (n1254,n1255,n1256);
and (n1255,n1184,n928);
and (n1256,n1178,n1080);
xor (n1257,n1258,n1175);
xor (n1258,n1170,n1173);
and (n1259,n1257,n1260);
or (n1260,n1261,n1267,n1281);
and (n1261,n1262,n1265);
xor (n1262,n1263,n1264);
wire s0n1263,s1n1263,notn1263;
or (n1263,s0n1263,s1n1263);
not(notn1263,n928);
and (s0n1263,notn1263,1'b0);
and (s1n1263,n928,n1190);
and (n1264,n1184,n1080);
xor (n1265,n1266,n1181);
xor (n1266,n1177,n1179);
and (n1267,n1265,n1268);
or (n1268,n1269,n1275,n1280);
and (n1269,n1270,n1273);
xor (n1270,n1271,n1272);
wire s0n1271,s1n1271,notn1271;
or (n1271,s0n1271,s1n1271);
not(notn1271,n928);
and (s0n1271,notn1271,1'b0);
and (s1n1271,n928,n1195);
wire s0n1272,s1n1272,notn1272;
or (n1272,s0n1272,s1n1272);
not(notn1272,n1080);
and (s0n1272,notn1272,1'b0);
and (s1n1272,n1080,n1190);
xor (n1273,n1274,n1187);
xor (n1274,n1183,n1185);
and (n1275,n1273,n1276);
and (n1276,n1277,n1278);
wire s0n1277,s1n1277,notn1277;
or (n1277,s0n1277,s1n1277);
not(notn1277,n1080);
and (s0n1277,notn1277,1'b0);
and (s1n1277,n1080,n1195);
xor (n1278,n1279,n1193);
xor (n1279,n1189,n1191);
and (n1280,n1270,n1276);
and (n1281,n1262,n1268);
and (n1282,n1254,n1260);
and (n1283,n1246,n1252);
and (n1284,n1238,n1244);
and (n1285,n1230,n1236);
and (n1286,n1222,n1228);
and (n1287,n1214,n1220);
and (n1288,n1207,n1212);
and (n1289,n1076,n1205);
xor (n1290,n1291,n1477);
wire s0n1291,s1n1291,notn1291;
or (n1291,s0n1291,s1n1291);
not(notn1291,n928);
and (s0n1291,notn1291,1'b0);
and (s1n1291,n928,n1292);
or (n1292,n1293,n1423,n1476);
and (n1293,n1294,n1306);
and (n1294,n587,n1295);
wire s0n1295,s1n1295,notn1295;
or (n1295,s0n1295,s1n1295);
not(notn1295,n568);
and (s0n1295,notn1295,n1296);
and (s1n1295,n568,n1298);
wire s0n1296,s1n1296,notn1296;
or (n1296,s0n1296,s1n1296);
not(notn1296,n15);
and (s0n1296,notn1296,1'b0);
and (s1n1296,n15,n1297);
or (n1298,1'b0,n1299,n1301,n1303,n1305);
and (n1299,n1300,n549);
and (n1301,n1302,n560);
and (n1303,n1304,n564);
and (n1305,n1297,n566);
and (n1306,n1307,n1308);
wire s0n1307,s1n1307,notn1307;
or (n1307,s0n1307,s1n1307);
not(notn1307,n644);
and (s0n1307,notn1307,1'b0);
and (s1n1307,n644,n1295);
or (n1308,n1309,n1323,n1422);
and (n1309,n1310,n1322);
wire s0n1310,s1n1310,notn1310;
or (n1310,s0n1310,s1n1310);
not(notn1310,n644);
and (s0n1310,notn1310,1'b0);
and (s1n1310,n644,n1311);
wire s0n1311,s1n1311,notn1311;
or (n1311,s0n1311,s1n1311);
not(notn1311,n568);
and (s0n1311,notn1311,n1312);
and (s1n1311,n568,n1314);
wire s0n1312,s1n1312,notn1312;
or (n1312,s0n1312,s1n1312);
not(notn1312,n15);
and (s0n1312,notn1312,1'b0);
and (s1n1312,n15,n1313);
or (n1314,1'b0,n1315,n1317,n1319,n1321);
and (n1315,n1316,n549);
and (n1317,n1318,n560);
and (n1319,n1320,n564);
and (n1321,n1313,n566);
wire s0n1322,s1n1322,notn1322;
or (n1322,s0n1322,s1n1322);
not(notn1322,n692);
and (s0n1322,notn1322,1'b0);
and (s1n1322,n692,n1295);
and (n1323,n1322,n1324);
or (n1324,n1325,n1339,n1421);
and (n1325,n1326,n1338);
wire s0n1326,s1n1326,notn1326;
or (n1326,s0n1326,s1n1326);
not(notn1326,n644);
and (s0n1326,notn1326,1'b0);
and (s1n1326,n644,n1327);
wire s0n1327,s1n1327,notn1327;
or (n1327,s0n1327,s1n1327);
not(notn1327,n568);
and (s0n1327,notn1327,n1328);
and (s1n1327,n568,n1330);
wire s0n1328,s1n1328,notn1328;
or (n1328,s0n1328,s1n1328);
not(notn1328,n15);
and (s0n1328,notn1328,1'b0);
and (s1n1328,n15,n1329);
or (n1330,1'b0,n1331,n1333,n1335,n1337);
and (n1331,n1332,n549);
and (n1333,n1334,n560);
and (n1335,n1336,n564);
and (n1337,n1329,n566);
wire s0n1338,s1n1338,notn1338;
or (n1338,s0n1338,s1n1338);
not(notn1338,n692);
and (s0n1338,notn1338,1'b0);
and (s1n1338,n692,n1311);
and (n1339,n1338,n1340);
or (n1340,n1341,n1355,n1420);
and (n1341,n1342,n1354);
wire s0n1342,s1n1342,notn1342;
or (n1342,s0n1342,s1n1342);
not(notn1342,n644);
and (s0n1342,notn1342,1'b0);
and (s1n1342,n644,n1343);
wire s0n1343,s1n1343,notn1343;
or (n1343,s0n1343,s1n1343);
not(notn1343,n568);
and (s0n1343,notn1343,n1344);
and (s1n1343,n568,n1346);
wire s0n1344,s1n1344,notn1344;
or (n1344,s0n1344,s1n1344);
not(notn1344,n15);
and (s0n1344,notn1344,1'b0);
and (s1n1344,n15,n1345);
or (n1346,1'b0,n1347,n1349,n1351,n1353);
and (n1347,n1348,n549);
and (n1349,n1350,n560);
and (n1351,n1352,n564);
and (n1353,n1345,n566);
wire s0n1354,s1n1354,notn1354;
or (n1354,s0n1354,s1n1354);
not(notn1354,n692);
and (s0n1354,notn1354,1'b0);
and (s1n1354,n692,n1327);
and (n1355,n1354,n1356);
or (n1356,n1357,n1371,n1419);
and (n1357,n1358,n1370);
wire s0n1358,s1n1358,notn1358;
or (n1358,s0n1358,s1n1358);
not(notn1358,n644);
and (s0n1358,notn1358,1'b0);
and (s1n1358,n644,n1359);
wire s0n1359,s1n1359,notn1359;
or (n1359,s0n1359,s1n1359);
not(notn1359,n568);
and (s0n1359,notn1359,n1360);
and (s1n1359,n568,n1362);
wire s0n1360,s1n1360,notn1360;
or (n1360,s0n1360,s1n1360);
not(notn1360,n15);
and (s0n1360,notn1360,1'b0);
and (s1n1360,n15,n1361);
or (n1362,1'b0,n1363,n1365,n1367,n1369);
and (n1363,n1364,n549);
and (n1365,n1366,n560);
and (n1367,n1368,n564);
and (n1369,n1361,n566);
wire s0n1370,s1n1370,notn1370;
or (n1370,s0n1370,s1n1370);
not(notn1370,n692);
and (s0n1370,notn1370,1'b0);
and (s1n1370,n692,n1343);
and (n1371,n1370,n1372);
or (n1372,n1373,n1387,n1389);
and (n1373,n1374,n1386);
wire s0n1374,s1n1374,notn1374;
or (n1374,s0n1374,s1n1374);
not(notn1374,n644);
and (s0n1374,notn1374,1'b0);
and (s1n1374,n644,n1375);
wire s0n1375,s1n1375,notn1375;
or (n1375,s0n1375,s1n1375);
not(notn1375,n568);
and (s0n1375,notn1375,n1376);
and (s1n1375,n568,n1378);
wire s0n1376,s1n1376,notn1376;
or (n1376,s0n1376,s1n1376);
not(notn1376,n15);
and (s0n1376,notn1376,1'b0);
and (s1n1376,n15,n1377);
or (n1378,1'b0,n1379,n1381,n1383,n1385);
and (n1379,n1380,n549);
and (n1381,n1382,n560);
and (n1383,n1384,n564);
and (n1385,n1377,n566);
wire s0n1386,s1n1386,notn1386;
or (n1386,s0n1386,s1n1386);
not(notn1386,n692);
and (s0n1386,notn1386,1'b0);
and (s1n1386,n692,n1359);
and (n1387,n1386,n1388);
or (n1388,n1389,n1404,n1405);
and (n1389,n1390,n1403);
not (n1390,n1391);
nand (n1391,n644,n1392);
wire s0n1392,s1n1392,notn1392;
or (n1392,s0n1392,s1n1392);
not(notn1392,n568);
and (s0n1392,notn1392,n1393);
and (s1n1392,n568,n1395);
wire s0n1393,s1n1393,notn1393;
or (n1393,s0n1393,s1n1393);
not(notn1393,n15);
and (s0n1393,notn1393,1'b0);
and (s1n1393,n15,n1394);
or (n1395,1'b0,n1396,n1398,n1400,n1402);
and (n1396,n1397,n549);
and (n1398,n1399,n560);
and (n1400,n1401,n564);
and (n1402,n1394,n566);
wire s0n1403,s1n1403,notn1403;
or (n1403,s0n1403,s1n1403);
not(notn1403,n692);
and (s0n1403,notn1403,1'b0);
and (s1n1403,n692,n1375);
and (n1404,n1403,n1405);
and (n1405,n1406,n1418);
wire s0n1406,s1n1406,notn1406;
or (n1406,s0n1406,s1n1406);
not(notn1406,n644);
and (s0n1406,notn1406,1'b0);
and (s1n1406,n644,n1407);
wire s0n1407,s1n1407,notn1407;
or (n1407,s0n1407,s1n1407);
not(notn1407,n568);
and (s0n1407,notn1407,n1408);
and (s1n1407,n568,n1410);
wire s0n1408,s1n1408,notn1408;
or (n1408,s0n1408,s1n1408);
not(notn1408,n15);
and (s0n1408,notn1408,1'b0);
and (s1n1408,n15,n1409);
or (n1410,1'b0,n1411,n1413,n1415,n1417);
and (n1411,n1412,n549);
and (n1413,n1414,n560);
and (n1415,n1416,n564);
and (n1417,n1409,n566);
wire s0n1418,s1n1418,notn1418;
or (n1418,s0n1418,s1n1418);
not(notn1418,n692);
and (s0n1418,notn1418,1'b0);
and (s1n1418,n692,n1392);
and (n1419,n1358,n1372);
and (n1420,n1342,n1356);
and (n1421,n1326,n1340);
and (n1422,n1310,n1324);
and (n1423,n1306,n1424);
or (n1424,n1425,n1429,n1475);
and (n1425,n1426,n1428);
not (n1426,n1427);
nand (n1427,n587,n1311);
xor (n1428,n1307,n1308);
and (n1429,n1428,n1430);
or (n1430,n1431,n1436,n1474);
and (n1431,n1432,n1434);
not (n1432,n1433);
nand (n1433,n587,n1327);
xor (n1434,n1435,n1324);
xor (n1435,n1310,n1322);
and (n1436,n1434,n1437);
or (n1437,n1438,n1443,n1473);
and (n1438,n1439,n1441);
not (n1439,n1440);
nand (n1440,n587,n1343);
xor (n1441,n1442,n1340);
xor (n1442,n1326,n1338);
and (n1443,n1441,n1444);
or (n1444,n1445,n1450,n1472);
and (n1445,n1446,n1448);
not (n1446,n1447);
nand (n1447,n587,n1359);
xor (n1448,n1449,n1356);
xor (n1449,n1342,n1354);
and (n1450,n1448,n1451);
or (n1451,n1452,n1457,n1471);
and (n1452,n1453,n1455);
not (n1453,n1454);
nand (n1454,n587,n1375);
xor (n1455,n1456,n1372);
xor (n1456,n1358,n1370);
and (n1457,n1455,n1458);
or (n1458,n1459,n1464,n1470);
and (n1459,n1460,n1462);
not (n1460,n1461);
nand (n1461,n587,n1392);
xor (n1462,n1463,n1388);
xor (n1463,n1374,n1386);
and (n1464,n1462,n1465);
and (n1465,n1466,n1468);
not (n1466,n1467);
nand (n1467,n587,n1407);
xor (n1468,n1469,n1405);
xor (n1469,n1390,n1403);
and (n1470,n1460,n1465);
and (n1471,n1453,n1458);
and (n1472,n1446,n1451);
and (n1473,n1439,n1444);
and (n1474,n1432,n1437);
and (n1475,n1426,n1430);
and (n1476,n1294,n1424);
or (n1477,n1478,n1633,n1718);
and (n1478,n1479,n1484);
xor (n1479,n1480,n1483);
wire s0n1480,s1n1480,notn1480;
or (n1480,s0n1480,s1n1480);
not(notn1480,n928);
and (s0n1480,notn1480,1'b0);
and (s1n1480,n928,n1481);
xor (n1481,n1482,n1424);
xor (n1482,n1294,n1306);
wire s0n1483,s1n1483,notn1483;
or (n1483,s0n1483,s1n1483);
not(notn1483,n1080);
and (s0n1483,notn1483,1'b0);
and (s1n1483,n1080,n1292);
and (n1484,n1485,n1486);
wire s0n1485,s1n1485,notn1485;
or (n1485,s0n1485,s1n1485);
not(notn1485,n1083);
and (s0n1485,notn1485,1'b0);
and (s1n1485,n1083,n1292);
or (n1486,n1487,n1490,n1632);
and (n1487,n1488,n1489);
wire s0n1488,s1n1488,notn1488;
or (n1488,s0n1488,s1n1488);
not(notn1488,n1083);
and (s0n1488,notn1488,1'b0);
and (s1n1488,n1083,n1481);
wire s0n1489,s1n1489,notn1489;
or (n1489,s0n1489,s1n1489);
not(notn1489,n1027);
and (s0n1489,notn1489,1'b0);
and (s1n1489,n1027,n1292);
and (n1490,n1489,n1491);
or (n1491,n1492,n1578,n1631);
and (n1492,n1493,n1577);
and (n1493,n1494,n1083);
xor (n1494,n1495,n1508);
xor (n1495,n1496,n1504);
nand (n1496,n1497,n1501);
or (n1497,n1498,n1500);
and (n1498,n1499,n1433);
not (n1499,n1322);
not (n1500,n1310);
or (n1501,n1502,n1503);
not (n1502,n1354);
not (n1503,n1294);
not (n1504,n1505);
xnor (n1505,n1506,n1507);
not (n1506,n1426);
not (n1507,n1307);
or (n1508,n1509,n1576);
and (n1509,n1510,n1522);
xor (n1510,n1511,n1516);
nor (n1511,n1512,n1514);
and (n1512,n1513,n1310);
xor (n1513,n1499,n1433);
and (n1514,n1515,n1500);
not (n1515,n1513);
nand (n1516,n1517,n1519,n1521);
or (n1517,n1433,n1518);
not (n1518,n1342);
or (n1519,n1440,n1520);
not (n1520,n1338);
not (n1521,n1325);
nand (n1522,n1523,n1575);
or (n1523,n1524,n1536);
not (n1524,n1525);
nand (n1525,n1526,n1528);
xor (n1526,n1442,n1527);
not (n1527,n1439);
not (n1528,n1529);
nand (n1529,n1530,n1533,n1535);
or (n1530,n1531,n1532);
not (n1531,n1386);
not (n1532,n1432);
or (n1533,n1527,n1534);
not (n1534,n1358);
not (n1535,n1341);
not (n1536,n1537);
or (n1537,n1538,n1574);
and (n1538,n1539,n1549);
xor (n1539,n1540,n1546);
nand (n1540,n1541,n1543,n1545);
or (n1541,n1440,n1542);
not (n1542,n1403);
or (n1543,n1447,n1544);
not (n1544,n1374);
not (n1545,n1357);
nand (n1546,n1547,n1548);
or (n1547,n1447,n1449);
nand (n1548,n1449,n1447);
or (n1549,n1550,n1573);
and (n1550,n1551,n1560);
xor (n1551,n1552,n1558);
nand (n1552,n1553,n1555,n1557);
not (n1553,n1554);
and (n1554,n1453,n1390);
or (n1555,n1447,n1556);
not (n1556,n1418);
not (n1557,n1373);
xnor (n1558,n1559,n1456);
not (n1559,n1453);
or (n1560,n1561,n1572);
and (n1561,n1562,n1568);
xor (n1562,n1563,n1564);
nor (n1563,n1467,n1542);
xnor (n1564,n1565,n1544);
nand (n1565,n1566,n1567);
or (n1566,n1460,n1531);
nand (n1567,n1460,n1531);
nand (n1568,n1569,n1571);
or (n1569,n1570,n1391);
xnor (n1570,n1542,n1467);
not (n1571,n1405);
and (n1572,n1563,n1564);
and (n1573,n1552,n1558);
and (n1574,n1540,n1546);
or (n1575,n1526,n1528);
and (n1576,n1511,n1516);
wire s0n1577,s1n1577,notn1577;
or (n1577,s0n1577,s1n1577);
not(notn1577,n1027);
and (s0n1577,notn1577,1'b0);
and (s1n1577,n1027,n1481);
and (n1578,n1577,n1579);
or (n1579,n1580,n1584,n1630);
and (n1580,n1581,n1583);
and (n1581,n1582,n1083);
xor (n1582,n1510,n1522);
wire s0n1583,s1n1583,notn1583;
or (n1583,s0n1583,s1n1583);
not(notn1583,n1027);
and (s0n1583,notn1583,1'b0);
and (s1n1583,n1027,n1494);
and (n1584,n1583,n1585);
or (n1585,n1586,n1591,n1629);
and (n1586,n1587,n1590);
wire s0n1587,s1n1587,notn1587;
or (n1587,s0n1587,s1n1587);
not(notn1587,n1083);
and (s0n1587,notn1587,1'b0);
and (s1n1587,n1083,n1588);
xor (n1588,n1589,n1444);
xor (n1589,n1439,n1441);
wire s0n1590,s1n1590,notn1590;
or (n1590,s0n1590,s1n1590);
not(notn1590,n1027);
and (s0n1590,notn1590,1'b0);
and (s1n1590,n1027,n1582);
and (n1591,n1590,n1592);
or (n1592,n1593,n1597,n1628);
and (n1593,n1594,n1596);
and (n1594,n1595,n1083);
xor (n1595,n1539,n1549);
wire s0n1596,s1n1596,notn1596;
or (n1596,s0n1596,s1n1596);
not(notn1596,n1027);
and (s0n1596,notn1596,1'b0);
and (s1n1596,n1027,n1588);
and (n1597,n1596,n1598);
or (n1598,n1599,n1603,n1627);
and (n1599,n1600,n1602);
and (n1600,n1601,n1083);
xor (n1601,n1551,n1560);
wire s0n1602,s1n1602,notn1602;
or (n1602,s0n1602,s1n1602);
not(notn1602,n1027);
and (s0n1602,notn1602,1'b0);
and (s1n1602,n1027,n1595);
and (n1603,n1602,n1604);
or (n1604,n1605,n1609,n1626);
and (n1605,n1606,n1608);
and (n1606,n1607,n1083);
xor (n1607,n1562,n1568);
wire s0n1608,s1n1608,notn1608;
or (n1608,s0n1608,s1n1608);
not(notn1608,n1027);
and (s0n1608,notn1608,1'b0);
and (s1n1608,n1027,n1601);
and (n1609,n1608,n1610);
or (n1610,n1611,n1615,n1617);
and (n1611,n1612,n1614);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n1083);
and (s0n1612,notn1612,1'b0);
and (s1n1612,n1083,n1613);
xor (n1613,n1466,n1468);
wire s0n1614,s1n1614,notn1614;
or (n1614,s0n1614,s1n1614);
not(notn1614,n1027);
and (s0n1614,notn1614,1'b0);
and (s1n1614,n1027,n1607);
and (n1615,n1614,n1616);
or (n1616,n1617,n1621,n1622);
and (n1617,n1618,n1620);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n1083);
and (s0n1618,notn1618,1'b0);
and (s1n1618,n1083,n1619);
xor (n1619,n1406,n1418);
wire s0n1620,s1n1620,notn1620;
or (n1620,s0n1620,s1n1620);
not(notn1620,n1027);
and (s0n1620,notn1620,1'b0);
and (s1n1620,n1027,n1613);
and (n1621,n1620,n1622);
and (n1622,n1623,n1625);
wire s0n1623,s1n1623,notn1623;
or (n1623,s0n1623,s1n1623);
not(notn1623,n1083);
and (s0n1623,notn1623,1'b0);
and (s1n1623,n1083,n1624);
wire s0n1624,s1n1624,notn1624;
or (n1624,s0n1624,s1n1624);
not(notn1624,n692);
and (s0n1624,notn1624,1'b0);
and (s1n1624,n692,n1407);
wire s0n1625,s1n1625,notn1625;
or (n1625,s0n1625,s1n1625);
not(notn1625,n1027);
and (s0n1625,notn1625,1'b0);
and (s1n1625,n1027,n1619);
and (n1626,n1606,n1610);
and (n1627,n1600,n1604);
and (n1628,n1594,n1598);
and (n1629,n1587,n1592);
and (n1630,n1581,n1585);
and (n1631,n1493,n1579);
and (n1632,n1488,n1491);
and (n1633,n1484,n1634);
or (n1634,n1635,n1640,n1717);
and (n1635,n1636,n1639);
xor (n1636,n1637,n1638);
and (n1637,n1494,n928);
wire s0n1638,s1n1638,notn1638;
or (n1638,s0n1638,s1n1638);
not(notn1638,n1080);
and (s0n1638,notn1638,1'b0);
and (s1n1638,n1080,n1481);
xor (n1639,n1485,n1486);
and (n1640,n1639,n1641);
or (n1641,n1642,n1648,n1716);
and (n1642,n1643,n1646);
xor (n1643,n1644,n1645);
and (n1644,n1582,n928);
and (n1645,n1494,n1080);
xor (n1646,n1647,n1491);
xor (n1647,n1488,n1489);
and (n1648,n1646,n1649);
or (n1649,n1650,n1656,n1715);
and (n1650,n1651,n1654);
xor (n1651,n1652,n1653);
wire s0n1652,s1n1652,notn1652;
or (n1652,s0n1652,s1n1652);
not(notn1652,n928);
and (s0n1652,notn1652,1'b0);
and (s1n1652,n928,n1588);
and (n1653,n1582,n1080);
xor (n1654,n1655,n1579);
xor (n1655,n1493,n1577);
and (n1656,n1654,n1657);
or (n1657,n1658,n1664,n1714);
and (n1658,n1659,n1662);
xor (n1659,n1660,n1661);
and (n1660,n1595,n928);
wire s0n1661,s1n1661,notn1661;
or (n1661,s0n1661,s1n1661);
not(notn1661,n1080);
and (s0n1661,notn1661,1'b0);
and (s1n1661,n1080,n1588);
xor (n1662,n1663,n1585);
xor (n1663,n1581,n1583);
and (n1664,n1662,n1665);
or (n1665,n1666,n1672,n1713);
and (n1666,n1667,n1670);
xor (n1667,n1668,n1669);
and (n1668,n1601,n928);
and (n1669,n1595,n1080);
xor (n1670,n1671,n1592);
xor (n1671,n1587,n1590);
and (n1672,n1670,n1673);
or (n1673,n1674,n1680,n1712);
and (n1674,n1675,n1678);
xor (n1675,n1676,n1677);
and (n1676,n1607,n928);
and (n1677,n1601,n1080);
xor (n1678,n1679,n1598);
xor (n1679,n1594,n1596);
and (n1680,n1678,n1681);
or (n1681,n1682,n1688,n1711);
and (n1682,n1683,n1686);
xor (n1683,n1684,n1685);
wire s0n1684,s1n1684,notn1684;
or (n1684,s0n1684,s1n1684);
not(notn1684,n928);
and (s0n1684,notn1684,1'b0);
and (s1n1684,n928,n1613);
and (n1685,n1607,n1080);
xor (n1686,n1687,n1604);
xor (n1687,n1600,n1602);
and (n1688,n1686,n1689);
or (n1689,n1690,n1696,n1710);
and (n1690,n1691,n1694);
xor (n1691,n1692,n1693);
and (n1692,n928,n1619);
wire s0n1693,s1n1693,notn1693;
or (n1693,s0n1693,s1n1693);
not(notn1693,n1080);
and (s0n1693,notn1693,1'b0);
and (s1n1693,n1080,n1613);
xor (n1694,n1695,n1610);
xor (n1695,n1606,n1608);
and (n1696,n1694,n1697);
or (n1697,n1698,n1704,n1709);
and (n1698,n1699,n1702);
xor (n1699,n1700,n1701);
wire s0n1700,s1n1700,notn1700;
or (n1700,s0n1700,s1n1700);
not(notn1700,n928);
and (s0n1700,notn1700,1'b0);
and (s1n1700,n928,n1624);
and (n1701,n1080,n1619);
xor (n1702,n1703,n1616);
xor (n1703,n1612,n1614);
and (n1704,n1702,n1705);
and (n1705,n1706,n1707);
wire s0n1706,s1n1706,notn1706;
or (n1706,s0n1706,s1n1706);
not(notn1706,n1080);
and (s0n1706,notn1706,1'b0);
and (s1n1706,n1080,n1624);
xor (n1707,n1708,n1622);
xor (n1708,n1618,n1620);
and (n1709,n1699,n1705);
and (n1710,n1691,n1697);
and (n1711,n1683,n1689);
and (n1712,n1675,n1681);
and (n1713,n1667,n1673);
and (n1714,n1659,n1665);
and (n1715,n1651,n1657);
and (n1716,n1643,n1649);
and (n1717,n1636,n1641);
and (n1718,n1479,n1634);
or (n1719,n1720,n1725,n1813);
and (n1720,n1721,n1723);
xor (n1721,n1722,n1205);
xor (n1722,n1076,n1081);
xor (n1723,n1724,n1634);
xor (n1724,n1479,n1484);
and (n1725,n1723,n1726);
or (n1726,n1727,n1732,n1812);
and (n1727,n1728,n1730);
xor (n1728,n1729,n1212);
xor (n1729,n1207,n1210);
xor (n1730,n1731,n1641);
xor (n1731,n1636,n1639);
and (n1732,n1730,n1733);
or (n1733,n1734,n1739,n1811);
and (n1734,n1735,n1737);
xor (n1735,n1736,n1220);
xor (n1736,n1214,n1217);
xor (n1737,n1738,n1649);
xor (n1738,n1643,n1646);
and (n1739,n1737,n1740);
or (n1740,n1741,n1746,n1810);
and (n1741,n1742,n1744);
xor (n1742,n1743,n1228);
xor (n1743,n1222,n1225);
xor (n1744,n1745,n1657);
xor (n1745,n1651,n1654);
and (n1746,n1744,n1747);
or (n1747,n1748,n1753,n1809);
and (n1748,n1749,n1751);
xor (n1749,n1750,n1236);
xor (n1750,n1230,n1233);
xor (n1751,n1752,n1665);
xor (n1752,n1659,n1662);
and (n1753,n1751,n1754);
or (n1754,n1755,n1760,n1808);
and (n1755,n1756,n1758);
xor (n1756,n1757,n1244);
xor (n1757,n1238,n1241);
xor (n1758,n1759,n1673);
xor (n1759,n1667,n1670);
and (n1760,n1758,n1761);
or (n1761,n1762,n1767,n1807);
and (n1762,n1763,n1765);
xor (n1763,n1764,n1252);
xor (n1764,n1246,n1249);
xor (n1765,n1766,n1681);
xor (n1766,n1675,n1678);
and (n1767,n1765,n1768);
or (n1768,n1769,n1774,n1806);
and (n1769,n1770,n1772);
xor (n1770,n1771,n1260);
xor (n1771,n1254,n1257);
xor (n1772,n1773,n1689);
xor (n1773,n1683,n1686);
and (n1774,n1772,n1775);
or (n1775,n1776,n1781,n1805);
and (n1776,n1777,n1779);
xor (n1777,n1778,n1268);
xor (n1778,n1262,n1265);
xor (n1779,n1780,n1697);
xor (n1780,n1691,n1694);
and (n1781,n1779,n1782);
or (n1782,n1783,n1788,n1804);
and (n1783,n1784,n1786);
xor (n1784,n1785,n1276);
xor (n1785,n1270,n1273);
xor (n1786,n1787,n1705);
xor (n1787,n1699,n1702);
and (n1788,n1786,n1789);
or (n1789,n1790,n1793,n1803);
and (n1790,n1791,n1792);
xor (n1791,n1277,n1278);
xor (n1792,n1706,n1707);
and (n1793,n1792,n1794);
or (n1794,n1795,n1798,n1802);
and (n1795,n1796,n1797);
xor (n1796,n1194,n1196);
xor (n1797,n1623,n1625);
and (n1798,n1797,n1799);
and (n1799,n1800,n1801);
wire s0n1800,s1n1800,notn1800;
or (n1800,s0n1800,s1n1800);
not(notn1800,n1027);
and (s0n1800,notn1800,1'b0);
and (s1n1800,n1027,n1195);
wire s0n1801,s1n1801,notn1801;
or (n1801,s0n1801,s1n1801);
not(notn1801,n1027);
and (s0n1801,notn1801,1'b0);
and (s1n1801,n1027,n1624);
and (n1802,n1796,n1799);
and (n1803,n1791,n1794);
and (n1804,n1784,n1789);
and (n1805,n1777,n1782);
and (n1806,n1770,n1775);
and (n1807,n1763,n1768);
and (n1808,n1756,n1761);
and (n1809,n1749,n1754);
and (n1810,n1742,n1747);
and (n1811,n1735,n1740);
and (n1812,n1728,n1733);
and (n1813,n1721,n1726);
xor (n1814,n1815,n2475);
xor (n1815,n1816,n2153);
or (n1816,n1817,n2085,n2152);
and (n1817,n1818,n2018);
and (n1818,n1819,n930);
xnor (n1819,n1820,n1833);
not (n1820,n1821);
and (n1821,n585,n1822);
wire s0n1822,s1n1822,notn1822;
or (n1822,s0n1822,s1n1822);
not(notn1822,n568);
and (s0n1822,notn1822,n1823);
and (s1n1822,n568,n1825);
wire s0n1823,s1n1823,notn1823;
or (n1823,s0n1823,s1n1823);
not(notn1823,n15);
and (s0n1823,notn1823,1'b0);
and (s1n1823,n15,n1824);
or (n1825,1'b0,n1826,n1828,n1830,n1832);
and (n1826,n1827,n549);
and (n1828,n1829,n560);
and (n1830,n1831,n564);
and (n1832,n1824,n566);
or (n1833,n1834,n1871);
and (n1834,n1835,n1872);
xor (n1835,n1836,n1850);
xor (n1836,n1837,n1838);
and (n1837,n756,n1822);
and (n1838,n585,n1839);
wire s0n1839,s1n1839,notn1839;
or (n1839,s0n1839,s1n1839);
not(notn1839,n568);
and (s0n1839,notn1839,n1840);
and (s1n1839,n568,n1842);
wire s0n1840,s1n1840,notn1840;
or (n1840,s0n1840,s1n1840);
not(notn1840,n15);
and (s0n1840,notn1840,1'b0);
and (s1n1840,n15,n1841);
or (n1842,1'b0,n1843,n1845,n1847,n1849);
and (n1843,n1844,n549);
and (n1845,n1846,n560);
and (n1847,n1848,n564);
and (n1849,n1841,n566);
or (n1850,n1851,n1871);
and (n1851,n1852,n1868);
xor (n1852,n1853,n1867);
xor (n1853,n1854,n1855);
and (n1854,n763,n1822);
and (n1855,n585,n1856);
wire s0n1856,s1n1856,notn1856;
or (n1856,s0n1856,s1n1856);
not(notn1856,n568);
and (s0n1856,notn1856,n1857);
and (s1n1856,n568,n1859);
wire s0n1857,s1n1857,notn1857;
or (n1857,s0n1857,s1n1857);
not(notn1857,n15);
and (s0n1857,notn1857,1'b0);
and (s1n1857,n15,n1858);
or (n1859,1'b0,n1860,n1862,n1864,n1866);
and (n1860,n1861,n549);
and (n1862,n1863,n560);
and (n1864,n1865,n564);
and (n1866,n1858,n566);
and (n1867,n756,n1839);
and (n1868,n1869,n1870);
and (n1869,n763,n1839);
wire s0n1870,s1n1870,notn1870;
or (n1870,s0n1870,s1n1870);
not(notn1870,n692);
and (s0n1870,notn1870,1'b0);
and (s1n1870,n692,n1822);
and (n1871,n1853,n1867);
or (n1872,n1873,n2017);
and (n1873,n1874,n1898);
xor (n1874,n1875,n1897);
or (n1875,n1876,n1896);
and (n1876,n1877,n1893);
xor (n1877,n1878,n1892);
xor (n1878,n1879,n1880);
xor (n1879,n1869,n1870);
and (n1880,n585,n1881);
wire s0n1881,s1n1881,notn1881;
or (n1881,s0n1881,s1n1881);
not(notn1881,n568);
and (s0n1881,notn1881,n1882);
and (s1n1881,n568,n1884);
wire s0n1882,s1n1882,notn1882;
or (n1882,s0n1882,s1n1882);
not(notn1882,n15);
and (s0n1882,notn1882,1'b0);
and (s1n1882,n15,n1883);
or (n1884,1'b0,n1885,n1887,n1889,n1891);
and (n1885,n1886,n549);
and (n1887,n1888,n560);
and (n1889,n1890,n564);
and (n1891,n1883,n566);
and (n1892,n756,n1856);
and (n1893,n1894,n1895);
wire s0n1894,s1n1894,notn1894;
or (n1894,s0n1894,s1n1894);
not(notn1894,n692);
and (s0n1894,notn1894,1'b0);
and (s1n1894,n692,n1839);
and (n1895,n763,n1856);
and (n1896,n1878,n1892);
xor (n1897,n1852,n1868);
or (n1898,n1899,n2016);
and (n1899,n1900,n1924);
xor (n1900,n1901,n1923);
or (n1901,n1902,n1922);
and (n1902,n1903,n1919);
xor (n1903,n1904,n1905);
and (n1904,n756,n1881);
xor (n1905,n1906,n1907);
xor (n1906,n1894,n1895);
and (n1907,n585,n1908);
wire s0n1908,s1n1908,notn1908;
or (n1908,s0n1908,s1n1908);
not(notn1908,n568);
and (s0n1908,notn1908,n1909);
and (s1n1908,n568,n1911);
wire s0n1909,s1n1909,notn1909;
or (n1909,s0n1909,s1n1909);
not(notn1909,n15);
and (s0n1909,notn1909,1'b0);
and (s1n1909,n15,n1910);
or (n1911,1'b0,n1912,n1914,n1916,n1918);
and (n1912,n1913,n549);
and (n1914,n1915,n560);
and (n1916,n1917,n564);
and (n1918,n1910,n566);
and (n1919,n1920,n1921);
wire s0n1920,s1n1920,notn1920;
or (n1920,s0n1920,s1n1920);
not(notn1920,n692);
and (s0n1920,notn1920,1'b0);
and (s1n1920,n692,n1856);
and (n1921,n763,n1881);
and (n1922,n1904,n1905);
xor (n1923,n1877,n1893);
or (n1924,n1925,n2015);
and (n1925,n1926,n1950);
xor (n1926,n1927,n1949);
or (n1927,n1928,n1948);
and (n1928,n1929,n1945);
xor (n1929,n1930,n1931);
and (n1930,n756,n1908);
xor (n1931,n1932,n1933);
xor (n1932,n1920,n1921);
and (n1933,n585,n1934);
wire s0n1934,s1n1934,notn1934;
or (n1934,s0n1934,s1n1934);
not(notn1934,n568);
and (s0n1934,notn1934,n1935);
and (s1n1934,n568,n1937);
wire s0n1935,s1n1935,notn1935;
or (n1935,s0n1935,s1n1935);
not(notn1935,n15);
and (s0n1935,notn1935,1'b0);
and (s1n1935,n15,n1936);
or (n1937,1'b0,n1938,n1940,n1942,n1944);
and (n1938,n1939,n549);
and (n1940,n1941,n560);
and (n1942,n1943,n564);
and (n1944,n1936,n566);
and (n1945,n1946,n1947);
and (n1946,n763,n1908);
wire s0n1947,s1n1947,notn1947;
or (n1947,s0n1947,s1n1947);
not(notn1947,n692);
and (s0n1947,notn1947,1'b0);
and (s1n1947,n692,n1881);
and (n1948,n1930,n1931);
xor (n1949,n1903,n1919);
or (n1950,n1951,n2014);
and (n1951,n1952,n1976);
xor (n1952,n1953,n1975);
or (n1953,n1954,n1974);
and (n1954,n1955,n1960);
xor (n1955,n1956,n1957);
and (n1956,n756,n1934);
and (n1957,n1958,n1959);
wire s0n1958,s1n1958,notn1958;
or (n1958,s0n1958,s1n1958);
not(notn1958,n692);
and (s0n1958,notn1958,1'b0);
and (s1n1958,n692,n1908);
and (n1959,n763,n1934);
xor (n1960,n1961,n1962);
xor (n1961,n1946,n1947);
and (n1962,n585,n1963);
wire s0n1963,s1n1963,notn1963;
or (n1963,s0n1963,s1n1963);
not(notn1963,n568);
and (s0n1963,notn1963,n1964);
and (s1n1963,n568,n1966);
wire s0n1964,s1n1964,notn1964;
or (n1964,s0n1964,s1n1964);
not(notn1964,n15);
and (s0n1964,notn1964,1'b0);
and (s1n1964,n15,n1965);
or (n1966,1'b0,n1967,n1969,n1971,n1973);
and (n1967,n1968,n549);
and (n1969,n1970,n560);
and (n1971,n1972,n564);
and (n1973,n1965,n566);
and (n1974,n1956,n1957);
xor (n1975,n1929,n1945);
or (n1976,n1977,n2013);
and (n1977,n1978,n1996);
xor (n1978,n1979,n1995);
and (n1979,n1980,n1994);
xor (n1980,n1981,n1993);
and (n1981,n585,n1982);
wire s0n1982,s1n1982,notn1982;
or (n1982,s0n1982,s1n1982);
not(notn1982,n568);
and (s0n1982,notn1982,n1983);
and (s1n1982,n568,n1985);
wire s0n1983,s1n1983,notn1983;
or (n1983,s0n1983,s1n1983);
not(notn1983,n15);
and (s0n1983,notn1983,1'b0);
and (s1n1983,n15,n1984);
or (n1985,1'b0,n1986,n1988,n1990,n1992);
and (n1986,n1987,n549);
and (n1988,n1989,n560);
and (n1990,n1991,n564);
and (n1992,n1984,n566);
and (n1993,n756,n1963);
xor (n1994,n1958,n1959);
xor (n1995,n1955,n1960);
or (n1996,n1997,n2012);
and (n1997,n1998,n2011);
xor (n1998,n1999,n2002);
and (n1999,n2000,n2001);
wire s0n2000,s1n2000,notn2000;
or (n2000,s0n2000,s1n2000);
not(notn2000,n692);
and (s0n2000,notn2000,1'b0);
and (s1n2000,n692,n1934);
and (n2001,n763,n1963);
or (n2002,n2003,n2010);
and (n2003,n2004,n2009);
xor (n2004,n2005,n2008);
and (n2005,n2006,n2007);
and (n2006,n763,n1982);
wire s0n2007,s1n2007,notn2007;
or (n2007,s0n2007,s1n2007);
not(notn2007,n692);
and (s0n2007,notn2007,1'b0);
and (s1n2007,n692,n1963);
xor (n2008,n2000,n2001);
and (n2009,n756,n1982);
and (n2010,n2005,n2008);
xor (n2011,n1980,n1994);
and (n2012,n1999,n2002);
and (n2013,n1979,n1995);
and (n2014,n1953,n1975);
and (n2015,n1927,n1949);
and (n2016,n1901,n1923);
and (n2017,n1875,n1897);
and (n2018,n2019,n2020);
and (n2019,n1819,n979);
or (n2020,n2021,n2025,n2084);
and (n2021,n2022,n2024);
and (n2022,n2023,n979);
xor (n2023,n1835,n1872);
and (n2024,n1819,n1027);
and (n2025,n2024,n2026);
or (n2026,n2027,n2031,n2083);
and (n2027,n2028,n2030);
and (n2028,n2029,n979);
xor (n2029,n1874,n1898);
and (n2030,n2023,n1027);
and (n2031,n2030,n2032);
or (n2032,n2033,n2037,n2082);
and (n2033,n2034,n2036);
and (n2034,n2035,n979);
xor (n2035,n1900,n1924);
and (n2036,n2029,n1027);
and (n2037,n2036,n2038);
or (n2038,n2039,n2043,n2081);
and (n2039,n2040,n2042);
and (n2040,n2041,n979);
xor (n2041,n1926,n1950);
and (n2042,n2035,n1027);
and (n2043,n2042,n2044);
or (n2044,n2045,n2049,n2080);
and (n2045,n2046,n2048);
and (n2046,n2047,n979);
xor (n2047,n1952,n1976);
and (n2048,n2041,n1027);
and (n2049,n2048,n2050);
or (n2050,n2051,n2055,n2079);
and (n2051,n2052,n2054);
and (n2052,n2053,n979);
xor (n2053,n1978,n1996);
and (n2054,n2047,n1027);
and (n2055,n2054,n2056);
or (n2056,n2057,n2061,n2078);
and (n2057,n2058,n2060);
and (n2058,n2059,n979);
xor (n2059,n1998,n2011);
and (n2060,n2053,n1027);
and (n2061,n2060,n2062);
or (n2062,n2063,n2067,n2069);
and (n2063,n2064,n2066);
and (n2064,n2065,n979);
xor (n2065,n2004,n2009);
and (n2066,n2059,n1027);
and (n2067,n2066,n2068);
or (n2068,n2069,n2073,n2074);
and (n2069,n2070,n2072);
and (n2070,n2071,n979);
xor (n2071,n2006,n2007);
and (n2072,n2065,n1027);
and (n2073,n2072,n2074);
and (n2074,n2075,n2077);
wire s0n2075,s1n2075,notn2075;
or (n2075,s0n2075,s1n2075);
not(notn2075,n979);
and (s0n2075,notn2075,1'b0);
and (s1n2075,n979,n2076);
wire s0n2076,s1n2076,notn2076;
or (n2076,s0n2076,s1n2076);
not(notn2076,n692);
and (s0n2076,notn2076,1'b0);
and (s1n2076,n692,n1982);
and (n2077,n2071,n1027);
and (n2078,n2058,n2062);
and (n2079,n2052,n2056);
and (n2080,n2046,n2050);
and (n2081,n2040,n2044);
and (n2082,n2034,n2038);
and (n2083,n2028,n2032);
and (n2084,n2022,n2026);
and (n2085,n2018,n2086);
or (n2086,n2087,n2090,n2151);
and (n2087,n2088,n2089);
and (n2088,n2023,n930);
xor (n2089,n2019,n2020);
and (n2090,n2089,n2091);
or (n2091,n2092,n2096,n2150);
and (n2092,n2093,n2094);
and (n2093,n2029,n930);
xor (n2094,n2095,n2026);
xor (n2095,n2022,n2024);
and (n2096,n2094,n2097);
or (n2097,n2098,n2102,n2149);
and (n2098,n2099,n2100);
and (n2099,n2035,n930);
xor (n2100,n2101,n2032);
xor (n2101,n2028,n2030);
and (n2102,n2100,n2103);
or (n2103,n2104,n2108,n2148);
and (n2104,n2105,n2106);
and (n2105,n2041,n930);
xor (n2106,n2107,n2038);
xor (n2107,n2034,n2036);
and (n2108,n2106,n2109);
or (n2109,n2110,n2114,n2147);
and (n2110,n2111,n2112);
and (n2111,n2047,n930);
xor (n2112,n2113,n2044);
xor (n2113,n2040,n2042);
and (n2114,n2112,n2115);
or (n2115,n2116,n2120,n2146);
and (n2116,n2117,n2118);
and (n2117,n2053,n930);
xor (n2118,n2119,n2050);
xor (n2119,n2046,n2048);
and (n2120,n2118,n2121);
or (n2121,n2122,n2126,n2145);
and (n2122,n2123,n2124);
and (n2123,n2059,n930);
xor (n2124,n2125,n2056);
xor (n2125,n2052,n2054);
and (n2126,n2124,n2127);
or (n2127,n2128,n2132,n2144);
and (n2128,n2129,n2130);
and (n2129,n2065,n930);
xor (n2130,n2131,n2062);
xor (n2131,n2058,n2060);
and (n2132,n2130,n2133);
or (n2133,n2134,n2138,n2143);
and (n2134,n2135,n2136);
and (n2135,n2071,n930);
xor (n2136,n2137,n2068);
xor (n2137,n2064,n2066);
and (n2138,n2136,n2139);
and (n2139,n2140,n2141);
wire s0n2140,s1n2140,notn2140;
or (n2140,s0n2140,s1n2140);
not(notn2140,n930);
and (s0n2140,notn2140,1'b0);
and (s1n2140,n930,n2076);
xor (n2141,n2142,n2074);
xor (n2142,n2070,n2072);
and (n2143,n2135,n2139);
and (n2144,n2129,n2133);
and (n2145,n2123,n2127);
and (n2146,n2117,n2121);
and (n2147,n2111,n2115);
and (n2148,n2105,n2109);
and (n2149,n2099,n2103);
and (n2150,n2093,n2097);
and (n2151,n2088,n2091);
and (n2152,n1818,n2086);
or (n2153,n2154,n2407,n2474);
and (n2154,n2155,n2333);
wire s0n2155,s1n2155,notn2155;
or (n2155,s0n2155,s1n2155);
not(notn2155,n930);
and (s0n2155,notn2155,1'b0);
and (s1n2155,n930,n2156);
or (n2156,n2157,n2286,n2332);
and (n2157,n2158,n2170);
wire s0n2158,s1n2158,notn2158;
or (n2158,s0n2158,s1n2158);
not(notn2158,n587);
and (s0n2158,notn2158,1'b0);
and (s1n2158,n587,n2159);
wire s0n2159,s1n2159,notn2159;
or (n2159,s0n2159,s1n2159);
not(notn2159,n568);
and (s0n2159,notn2159,n2160);
and (s1n2159,n568,n2162);
wire s0n2160,s1n2160,notn2160;
or (n2160,s0n2160,s1n2160);
not(notn2160,n15);
and (s0n2160,notn2160,1'b0);
and (s1n2160,n15,n2161);
or (n2162,1'b0,n2163,n2165,n2167,n2169);
and (n2163,n2164,n549);
and (n2165,n2166,n560);
and (n2167,n2168,n564);
and (n2169,n2161,n566);
and (n2170,n2171,n2172);
wire s0n2171,s1n2171,notn2171;
or (n2171,s0n2171,s1n2171);
not(notn2171,n644);
and (s0n2171,notn2171,1'b0);
and (s1n2171,n644,n2159);
or (n2172,n2173,n2187,n2285);
and (n2173,n2174,n2186);
wire s0n2174,s1n2174,notn2174;
or (n2174,s0n2174,s1n2174);
not(notn2174,n644);
and (s0n2174,notn2174,1'b0);
and (s1n2174,n644,n2175);
wire s0n2175,s1n2175,notn2175;
or (n2175,s0n2175,s1n2175);
not(notn2175,n568);
and (s0n2175,notn2175,n2176);
and (s1n2175,n568,n2178);
wire s0n2176,s1n2176,notn2176;
or (n2176,s0n2176,s1n2176);
not(notn2176,n15);
and (s0n2176,notn2176,1'b0);
and (s1n2176,n15,n2177);
or (n2178,1'b0,n2179,n2181,n2183,n2185);
and (n2179,n2180,n549);
and (n2181,n2182,n560);
and (n2183,n2184,n564);
and (n2185,n2177,n566);
wire s0n2186,s1n2186,notn2186;
or (n2186,s0n2186,s1n2186);
not(notn2186,n692);
and (s0n2186,notn2186,1'b0);
and (s1n2186,n692,n2159);
and (n2187,n2186,n2188);
or (n2188,n2189,n2203,n2284);
and (n2189,n2190,n2202);
wire s0n2190,s1n2190,notn2190;
or (n2190,s0n2190,s1n2190);
not(notn2190,n644);
and (s0n2190,notn2190,1'b0);
and (s1n2190,n644,n2191);
wire s0n2191,s1n2191,notn2191;
or (n2191,s0n2191,s1n2191);
not(notn2191,n568);
and (s0n2191,notn2191,n2192);
and (s1n2191,n568,n2194);
wire s0n2192,s1n2192,notn2192;
or (n2192,s0n2192,s1n2192);
not(notn2192,n15);
and (s0n2192,notn2192,1'b0);
and (s1n2192,n15,n2193);
or (n2194,1'b0,n2195,n2197,n2199,n2201);
and (n2195,n2196,n549);
and (n2197,n2198,n560);
and (n2199,n2200,n564);
and (n2201,n2193,n566);
wire s0n2202,s1n2202,notn2202;
or (n2202,s0n2202,s1n2202);
not(notn2202,n692);
and (s0n2202,notn2202,1'b0);
and (s1n2202,n692,n2175);
and (n2203,n2202,n2204);
or (n2204,n2205,n2219,n2283);
and (n2205,n2206,n2218);
wire s0n2206,s1n2206,notn2206;
or (n2206,s0n2206,s1n2206);
not(notn2206,n644);
and (s0n2206,notn2206,1'b0);
and (s1n2206,n644,n2207);
wire s0n2207,s1n2207,notn2207;
or (n2207,s0n2207,s1n2207);
not(notn2207,n568);
and (s0n2207,notn2207,n2208);
and (s1n2207,n568,n2210);
wire s0n2208,s1n2208,notn2208;
or (n2208,s0n2208,s1n2208);
not(notn2208,n15);
and (s0n2208,notn2208,1'b0);
and (s1n2208,n15,n2209);
or (n2210,1'b0,n2211,n2213,n2215,n2217);
and (n2211,n2212,n549);
and (n2213,n2214,n560);
and (n2215,n2216,n564);
and (n2217,n2209,n566);
wire s0n2218,s1n2218,notn2218;
or (n2218,s0n2218,s1n2218);
not(notn2218,n692);
and (s0n2218,notn2218,1'b0);
and (s1n2218,n692,n2191);
and (n2219,n2218,n2220);
or (n2220,n2221,n2235,n2282);
and (n2221,n2222,n2234);
wire s0n2222,s1n2222,notn2222;
or (n2222,s0n2222,s1n2222);
not(notn2222,n644);
and (s0n2222,notn2222,1'b0);
and (s1n2222,n644,n2223);
wire s0n2223,s1n2223,notn2223;
or (n2223,s0n2223,s1n2223);
not(notn2223,n568);
and (s0n2223,notn2223,n2224);
and (s1n2223,n568,n2226);
wire s0n2224,s1n2224,notn2224;
or (n2224,s0n2224,s1n2224);
not(notn2224,n15);
and (s0n2224,notn2224,1'b0);
and (s1n2224,n15,n2225);
or (n2226,1'b0,n2227,n2229,n2231,n2233);
and (n2227,n2228,n549);
and (n2229,n2230,n560);
and (n2231,n2232,n564);
and (n2233,n2225,n566);
wire s0n2234,s1n2234,notn2234;
or (n2234,s0n2234,s1n2234);
not(notn2234,n692);
and (s0n2234,notn2234,1'b0);
and (s1n2234,n692,n2207);
and (n2235,n2234,n2236);
or (n2236,n2237,n2251,n2253);
and (n2237,n2238,n2250);
wire s0n2238,s1n2238,notn2238;
or (n2238,s0n2238,s1n2238);
not(notn2238,n644);
and (s0n2238,notn2238,1'b0);
and (s1n2238,n644,n2239);
wire s0n2239,s1n2239,notn2239;
or (n2239,s0n2239,s1n2239);
not(notn2239,n568);
and (s0n2239,notn2239,n2240);
and (s1n2239,n568,n2242);
wire s0n2240,s1n2240,notn2240;
or (n2240,s0n2240,s1n2240);
not(notn2240,n15);
and (s0n2240,notn2240,1'b0);
and (s1n2240,n15,n2241);
or (n2242,1'b0,n2243,n2245,n2247,n2249);
and (n2243,n2244,n549);
and (n2245,n2246,n560);
and (n2247,n2248,n564);
and (n2249,n2241,n566);
wire s0n2250,s1n2250,notn2250;
or (n2250,s0n2250,s1n2250);
not(notn2250,n692);
and (s0n2250,notn2250,1'b0);
and (s1n2250,n692,n2223);
and (n2251,n2250,n2252);
or (n2252,n2253,n2267,n2268);
and (n2253,n2254,n2266);
wire s0n2254,s1n2254,notn2254;
or (n2254,s0n2254,s1n2254);
not(notn2254,n644);
and (s0n2254,notn2254,1'b0);
and (s1n2254,n644,n2255);
wire s0n2255,s1n2255,notn2255;
or (n2255,s0n2255,s1n2255);
not(notn2255,n568);
and (s0n2255,notn2255,n2256);
and (s1n2255,n568,n2258);
wire s0n2256,s1n2256,notn2256;
or (n2256,s0n2256,s1n2256);
not(notn2256,n15);
and (s0n2256,notn2256,1'b0);
and (s1n2256,n15,n2257);
or (n2258,1'b0,n2259,n2261,n2263,n2265);
and (n2259,n2260,n549);
and (n2261,n2262,n560);
and (n2263,n2264,n564);
and (n2265,n2257,n566);
wire s0n2266,s1n2266,notn2266;
or (n2266,s0n2266,s1n2266);
not(notn2266,n692);
and (s0n2266,notn2266,1'b0);
and (s1n2266,n692,n2239);
and (n2267,n2266,n2268);
and (n2268,n2269,n2281);
wire s0n2269,s1n2269,notn2269;
or (n2269,s0n2269,s1n2269);
not(notn2269,n644);
and (s0n2269,notn2269,1'b0);
and (s1n2269,n644,n2270);
wire s0n2270,s1n2270,notn2270;
or (n2270,s0n2270,s1n2270);
not(notn2270,n568);
and (s0n2270,notn2270,n2271);
and (s1n2270,n568,n2273);
wire s0n2271,s1n2271,notn2271;
or (n2271,s0n2271,s1n2271);
not(notn2271,n15);
and (s0n2271,notn2271,1'b0);
and (s1n2271,n15,n2272);
or (n2273,1'b0,n2274,n2276,n2278,n2280);
and (n2274,n2275,n549);
and (n2276,n2277,n560);
and (n2278,n2279,n564);
and (n2280,n2272,n566);
wire s0n2281,s1n2281,notn2281;
or (n2281,s0n2281,s1n2281);
not(notn2281,n692);
and (s0n2281,notn2281,1'b0);
and (s1n2281,n692,n2255);
and (n2282,n2222,n2236);
and (n2283,n2206,n2220);
and (n2284,n2190,n2204);
and (n2285,n2174,n2188);
and (n2286,n2170,n2287);
or (n2287,n2288,n2291,n2331);
and (n2288,n2289,n2290);
wire s0n2289,s1n2289,notn2289;
or (n2289,s0n2289,s1n2289);
not(notn2289,n587);
and (s0n2289,notn2289,1'b0);
and (s1n2289,n587,n2175);
xor (n2290,n2171,n2172);
and (n2291,n2290,n2292);
or (n2292,n2293,n2297,n2330);
and (n2293,n2294,n2295);
wire s0n2294,s1n2294,notn2294;
or (n2294,s0n2294,s1n2294);
not(notn2294,n587);
and (s0n2294,notn2294,1'b0);
and (s1n2294,n587,n2191);
xor (n2295,n2296,n2188);
xor (n2296,n2174,n2186);
and (n2297,n2295,n2298);
or (n2298,n2299,n2303,n2329);
and (n2299,n2300,n2301);
wire s0n2300,s1n2300,notn2300;
or (n2300,s0n2300,s1n2300);
not(notn2300,n587);
and (s0n2300,notn2300,1'b0);
and (s1n2300,n587,n2207);
xor (n2301,n2302,n2204);
xor (n2302,n2190,n2202);
and (n2303,n2301,n2304);
or (n2304,n2305,n2309,n2328);
and (n2305,n2306,n2307);
wire s0n2306,s1n2306,notn2306;
or (n2306,s0n2306,s1n2306);
not(notn2306,n587);
and (s0n2306,notn2306,1'b0);
and (s1n2306,n587,n2223);
xor (n2307,n2308,n2220);
xor (n2308,n2206,n2218);
and (n2309,n2307,n2310);
or (n2310,n2311,n2315,n2327);
and (n2311,n2312,n2313);
wire s0n2312,s1n2312,notn2312;
or (n2312,s0n2312,s1n2312);
not(notn2312,n587);
and (s0n2312,notn2312,1'b0);
and (s1n2312,n587,n2239);
xor (n2313,n2314,n2236);
xor (n2314,n2222,n2234);
and (n2315,n2313,n2316);
or (n2316,n2317,n2321,n2326);
and (n2317,n2318,n2319);
wire s0n2318,s1n2318,notn2318;
or (n2318,s0n2318,s1n2318);
not(notn2318,n587);
and (s0n2318,notn2318,1'b0);
and (s1n2318,n587,n2255);
xor (n2319,n2320,n2252);
xor (n2320,n2238,n2250);
and (n2321,n2319,n2322);
and (n2322,n2323,n2324);
wire s0n2323,s1n2323,notn2323;
or (n2323,s0n2323,s1n2323);
not(notn2323,n587);
and (s0n2323,notn2323,1'b0);
and (s1n2323,n587,n2270);
xor (n2324,n2325,n2268);
xor (n2325,n2254,n2266);
and (n2326,n2318,n2322);
and (n2327,n2312,n2316);
and (n2328,n2306,n2310);
and (n2329,n2300,n2304);
and (n2330,n2294,n2298);
and (n2331,n2289,n2292);
and (n2332,n2158,n2287);
and (n2333,n2334,n2335);
wire s0n2334,s1n2334,notn2334;
or (n2334,s0n2334,s1n2334);
not(notn2334,n979);
and (s0n2334,notn2334,1'b0);
and (s1n2334,n979,n2156);
or (n2335,n2336,n2341,n2406);
and (n2336,n2337,n2340);
wire s0n2337,s1n2337,notn2337;
or (n2337,s0n2337,s1n2337);
not(notn2337,n979);
and (s0n2337,notn2337,1'b0);
and (s1n2337,n979,n2338);
xor (n2338,n2339,n2287);
xor (n2339,n2158,n2170);
wire s0n2340,s1n2340,notn2340;
or (n2340,s0n2340,s1n2340);
not(notn2340,n1027);
and (s0n2340,notn2340,1'b0);
and (s1n2340,n1027,n2156);
and (n2341,n2340,n2342);
or (n2342,n2343,n2348,n2405);
and (n2343,n2344,n2347);
wire s0n2344,s1n2344,notn2344;
or (n2344,s0n2344,s1n2344);
not(notn2344,n979);
and (s0n2344,notn2344,1'b0);
and (s1n2344,n979,n2345);
xor (n2345,n2346,n2292);
xor (n2346,n2289,n2290);
wire s0n2347,s1n2347,notn2347;
or (n2347,s0n2347,s1n2347);
not(notn2347,n1027);
and (s0n2347,notn2347,1'b0);
and (s1n2347,n1027,n2338);
and (n2348,n2347,n2349);
or (n2349,n2350,n2355,n2404);
and (n2350,n2351,n2354);
wire s0n2351,s1n2351,notn2351;
or (n2351,s0n2351,s1n2351);
not(notn2351,n979);
and (s0n2351,notn2351,1'b0);
and (s1n2351,n979,n2352);
xor (n2352,n2353,n2298);
xor (n2353,n2294,n2295);
wire s0n2354,s1n2354,notn2354;
or (n2354,s0n2354,s1n2354);
not(notn2354,n1027);
and (s0n2354,notn2354,1'b0);
and (s1n2354,n1027,n2345);
and (n2355,n2354,n2356);
or (n2356,n2357,n2362,n2403);
and (n2357,n2358,n2361);
wire s0n2358,s1n2358,notn2358;
or (n2358,s0n2358,s1n2358);
not(notn2358,n979);
and (s0n2358,notn2358,1'b0);
and (s1n2358,n979,n2359);
xor (n2359,n2360,n2304);
xor (n2360,n2300,n2301);
wire s0n2361,s1n2361,notn2361;
or (n2361,s0n2361,s1n2361);
not(notn2361,n1027);
and (s0n2361,notn2361,1'b0);
and (s1n2361,n1027,n2352);
and (n2362,n2361,n2363);
or (n2363,n2364,n2369,n2402);
and (n2364,n2365,n2368);
wire s0n2365,s1n2365,notn2365;
or (n2365,s0n2365,s1n2365);
not(notn2365,n979);
and (s0n2365,notn2365,1'b0);
and (s1n2365,n979,n2366);
xor (n2366,n2367,n2310);
xor (n2367,n2306,n2307);
wire s0n2368,s1n2368,notn2368;
or (n2368,s0n2368,s1n2368);
not(notn2368,n1027);
and (s0n2368,notn2368,1'b0);
and (s1n2368,n1027,n2359);
and (n2369,n2368,n2370);
or (n2370,n2371,n2376,n2401);
and (n2371,n2372,n2375);
wire s0n2372,s1n2372,notn2372;
or (n2372,s0n2372,s1n2372);
not(notn2372,n979);
and (s0n2372,notn2372,1'b0);
and (s1n2372,n979,n2373);
xor (n2373,n2374,n2316);
xor (n2374,n2312,n2313);
wire s0n2375,s1n2375,notn2375;
or (n2375,s0n2375,s1n2375);
not(notn2375,n1027);
and (s0n2375,notn2375,1'b0);
and (s1n2375,n1027,n2366);
and (n2376,n2375,n2377);
or (n2377,n2378,n2383,n2400);
and (n2378,n2379,n2382);
wire s0n2379,s1n2379,notn2379;
or (n2379,s0n2379,s1n2379);
not(notn2379,n979);
and (s0n2379,notn2379,1'b0);
and (s1n2379,n979,n2380);
xor (n2380,n2381,n2322);
xor (n2381,n2318,n2319);
wire s0n2382,s1n2382,notn2382;
or (n2382,s0n2382,s1n2382);
not(notn2382,n1027);
and (s0n2382,notn2382,1'b0);
and (s1n2382,n1027,n2373);
and (n2383,n2382,n2384);
or (n2384,n2385,n2389,n2391);
and (n2385,n2386,n2388);
wire s0n2386,s1n2386,notn2386;
or (n2386,s0n2386,s1n2386);
not(notn2386,n979);
and (s0n2386,notn2386,1'b0);
and (s1n2386,n979,n2387);
xor (n2387,n2323,n2324);
wire s0n2388,s1n2388,notn2388;
or (n2388,s0n2388,s1n2388);
not(notn2388,n1027);
and (s0n2388,notn2388,1'b0);
and (s1n2388,n1027,n2380);
and (n2389,n2388,n2390);
or (n2390,n2391,n2395,n2396);
and (n2391,n2392,n2394);
wire s0n2392,s1n2392,notn2392;
or (n2392,s0n2392,s1n2392);
not(notn2392,n979);
and (s0n2392,notn2392,1'b0);
and (s1n2392,n979,n2393);
xor (n2393,n2269,n2281);
wire s0n2394,s1n2394,notn2394;
or (n2394,s0n2394,s1n2394);
not(notn2394,n1027);
and (s0n2394,notn2394,1'b0);
and (s1n2394,n1027,n2387);
and (n2395,n2394,n2396);
and (n2396,n2397,n2399);
wire s0n2397,s1n2397,notn2397;
or (n2397,s0n2397,s1n2397);
not(notn2397,n979);
and (s0n2397,notn2397,1'b0);
and (s1n2397,n979,n2398);
wire s0n2398,s1n2398,notn2398;
or (n2398,s0n2398,s1n2398);
not(notn2398,n692);
and (s0n2398,notn2398,1'b0);
and (s1n2398,n692,n2270);
wire s0n2399,s1n2399,notn2399;
or (n2399,s0n2399,s1n2399);
not(notn2399,n1027);
and (s0n2399,notn2399,1'b0);
and (s1n2399,n1027,n2393);
and (n2400,n2379,n2384);
and (n2401,n2372,n2377);
and (n2402,n2365,n2370);
and (n2403,n2358,n2363);
and (n2404,n2351,n2356);
and (n2405,n2344,n2349);
and (n2406,n2337,n2342);
and (n2407,n2333,n2408);
or (n2408,n2409,n2412,n2473);
and (n2409,n2410,n2411);
wire s0n2410,s1n2410,notn2410;
or (n2410,s0n2410,s1n2410);
not(notn2410,n930);
and (s0n2410,notn2410,1'b0);
and (s1n2410,n930,n2338);
xor (n2411,n2334,n2335);
and (n2412,n2411,n2413);
or (n2413,n2414,n2418,n2472);
and (n2414,n2415,n2416);
wire s0n2415,s1n2415,notn2415;
or (n2415,s0n2415,s1n2415);
not(notn2415,n930);
and (s0n2415,notn2415,1'b0);
and (s1n2415,n930,n2345);
xor (n2416,n2417,n2342);
xor (n2417,n2337,n2340);
and (n2418,n2416,n2419);
or (n2419,n2420,n2424,n2471);
and (n2420,n2421,n2422);
wire s0n2421,s1n2421,notn2421;
or (n2421,s0n2421,s1n2421);
not(notn2421,n930);
and (s0n2421,notn2421,1'b0);
and (s1n2421,n930,n2352);
xor (n2422,n2423,n2349);
xor (n2423,n2344,n2347);
and (n2424,n2422,n2425);
or (n2425,n2426,n2430,n2470);
and (n2426,n2427,n2428);
wire s0n2427,s1n2427,notn2427;
or (n2427,s0n2427,s1n2427);
not(notn2427,n930);
and (s0n2427,notn2427,1'b0);
and (s1n2427,n930,n2359);
xor (n2428,n2429,n2356);
xor (n2429,n2351,n2354);
and (n2430,n2428,n2431);
or (n2431,n2432,n2436,n2469);
and (n2432,n2433,n2434);
wire s0n2433,s1n2433,notn2433;
or (n2433,s0n2433,s1n2433);
not(notn2433,n930);
and (s0n2433,notn2433,1'b0);
and (s1n2433,n930,n2366);
xor (n2434,n2435,n2363);
xor (n2435,n2358,n2361);
and (n2436,n2434,n2437);
or (n2437,n2438,n2442,n2468);
and (n2438,n2439,n2440);
wire s0n2439,s1n2439,notn2439;
or (n2439,s0n2439,s1n2439);
not(notn2439,n930);
and (s0n2439,notn2439,1'b0);
and (s1n2439,n930,n2373);
xor (n2440,n2441,n2370);
xor (n2441,n2365,n2368);
and (n2442,n2440,n2443);
or (n2443,n2444,n2448,n2467);
and (n2444,n2445,n2446);
wire s0n2445,s1n2445,notn2445;
or (n2445,s0n2445,s1n2445);
not(notn2445,n930);
and (s0n2445,notn2445,1'b0);
and (s1n2445,n930,n2380);
xor (n2446,n2447,n2377);
xor (n2447,n2372,n2375);
and (n2448,n2446,n2449);
or (n2449,n2450,n2454,n2466);
and (n2450,n2451,n2452);
wire s0n2451,s1n2451,notn2451;
or (n2451,s0n2451,s1n2451);
not(notn2451,n930);
and (s0n2451,notn2451,1'b0);
and (s1n2451,n930,n2387);
xor (n2452,n2453,n2384);
xor (n2453,n2379,n2382);
and (n2454,n2452,n2455);
or (n2455,n2456,n2460,n2465);
and (n2456,n2457,n2458);
wire s0n2457,s1n2457,notn2457;
or (n2457,s0n2457,s1n2457);
not(notn2457,n930);
and (s0n2457,notn2457,1'b0);
and (s1n2457,n930,n2393);
xor (n2458,n2459,n2390);
xor (n2459,n2386,n2388);
and (n2460,n2458,n2461);
and (n2461,n2462,n2463);
wire s0n2462,s1n2462,notn2462;
or (n2462,s0n2462,s1n2462);
not(notn2462,n930);
and (s0n2462,notn2462,1'b0);
and (s1n2462,n930,n2398);
xor (n2463,n2464,n2396);
xor (n2464,n2392,n2394);
and (n2465,n2457,n2461);
and (n2466,n2451,n2455);
and (n2467,n2445,n2449);
and (n2468,n2439,n2443);
and (n2469,n2433,n2437);
and (n2470,n2427,n2431);
and (n2471,n2421,n2425);
and (n2472,n2415,n2419);
and (n2473,n2410,n2413);
and (n2474,n2155,n2408);
or (n2475,n2476,n2481,n2569);
and (n2476,n2477,n2479);
xor (n2477,n2478,n2086);
xor (n2478,n1818,n2018);
xor (n2479,n2480,n2408);
xor (n2480,n2155,n2333);
and (n2481,n2479,n2482);
or (n2482,n2483,n2488,n2568);
and (n2483,n2484,n2486);
xor (n2484,n2485,n2091);
xor (n2485,n2088,n2089);
xor (n2486,n2487,n2413);
xor (n2487,n2410,n2411);
and (n2488,n2486,n2489);
or (n2489,n2490,n2495,n2567);
and (n2490,n2491,n2493);
xor (n2491,n2492,n2097);
xor (n2492,n2093,n2094);
xor (n2493,n2494,n2419);
xor (n2494,n2415,n2416);
and (n2495,n2493,n2496);
or (n2496,n2497,n2502,n2566);
and (n2497,n2498,n2500);
xor (n2498,n2499,n2103);
xor (n2499,n2099,n2100);
xor (n2500,n2501,n2425);
xor (n2501,n2421,n2422);
and (n2502,n2500,n2503);
or (n2503,n2504,n2509,n2565);
and (n2504,n2505,n2507);
xor (n2505,n2506,n2109);
xor (n2506,n2105,n2106);
xor (n2507,n2508,n2431);
xor (n2508,n2427,n2428);
and (n2509,n2507,n2510);
or (n2510,n2511,n2516,n2564);
and (n2511,n2512,n2514);
xor (n2512,n2513,n2115);
xor (n2513,n2111,n2112);
xor (n2514,n2515,n2437);
xor (n2515,n2433,n2434);
and (n2516,n2514,n2517);
or (n2517,n2518,n2523,n2563);
and (n2518,n2519,n2521);
xor (n2519,n2520,n2121);
xor (n2520,n2117,n2118);
xor (n2521,n2522,n2443);
xor (n2522,n2439,n2440);
and (n2523,n2521,n2524);
or (n2524,n2525,n2530,n2562);
and (n2525,n2526,n2528);
xor (n2526,n2527,n2127);
xor (n2527,n2123,n2124);
xor (n2528,n2529,n2449);
xor (n2529,n2445,n2446);
and (n2530,n2528,n2531);
or (n2531,n2532,n2537,n2561);
and (n2532,n2533,n2535);
xor (n2533,n2534,n2133);
xor (n2534,n2129,n2130);
xor (n2535,n2536,n2455);
xor (n2536,n2451,n2452);
and (n2537,n2535,n2538);
or (n2538,n2539,n2544,n2560);
and (n2539,n2540,n2542);
xor (n2540,n2541,n2139);
xor (n2541,n2135,n2136);
xor (n2542,n2543,n2461);
xor (n2543,n2457,n2458);
and (n2544,n2542,n2545);
or (n2545,n2546,n2549,n2559);
and (n2546,n2547,n2548);
xor (n2547,n2140,n2141);
xor (n2548,n2462,n2463);
and (n2549,n2548,n2550);
or (n2550,n2551,n2554,n2558);
and (n2551,n2552,n2553);
xor (n2552,n2075,n2077);
xor (n2553,n2397,n2399);
and (n2554,n2553,n2555);
and (n2555,n2556,n2557);
wire s0n2556,s1n2556,notn2556;
or (n2556,s0n2556,s1n2556);
not(notn2556,n1027);
and (s0n2556,notn2556,1'b0);
and (s1n2556,n1027,n2076);
wire s0n2557,s1n2557,notn2557;
or (n2557,s0n2557,s1n2557);
not(notn2557,n1027);
and (s0n2557,notn2557,1'b0);
and (s1n2557,n1027,n2398);
and (n2558,n2552,n2555);
and (n2559,n2547,n2550);
and (n2560,n2540,n2545);
and (n2561,n2533,n2538);
and (n2562,n2526,n2531);
and (n2563,n2519,n2524);
and (n2564,n2512,n2517);
and (n2565,n2505,n2510);
and (n2566,n2498,n2503);
and (n2567,n2491,n2496);
and (n2568,n2484,n2489);
and (n2569,n2477,n2482);
or (n2570,n2571,n2576,n2668);
and (n2571,n2572,n2574);
xor (n2572,n2573,n1726);
xor (n2573,n1721,n1723);
xor (n2574,n2575,n2482);
xor (n2575,n2477,n2479);
and (n2576,n2574,n2577);
or (n2577,n2578,n2583,n2667);
and (n2578,n2579,n2581);
xor (n2579,n2580,n1733);
xor (n2580,n1728,n1730);
xor (n2581,n2582,n2489);
xor (n2582,n2484,n2486);
and (n2583,n2581,n2584);
or (n2584,n2585,n2590,n2666);
and (n2585,n2586,n2588);
xor (n2586,n2587,n1740);
xor (n2587,n1735,n1737);
xor (n2588,n2589,n2496);
xor (n2589,n2491,n2493);
and (n2590,n2588,n2591);
or (n2591,n2592,n2597,n2665);
and (n2592,n2593,n2595);
xor (n2593,n2594,n1747);
xor (n2594,n1742,n1744);
xor (n2595,n2596,n2503);
xor (n2596,n2498,n2500);
and (n2597,n2595,n2598);
or (n2598,n2599,n2604,n2664);
and (n2599,n2600,n2602);
xor (n2600,n2601,n1754);
xor (n2601,n1749,n1751);
xor (n2602,n2603,n2510);
xor (n2603,n2505,n2507);
and (n2604,n2602,n2605);
or (n2605,n2606,n2611,n2663);
and (n2606,n2607,n2609);
xor (n2607,n2608,n1761);
xor (n2608,n1756,n1758);
xor (n2609,n2610,n2517);
xor (n2610,n2512,n2514);
and (n2611,n2609,n2612);
or (n2612,n2613,n2618,n2662);
and (n2613,n2614,n2616);
xor (n2614,n2615,n1768);
xor (n2615,n1763,n1765);
xor (n2616,n2617,n2524);
xor (n2617,n2519,n2521);
and (n2618,n2616,n2619);
or (n2619,n2620,n2625,n2661);
and (n2620,n2621,n2623);
xor (n2621,n2622,n1775);
xor (n2622,n1770,n1772);
xor (n2623,n2624,n2531);
xor (n2624,n2526,n2528);
and (n2625,n2623,n2626);
or (n2626,n2627,n2632,n2660);
and (n2627,n2628,n2630);
xor (n2628,n2629,n1782);
xor (n2629,n1777,n1779);
xor (n2630,n2631,n2538);
xor (n2631,n2533,n2535);
and (n2632,n2630,n2633);
or (n2633,n2634,n2639,n2659);
and (n2634,n2635,n2637);
xor (n2635,n2636,n1789);
xor (n2636,n1784,n1786);
xor (n2637,n2638,n2545);
xor (n2638,n2540,n2542);
and (n2639,n2637,n2640);
or (n2640,n2641,n2646,n2658);
and (n2641,n2642,n2644);
xor (n2642,n2643,n1794);
xor (n2643,n1791,n1792);
xor (n2644,n2645,n2550);
xor (n2645,n2547,n2548);
and (n2646,n2644,n2647);
or (n2647,n2648,n2653,n2657);
and (n2648,n2649,n2651);
xor (n2649,n2650,n1799);
xor (n2650,n1796,n1797);
xor (n2651,n2652,n2555);
xor (n2652,n2552,n2553);
and (n2653,n2651,n2654);
and (n2654,n2655,n2656);
xor (n2655,n1800,n1801);
xor (n2656,n2556,n2557);
and (n2657,n2649,n2654);
and (n2658,n2642,n2647);
and (n2659,n2635,n2640);
and (n2660,n2628,n2633);
and (n2661,n2621,n2626);
and (n2662,n2614,n2619);
and (n2663,n2607,n2612);
and (n2664,n2600,n2605);
and (n2665,n2593,n2598);
and (n2666,n2586,n2591);
and (n2667,n2579,n2584);
and (n2668,n2572,n2577);
and (n2669,n2670,n2672);
xor (n2670,n2671,n2577);
xor (n2671,n2572,n2574);
and (n2672,n2673,n2675);
xor (n2673,n2674,n2584);
xor (n2674,n2579,n2581);
and (n2675,n2676,n2678);
xor (n2676,n2677,n2591);
xor (n2677,n2586,n2588);
and (n2678,n2679,n2681);
xor (n2679,n2680,n2598);
xor (n2680,n2593,n2595);
and (n2681,n2682,n2684);
xor (n2682,n2683,n2605);
xor (n2683,n2600,n2602);
and (n2684,n2685,n2687);
xor (n2685,n2686,n2612);
xor (n2686,n2607,n2609);
and (n2687,n2688,n2690);
xor (n2688,n2689,n2619);
xor (n2689,n2614,n2616);
xor (n2690,n2691,n2626);
xor (n2691,n2621,n2623);
wire s0n2692,s1n2692,notn2692;
or (n2692,s0n2692,s1n2692);
not(notn2692,n2747);
and (s0n2692,notn2692,n2693);
and (s1n2692,n2747,n2699);
wire s0n2693,s1n2693,notn2693;
or (n2693,s0n2693,s1n2693);
not(notn2693,n2697);
and (s0n2693,notn2693,1'b0);
and (s1n2693,n2697,n2694);
wire s0n2694,s1n2694,notn2694;
or (n2694,s0n2694,s1n2694);
not(notn2694,n570);
and (s0n2694,notn2694,n555);
and (s1n2694,n570,n2695);
wire s0n2695,s1n2695,notn2695;
or (n2695,s0n2695,s1n2695);
not(notn2695,n2696);
and (s0n2695,notn2695,1'b0);
and (s1n2695,n2696,n14);
or (n2696,n551,n552,n553,n554);
and (n2697,n2698,n928);
and (n2698,n33,n585);
or (n2699,1'b0,n2700,n2712,n2724,n2736);
and (n2700,n2701,n2710);
or (n2701,1'b0,n2702,n2704,n2706,n2708);
and (n2702,n2703,n549);
and (n2704,n2705,n560);
and (n2706,n2707,n564);
and (n2708,n2709,n566);
and (n2710,n583,n2711);
and (n2711,n569,n20);
and (n2712,n2713,n2722);
or (n2713,1'b0,n2714,n2716,n2718,n2720);
and (n2714,n2715,n549);
and (n2716,n2717,n560);
and (n2718,n2719,n564);
and (n2720,n2721,n566);
and (n2722,n583,n2723);
and (n2723,n569,n25);
and (n2724,n2725,n2734);
or (n2725,1'b0,n2726,n2728,n2730,n2732);
and (n2726,n2727,n549);
and (n2728,n2729,n560);
and (n2730,n2731,n564);
and (n2732,n2733,n566);
and (n2734,n583,n2735);
and (n2735,n569,n29);
and (n2736,n2737,n2744);
or (n2737,1'b0,n2738,n2740,n2742,n2743);
and (n2738,n2739,n549);
and (n2740,n2741,n560);
and (n2742,n2164,n564);
and (n2743,n1827,n566);
and (n2744,n583,n2745);
or (n2745,n570,n2746);
and (n2746,n569,n32);
and (n2747,n583,n2748);
nor (n2748,n2749,n2792,n2818,n2844);
wire s0n2749,s1n2749,notn2749;
or (n2749,s0n2749,s1n2749);
not(notn2749,n583);
and (s0n2749,notn2749,1'b0);
and (s1n2749,n583,n2750);
wire s0n2750,s1n2750,notn2750;
or (n2750,s0n2750,s1n2750);
not(notn2750,n583);
and (s0n2750,notn2750,n1027);
and (s1n2750,n583,n2751);
wire s0n2751,s1n2751,notn2751;
or (n2751,s0n2751,s1n2751);
not(notn2751,n641);
and (s0n2751,notn2751,n2752);
and (s1n2751,n641,n1065);
wire s0n2752,s1n2752,notn2752;
or (n2752,s0n2752,s1n2752);
not(notn2752,n570);
and (s0n2752,notn2752,n2753);
and (s1n2752,n570,n2758);
or (n2753,n2754,n2755,n2756,n2757);
and (n2754,n1032,n573);
and (n2755,n1043,n577);
and (n2756,n1054,n580);
and (n2757,n1065,n582);
or (n2758,1'b0,n2759,n2761,n2763,n2766,n2768,n2770,n2772,n2774,n2776,n2778,n2780,n2782,n2784,n2786,n2788,n2790);
and (n2759,n1035,n2760);
and (n2760,n21,n22,n574,n575,n584);
and (n2761,n1037,n2762);
and (n2762,n26,n22,n574,n575,n584);
and (n2763,n1039,n2764);
and (n2764,n21,n2765,n574,n575,n584);
not (n2765,n22);
and (n2766,n1032,n2767);
and (n2767,n26,n2765,n574,n575,n584);
and (n2768,n1046,n2769);
and (n2769,n21,n22,n578,n575,n584);
and (n2770,n1048,n2771);
and (n2771,n26,n22,n578,n575,n584);
and (n2772,n1050,n2773);
and (n2773,n21,n2765,n578,n575,n584);
and (n2774,n1043,n2775);
and (n2775,n26,n2765,n578,n575,n584);
and (n2776,n1057,n2777);
nor (n2777,n26,n2765,n578,n575,n548);
and (n2778,n1059,n2779);
nor (n2779,n21,n2765,n578,n575,n548);
and (n2780,n1061,n2781);
nor (n2781,n26,n22,n578,n575,n548);
and (n2782,n1054,n2783);
nor (n2783,n21,n22,n578,n575,n548);
and (n2784,n1068,n2785);
nor (n2785,n26,n2765,n574,n575,n548);
and (n2786,n1070,n2787);
nor (n2787,n21,n2765,n574,n575,n548);
and (n2788,n1072,n2789);
nor (n2789,n26,n22,n574,n575,n548);
and (n2790,n1065,n2791);
nor (n2791,n21,n22,n574,n575,n548);
wire s0n2792,s1n2792,notn2792;
or (n2792,s0n2792,s1n2792);
not(notn2792,n583);
and (s0n2792,notn2792,1'b0);
and (s1n2792,n583,n2793);
wire s0n2793,s1n2793,notn2793;
or (n2793,s0n2793,s1n2793);
not(notn2793,n583);
and (s0n2793,notn2793,n979);
and (s1n2793,n583,n2794);
wire s0n2794,s1n2794,notn2794;
or (n2794,s0n2794,s1n2794);
not(notn2794,n641);
and (s0n2794,notn2794,n2795);
and (s1n2794,n641,n1017);
wire s0n2795,s1n2795,notn2795;
or (n2795,s0n2795,s1n2795);
not(notn2795,n570);
and (s0n2795,notn2795,n2796);
and (s1n2795,n570,n2801);
or (n2796,n2797,n2798,n2799,n2800);
and (n2797,n984,n573);
and (n2798,n995,n577);
and (n2799,n1006,n580);
and (n2800,n1017,n582);
or (n2801,1'b0,n2802,n2803,n2804,n2805,n2806,n2807,n2808,n2809,n2810,n2811,n2812,n2813,n2814,n2815,n2816,n2817);
and (n2802,n987,n2760);
and (n2803,n989,n2762);
and (n2804,n991,n2764);
and (n2805,n984,n2767);
and (n2806,n998,n2769);
and (n2807,n1000,n2771);
and (n2808,n1002,n2773);
and (n2809,n995,n2775);
and (n2810,n1009,n2777);
and (n2811,n1011,n2779);
and (n2812,n1013,n2781);
and (n2813,n1006,n2783);
and (n2814,n1020,n2785);
and (n2815,n1022,n2787);
and (n2816,n1024,n2789);
and (n2817,n1017,n2791);
wire s0n2818,s1n2818,notn2818;
or (n2818,s0n2818,s1n2818);
not(notn2818,n583);
and (s0n2818,notn2818,1'b0);
and (s1n2818,n583,n2819);
wire s0n2819,s1n2819,notn2819;
or (n2819,s0n2819,s1n2819);
not(notn2819,n583);
and (s0n2819,notn2819,n692);
and (s1n2819,n583,n2820);
wire s0n2820,s1n2820,notn2820;
or (n2820,s0n2820,s1n2820);
not(notn2820,n641);
and (s0n2820,notn2820,n2821);
and (s1n2820,n641,n730);
wire s0n2821,s1n2821,notn2821;
or (n2821,s0n2821,s1n2821);
not(notn2821,n570);
and (s0n2821,notn2821,n2822);
and (s1n2821,n570,n2827);
or (n2822,n2823,n2824,n2825,n2826);
and (n2823,n697,n573);
and (n2824,n708,n577);
and (n2825,n719,n580);
and (n2826,n730,n582);
or (n2827,1'b0,n2828,n2829,n2830,n2831,n2832,n2833,n2834,n2835,n2836,n2837,n2838,n2839,n2840,n2841,n2842,n2843);
and (n2828,n700,n2760);
and (n2829,n702,n2762);
and (n2830,n704,n2764);
and (n2831,n697,n2767);
and (n2832,n711,n2769);
and (n2833,n713,n2771);
and (n2834,n715,n2773);
and (n2835,n708,n2775);
and (n2836,n722,n2777);
and (n2837,n724,n2779);
and (n2838,n726,n2781);
and (n2839,n719,n2783);
and (n2840,n733,n2785);
and (n2841,n735,n2787);
and (n2842,n737,n2789);
and (n2843,n730,n2791);
wire s0n2844,s1n2844,notn2844;
or (n2844,s0n2844,s1n2844);
not(notn2844,n583);
and (s0n2844,notn2844,1'b0);
and (s1n2844,n583,n2845);
wire s0n2845,s1n2845,notn2845;
or (n2845,s0n2845,s1n2845);
not(notn2845,n583);
and (s0n2845,notn2845,n644);
and (s1n2845,n583,n2846);
wire s0n2846,s1n2846,notn2846;
or (n2846,s0n2846,s1n2846);
not(notn2846,n641);
and (s0n2846,notn2846,n2847);
and (s1n2846,n641,n682);
wire s0n2847,s1n2847,notn2847;
or (n2847,s0n2847,s1n2847);
not(notn2847,n570);
and (s0n2847,notn2847,n2848);
and (s1n2847,n570,n2853);
or (n2848,n2849,n2850,n2851,n2852);
and (n2849,n649,n573);
and (n2850,n660,n577);
and (n2851,n671,n580);
and (n2852,n682,n582);
or (n2853,1'b0,n2854,n2855,n2856,n2857,n2858,n2859,n2860,n2861,n2862,n2863,n2864,n2865,n2866,n2867,n2868,n2869);
and (n2854,n652,n2760);
and (n2855,n654,n2762);
and (n2856,n656,n2764);
and (n2857,n649,n2767);
and (n2858,n663,n2769);
and (n2859,n665,n2771);
and (n2860,n667,n2773);
and (n2861,n660,n2775);
and (n2862,n674,n2777);
and (n2863,n676,n2779);
and (n2864,n678,n2781);
and (n2865,n671,n2783);
and (n2866,n685,n2785);
and (n2867,n687,n2787);
and (n2868,n689,n2789);
and (n2869,n682,n2791);
or (n2870,n2871,n2874,n2692);
and (n2871,n2872,n8859);
wire s0n2872,s1n2872,notn2872;
or (n2872,s0n2872,s1n2872);
not(notn2872,n5024);
and (s0n2872,notn2872,1'b0);
and (s1n2872,n5024,n2873);
or (n2873,1'b0,n2874,n8846,n8856,n8857,n8858);
and (n2874,n2875,n2899);
wire s0n2875,s1n2875,notn2875;
or (n2875,s0n2875,s1n2875);
not(notn2875,n2894);
and (s0n2875,notn2875,1'b0);
and (s1n2875,n2894,n2876);
xor (n2876,n2877,n8824);
or (n2877,n2878,n8050,n8823);
and (n2878,n2879,n5005);
or (n2879,1'b0,n2880,n2891,n2902,n4941);
and (n2880,n2881,n2885);
wire s0n2881,s1n2881,notn2881;
or (n2881,s0n2881,s1n2881);
not(notn2881,n2883);
and (s0n2881,notn2881,1'b0);
and (s1n2881,n2883,n2882);
and (n2883,n2884,n2696);
nand (n2884,n551,n561,n553,n567);
or (n2885,n2886,n2889);
nor (n2886,n2887,n2792,n2818,n2888);
not (n2887,n2749);
not (n2888,n2844);
and (n2889,n2749,n2792,n2890,n2844);
not (n2890,n2818);
and (n2891,n2892,n2899);
wire s0n2892,s1n2892,notn2892;
or (n2892,s0n2892,s1n2892);
not(notn2892,n2894);
and (s0n2892,notn2892,1'b0);
and (s1n2892,n2894,n2893);
or (n2894,n2895,n549);
or (n2895,n2896,n564);
or (n2896,n2897,n2898);
and (n2897,n551,n552,n553,n567);
not (n2898,n2884);
or (n2899,n2900,n2901);
and (n2900,n2887,n2792,n2818,n2888);
and (n2901,n2887,n2792,n2818,n2844);
and (n2902,n2903,n4938);
wire s0n2903,s1n2903,notn2903;
or (n2903,s0n2903,s1n2903);
not(notn2903,n4933);
and (s0n2903,notn2903,n2904);
and (s1n2903,n4933,1'b0);
wire s0n2904,s1n2904,notn2904;
or (n2904,s0n2904,s1n2904);
not(notn2904,n4928);
and (s0n2904,notn2904,n2905);
and (s1n2904,n4928,1'b1);
wire s0n2905,s1n2905,notn2905;
or (n2905,s0n2905,s1n2905);
not(notn2905,n4916);
and (s0n2905,notn2905,1'b0);
and (s1n2905,n4916,n2906);
xor (n2906,n2907,n4893);
xor (n2907,n2908,n4840);
xor (n2908,n2909,n4402);
xor (n2909,n2910,n4400);
xor (n2910,n2911,n4370);
not (n2911,n2912);
or (n2912,n2913,n3784);
or (n2913,n2914,n3043,n3783);
and (n2914,n2915,n3012);
or (n2915,1'b0,n2916,n2970,n2984,n2998);
and (n2916,n2917,n2710);
or (n2917,1'b0,n2918,n2944,n2952,n2961);
and (n2918,n2919,n2924);
wire s0n2919,s1n2919,notn2919;
or (n2919,s0n2919,s1n2919);
not(notn2919,n2921);
and (s0n2919,notn2919,n2703);
and (s1n2919,n2921,n2920);
or (n2921,n2922,n2923);
and (n2922,n2749,n2792,n2818,n2888);
and (n2923,n2749,n2792,n2818,n2844);
or (n2924,n2925,n2943);
or (n2925,n2926,n2939);
and (n2926,n2927,n549);
or (n2927,n2928,n2923);
or (n2928,n2929,n2922);
or (n2929,n2930,n2938);
or (n2930,n2931,n2937);
or (n2931,n2932,n2936);
or (n2932,n2933,n2934);
nor (n2933,n2749,n2792,n2818,n2888);
and (n2934,n2887,n2935,n2818,n2888);
not (n2935,n2792);
and (n2936,n2887,n2935,n2818,n2844);
and (n2937,n2749,n2935,n2818,n2888);
and (n2938,n2749,n2935,n2818,n2844);
and (n2939,n2940,n560);
or (n2940,n2941,n2889);
or (n2941,n2942,n2886);
nor (n2942,n2749,n2935,n2818,n2888);
and (n2943,n2899,n560);
and (n2944,n2945,n2947);
wire s0n2945,s1n2945,notn2945;
or (n2945,s0n2945,s1n2945);
not(notn2945,n2921);
and (s0n2945,notn2945,n2705);
and (s1n2945,n2921,n2946);
or (n2947,n2948,n2951);
or (n2948,n2949,n2950);
and (n2949,n2927,n560);
and (n2950,n2940,n564);
and (n2951,n2899,n566);
and (n2952,n2953,n2955);
wire s0n2953,s1n2953,notn2953;
or (n2953,s0n2953,s1n2953);
not(notn2953,n2921);
and (s0n2953,notn2953,n2707);
and (s1n2953,n2921,n2954);
or (n2955,n2956,n2959);
or (n2956,n2957,n2958);
and (n2957,n2927,n564);
and (n2958,n2940,n566);
and (n2959,n2899,n2960);
and (n2960,n550,n552,n553,n567);
and (n2961,n2962,n2964);
wire s0n2962,s1n2962,notn2962;
or (n2962,s0n2962,s1n2962);
not(notn2962,n2921);
and (s0n2962,notn2962,n2709);
and (s1n2962,n2921,n2963);
or (n2964,n2965,n2968);
or (n2965,n2966,n2967);
and (n2966,n2927,n566);
and (n2967,n2940,n2898);
and (n2968,n2899,n2969);
nor (n2969,n551,n552,n553,n567);
and (n2970,n2971,n2722);
or (n2971,1'b0,n2972,n2975,n2978,n2981);
and (n2972,n2973,n2924);
wire s0n2973,s1n2973,notn2973;
or (n2973,s0n2973,s1n2973);
not(notn2973,n2921);
and (s0n2973,notn2973,n2715);
and (s1n2973,n2921,n2974);
and (n2975,n2976,n2947);
wire s0n2976,s1n2976,notn2976;
or (n2976,s0n2976,s1n2976);
not(notn2976,n2921);
and (s0n2976,notn2976,n2717);
and (s1n2976,n2921,n2977);
and (n2978,n2979,n2955);
wire s0n2979,s1n2979,notn2979;
or (n2979,s0n2979,s1n2979);
not(notn2979,n2921);
and (s0n2979,notn2979,n2719);
and (s1n2979,n2921,n2980);
and (n2981,n2982,n2964);
wire s0n2982,s1n2982,notn2982;
or (n2982,s0n2982,s1n2982);
not(notn2982,n2921);
and (s0n2982,notn2982,n2721);
and (s1n2982,n2921,n2983);
and (n2984,n2985,n2734);
or (n2985,1'b0,n2986,n2989,n2992,n2995);
and (n2986,n2987,n2924);
wire s0n2987,s1n2987,notn2987;
or (n2987,s0n2987,s1n2987);
not(notn2987,n2921);
and (s0n2987,notn2987,n2727);
and (s1n2987,n2921,n2988);
and (n2989,n2990,n2947);
wire s0n2990,s1n2990,notn2990;
or (n2990,s0n2990,s1n2990);
not(notn2990,n2921);
and (s0n2990,notn2990,n2729);
and (s1n2990,n2921,n2991);
and (n2992,n2993,n2955);
wire s0n2993,s1n2993,notn2993;
or (n2993,s0n2993,s1n2993);
not(notn2993,n2921);
and (s0n2993,notn2993,n2731);
and (s1n2993,n2921,n2994);
and (n2995,n2996,n2964);
wire s0n2996,s1n2996,notn2996;
or (n2996,s0n2996,s1n2996);
not(notn2996,n2921);
and (s0n2996,notn2996,n2733);
and (s1n2996,n2921,n2997);
and (n2998,n2999,n2744);
or (n2999,1'b0,n3000,n3003,n3006,n3009);
and (n3000,n3001,n2924);
wire s0n3001,s1n3001,notn3001;
or (n3001,s0n3001,s1n3001);
not(notn3001,n2921);
and (s0n3001,notn3001,n2739);
and (s1n3001,n2921,n3002);
and (n3003,n3004,n2947);
wire s0n3004,s1n3004,notn3004;
or (n3004,s0n3004,s1n3004);
not(notn3004,n2921);
and (s0n3004,notn3004,n2741);
and (s1n3004,n2921,n3005);
and (n3006,n3007,n2955);
wire s0n3007,s1n3007,notn3007;
or (n3007,s0n3007,s1n3007);
not(notn3007,n2921);
and (s0n3007,notn3007,n2164);
and (s1n3007,n2921,n3008);
and (n3009,n3010,n2964);
wire s0n3010,s1n3010,notn3010;
or (n3010,s0n3010,s1n3010);
not(notn3010,n2921);
and (s0n3010,notn3010,n1827);
and (s1n3010,n2921,n3011);
or (n3012,1'b0,n3013,n3022,n3028,n3037);
and (n3013,n3014,n2710);
or (n3014,1'b0,n3015,n3019,n3020,n3021);
and (n3015,n3016,n2924);
wire s0n3016,s1n3016,notn3016;
or (n3016,s0n3016,s1n3016);
not(notn3016,n2921);
and (s0n3016,notn3016,n3017);
and (s1n3016,n2921,n3018);
and (n3019,n2919,n2947);
and (n3020,n2945,n2955);
and (n3021,n2953,n2964);
and (n3022,n3023,n2722);
or (n3023,1'b0,n3024,n3025,n3026,n3027);
and (n3024,n2962,n2924);
and (n3025,n2973,n2947);
and (n3026,n2976,n2955);
and (n3027,n2979,n2964);
and (n3028,n3029,n2734);
or (n3029,1'b0,n3030,n3034,n3035,n3036);
and (n3030,n3031,n2924);
wire s0n3031,s1n3031,notn3031;
or (n3031,s0n3031,s1n3031);
not(notn3031,n2921);
and (s0n3031,notn3031,n3032);
and (s1n3031,n2921,n3033);
and (n3034,n2987,n2947);
and (n3035,n2990,n2955);
and (n3036,n2993,n2964);
and (n3037,n3038,n2744);
or (n3038,1'b0,n3039,n3040,n3041,n3042);
and (n3039,n2996,n2924);
and (n3040,n3001,n2947);
and (n3041,n3004,n2955);
and (n3042,n3007,n2964);
and (n3043,n3012,n3044);
or (n3044,n3045,n3148,n3782);
and (n3045,n3046,n3117);
or (n3046,1'b0,n3047,n3065,n3083,n3101);
and (n3047,n3048,n2710);
or (n3048,1'b0,n3049,n3053,n3057,n3061);
and (n3049,n3050,n2924);
wire s0n3050,s1n3050,notn3050;
or (n3050,s0n3050,s1n3050);
not(notn3050,n2921);
and (s0n3050,notn3050,n3051);
and (s1n3050,n2921,n3052);
and (n3053,n3054,n2947);
wire s0n3054,s1n3054,notn3054;
or (n3054,s0n3054,s1n3054);
not(notn3054,n2921);
and (s0n3054,notn3054,n3055);
and (s1n3054,n2921,n3056);
and (n3057,n3058,n2955);
wire s0n3058,s1n3058,notn3058;
or (n3058,s0n3058,s1n3058);
not(notn3058,n2921);
and (s0n3058,notn3058,n3059);
and (s1n3058,n2921,n3060);
and (n3061,n3062,n2964);
wire s0n3062,s1n3062,notn3062;
or (n3062,s0n3062,s1n3062);
not(notn3062,n2921);
and (s0n3062,notn3062,n3063);
and (s1n3062,n2921,n3064);
and (n3065,n3066,n2722);
or (n3066,1'b0,n3067,n3071,n3075,n3079);
and (n3067,n3068,n2924);
wire s0n3068,s1n3068,notn3068;
or (n3068,s0n3068,s1n3068);
not(notn3068,n2921);
and (s0n3068,notn3068,n3069);
and (s1n3068,n2921,n3070);
and (n3071,n3072,n2947);
wire s0n3072,s1n3072,notn3072;
or (n3072,s0n3072,s1n3072);
not(notn3072,n2921);
and (s0n3072,notn3072,n3073);
and (s1n3072,n2921,n3074);
and (n3075,n3076,n2955);
wire s0n3076,s1n3076,notn3076;
or (n3076,s0n3076,s1n3076);
not(notn3076,n2921);
and (s0n3076,notn3076,n3077);
and (s1n3076,n2921,n3078);
and (n3079,n3080,n2964);
wire s0n3080,s1n3080,notn3080;
or (n3080,s0n3080,s1n3080);
not(notn3080,n2921);
and (s0n3080,notn3080,n3081);
and (s1n3080,n2921,n3082);
and (n3083,n3084,n2734);
or (n3084,1'b0,n3085,n3089,n3093,n3097);
and (n3085,n3086,n2924);
wire s0n3086,s1n3086,notn3086;
or (n3086,s0n3086,s1n3086);
not(notn3086,n2921);
and (s0n3086,notn3086,n3087);
and (s1n3086,n2921,n3088);
and (n3089,n3090,n2947);
wire s0n3090,s1n3090,notn3090;
or (n3090,s0n3090,s1n3090);
not(notn3090,n2921);
and (s0n3090,notn3090,n3091);
and (s1n3090,n2921,n3092);
and (n3093,n3094,n2955);
wire s0n3094,s1n3094,notn3094;
or (n3094,s0n3094,s1n3094);
not(notn3094,n2921);
and (s0n3094,notn3094,n3095);
and (s1n3094,n2921,n3096);
and (n3097,n3098,n2964);
wire s0n3098,s1n3098,notn3098;
or (n3098,s0n3098,s1n3098);
not(notn3098,n2921);
and (s0n3098,notn3098,n3099);
and (s1n3098,n2921,n3100);
and (n3101,n3102,n2744);
or (n3102,1'b0,n3103,n3107,n3111,n3114);
and (n3103,n3104,n2924);
wire s0n3104,s1n3104,notn3104;
or (n3104,s0n3104,s1n3104);
not(notn3104,n2921);
and (s0n3104,notn3104,n3105);
and (s1n3104,n2921,n3106);
and (n3107,n3108,n2947);
wire s0n3108,s1n3108,notn3108;
or (n3108,s0n3108,s1n3108);
not(notn3108,n2921);
and (s0n3108,notn3108,n3109);
and (s1n3108,n2921,n3110);
and (n3111,n3112,n2955);
wire s0n3112,s1n3112,notn3112;
or (n3112,s0n3112,s1n3112);
not(notn3112,n2921);
and (s0n3112,notn3112,n2180);
and (s1n3112,n2921,n3113);
and (n3114,n3115,n2964);
wire s0n3115,s1n3115,notn3115;
or (n3115,s0n3115,s1n3115);
not(notn3115,n2921);
and (s0n3115,notn3115,n1844);
and (s1n3115,n2921,n3116);
or (n3117,1'b0,n3118,n3127,n3133,n3142);
and (n3118,n3119,n2710);
or (n3119,1'b0,n3120,n3124,n3125,n3126);
and (n3120,n3121,n2924);
wire s0n3121,s1n3121,notn3121;
or (n3121,s0n3121,s1n3121);
not(notn3121,n2921);
and (s0n3121,notn3121,n3122);
and (s1n3121,n2921,n3123);
and (n3124,n3050,n2947);
and (n3125,n3054,n2955);
and (n3126,n3058,n2964);
and (n3127,n3128,n2722);
or (n3128,1'b0,n3129,n3130,n3131,n3132);
and (n3129,n3062,n2924);
and (n3130,n3068,n2947);
and (n3131,n3072,n2955);
and (n3132,n3076,n2964);
and (n3133,n3134,n2734);
or (n3134,1'b0,n3135,n3139,n3140,n3141);
and (n3135,n3136,n2924);
wire s0n3136,s1n3136,notn3136;
or (n3136,s0n3136,s1n3136);
not(notn3136,n2921);
and (s0n3136,notn3136,n3137);
and (s1n3136,n2921,n3138);
and (n3139,n3086,n2947);
and (n3140,n3090,n2955);
and (n3141,n3094,n2964);
and (n3142,n3143,n2744);
or (n3143,1'b0,n3144,n3145,n3146,n3147);
and (n3144,n3098,n2924);
and (n3145,n3104,n2947);
and (n3146,n3108,n2955);
and (n3147,n3112,n2964);
and (n3148,n3117,n3149);
or (n3149,n3150,n3253,n3781);
and (n3150,n3151,n3222);
or (n3151,1'b0,n3152,n3170,n3188,n3206);
and (n3152,n3153,n2710);
or (n3153,1'b0,n3154,n3158,n3162,n3166);
and (n3154,n3155,n2924);
wire s0n3155,s1n3155,notn3155;
or (n3155,s0n3155,s1n3155);
not(notn3155,n2921);
and (s0n3155,notn3155,n3156);
and (s1n3155,n2921,n3157);
and (n3158,n3159,n2947);
wire s0n3159,s1n3159,notn3159;
or (n3159,s0n3159,s1n3159);
not(notn3159,n2921);
and (s0n3159,notn3159,n3160);
and (s1n3159,n2921,n3161);
and (n3162,n3163,n2955);
wire s0n3163,s1n3163,notn3163;
or (n3163,s0n3163,s1n3163);
not(notn3163,n2921);
and (s0n3163,notn3163,n3164);
and (s1n3163,n2921,n3165);
and (n3166,n3167,n2964);
wire s0n3167,s1n3167,notn3167;
or (n3167,s0n3167,s1n3167);
not(notn3167,n2921);
and (s0n3167,notn3167,n3168);
and (s1n3167,n2921,n3169);
and (n3170,n3171,n2722);
or (n3171,1'b0,n3172,n3176,n3180,n3184);
and (n3172,n3173,n2924);
wire s0n3173,s1n3173,notn3173;
or (n3173,s0n3173,s1n3173);
not(notn3173,n2921);
and (s0n3173,notn3173,n3174);
and (s1n3173,n2921,n3175);
and (n3176,n3177,n2947);
wire s0n3177,s1n3177,notn3177;
or (n3177,s0n3177,s1n3177);
not(notn3177,n2921);
and (s0n3177,notn3177,n3178);
and (s1n3177,n2921,n3179);
and (n3180,n3181,n2955);
wire s0n3181,s1n3181,notn3181;
or (n3181,s0n3181,s1n3181);
not(notn3181,n2921);
and (s0n3181,notn3181,n3182);
and (s1n3181,n2921,n3183);
and (n3184,n3185,n2964);
wire s0n3185,s1n3185,notn3185;
or (n3185,s0n3185,s1n3185);
not(notn3185,n2921);
and (s0n3185,notn3185,n3186);
and (s1n3185,n2921,n3187);
and (n3188,n3189,n2734);
or (n3189,1'b0,n3190,n3194,n3198,n3202);
and (n3190,n3191,n2924);
wire s0n3191,s1n3191,notn3191;
or (n3191,s0n3191,s1n3191);
not(notn3191,n2921);
and (s0n3191,notn3191,n3192);
and (s1n3191,n2921,n3193);
and (n3194,n3195,n2947);
wire s0n3195,s1n3195,notn3195;
or (n3195,s0n3195,s1n3195);
not(notn3195,n2921);
and (s0n3195,notn3195,n3196);
and (s1n3195,n2921,n3197);
and (n3198,n3199,n2955);
wire s0n3199,s1n3199,notn3199;
or (n3199,s0n3199,s1n3199);
not(notn3199,n2921);
and (s0n3199,notn3199,n3200);
and (s1n3199,n2921,n3201);
and (n3202,n3203,n2964);
wire s0n3203,s1n3203,notn3203;
or (n3203,s0n3203,s1n3203);
not(notn3203,n2921);
and (s0n3203,notn3203,n3204);
and (s1n3203,n2921,n3205);
and (n3206,n3207,n2744);
or (n3207,1'b0,n3208,n3212,n3216,n3219);
and (n3208,n3209,n2924);
wire s0n3209,s1n3209,notn3209;
or (n3209,s0n3209,s1n3209);
not(notn3209,n2921);
and (s0n3209,notn3209,n3210);
and (s1n3209,n2921,n3211);
and (n3212,n3213,n2947);
wire s0n3213,s1n3213,notn3213;
or (n3213,s0n3213,s1n3213);
not(notn3213,n2921);
and (s0n3213,notn3213,n3214);
and (s1n3213,n2921,n3215);
and (n3216,n3217,n2955);
wire s0n3217,s1n3217,notn3217;
or (n3217,s0n3217,s1n3217);
not(notn3217,n2921);
and (s0n3217,notn3217,n2196);
and (s1n3217,n2921,n3218);
and (n3219,n3220,n2964);
wire s0n3220,s1n3220,notn3220;
or (n3220,s0n3220,s1n3220);
not(notn3220,n2921);
and (s0n3220,notn3220,n1861);
and (s1n3220,n2921,n3221);
or (n3222,1'b0,n3223,n3232,n3238,n3247);
and (n3223,n3224,n2710);
or (n3224,1'b0,n3225,n3229,n3230,n3231);
and (n3225,n3226,n2924);
wire s0n3226,s1n3226,notn3226;
or (n3226,s0n3226,s1n3226);
not(notn3226,n2921);
and (s0n3226,notn3226,n3227);
and (s1n3226,n2921,n3228);
and (n3229,n3155,n2947);
and (n3230,n3159,n2955);
and (n3231,n3163,n2964);
and (n3232,n3233,n2722);
or (n3233,1'b0,n3234,n3235,n3236,n3237);
and (n3234,n3167,n2924);
and (n3235,n3173,n2947);
and (n3236,n3177,n2955);
and (n3237,n3181,n2964);
and (n3238,n3239,n2734);
or (n3239,1'b0,n3240,n3244,n3245,n3246);
and (n3240,n3241,n2924);
wire s0n3241,s1n3241,notn3241;
or (n3241,s0n3241,s1n3241);
not(notn3241,n2921);
and (s0n3241,notn3241,n3242);
and (s1n3241,n2921,n3243);
and (n3244,n3191,n2947);
and (n3245,n3195,n2955);
and (n3246,n3199,n2964);
and (n3247,n3248,n2744);
or (n3248,1'b0,n3249,n3250,n3251,n3252);
and (n3249,n3203,n2924);
and (n3250,n3209,n2947);
and (n3251,n3213,n2955);
and (n3252,n3217,n2964);
and (n3253,n3222,n3254);
or (n3254,n3255,n3358,n3780);
and (n3255,n3256,n3327);
or (n3256,1'b0,n3257,n3275,n3293,n3311);
and (n3257,n3258,n2710);
or (n3258,1'b0,n3259,n3263,n3267,n3271);
and (n3259,n3260,n2924);
wire s0n3260,s1n3260,notn3260;
or (n3260,s0n3260,s1n3260);
not(notn3260,n2921);
and (s0n3260,notn3260,n3261);
and (s1n3260,n2921,n3262);
and (n3263,n3264,n2947);
wire s0n3264,s1n3264,notn3264;
or (n3264,s0n3264,s1n3264);
not(notn3264,n2921);
and (s0n3264,notn3264,n3265);
and (s1n3264,n2921,n3266);
and (n3267,n3268,n2955);
wire s0n3268,s1n3268,notn3268;
or (n3268,s0n3268,s1n3268);
not(notn3268,n2921);
and (s0n3268,notn3268,n3269);
and (s1n3268,n2921,n3270);
and (n3271,n3272,n2964);
wire s0n3272,s1n3272,notn3272;
or (n3272,s0n3272,s1n3272);
not(notn3272,n2921);
and (s0n3272,notn3272,n3273);
and (s1n3272,n2921,n3274);
and (n3275,n3276,n2722);
or (n3276,1'b0,n3277,n3281,n3285,n3289);
and (n3277,n3278,n2924);
wire s0n3278,s1n3278,notn3278;
or (n3278,s0n3278,s1n3278);
not(notn3278,n2921);
and (s0n3278,notn3278,n3279);
and (s1n3278,n2921,n3280);
and (n3281,n3282,n2947);
wire s0n3282,s1n3282,notn3282;
or (n3282,s0n3282,s1n3282);
not(notn3282,n2921);
and (s0n3282,notn3282,n3283);
and (s1n3282,n2921,n3284);
and (n3285,n3286,n2955);
wire s0n3286,s1n3286,notn3286;
or (n3286,s0n3286,s1n3286);
not(notn3286,n2921);
and (s0n3286,notn3286,n3287);
and (s1n3286,n2921,n3288);
and (n3289,n3290,n2964);
wire s0n3290,s1n3290,notn3290;
or (n3290,s0n3290,s1n3290);
not(notn3290,n2921);
and (s0n3290,notn3290,n3291);
and (s1n3290,n2921,n3292);
and (n3293,n3294,n2734);
or (n3294,1'b0,n3295,n3299,n3303,n3307);
and (n3295,n3296,n2924);
wire s0n3296,s1n3296,notn3296;
or (n3296,s0n3296,s1n3296);
not(notn3296,n2921);
and (s0n3296,notn3296,n3297);
and (s1n3296,n2921,n3298);
and (n3299,n3300,n2947);
wire s0n3300,s1n3300,notn3300;
or (n3300,s0n3300,s1n3300);
not(notn3300,n2921);
and (s0n3300,notn3300,n3301);
and (s1n3300,n2921,n3302);
and (n3303,n3304,n2955);
wire s0n3304,s1n3304,notn3304;
or (n3304,s0n3304,s1n3304);
not(notn3304,n2921);
and (s0n3304,notn3304,n3305);
and (s1n3304,n2921,n3306);
and (n3307,n3308,n2964);
wire s0n3308,s1n3308,notn3308;
or (n3308,s0n3308,s1n3308);
not(notn3308,n2921);
and (s0n3308,notn3308,n3309);
and (s1n3308,n2921,n3310);
and (n3311,n3312,n2744);
or (n3312,1'b0,n3313,n3317,n3321,n3324);
and (n3313,n3314,n2924);
wire s0n3314,s1n3314,notn3314;
or (n3314,s0n3314,s1n3314);
not(notn3314,n2921);
and (s0n3314,notn3314,n3315);
and (s1n3314,n2921,n3316);
and (n3317,n3318,n2947);
wire s0n3318,s1n3318,notn3318;
or (n3318,s0n3318,s1n3318);
not(notn3318,n2921);
and (s0n3318,notn3318,n3319);
and (s1n3318,n2921,n3320);
and (n3321,n3322,n2955);
wire s0n3322,s1n3322,notn3322;
or (n3322,s0n3322,s1n3322);
not(notn3322,n2921);
and (s0n3322,notn3322,n2212);
and (s1n3322,n2921,n3323);
and (n3324,n3325,n2964);
wire s0n3325,s1n3325,notn3325;
or (n3325,s0n3325,s1n3325);
not(notn3325,n2921);
and (s0n3325,notn3325,n1886);
and (s1n3325,n2921,n3326);
or (n3327,1'b0,n3328,n3337,n3343,n3352);
and (n3328,n3329,n2710);
or (n3329,1'b0,n3330,n3334,n3335,n3336);
and (n3330,n3331,n2924);
wire s0n3331,s1n3331,notn3331;
or (n3331,s0n3331,s1n3331);
not(notn3331,n2921);
and (s0n3331,notn3331,n3332);
and (s1n3331,n2921,n3333);
and (n3334,n3260,n2947);
and (n3335,n3264,n2955);
and (n3336,n3268,n2964);
and (n3337,n3338,n2722);
or (n3338,1'b0,n3339,n3340,n3341,n3342);
and (n3339,n3272,n2924);
and (n3340,n3278,n2947);
and (n3341,n3282,n2955);
and (n3342,n3286,n2964);
and (n3343,n3344,n2734);
or (n3344,1'b0,n3345,n3349,n3350,n3351);
and (n3345,n3346,n2924);
wire s0n3346,s1n3346,notn3346;
or (n3346,s0n3346,s1n3346);
not(notn3346,n2921);
and (s0n3346,notn3346,n3347);
and (s1n3346,n2921,n3348);
and (n3349,n3296,n2947);
and (n3350,n3300,n2955);
and (n3351,n3304,n2964);
and (n3352,n3353,n2744);
or (n3353,1'b0,n3354,n3355,n3356,n3357);
and (n3354,n3308,n2924);
and (n3355,n3314,n2947);
and (n3356,n3318,n2955);
and (n3357,n3322,n2964);
and (n3358,n3327,n3359);
or (n3359,n3360,n3463,n3779);
and (n3360,n3361,n3432);
or (n3361,1'b0,n3362,n3380,n3398,n3416);
and (n3362,n3363,n2710);
or (n3363,1'b0,n3364,n3368,n3372,n3376);
and (n3364,n3365,n2924);
wire s0n3365,s1n3365,notn3365;
or (n3365,s0n3365,s1n3365);
not(notn3365,n2921);
and (s0n3365,notn3365,n3366);
and (s1n3365,n2921,n3367);
and (n3368,n3369,n2947);
wire s0n3369,s1n3369,notn3369;
or (n3369,s0n3369,s1n3369);
not(notn3369,n2921);
and (s0n3369,notn3369,n3370);
and (s1n3369,n2921,n3371);
and (n3372,n3373,n2955);
wire s0n3373,s1n3373,notn3373;
or (n3373,s0n3373,s1n3373);
not(notn3373,n2921);
and (s0n3373,notn3373,n3374);
and (s1n3373,n2921,n3375);
and (n3376,n3377,n2964);
wire s0n3377,s1n3377,notn3377;
or (n3377,s0n3377,s1n3377);
not(notn3377,n2921);
and (s0n3377,notn3377,n3378);
and (s1n3377,n2921,n3379);
and (n3380,n3381,n2722);
or (n3381,1'b0,n3382,n3386,n3390,n3394);
and (n3382,n3383,n2924);
wire s0n3383,s1n3383,notn3383;
or (n3383,s0n3383,s1n3383);
not(notn3383,n2921);
and (s0n3383,notn3383,n3384);
and (s1n3383,n2921,n3385);
and (n3386,n3387,n2947);
wire s0n3387,s1n3387,notn3387;
or (n3387,s0n3387,s1n3387);
not(notn3387,n2921);
and (s0n3387,notn3387,n3388);
and (s1n3387,n2921,n3389);
and (n3390,n3391,n2955);
wire s0n3391,s1n3391,notn3391;
or (n3391,s0n3391,s1n3391);
not(notn3391,n2921);
and (s0n3391,notn3391,n3392);
and (s1n3391,n2921,n3393);
and (n3394,n3395,n2964);
wire s0n3395,s1n3395,notn3395;
or (n3395,s0n3395,s1n3395);
not(notn3395,n2921);
and (s0n3395,notn3395,n3396);
and (s1n3395,n2921,n3397);
and (n3398,n3399,n2734);
or (n3399,1'b0,n3400,n3404,n3408,n3412);
and (n3400,n3401,n2924);
wire s0n3401,s1n3401,notn3401;
or (n3401,s0n3401,s1n3401);
not(notn3401,n2921);
and (s0n3401,notn3401,n3402);
and (s1n3401,n2921,n3403);
and (n3404,n3405,n2947);
wire s0n3405,s1n3405,notn3405;
or (n3405,s0n3405,s1n3405);
not(notn3405,n2921);
and (s0n3405,notn3405,n3406);
and (s1n3405,n2921,n3407);
and (n3408,n3409,n2955);
wire s0n3409,s1n3409,notn3409;
or (n3409,s0n3409,s1n3409);
not(notn3409,n2921);
and (s0n3409,notn3409,n3410);
and (s1n3409,n2921,n3411);
and (n3412,n3413,n2964);
wire s0n3413,s1n3413,notn3413;
or (n3413,s0n3413,s1n3413);
not(notn3413,n2921);
and (s0n3413,notn3413,n3414);
and (s1n3413,n2921,n3415);
and (n3416,n3417,n2744);
or (n3417,1'b0,n3418,n3422,n3426,n3429);
and (n3418,n3419,n2924);
wire s0n3419,s1n3419,notn3419;
or (n3419,s0n3419,s1n3419);
not(notn3419,n2921);
and (s0n3419,notn3419,n3420);
and (s1n3419,n2921,n3421);
and (n3422,n3423,n2947);
wire s0n3423,s1n3423,notn3423;
or (n3423,s0n3423,s1n3423);
not(notn3423,n2921);
and (s0n3423,notn3423,n3424);
and (s1n3423,n2921,n3425);
and (n3426,n3427,n2955);
wire s0n3427,s1n3427,notn3427;
or (n3427,s0n3427,s1n3427);
not(notn3427,n2921);
and (s0n3427,notn3427,n2228);
and (s1n3427,n2921,n3428);
and (n3429,n3430,n2964);
wire s0n3430,s1n3430,notn3430;
or (n3430,s0n3430,s1n3430);
not(notn3430,n2921);
and (s0n3430,notn3430,n1913);
and (s1n3430,n2921,n3431);
or (n3432,1'b0,n3433,n3442,n3448,n3457);
and (n3433,n3434,n2710);
or (n3434,1'b0,n3435,n3439,n3440,n3441);
and (n3435,n3436,n2924);
wire s0n3436,s1n3436,notn3436;
or (n3436,s0n3436,s1n3436);
not(notn3436,n2921);
and (s0n3436,notn3436,n3437);
and (s1n3436,n2921,n3438);
and (n3439,n3365,n2947);
and (n3440,n3369,n2955);
and (n3441,n3373,n2964);
and (n3442,n3443,n2722);
or (n3443,1'b0,n3444,n3445,n3446,n3447);
and (n3444,n3377,n2924);
and (n3445,n3383,n2947);
and (n3446,n3387,n2955);
and (n3447,n3391,n2964);
and (n3448,n3449,n2734);
or (n3449,1'b0,n3450,n3454,n3455,n3456);
and (n3450,n3451,n2924);
wire s0n3451,s1n3451,notn3451;
or (n3451,s0n3451,s1n3451);
not(notn3451,n2921);
and (s0n3451,notn3451,n3452);
and (s1n3451,n2921,n3453);
and (n3454,n3401,n2947);
and (n3455,n3405,n2955);
and (n3456,n3409,n2964);
and (n3457,n3458,n2744);
or (n3458,1'b0,n3459,n3460,n3461,n3462);
and (n3459,n3413,n2924);
and (n3460,n3419,n2947);
and (n3461,n3423,n2955);
and (n3462,n3427,n2964);
and (n3463,n3432,n3464);
or (n3464,n3465,n3568,n3778);
and (n3465,n3466,n3537);
or (n3466,1'b0,n3467,n3485,n3503,n3521);
and (n3467,n3468,n2710);
or (n3468,1'b0,n3469,n3473,n3477,n3481);
and (n3469,n3470,n2924);
wire s0n3470,s1n3470,notn3470;
or (n3470,s0n3470,s1n3470);
not(notn3470,n2921);
and (s0n3470,notn3470,n3471);
and (s1n3470,n2921,n3472);
and (n3473,n3474,n2947);
wire s0n3474,s1n3474,notn3474;
or (n3474,s0n3474,s1n3474);
not(notn3474,n2921);
and (s0n3474,notn3474,n3475);
and (s1n3474,n2921,n3476);
and (n3477,n3478,n2955);
wire s0n3478,s1n3478,notn3478;
or (n3478,s0n3478,s1n3478);
not(notn3478,n2921);
and (s0n3478,notn3478,n3479);
and (s1n3478,n2921,n3480);
and (n3481,n3482,n2964);
wire s0n3482,s1n3482,notn3482;
or (n3482,s0n3482,s1n3482);
not(notn3482,n2921);
and (s0n3482,notn3482,n3483);
and (s1n3482,n2921,n3484);
and (n3485,n3486,n2722);
or (n3486,1'b0,n3487,n3491,n3495,n3499);
and (n3487,n3488,n2924);
wire s0n3488,s1n3488,notn3488;
or (n3488,s0n3488,s1n3488);
not(notn3488,n2921);
and (s0n3488,notn3488,n3489);
and (s1n3488,n2921,n3490);
and (n3491,n3492,n2947);
wire s0n3492,s1n3492,notn3492;
or (n3492,s0n3492,s1n3492);
not(notn3492,n2921);
and (s0n3492,notn3492,n3493);
and (s1n3492,n2921,n3494);
and (n3495,n3496,n2955);
wire s0n3496,s1n3496,notn3496;
or (n3496,s0n3496,s1n3496);
not(notn3496,n2921);
and (s0n3496,notn3496,n3497);
and (s1n3496,n2921,n3498);
and (n3499,n3500,n2964);
wire s0n3500,s1n3500,notn3500;
or (n3500,s0n3500,s1n3500);
not(notn3500,n2921);
and (s0n3500,notn3500,n3501);
and (s1n3500,n2921,n3502);
and (n3503,n3504,n2734);
or (n3504,1'b0,n3505,n3509,n3513,n3517);
and (n3505,n3506,n2924);
wire s0n3506,s1n3506,notn3506;
or (n3506,s0n3506,s1n3506);
not(notn3506,n2921);
and (s0n3506,notn3506,n3507);
and (s1n3506,n2921,n3508);
and (n3509,n3510,n2947);
wire s0n3510,s1n3510,notn3510;
or (n3510,s0n3510,s1n3510);
not(notn3510,n2921);
and (s0n3510,notn3510,n3511);
and (s1n3510,n2921,n3512);
and (n3513,n3514,n2955);
wire s0n3514,s1n3514,notn3514;
or (n3514,s0n3514,s1n3514);
not(notn3514,n2921);
and (s0n3514,notn3514,n3515);
and (s1n3514,n2921,n3516);
and (n3517,n3518,n2964);
wire s0n3518,s1n3518,notn3518;
or (n3518,s0n3518,s1n3518);
not(notn3518,n2921);
and (s0n3518,notn3518,n3519);
and (s1n3518,n2921,n3520);
and (n3521,n3522,n2744);
or (n3522,1'b0,n3523,n3527,n3531,n3534);
and (n3523,n3524,n2924);
wire s0n3524,s1n3524,notn3524;
or (n3524,s0n3524,s1n3524);
not(notn3524,n2921);
and (s0n3524,notn3524,n3525);
and (s1n3524,n2921,n3526);
and (n3527,n3528,n2947);
wire s0n3528,s1n3528,notn3528;
or (n3528,s0n3528,s1n3528);
not(notn3528,n2921);
and (s0n3528,notn3528,n3529);
and (s1n3528,n2921,n3530);
and (n3531,n3532,n2955);
wire s0n3532,s1n3532,notn3532;
or (n3532,s0n3532,s1n3532);
not(notn3532,n2921);
and (s0n3532,notn3532,n2244);
and (s1n3532,n2921,n3533);
and (n3534,n3535,n2964);
wire s0n3535,s1n3535,notn3535;
or (n3535,s0n3535,s1n3535);
not(notn3535,n2921);
and (s0n3535,notn3535,n1939);
and (s1n3535,n2921,n3536);
or (n3537,1'b0,n3538,n3547,n3553,n3562);
and (n3538,n3539,n2710);
or (n3539,1'b0,n3540,n3544,n3545,n3546);
and (n3540,n3541,n2924);
wire s0n3541,s1n3541,notn3541;
or (n3541,s0n3541,s1n3541);
not(notn3541,n2921);
and (s0n3541,notn3541,n3542);
and (s1n3541,n2921,n3543);
and (n3544,n3470,n2947);
and (n3545,n3474,n2955);
and (n3546,n3478,n2964);
and (n3547,n3548,n2722);
or (n3548,1'b0,n3549,n3550,n3551,n3552);
and (n3549,n3482,n2924);
and (n3550,n3488,n2947);
and (n3551,n3492,n2955);
and (n3552,n3496,n2964);
and (n3553,n3554,n2734);
or (n3554,1'b0,n3555,n3559,n3560,n3561);
and (n3555,n3556,n2924);
wire s0n3556,s1n3556,notn3556;
or (n3556,s0n3556,s1n3556);
not(notn3556,n2921);
and (s0n3556,notn3556,n3557);
and (s1n3556,n2921,n3558);
and (n3559,n3506,n2947);
and (n3560,n3510,n2955);
and (n3561,n3514,n2964);
and (n3562,n3563,n2744);
or (n3563,1'b0,n3564,n3565,n3566,n3567);
and (n3564,n3518,n2924);
and (n3565,n3524,n2947);
and (n3566,n3528,n2955);
and (n3567,n3532,n2964);
and (n3568,n3537,n3569);
or (n3569,n3570,n3673,n3777);
and (n3570,n3571,n3642);
or (n3571,1'b0,n3572,n3590,n3608,n3626);
and (n3572,n3573,n2710);
or (n3573,1'b0,n3574,n3578,n3582,n3586);
and (n3574,n3575,n2924);
wire s0n3575,s1n3575,notn3575;
or (n3575,s0n3575,s1n3575);
not(notn3575,n2921);
and (s0n3575,notn3575,n3576);
and (s1n3575,n2921,n3577);
and (n3578,n3579,n2947);
wire s0n3579,s1n3579,notn3579;
or (n3579,s0n3579,s1n3579);
not(notn3579,n2921);
and (s0n3579,notn3579,n3580);
and (s1n3579,n2921,n3581);
and (n3582,n3583,n2955);
wire s0n3583,s1n3583,notn3583;
or (n3583,s0n3583,s1n3583);
not(notn3583,n2921);
and (s0n3583,notn3583,n3584);
and (s1n3583,n2921,n3585);
and (n3586,n3587,n2964);
wire s0n3587,s1n3587,notn3587;
or (n3587,s0n3587,s1n3587);
not(notn3587,n2921);
and (s0n3587,notn3587,n3588);
and (s1n3587,n2921,n3589);
and (n3590,n3591,n2722);
or (n3591,1'b0,n3592,n3596,n3600,n3604);
and (n3592,n3593,n2924);
wire s0n3593,s1n3593,notn3593;
or (n3593,s0n3593,s1n3593);
not(notn3593,n2921);
and (s0n3593,notn3593,n3594);
and (s1n3593,n2921,n3595);
and (n3596,n3597,n2947);
wire s0n3597,s1n3597,notn3597;
or (n3597,s0n3597,s1n3597);
not(notn3597,n2921);
and (s0n3597,notn3597,n3598);
and (s1n3597,n2921,n3599);
and (n3600,n3601,n2955);
wire s0n3601,s1n3601,notn3601;
or (n3601,s0n3601,s1n3601);
not(notn3601,n2921);
and (s0n3601,notn3601,n3602);
and (s1n3601,n2921,n3603);
and (n3604,n3605,n2964);
wire s0n3605,s1n3605,notn3605;
or (n3605,s0n3605,s1n3605);
not(notn3605,n2921);
and (s0n3605,notn3605,n3606);
and (s1n3605,n2921,n3607);
and (n3608,n3609,n2734);
or (n3609,1'b0,n3610,n3614,n3618,n3622);
and (n3610,n3611,n2924);
wire s0n3611,s1n3611,notn3611;
or (n3611,s0n3611,s1n3611);
not(notn3611,n2921);
and (s0n3611,notn3611,n3612);
and (s1n3611,n2921,n3613);
and (n3614,n3615,n2947);
wire s0n3615,s1n3615,notn3615;
or (n3615,s0n3615,s1n3615);
not(notn3615,n2921);
and (s0n3615,notn3615,n3616);
and (s1n3615,n2921,n3617);
and (n3618,n3619,n2955);
wire s0n3619,s1n3619,notn3619;
or (n3619,s0n3619,s1n3619);
not(notn3619,n2921);
and (s0n3619,notn3619,n3620);
and (s1n3619,n2921,n3621);
and (n3622,n3623,n2964);
wire s0n3623,s1n3623,notn3623;
or (n3623,s0n3623,s1n3623);
not(notn3623,n2921);
and (s0n3623,notn3623,n3624);
and (s1n3623,n2921,n3625);
and (n3626,n3627,n2744);
or (n3627,1'b0,n3628,n3632,n3636,n3639);
and (n3628,n3629,n2924);
wire s0n3629,s1n3629,notn3629;
or (n3629,s0n3629,s1n3629);
not(notn3629,n2921);
and (s0n3629,notn3629,n3630);
and (s1n3629,n2921,n3631);
and (n3632,n3633,n2947);
wire s0n3633,s1n3633,notn3633;
or (n3633,s0n3633,s1n3633);
not(notn3633,n2921);
and (s0n3633,notn3633,n3634);
and (s1n3633,n2921,n3635);
and (n3636,n3637,n2955);
wire s0n3637,s1n3637,notn3637;
or (n3637,s0n3637,s1n3637);
not(notn3637,n2921);
and (s0n3637,notn3637,n2260);
and (s1n3637,n2921,n3638);
and (n3639,n3640,n2964);
wire s0n3640,s1n3640,notn3640;
or (n3640,s0n3640,s1n3640);
not(notn3640,n2921);
and (s0n3640,notn3640,n1968);
and (s1n3640,n2921,n3641);
or (n3642,1'b0,n3643,n3652,n3658,n3667);
and (n3643,n3644,n2710);
or (n3644,1'b0,n3645,n3649,n3650,n3651);
and (n3645,n3646,n2924);
wire s0n3646,s1n3646,notn3646;
or (n3646,s0n3646,s1n3646);
not(notn3646,n2921);
and (s0n3646,notn3646,n3647);
and (s1n3646,n2921,n3648);
and (n3649,n3575,n2947);
and (n3650,n3579,n2955);
and (n3651,n3583,n2964);
and (n3652,n3653,n2722);
or (n3653,1'b0,n3654,n3655,n3656,n3657);
and (n3654,n3587,n2924);
and (n3655,n3593,n2947);
and (n3656,n3597,n2955);
and (n3657,n3601,n2964);
and (n3658,n3659,n2734);
or (n3659,1'b0,n3660,n3664,n3665,n3666);
and (n3660,n3661,n2924);
wire s0n3661,s1n3661,notn3661;
or (n3661,s0n3661,s1n3661);
not(notn3661,n2921);
and (s0n3661,notn3661,n3662);
and (s1n3661,n2921,n3663);
and (n3664,n3611,n2947);
and (n3665,n3615,n2955);
and (n3666,n3619,n2964);
and (n3667,n3668,n2744);
or (n3668,1'b0,n3669,n3670,n3671,n3672);
and (n3669,n3623,n2924);
and (n3670,n3629,n2947);
and (n3671,n3633,n2955);
and (n3672,n3637,n2964);
and (n3673,n3642,n3674);
and (n3674,n3675,n3746);
or (n3675,1'b0,n3676,n3694,n3712,n3730);
and (n3676,n3677,n2710);
or (n3677,1'b0,n3678,n3682,n3686,n3690);
and (n3678,n3679,n2924);
wire s0n3679,s1n3679,notn3679;
or (n3679,s0n3679,s1n3679);
not(notn3679,n2921);
and (s0n3679,notn3679,n3680);
and (s1n3679,n2921,n3681);
and (n3682,n3683,n2947);
wire s0n3683,s1n3683,notn3683;
or (n3683,s0n3683,s1n3683);
not(notn3683,n2921);
and (s0n3683,notn3683,n3684);
and (s1n3683,n2921,n3685);
and (n3686,n3687,n2955);
wire s0n3687,s1n3687,notn3687;
or (n3687,s0n3687,s1n3687);
not(notn3687,n2921);
and (s0n3687,notn3687,n3688);
and (s1n3687,n2921,n3689);
and (n3690,n3691,n2964);
wire s0n3691,s1n3691,notn3691;
or (n3691,s0n3691,s1n3691);
not(notn3691,n2921);
and (s0n3691,notn3691,n3692);
and (s1n3691,n2921,n3693);
and (n3694,n3695,n2722);
or (n3695,1'b0,n3696,n3700,n3704,n3708);
and (n3696,n3697,n2924);
wire s0n3697,s1n3697,notn3697;
or (n3697,s0n3697,s1n3697);
not(notn3697,n2921);
and (s0n3697,notn3697,n3698);
and (s1n3697,n2921,n3699);
and (n3700,n3701,n2947);
wire s0n3701,s1n3701,notn3701;
or (n3701,s0n3701,s1n3701);
not(notn3701,n2921);
and (s0n3701,notn3701,n3702);
and (s1n3701,n2921,n3703);
and (n3704,n3705,n2955);
wire s0n3705,s1n3705,notn3705;
or (n3705,s0n3705,s1n3705);
not(notn3705,n2921);
and (s0n3705,notn3705,n3706);
and (s1n3705,n2921,n3707);
and (n3708,n3709,n2964);
wire s0n3709,s1n3709,notn3709;
or (n3709,s0n3709,s1n3709);
not(notn3709,n2921);
and (s0n3709,notn3709,n3710);
and (s1n3709,n2921,n3711);
and (n3712,n3713,n2734);
or (n3713,1'b0,n3714,n3718,n3722,n3726);
and (n3714,n3715,n2924);
wire s0n3715,s1n3715,notn3715;
or (n3715,s0n3715,s1n3715);
not(notn3715,n2921);
and (s0n3715,notn3715,n3716);
and (s1n3715,n2921,n3717);
and (n3718,n3719,n2947);
wire s0n3719,s1n3719,notn3719;
or (n3719,s0n3719,s1n3719);
not(notn3719,n2921);
and (s0n3719,notn3719,n3720);
and (s1n3719,n2921,n3721);
and (n3722,n3723,n2955);
wire s0n3723,s1n3723,notn3723;
or (n3723,s0n3723,s1n3723);
not(notn3723,n2921);
and (s0n3723,notn3723,n3724);
and (s1n3723,n2921,n3725);
and (n3726,n3727,n2964);
wire s0n3727,s1n3727,notn3727;
or (n3727,s0n3727,s1n3727);
not(notn3727,n2921);
and (s0n3727,notn3727,n3728);
and (s1n3727,n2921,n3729);
and (n3730,n3731,n2744);
or (n3731,1'b0,n3732,n3736,n3740,n3743);
and (n3732,n3733,n2924);
wire s0n3733,s1n3733,notn3733;
or (n3733,s0n3733,s1n3733);
not(notn3733,n2921);
and (s0n3733,notn3733,n3734);
and (s1n3733,n2921,n3735);
and (n3736,n3737,n2947);
wire s0n3737,s1n3737,notn3737;
or (n3737,s0n3737,s1n3737);
not(notn3737,n2921);
and (s0n3737,notn3737,n3738);
and (s1n3737,n2921,n3739);
and (n3740,n3741,n2955);
wire s0n3741,s1n3741,notn3741;
or (n3741,s0n3741,s1n3741);
not(notn3741,n2921);
and (s0n3741,notn3741,n2275);
and (s1n3741,n2921,n3742);
and (n3743,n3744,n2964);
wire s0n3744,s1n3744,notn3744;
or (n3744,s0n3744,s1n3744);
not(notn3744,n2921);
and (s0n3744,notn3744,n1987);
and (s1n3744,n2921,n3745);
or (n3746,1'b0,n3747,n3756,n3762,n3771);
and (n3747,n3748,n2710);
or (n3748,1'b0,n3749,n3753,n3754,n3755);
and (n3749,n3750,n2924);
wire s0n3750,s1n3750,notn3750;
or (n3750,s0n3750,s1n3750);
not(notn3750,n2921);
and (s0n3750,notn3750,n3751);
and (s1n3750,n2921,n3752);
and (n3753,n3679,n2947);
and (n3754,n3683,n2955);
and (n3755,n3687,n2964);
and (n3756,n3757,n2722);
or (n3757,1'b0,n3758,n3759,n3760,n3761);
and (n3758,n3691,n2924);
and (n3759,n3697,n2947);
and (n3760,n3701,n2955);
and (n3761,n3705,n2964);
and (n3762,n3763,n2734);
or (n3763,1'b0,n3764,n3768,n3769,n3770);
and (n3764,n3765,n2924);
wire s0n3765,s1n3765,notn3765;
or (n3765,s0n3765,s1n3765);
not(notn3765,n2921);
and (s0n3765,notn3765,n3766);
and (s1n3765,n2921,n3767);
and (n3768,n3715,n2947);
and (n3769,n3719,n2955);
and (n3770,n3723,n2964);
and (n3771,n3772,n2744);
or (n3772,1'b0,n3773,n3774,n3775,n3776);
and (n3773,n3727,n2924);
and (n3774,n3733,n2947);
and (n3775,n3737,n2955);
and (n3776,n3741,n2964);
and (n3777,n3571,n3674);
and (n3778,n3466,n3569);
and (n3779,n3361,n3464);
and (n3780,n3256,n3359);
and (n3781,n3151,n3254);
and (n3782,n3046,n3149);
and (n3783,n2915,n3044);
or (n3784,n3785,n3787);
xor (n3785,n3786,n3044);
xor (n3786,n2915,n3012);
or (n3787,n3788,n4318,n4369);
and (n3788,n3789,n3791);
xor (n3789,n3790,n3149);
xor (n3790,n3046,n3117);
not (n3791,n3792);
or (n3792,n3793,n3855,n4317);
and (n3793,n3794,n3824);
or (n3794,1'b0,n3795,n3801,n3810,n3816);
and (n3795,n3796,n2710);
or (n3796,1'b0,n3797,n3798,n3799,n3800);
and (n3797,n2945,n2924);
and (n3798,n2953,n2947);
and (n3799,n2962,n2955);
and (n3800,n2973,n2964);
and (n3801,n3802,n2722);
or (n3802,1'b0,n3803,n3804,n3805,n3806);
and (n3803,n2976,n2924);
and (n3804,n2979,n2947);
and (n3805,n2982,n2955);
and (n3806,n3807,n2964);
wire s0n3807,s1n3807,notn3807;
or (n3807,s0n3807,s1n3807);
not(notn3807,n2921);
and (s0n3807,notn3807,n3808);
and (s1n3807,n2921,n3809);
and (n3810,n3811,n2734);
or (n3811,1'b0,n3812,n3813,n3814,n3815);
and (n3812,n2990,n2924);
and (n3813,n2993,n2947);
and (n3814,n2996,n2955);
and (n3815,n3001,n2964);
and (n3816,n3817,n2744);
or (n3817,1'b0,n3818,n3819,n3820,n3821);
and (n3818,n3004,n2924);
and (n3819,n3007,n2947);
and (n3820,n3010,n2955);
and (n3821,n3822,n2964);
wire s0n3822,s1n3822,notn3822;
or (n3822,s0n3822,s1n3822);
not(notn3822,n2921);
and (s0n3822,notn3822,n2166);
and (s1n3822,n2921,n3823);
or (n3824,1'b0,n3825,n3834,n3840,n3849);
and (n3825,n3826,n2710);
or (n3826,1'b0,n3827,n3831,n3832,n3833);
and (n3827,n3828,n2924);
wire s0n3828,s1n3828,notn3828;
or (n3828,s0n3828,s1n3828);
not(notn3828,n2921);
and (s0n3828,notn3828,n3829);
and (s1n3828,n2921,n3830);
and (n3831,n3016,n2947);
and (n3832,n2919,n2955);
and (n3833,n2945,n2964);
and (n3834,n3835,n2722);
or (n3835,1'b0,n3836,n3837,n3838,n3839);
and (n3836,n2953,n2924);
and (n3837,n2962,n2947);
and (n3838,n2973,n2955);
and (n3839,n2976,n2964);
and (n3840,n3841,n2734);
or (n3841,1'b0,n3842,n3846,n3847,n3848);
and (n3842,n3843,n2924);
wire s0n3843,s1n3843,notn3843;
or (n3843,s0n3843,s1n3843);
not(notn3843,n2921);
and (s0n3843,notn3843,n3844);
and (s1n3843,n2921,n3845);
and (n3846,n3031,n2947);
and (n3847,n2987,n2955);
and (n3848,n2990,n2964);
and (n3849,n3850,n2744);
or (n3850,1'b0,n3851,n3852,n3853,n3854);
and (n3851,n2993,n2924);
and (n3852,n2996,n2947);
and (n3853,n3001,n2955);
and (n3854,n3004,n2964);
and (n3855,n3824,n3856);
or (n3856,n3857,n3919,n4316);
and (n3857,n3858,n3888);
or (n3858,1'b0,n3859,n3865,n3874,n3880);
and (n3859,n3860,n2710);
or (n3860,1'b0,n3861,n3862,n3863,n3864);
and (n3861,n3054,n2924);
and (n3862,n3058,n2947);
and (n3863,n3062,n2955);
and (n3864,n3068,n2964);
and (n3865,n3866,n2722);
or (n3866,1'b0,n3867,n3868,n3869,n3870);
and (n3867,n3072,n2924);
and (n3868,n3076,n2947);
and (n3869,n3080,n2955);
and (n3870,n3871,n2964);
wire s0n3871,s1n3871,notn3871;
or (n3871,s0n3871,s1n3871);
not(notn3871,n2921);
and (s0n3871,notn3871,n3872);
and (s1n3871,n2921,n3873);
and (n3874,n3875,n2734);
or (n3875,1'b0,n3876,n3877,n3878,n3879);
and (n3876,n3090,n2924);
and (n3877,n3094,n2947);
and (n3878,n3098,n2955);
and (n3879,n3104,n2964);
and (n3880,n3881,n2744);
or (n3881,1'b0,n3882,n3883,n3884,n3885);
and (n3882,n3108,n2924);
and (n3883,n3112,n2947);
and (n3884,n3115,n2955);
and (n3885,n3886,n2964);
wire s0n3886,s1n3886,notn3886;
or (n3886,s0n3886,s1n3886);
not(notn3886,n2921);
and (s0n3886,notn3886,n2182);
and (s1n3886,n2921,n3887);
or (n3888,1'b0,n3889,n3898,n3904,n3913);
and (n3889,n3890,n2710);
or (n3890,1'b0,n3891,n3895,n3896,n3897);
and (n3891,n3892,n2924);
wire s0n3892,s1n3892,notn3892;
or (n3892,s0n3892,s1n3892);
not(notn3892,n2921);
and (s0n3892,notn3892,n3893);
and (s1n3892,n2921,n3894);
and (n3895,n3121,n2947);
and (n3896,n3050,n2955);
and (n3897,n3054,n2964);
and (n3898,n3899,n2722);
or (n3899,1'b0,n3900,n3901,n3902,n3903);
and (n3900,n3058,n2924);
and (n3901,n3062,n2947);
and (n3902,n3068,n2955);
and (n3903,n3072,n2964);
and (n3904,n3905,n2734);
or (n3905,1'b0,n3906,n3910,n3911,n3912);
and (n3906,n3907,n2924);
wire s0n3907,s1n3907,notn3907;
or (n3907,s0n3907,s1n3907);
not(notn3907,n2921);
and (s0n3907,notn3907,n3908);
and (s1n3907,n2921,n3909);
and (n3910,n3136,n2947);
and (n3911,n3086,n2955);
and (n3912,n3090,n2964);
and (n3913,n3914,n2744);
or (n3914,1'b0,n3915,n3916,n3917,n3918);
and (n3915,n3094,n2924);
and (n3916,n3098,n2947);
and (n3917,n3104,n2955);
and (n3918,n3108,n2964);
and (n3919,n3888,n3920);
or (n3920,n3921,n3983,n4315);
and (n3921,n3922,n3952);
or (n3922,1'b0,n3923,n3929,n3938,n3944);
and (n3923,n3924,n2710);
or (n3924,1'b0,n3925,n3926,n3927,n3928);
and (n3925,n3159,n2924);
and (n3926,n3163,n2947);
and (n3927,n3167,n2955);
and (n3928,n3173,n2964);
and (n3929,n3930,n2722);
or (n3930,1'b0,n3931,n3932,n3933,n3934);
and (n3931,n3177,n2924);
and (n3932,n3181,n2947);
and (n3933,n3185,n2955);
and (n3934,n3935,n2964);
wire s0n3935,s1n3935,notn3935;
or (n3935,s0n3935,s1n3935);
not(notn3935,n2921);
and (s0n3935,notn3935,n3936);
and (s1n3935,n2921,n3937);
and (n3938,n3939,n2734);
or (n3939,1'b0,n3940,n3941,n3942,n3943);
and (n3940,n3195,n2924);
and (n3941,n3199,n2947);
and (n3942,n3203,n2955);
and (n3943,n3209,n2964);
and (n3944,n3945,n2744);
or (n3945,1'b0,n3946,n3947,n3948,n3949);
and (n3946,n3213,n2924);
and (n3947,n3217,n2947);
and (n3948,n3220,n2955);
and (n3949,n3950,n2964);
wire s0n3950,s1n3950,notn3950;
or (n3950,s0n3950,s1n3950);
not(notn3950,n2921);
and (s0n3950,notn3950,n2198);
and (s1n3950,n2921,n3951);
or (n3952,1'b0,n3953,n3962,n3968,n3977);
and (n3953,n3954,n2710);
or (n3954,1'b0,n3955,n3959,n3960,n3961);
and (n3955,n3956,n2924);
wire s0n3956,s1n3956,notn3956;
or (n3956,s0n3956,s1n3956);
not(notn3956,n2921);
and (s0n3956,notn3956,n3957);
and (s1n3956,n2921,n3958);
and (n3959,n3226,n2947);
and (n3960,n3155,n2955);
and (n3961,n3159,n2964);
and (n3962,n3963,n2722);
or (n3963,1'b0,n3964,n3965,n3966,n3967);
and (n3964,n3163,n2924);
and (n3965,n3167,n2947);
and (n3966,n3173,n2955);
and (n3967,n3177,n2964);
and (n3968,n3969,n2734);
or (n3969,1'b0,n3970,n3974,n3975,n3976);
and (n3970,n3971,n2924);
wire s0n3971,s1n3971,notn3971;
or (n3971,s0n3971,s1n3971);
not(notn3971,n2921);
and (s0n3971,notn3971,n3972);
and (s1n3971,n2921,n3973);
and (n3974,n3241,n2947);
and (n3975,n3191,n2955);
and (n3976,n3195,n2964);
and (n3977,n3978,n2744);
or (n3978,1'b0,n3979,n3980,n3981,n3982);
and (n3979,n3199,n2924);
and (n3980,n3203,n2947);
and (n3981,n3209,n2955);
and (n3982,n3213,n2964);
and (n3983,n3952,n3984);
or (n3984,n3985,n4047,n4314);
and (n3985,n3986,n4016);
or (n3986,1'b0,n3987,n3993,n4002,n4008);
and (n3987,n3988,n2710);
or (n3988,1'b0,n3989,n3990,n3991,n3992);
and (n3989,n3264,n2924);
and (n3990,n3268,n2947);
and (n3991,n3272,n2955);
and (n3992,n3278,n2964);
and (n3993,n3994,n2722);
or (n3994,1'b0,n3995,n3996,n3997,n3998);
and (n3995,n3282,n2924);
and (n3996,n3286,n2947);
and (n3997,n3290,n2955);
and (n3998,n3999,n2964);
wire s0n3999,s1n3999,notn3999;
or (n3999,s0n3999,s1n3999);
not(notn3999,n2921);
and (s0n3999,notn3999,n4000);
and (s1n3999,n2921,n4001);
and (n4002,n4003,n2734);
or (n4003,1'b0,n4004,n4005,n4006,n4007);
and (n4004,n3300,n2924);
and (n4005,n3304,n2947);
and (n4006,n3308,n2955);
and (n4007,n3314,n2964);
and (n4008,n4009,n2744);
or (n4009,1'b0,n4010,n4011,n4012,n4013);
and (n4010,n3318,n2924);
and (n4011,n3322,n2947);
and (n4012,n3325,n2955);
and (n4013,n4014,n2964);
wire s0n4014,s1n4014,notn4014;
or (n4014,s0n4014,s1n4014);
not(notn4014,n2921);
and (s0n4014,notn4014,n2214);
and (s1n4014,n2921,n4015);
or (n4016,1'b0,n4017,n4026,n4032,n4041);
and (n4017,n4018,n2710);
or (n4018,1'b0,n4019,n4023,n4024,n4025);
and (n4019,n4020,n2924);
wire s0n4020,s1n4020,notn4020;
or (n4020,s0n4020,s1n4020);
not(notn4020,n2921);
and (s0n4020,notn4020,n4021);
and (s1n4020,n2921,n4022);
and (n4023,n3331,n2947);
and (n4024,n3260,n2955);
and (n4025,n3264,n2964);
and (n4026,n4027,n2722);
or (n4027,1'b0,n4028,n4029,n4030,n4031);
and (n4028,n3268,n2924);
and (n4029,n3272,n2947);
and (n4030,n3278,n2955);
and (n4031,n3282,n2964);
and (n4032,n4033,n2734);
or (n4033,1'b0,n4034,n4038,n4039,n4040);
and (n4034,n4035,n2924);
wire s0n4035,s1n4035,notn4035;
or (n4035,s0n4035,s1n4035);
not(notn4035,n2921);
and (s0n4035,notn4035,n4036);
and (s1n4035,n2921,n4037);
and (n4038,n3346,n2947);
and (n4039,n3296,n2955);
and (n4040,n3300,n2964);
and (n4041,n4042,n2744);
or (n4042,1'b0,n4043,n4044,n4045,n4046);
and (n4043,n3304,n2924);
and (n4044,n3308,n2947);
and (n4045,n3314,n2955);
and (n4046,n3318,n2964);
and (n4047,n4016,n4048);
or (n4048,n4049,n4114,n4313);
and (n4049,n4050,n4081);
or (n4050,1'b0,n4051,n4058,n4067,n4073);
not (n4051,n4052);
nand (n4052,n4053,n2710);
or (n4053,1'b0,n4054,n4055,n4056,n4057);
and (n4054,n3369,n2924);
and (n4055,n3373,n2947);
and (n4056,n3377,n2955);
and (n4057,n3383,n2964);
and (n4058,n4059,n2722);
or (n4059,1'b0,n4060,n4061,n4062,n4063);
and (n4060,n3387,n2924);
and (n4061,n3391,n2947);
and (n4062,n3395,n2955);
and (n4063,n4064,n2964);
wire s0n4064,s1n4064,notn4064;
or (n4064,s0n4064,s1n4064);
not(notn4064,n2921);
and (s0n4064,notn4064,n4065);
and (s1n4064,n2921,n4066);
and (n4067,n4068,n2734);
or (n4068,1'b0,n4069,n4070,n4071,n4072);
and (n4069,n3405,n2924);
and (n4070,n3409,n2947);
and (n4071,n3413,n2955);
and (n4072,n3419,n2964);
and (n4073,n4074,n2744);
or (n4074,1'b0,n4075,n4076,n4077,n4078);
and (n4075,n3423,n2924);
and (n4076,n3427,n2947);
and (n4077,n3430,n2955);
and (n4078,n4079,n2964);
wire s0n4079,s1n4079,notn4079;
or (n4079,s0n4079,s1n4079);
not(notn4079,n2921);
and (s0n4079,notn4079,n2230);
and (s1n4079,n2921,n4080);
or (n4081,1'b0,n4082,n4091,n4098,n4107);
and (n4082,n4083,n2710);
or (n4083,1'b0,n4084,n4088,n4089,n4090);
and (n4084,n4085,n2924);
wire s0n4085,s1n4085,notn4085;
or (n4085,s0n4085,s1n4085);
not(notn4085,n2921);
and (s0n4085,notn4085,n4086);
and (s1n4085,n2921,n4087);
and (n4088,n3436,n2947);
and (n4089,n3365,n2955);
and (n4090,n3369,n2964);
not (n4091,n4092);
nand (n4092,n4093,n2722);
or (n4093,1'b0,n4094,n4095,n4096,n4097);
and (n4094,n3373,n2924);
and (n4095,n3377,n2947);
and (n4096,n3383,n2955);
and (n4097,n3387,n2964);
and (n4098,n4099,n2734);
or (n4099,1'b0,n4100,n4104,n4105,n4106);
and (n4100,n4101,n2924);
wire s0n4101,s1n4101,notn4101;
or (n4101,s0n4101,s1n4101);
not(notn4101,n2921);
and (s0n4101,notn4101,n4102);
and (s1n4101,n2921,n4103);
and (n4104,n3451,n2947);
and (n4105,n3401,n2955);
and (n4106,n3405,n2964);
not (n4107,n4108);
nand (n4108,n4109,n2744);
or (n4109,1'b0,n4110,n4111,n4112,n4113);
and (n4110,n3409,n2924);
and (n4111,n3413,n2947);
and (n4112,n3419,n2955);
and (n4113,n3423,n2964);
and (n4114,n4081,n4115);
or (n4115,n4116,n4180,n4312);
and (n4116,n4117,n4149);
or (n4117,1'b0,n4118,n4125,n4134,n4141);
not (n4118,n4119);
nand (n4119,n4120,n2710);
or (n4120,1'b0,n4121,n4122,n4123,n4124);
and (n4121,n3474,n2924);
and (n4122,n3478,n2947);
and (n4123,n3482,n2955);
and (n4124,n3488,n2964);
and (n4125,n4126,n2722);
or (n4126,1'b0,n4127,n4128,n4129,n4130);
and (n4127,n3492,n2924);
and (n4128,n3496,n2947);
and (n4129,n3500,n2955);
and (n4130,n4131,n2964);
wire s0n4131,s1n4131,notn4131;
or (n4131,s0n4131,s1n4131);
not(notn4131,n2921);
and (s0n4131,notn4131,n4132);
and (s1n4131,n2921,n4133);
not (n4134,n4135);
nand (n4135,n4136,n2734);
or (n4136,1'b0,n4137,n4138,n4139,n4140);
and (n4137,n3510,n2924);
and (n4138,n3514,n2947);
and (n4139,n3518,n2955);
and (n4140,n3524,n2964);
and (n4141,n4142,n2744);
or (n4142,1'b0,n4143,n4144,n4145,n4146);
and (n4143,n3528,n2924);
and (n4144,n3532,n2947);
and (n4145,n3535,n2955);
and (n4146,n4147,n2964);
wire s0n4147,s1n4147,notn4147;
or (n4147,s0n4147,s1n4147);
not(notn4147,n2921);
and (s0n4147,notn4147,n2246);
and (s1n4147,n2921,n4148);
or (n4149,1'b0,n4150,n4159,n4165,n4174);
and (n4150,n4151,n2710);
or (n4151,1'b0,n4152,n4156,n4157,n4158);
and (n4152,n4153,n2924);
wire s0n4153,s1n4153,notn4153;
or (n4153,s0n4153,s1n4153);
not(notn4153,n2921);
and (s0n4153,notn4153,n4154);
and (s1n4153,n2921,n4155);
and (n4156,n3541,n2947);
and (n4157,n3470,n2955);
and (n4158,n3474,n2964);
and (n4159,n4160,n2722);
or (n4160,1'b0,n4161,n4162,n4163,n4164);
and (n4161,n3478,n2924);
and (n4162,n3482,n2947);
and (n4163,n3488,n2955);
and (n4164,n3492,n2964);
and (n4165,n4166,n2734);
or (n4166,1'b0,n4167,n4171,n4172,n4173);
and (n4167,n4168,n2924);
wire s0n4168,s1n4168,notn4168;
or (n4168,s0n4168,s1n4168);
not(notn4168,n2921);
and (s0n4168,notn4168,n4169);
and (s1n4168,n2921,n4170);
and (n4171,n3556,n2947);
and (n4172,n3506,n2955);
and (n4173,n3510,n2964);
and (n4174,n4175,n2744);
or (n4175,1'b0,n4176,n4177,n4178,n4179);
and (n4176,n3514,n2924);
and (n4177,n3518,n2947);
and (n4178,n3524,n2955);
and (n4179,n3528,n2964);
and (n4180,n4149,n4181);
or (n4181,n4182,n4244,n4311);
and (n4182,n4183,n4213);
or (n4183,1'b0,n4184,n4190,n4199,n4205);
and (n4184,n4185,n2710);
or (n4185,1'b0,n4186,n4187,n4188,n4189);
and (n4186,n3579,n2924);
and (n4187,n3583,n2947);
and (n4188,n3587,n2955);
and (n4189,n3593,n2964);
and (n4190,n4191,n2722);
or (n4191,1'b0,n4192,n4193,n4194,n4195);
and (n4192,n3597,n2924);
and (n4193,n3601,n2947);
and (n4194,n3605,n2955);
and (n4195,n4196,n2964);
wire s0n4196,s1n4196,notn4196;
or (n4196,s0n4196,s1n4196);
not(notn4196,n2921);
and (s0n4196,notn4196,n4197);
and (s1n4196,n2921,n4198);
and (n4199,n4200,n2734);
or (n4200,1'b0,n4201,n4202,n4203,n4204);
and (n4201,n3615,n2924);
and (n4202,n3619,n2947);
and (n4203,n3623,n2955);
and (n4204,n3629,n2964);
and (n4205,n4206,n2744);
or (n4206,1'b0,n4207,n4208,n4209,n4210);
and (n4207,n3633,n2924);
and (n4208,n3637,n2947);
and (n4209,n3640,n2955);
and (n4210,n4211,n2964);
wire s0n4211,s1n4211,notn4211;
or (n4211,s0n4211,s1n4211);
not(notn4211,n2921);
and (s0n4211,notn4211,n2262);
and (s1n4211,n2921,n4212);
or (n4213,1'b0,n4214,n4223,n4229,n4238);
and (n4214,n4215,n2710);
or (n4215,1'b0,n4216,n4220,n4221,n4222);
and (n4216,n4217,n2924);
wire s0n4217,s1n4217,notn4217;
or (n4217,s0n4217,s1n4217);
not(notn4217,n2921);
and (s0n4217,notn4217,n4218);
and (s1n4217,n2921,n4219);
and (n4220,n3646,n2947);
and (n4221,n3575,n2955);
and (n4222,n3579,n2964);
and (n4223,n4224,n2722);
or (n4224,1'b0,n4225,n4226,n4227,n4228);
and (n4225,n3583,n2924);
and (n4226,n3587,n2947);
and (n4227,n3593,n2955);
and (n4228,n3597,n2964);
and (n4229,n4230,n2734);
or (n4230,1'b0,n4231,n4235,n4236,n4237);
and (n4231,n4232,n2924);
wire s0n4232,s1n4232,notn4232;
or (n4232,s0n4232,s1n4232);
not(notn4232,n2921);
and (s0n4232,notn4232,n4233);
and (s1n4232,n2921,n4234);
and (n4235,n3661,n2947);
and (n4236,n3611,n2955);
and (n4237,n3615,n2964);
and (n4238,n4239,n2744);
or (n4239,1'b0,n4240,n4241,n4242,n4243);
and (n4240,n3619,n2924);
and (n4241,n3623,n2947);
and (n4242,n3629,n2955);
and (n4243,n3633,n2964);
and (n4244,n4213,n4245);
and (n4245,n4246,n4278);
or (n4246,1'b0,n4247,n4254,n4263,n4270);
not (n4247,n4248);
nand (n4248,n4249,n2710);
or (n4249,1'b0,n4250,n4251,n4252,n4253);
and (n4250,n3683,n2924);
and (n4251,n3687,n2947);
and (n4252,n3691,n2955);
and (n4253,n3697,n2964);
and (n4254,n4255,n2722);
or (n4255,1'b0,n4256,n4257,n4258,n4259);
and (n4256,n3701,n2924);
and (n4257,n3705,n2947);
and (n4258,n3709,n2955);
and (n4259,n4260,n2964);
wire s0n4260,s1n4260,notn4260;
or (n4260,s0n4260,s1n4260);
not(notn4260,n2921);
and (s0n4260,notn4260,n4261);
and (s1n4260,n2921,n4262);
not (n4263,n4264);
nand (n4264,n4265,n2734);
or (n4265,1'b0,n4266,n4267,n4268,n4269);
and (n4266,n3719,n2924);
and (n4267,n3723,n2947);
and (n4268,n3727,n2955);
and (n4269,n3733,n2964);
and (n4270,n4271,n2744);
or (n4271,1'b0,n4272,n4273,n4274,n4275);
and (n4272,n3737,n2924);
and (n4273,n3741,n2947);
and (n4274,n3744,n2955);
and (n4275,n4276,n2964);
wire s0n4276,s1n4276,notn4276;
or (n4276,s0n4276,s1n4276);
not(notn4276,n2921);
and (s0n4276,notn4276,n2277);
and (s1n4276,n2921,n4277);
or (n4278,1'b0,n4279,n4288,n4295,n4304);
and (n4279,n4280,n2710);
or (n4280,1'b0,n4281,n4285,n4286,n4287);
and (n4281,n4282,n2924);
wire s0n4282,s1n4282,notn4282;
or (n4282,s0n4282,s1n4282);
not(notn4282,n2921);
and (s0n4282,notn4282,n4283);
and (s1n4282,n2921,n4284);
and (n4285,n3750,n2947);
and (n4286,n3679,n2955);
and (n4287,n3683,n2964);
not (n4288,n4289);
nand (n4289,n4290,n2722);
or (n4290,1'b0,n4291,n4292,n4293,n4294);
and (n4291,n3687,n2924);
and (n4292,n3691,n2947);
and (n4293,n3697,n2955);
and (n4294,n3701,n2964);
and (n4295,n4296,n2734);
or (n4296,1'b0,n4297,n4301,n4302,n4303);
and (n4297,n4298,n2924);
wire s0n4298,s1n4298,notn4298;
or (n4298,s0n4298,s1n4298);
not(notn4298,n2921);
and (s0n4298,notn4298,n4299);
and (s1n4298,n2921,n4300);
and (n4301,n3765,n2947);
and (n4302,n3715,n2955);
and (n4303,n3719,n2964);
not (n4304,n4305);
nand (n4305,n4306,n2744);
or (n4306,1'b0,n4307,n4308,n4309,n4310);
and (n4307,n3723,n2924);
and (n4308,n3727,n2947);
and (n4309,n3733,n2955);
and (n4310,n3737,n2964);
and (n4311,n4183,n4245);
and (n4312,n4117,n4181);
and (n4313,n4050,n4115);
and (n4314,n3986,n4048);
and (n4315,n3922,n3984);
and (n4316,n3858,n3920);
and (n4317,n3794,n3856);
and (n4318,n3791,n4319);
or (n4319,n4320,n4326,n4368);
and (n4320,n4321,n4323);
xor (n4321,n4322,n3254);
xor (n4322,n3151,n3222);
not (n4323,n4324);
xor (n4324,n4325,n3856);
xor (n4325,n3794,n3824);
and (n4326,n4323,n4327);
or (n4327,n4328,n4334,n4367);
and (n4328,n4329,n4331);
xor (n4329,n4330,n3359);
xor (n4330,n3256,n3327);
not (n4331,n4332);
xor (n4332,n4333,n3920);
xor (n4333,n3858,n3888);
and (n4334,n4331,n4335);
or (n4335,n4336,n4342,n4366);
and (n4336,n4337,n4339);
xor (n4337,n4338,n3464);
xor (n4338,n3361,n3432);
not (n4339,n4340);
xor (n4340,n4341,n3984);
xor (n4341,n3922,n3952);
and (n4342,n4339,n4343);
or (n4343,n4344,n4350,n4365);
and (n4344,n4345,n4347);
xor (n4345,n4346,n3569);
xor (n4346,n3466,n3537);
not (n4347,n4348);
xor (n4348,n4349,n4048);
xor (n4349,n3986,n4016);
and (n4350,n4347,n4351);
or (n4351,n4352,n4358,n4364);
and (n4352,n4353,n4355);
xor (n4353,n4354,n3674);
xor (n4354,n3571,n3642);
not (n4355,n4356);
xor (n4356,n4357,n4115);
xor (n4357,n4050,n4081);
and (n4358,n4355,n4359);
and (n4359,n4360,n4361);
xor (n4360,n3675,n3746);
not (n4361,n4362);
xor (n4362,n4363,n4181);
xor (n4363,n4117,n4149);
and (n4364,n4353,n4359);
and (n4365,n4345,n4351);
and (n4366,n4337,n4343);
and (n4367,n4329,n4335);
and (n4368,n4321,n4327);
and (n4369,n3789,n4319);
and (n4370,n4371,n4372);
xnor (n4371,n2913,n3784);
and (n4372,n4373,n4374);
xnor (n4373,n3785,n3787);
and (n4374,n4375,n4377);
xor (n4375,n4376,n4319);
xor (n4376,n3789,n3791);
and (n4377,n4378,n4380);
xor (n4378,n4379,n4327);
xor (n4379,n4321,n4323);
and (n4380,n4381,n4383);
xor (n4381,n4382,n4335);
xor (n4382,n4329,n4331);
and (n4383,n4384,n4386);
xor (n4384,n4385,n4343);
xor (n4385,n4337,n4339);
and (n4386,n4387,n4389);
xor (n4387,n4388,n4351);
xor (n4388,n4345,n4347);
and (n4389,n4390,n4392);
xor (n4390,n4391,n4359);
xor (n4391,n4353,n4355);
and (n4392,n4393,n4394);
xor (n4393,n4360,n4361);
and (n4394,n4395,n4398);
not (n4395,n4396);
xor (n4396,n4397,n4245);
xor (n4397,n4183,n4213);
not (n4398,n4399);
xor (n4399,n4246,n4278);
and (n4400,n2910,n4401);
and (n4401,n4402,n4403);
xor (n4402,n4371,n4372);
and (n4403,n4404,n4405);
xor (n4404,n4373,n4374);
or (n4405,n4406,n4787,n4839);
and (n4406,n4407,n4786);
or (n4407,n4408,n4453,n4785);
and (n4408,n4409,n4430);
or (n4409,1'b0,n4410,n4411,n4420,n4422);
and (n4410,n3835,n2710);
and (n4411,n4412,n2722);
or (n4412,1'b0,n4413,n4414,n4415,n4416);
and (n4413,n2979,n2924);
and (n4414,n2982,n2947);
and (n4415,n3807,n2955);
and (n4416,n4417,n2964);
wire s0n4417,s1n4417,notn4417;
or (n4417,s0n4417,s1n4417);
not(notn4417,n2921);
and (s0n4417,notn4417,n4418);
and (s1n4417,n2921,n4419);
not (n4420,n4421);
nand (n4421,n3850,n2734);
and (n4422,n4423,n2744);
or (n4423,1'b0,n4424,n4425,n4426,n4427);
and (n4424,n3007,n2924);
and (n4425,n3010,n2947);
and (n4426,n3822,n2955);
and (n4427,n4428,n2964);
wire s0n4428,s1n4428,notn4428;
or (n4428,s0n4428,s1n4428);
not(notn4428,n2921);
and (s0n4428,notn4428,n1829);
and (s1n4428,n2921,n4429);
or (n4430,1'b0,n4431,n4440,n4442,n4451);
and (n4431,n4432,n2710);
or (n4432,1'b0,n4433,n4437,n4438,n4439);
and (n4433,n4434,n2924);
wire s0n4434,s1n4434,notn4434;
or (n4434,s0n4434,s1n4434);
not(notn4434,n2921);
and (s0n4434,notn4434,n4435);
and (s1n4434,n2921,n4436);
and (n4437,n3828,n2947);
and (n4438,n3016,n2955);
and (n4439,n2919,n2964);
not (n4440,n4441);
nand (n4441,n3796,n2722);
and (n4442,n4443,n2734);
or (n4443,1'b0,n4444,n4448,n4449,n4450);
and (n4444,n4445,n2924);
wire s0n4445,s1n4445,notn4445;
or (n4445,s0n4445,s1n4445);
not(notn4445,n2921);
and (s0n4445,notn4445,n4446);
and (s1n4445,n2921,n4447);
and (n4448,n3843,n2947);
and (n4449,n3031,n2955);
and (n4450,n2987,n2964);
not (n4451,n4452);
nand (n4452,n3811,n2744);
and (n4453,n4430,n4454);
or (n4454,n4455,n4500,n4784);
and (n4455,n4456,n4477);
or (n4456,1'b0,n4457,n4458,n4467,n4469);
and (n4457,n3899,n2710);
and (n4458,n4459,n2722);
or (n4459,1'b0,n4460,n4461,n4462,n4463);
and (n4460,n3076,n2924);
and (n4461,n3080,n2947);
and (n4462,n3871,n2955);
and (n4463,n4464,n2964);
wire s0n4464,s1n4464,notn4464;
or (n4464,s0n4464,s1n4464);
not(notn4464,n2921);
and (s0n4464,notn4464,n4465);
and (s1n4464,n2921,n4466);
not (n4467,n4468);
nand (n4468,n3914,n2734);
and (n4469,n4470,n2744);
or (n4470,1'b0,n4471,n4472,n4473,n4474);
and (n4471,n3112,n2924);
and (n4472,n3115,n2947);
and (n4473,n3886,n2955);
and (n4474,n4475,n2964);
wire s0n4475,s1n4475,notn4475;
or (n4475,s0n4475,s1n4475);
not(notn4475,n2921);
and (s0n4475,notn4475,n1846);
and (s1n4475,n2921,n4476);
or (n4477,1'b0,n4478,n4487,n4489,n4498);
and (n4478,n4479,n2710);
or (n4479,1'b0,n4480,n4484,n4485,n4486);
and (n4480,n4481,n2924);
wire s0n4481,s1n4481,notn4481;
or (n4481,s0n4481,s1n4481);
not(notn4481,n2921);
and (s0n4481,notn4481,n4482);
and (s1n4481,n2921,n4483);
and (n4484,n3892,n2947);
and (n4485,n3121,n2955);
and (n4486,n3050,n2964);
not (n4487,n4488);
nand (n4488,n3860,n2722);
and (n4489,n4490,n2734);
or (n4490,1'b0,n4491,n4495,n4496,n4497);
and (n4491,n4492,n2924);
wire s0n4492,s1n4492,notn4492;
or (n4492,s0n4492,s1n4492);
not(notn4492,n2921);
and (s0n4492,notn4492,n4493);
and (s1n4492,n2921,n4494);
and (n4495,n3907,n2947);
and (n4496,n3136,n2955);
and (n4497,n3086,n2964);
not (n4498,n4499);
nand (n4499,n3875,n2744);
and (n4500,n4477,n4501);
or (n4501,n4502,n4547,n4783);
and (n4502,n4503,n4524);
or (n4503,1'b0,n4504,n4505,n4514,n4516);
and (n4504,n3963,n2710);
and (n4505,n4506,n2722);
or (n4506,1'b0,n4507,n4508,n4509,n4510);
and (n4507,n3181,n2924);
and (n4508,n3185,n2947);
and (n4509,n3935,n2955);
and (n4510,n4511,n2964);
wire s0n4511,s1n4511,notn4511;
or (n4511,s0n4511,s1n4511);
not(notn4511,n2921);
and (s0n4511,notn4511,n4512);
and (s1n4511,n2921,n4513);
not (n4514,n4515);
nand (n4515,n3978,n2734);
and (n4516,n4517,n2744);
or (n4517,1'b0,n4518,n4519,n4520,n4521);
and (n4518,n3217,n2924);
and (n4519,n3220,n2947);
and (n4520,n3950,n2955);
and (n4521,n4522,n2964);
wire s0n4522,s1n4522,notn4522;
or (n4522,s0n4522,s1n4522);
not(notn4522,n2921);
and (s0n4522,notn4522,n1863);
and (s1n4522,n2921,n4523);
or (n4524,1'b0,n4525,n4534,n4536,n4545);
and (n4525,n4526,n2710);
or (n4526,1'b0,n4527,n4531,n4532,n4533);
and (n4527,n4528,n2924);
wire s0n4528,s1n4528,notn4528;
or (n4528,s0n4528,s1n4528);
not(notn4528,n2921);
and (s0n4528,notn4528,n4529);
and (s1n4528,n2921,n4530);
and (n4531,n3956,n2947);
and (n4532,n3226,n2955);
and (n4533,n3155,n2964);
not (n4534,n4535);
nand (n4535,n3924,n2722);
and (n4536,n4537,n2734);
or (n4537,1'b0,n4538,n4542,n4543,n4544);
and (n4538,n4539,n2924);
wire s0n4539,s1n4539,notn4539;
or (n4539,s0n4539,s1n4539);
not(notn4539,n2921);
and (s0n4539,notn4539,n4540);
and (s1n4539,n2921,n4541);
and (n4542,n3971,n2947);
and (n4543,n3241,n2955);
and (n4544,n3191,n2964);
not (n4545,n4546);
nand (n4546,n3939,n2744);
and (n4547,n4524,n4548);
or (n4548,n4549,n4594,n4782);
and (n4549,n4550,n4571);
or (n4550,1'b0,n4551,n4552,n4561,n4563);
and (n4551,n4027,n2710);
and (n4552,n4553,n2722);
or (n4553,1'b0,n4554,n4555,n4556,n4557);
and (n4554,n3286,n2924);
and (n4555,n3290,n2947);
and (n4556,n3999,n2955);
and (n4557,n4558,n2964);
wire s0n4558,s1n4558,notn4558;
or (n4558,s0n4558,s1n4558);
not(notn4558,n2921);
and (s0n4558,notn4558,n4559);
and (s1n4558,n2921,n4560);
not (n4561,n4562);
nand (n4562,n4042,n2734);
and (n4563,n4564,n2744);
or (n4564,1'b0,n4565,n4566,n4567,n4568);
and (n4565,n3322,n2924);
and (n4566,n3325,n2947);
and (n4567,n4014,n2955);
and (n4568,n4569,n2964);
wire s0n4569,s1n4569,notn4569;
or (n4569,s0n4569,s1n4569);
not(notn4569,n2921);
and (s0n4569,notn4569,n1888);
and (s1n4569,n2921,n4570);
or (n4571,1'b0,n4572,n4581,n4583,n4592);
and (n4572,n4573,n2710);
or (n4573,1'b0,n4574,n4578,n4579,n4580);
and (n4574,n4575,n2924);
wire s0n4575,s1n4575,notn4575;
or (n4575,s0n4575,s1n4575);
not(notn4575,n2921);
and (s0n4575,notn4575,n4576);
and (s1n4575,n2921,n4577);
and (n4578,n4020,n2947);
and (n4579,n3331,n2955);
and (n4580,n3260,n2964);
not (n4581,n4582);
nand (n4582,n3988,n2722);
and (n4583,n4584,n2734);
or (n4584,1'b0,n4585,n4589,n4590,n4591);
and (n4585,n4586,n2924);
wire s0n4586,s1n4586,notn4586;
or (n4586,s0n4586,s1n4586);
not(notn4586,n2921);
and (s0n4586,notn4586,n4587);
and (s1n4586,n2921,n4588);
and (n4589,n4035,n2947);
and (n4590,n3346,n2955);
and (n4591,n3296,n2964);
not (n4592,n4593);
nand (n4593,n4003,n2744);
and (n4594,n4571,n4595);
or (n4595,n4596,n4639,n4781);
and (n4596,n4597,n4618);
or (n4597,1'b0,n4598,n4599,n4608,n4610);
and (n4598,n4093,n2710);
and (n4599,n4600,n2722);
or (n4600,1'b0,n4601,n4602,n4603,n4604);
and (n4601,n3391,n2924);
and (n4602,n3395,n2947);
and (n4603,n4064,n2955);
and (n4604,n4605,n2964);
wire s0n4605,s1n4605,notn4605;
or (n4605,s0n4605,s1n4605);
not(notn4605,n2921);
and (s0n4605,notn4605,n4606);
and (s1n4605,n2921,n4607);
not (n4608,n4609);
nand (n4609,n4109,n2734);
and (n4610,n4611,n2744);
or (n4611,1'b0,n4612,n4613,n4614,n4615);
and (n4612,n3427,n2924);
and (n4613,n3430,n2947);
and (n4614,n4079,n2955);
and (n4615,n4616,n2964);
wire s0n4616,s1n4616,notn4616;
or (n4616,s0n4616,s1n4616);
not(notn4616,n2921);
and (s0n4616,notn4616,n1915);
and (s1n4616,n2921,n4617);
or (n4618,1'b0,n4619,n4628,n4629,n4638);
and (n4619,n4620,n2710);
or (n4620,1'b0,n4621,n4625,n4626,n4627);
and (n4621,n4622,n2924);
wire s0n4622,s1n4622,notn4622;
or (n4622,s0n4622,s1n4622);
not(notn4622,n2921);
and (s0n4622,notn4622,n4623);
and (s1n4622,n2921,n4624);
and (n4625,n4085,n2947);
and (n4626,n3436,n2955);
and (n4627,n3365,n2964);
and (n4628,n4053,n2722);
and (n4629,n4630,n2734);
or (n4630,1'b0,n4631,n4635,n4636,n4637);
and (n4631,n4632,n2924);
wire s0n4632,s1n4632,notn4632;
or (n4632,s0n4632,s1n4632);
not(notn4632,n2921);
and (s0n4632,notn4632,n4633);
and (s1n4632,n2921,n4634);
and (n4635,n4101,n2947);
and (n4636,n3451,n2955);
and (n4637,n3401,n2964);
and (n4638,n4068,n2744);
and (n4639,n4618,n4640);
or (n4640,n4641,n4686,n4780);
and (n4641,n4642,n4663);
or (n4642,1'b0,n4643,n4644,n4653,n4655);
and (n4643,n4160,n2710);
and (n4644,n4645,n2722);
or (n4645,1'b0,n4646,n4647,n4648,n4649);
and (n4646,n3496,n2924);
and (n4647,n3500,n2947);
and (n4648,n4131,n2955);
and (n4649,n4650,n2964);
wire s0n4650,s1n4650,notn4650;
or (n4650,s0n4650,s1n4650);
not(notn4650,n2921);
and (s0n4650,notn4650,n4651);
and (s1n4650,n2921,n4652);
not (n4653,n4654);
nand (n4654,n4175,n2734);
and (n4655,n4656,n2744);
or (n4656,1'b0,n4657,n4658,n4659,n4660);
and (n4657,n3532,n2924);
and (n4658,n3535,n2947);
and (n4659,n4147,n2955);
and (n4660,n4661,n2964);
wire s0n4661,s1n4661,notn4661;
or (n4661,s0n4661,s1n4661);
not(notn4661,n2921);
and (s0n4661,notn4661,n1941);
and (s1n4661,n2921,n4662);
or (n4663,1'b0,n4664,n4673,n4675,n4684);
and (n4664,n4665,n2710);
or (n4665,1'b0,n4666,n4670,n4671,n4672);
and (n4666,n4667,n2924);
wire s0n4667,s1n4667,notn4667;
or (n4667,s0n4667,s1n4667);
not(notn4667,n2921);
and (s0n4667,notn4667,n4668);
and (s1n4667,n2921,n4669);
and (n4670,n4153,n2947);
and (n4671,n3541,n2955);
and (n4672,n3470,n2964);
not (n4673,n4674);
nand (n4674,n4120,n2722);
and (n4675,n4676,n2734);
or (n4676,1'b0,n4677,n4681,n4682,n4683);
and (n4677,n4678,n2924);
wire s0n4678,s1n4678,notn4678;
or (n4678,s0n4678,s1n4678);
not(notn4678,n2921);
and (s0n4678,notn4678,n4679);
and (s1n4678,n2921,n4680);
and (n4681,n4168,n2947);
and (n4682,n3556,n2955);
and (n4683,n3506,n2964);
not (n4684,n4685);
nand (n4685,n4136,n2744);
and (n4686,n4663,n4687);
or (n4687,n4688,n4733,n4779);
and (n4688,n4689,n4710);
or (n4689,1'b0,n4690,n4691,n4700,n4702);
and (n4690,n4224,n2710);
and (n4691,n4692,n2722);
or (n4692,1'b0,n4693,n4694,n4695,n4696);
and (n4693,n3601,n2924);
and (n4694,n3605,n2947);
and (n4695,n4196,n2955);
and (n4696,n4697,n2964);
wire s0n4697,s1n4697,notn4697;
or (n4697,s0n4697,s1n4697);
not(notn4697,n2921);
and (s0n4697,notn4697,n4698);
and (s1n4697,n2921,n4699);
not (n4700,n4701);
nand (n4701,n4239,n2734);
and (n4702,n4703,n2744);
or (n4703,1'b0,n4704,n4705,n4706,n4707);
and (n4704,n3637,n2924);
and (n4705,n3640,n2947);
and (n4706,n4211,n2955);
and (n4707,n4708,n2964);
wire s0n4708,s1n4708,notn4708;
or (n4708,s0n4708,s1n4708);
not(notn4708,n2921);
and (s0n4708,notn4708,n1970);
and (s1n4708,n2921,n4709);
or (n4710,1'b0,n4711,n4720,n4722,n4731);
and (n4711,n4712,n2710);
or (n4712,1'b0,n4713,n4717,n4718,n4719);
and (n4713,n4714,n2924);
wire s0n4714,s1n4714,notn4714;
or (n4714,s0n4714,s1n4714);
not(notn4714,n2921);
and (s0n4714,notn4714,n4715);
and (s1n4714,n2921,n4716);
and (n4717,n4217,n2947);
and (n4718,n3646,n2955);
and (n4719,n3575,n2964);
not (n4720,n4721);
nand (n4721,n4185,n2722);
and (n4722,n4723,n2734);
or (n4723,1'b0,n4724,n4728,n4729,n4730);
and (n4724,n4725,n2924);
wire s0n4725,s1n4725,notn4725;
or (n4725,s0n4725,s1n4725);
not(notn4725,n2921);
and (s0n4725,notn4725,n4726);
and (s1n4725,n2921,n4727);
and (n4728,n4232,n2947);
and (n4729,n3661,n2955);
and (n4730,n3611,n2964);
not (n4731,n4732);
nand (n4732,n4200,n2744);
and (n4733,n4710,n4734);
and (n4734,n4735,n4756);
or (n4735,1'b0,n4736,n4737,n4746,n4748);
and (n4736,n4290,n2710);
and (n4737,n4738,n2722);
or (n4738,1'b0,n4739,n4740,n4741,n4742);
and (n4739,n3705,n2924);
and (n4740,n3709,n2947);
and (n4741,n4260,n2955);
and (n4742,n4743,n2964);
wire s0n4743,s1n4743,notn4743;
or (n4743,s0n4743,s1n4743);
not(notn4743,n2921);
and (s0n4743,notn4743,n4744);
and (s1n4743,n2921,n4745);
not (n4746,n4747);
nand (n4747,n4306,n2734);
and (n4748,n4749,n2744);
or (n4749,1'b0,n4750,n4751,n4752,n4753);
and (n4750,n3741,n2924);
and (n4751,n3744,n2947);
and (n4752,n4276,n2955);
and (n4753,n4754,n2964);
wire s0n4754,s1n4754,notn4754;
or (n4754,s0n4754,s1n4754);
not(notn4754,n2921);
and (s0n4754,notn4754,n1989);
and (s1n4754,n2921,n4755);
or (n4756,1'b0,n4757,n4766,n4768,n4777);
and (n4757,n4758,n2710);
or (n4758,1'b0,n4759,n4763,n4764,n4765);
and (n4759,n4760,n2924);
wire s0n4760,s1n4760,notn4760;
or (n4760,s0n4760,s1n4760);
not(notn4760,n2921);
and (s0n4760,notn4760,n4761);
and (s1n4760,n2921,n4762);
and (n4763,n4282,n2947);
and (n4764,n3750,n2955);
and (n4765,n3679,n2964);
not (n4766,n4767);
nand (n4767,n4249,n2722);
and (n4768,n4769,n2734);
or (n4769,1'b0,n4770,n4774,n4775,n4776);
and (n4770,n4771,n2924);
wire s0n4771,s1n4771,notn4771;
or (n4771,s0n4771,s1n4771);
not(notn4771,n2921);
and (s0n4771,notn4771,n4772);
and (s1n4771,n2921,n4773);
and (n4774,n4298,n2947);
and (n4775,n3765,n2955);
and (n4776,n3715,n2964);
not (n4777,n4778);
nand (n4778,n4265,n2744);
and (n4779,n4689,n4734);
and (n4780,n4642,n4687);
and (n4781,n4597,n4640);
and (n4782,n4550,n4595);
and (n4783,n4503,n4548);
and (n4784,n4456,n4501);
and (n4785,n4409,n4454);
xor (n4786,n4375,n4377);
and (n4787,n4786,n4788);
or (n4788,n4789,n4793,n4838);
and (n4789,n4790,n4792);
xor (n4790,n4791,n4454);
xor (n4791,n4409,n4430);
xor (n4792,n4378,n4380);
and (n4793,n4792,n4794);
or (n4794,n4795,n4799,n4837);
and (n4795,n4796,n4798);
xor (n4796,n4797,n4501);
xor (n4797,n4456,n4477);
xor (n4798,n4381,n4383);
and (n4799,n4798,n4800);
or (n4800,n4801,n4805,n4836);
and (n4801,n4802,n4804);
xor (n4802,n4803,n4548);
xor (n4803,n4503,n4524);
xor (n4804,n4384,n4386);
and (n4805,n4804,n4806);
or (n4806,n4807,n4811,n4835);
and (n4807,n4808,n4810);
xor (n4808,n4809,n4595);
xor (n4809,n4550,n4571);
xor (n4810,n4387,n4389);
and (n4811,n4810,n4812);
or (n4812,n4813,n4817,n4834);
and (n4813,n4814,n4816);
xor (n4814,n4815,n4640);
xor (n4815,n4597,n4618);
xor (n4816,n4390,n4392);
and (n4817,n4816,n4818);
or (n4818,n4819,n4823,n4833);
and (n4819,n4820,n4822);
xor (n4820,n4821,n4687);
xor (n4821,n4642,n4663);
xor (n4822,n4393,n4394);
and (n4823,n4822,n4824);
or (n4824,n4825,n4829,n4832);
and (n4825,n4826,n4828);
xor (n4826,n4827,n4734);
xor (n4827,n4689,n4710);
xor (n4828,n4395,n4398);
and (n4829,n4828,n4830);
and (n4830,n4831,n4399);
xor (n4831,n4735,n4756);
and (n4832,n4826,n4830);
and (n4833,n4820,n4824);
and (n4834,n4814,n4818);
and (n4835,n4808,n4812);
and (n4836,n4802,n4806);
and (n4837,n4796,n4800);
and (n4838,n4790,n4794);
and (n4839,n4407,n4788);
or (n4840,n4841,n4842,n4892);
xor (n4841,n2910,n4401);
and (n4842,n4404,n4843);
or (n4843,n4844,n4846,n4891);
and (n4844,n4845,n4786);
xor (n4845,n4402,n4403);
and (n4846,n4786,n4847);
or (n4847,n4848,n4850,n4890);
and (n4848,n4849,n4792);
xor (n4849,n4404,n4405);
and (n4850,n4792,n4851);
or (n4851,n4852,n4855,n4889);
and (n4852,n4853,n4798);
xor (n4853,n4854,n4788);
xor (n4854,n4407,n4786);
and (n4855,n4798,n4856);
or (n4856,n4857,n4860,n4888);
and (n4857,n4858,n4804);
xor (n4858,n4859,n4794);
xor (n4859,n4790,n4792);
and (n4860,n4804,n4861);
or (n4861,n4862,n4865,n4887);
and (n4862,n4863,n4810);
xor (n4863,n4864,n4800);
xor (n4864,n4796,n4798);
and (n4865,n4810,n4866);
or (n4866,n4867,n4870,n4886);
and (n4867,n4868,n4816);
xor (n4868,n4869,n4806);
xor (n4869,n4802,n4804);
and (n4870,n4816,n4871);
or (n4871,n4872,n4875,n4885);
and (n4872,n4873,n4822);
xor (n4873,n4874,n4812);
xor (n4874,n4808,n4810);
and (n4875,n4822,n4876);
or (n4876,n4877,n4880,n4884);
and (n4877,n4878,n4828);
xor (n4878,n4879,n4818);
xor (n4879,n4814,n4816);
and (n4880,n4828,n4881);
and (n4881,n4882,n4399);
xor (n4882,n4883,n4824);
xor (n4883,n4820,n4822);
and (n4884,n4878,n4881);
and (n4885,n4873,n4876);
and (n4886,n4868,n4871);
and (n4887,n4863,n4866);
and (n4888,n4858,n4861);
and (n4889,n4853,n4856);
and (n4890,n4849,n4851);
and (n4891,n4845,n4847);
and (n4892,n4841,n4843);
and (n4893,n4894,n4896);
xor (n4894,n4895,n4843);
xor (n4895,n4841,n4404);
and (n4896,n4897,n4899);
xor (n4897,n4898,n4847);
xor (n4898,n4845,n4786);
and (n4899,n4900,n4902);
xor (n4900,n4901,n4851);
xor (n4901,n4849,n4792);
and (n4902,n4903,n4905);
xor (n4903,n4904,n4856);
xor (n4904,n4853,n4798);
and (n4905,n4906,n4908);
xor (n4906,n4907,n4861);
xor (n4907,n4858,n4804);
and (n4908,n4909,n4911);
xor (n4909,n4910,n4866);
xor (n4910,n4863,n4810);
and (n4911,n4912,n4914);
xor (n4912,n4913,n4871);
xor (n4913,n4868,n4816);
xor (n4914,n4915,n4876);
xor (n4915,n4873,n4822);
and (n4916,n4917,n4927);
and (n4917,n4918,n4926);
and (n4918,n4919,n4925);
and (n4919,n4920,n4924);
and (n4920,n4921,n4923);
and (n4921,n2696,n4922);
not (n4922,n2748);
not (n4923,n2900);
not (n4924,n2942);
not (n4925,n2901);
or (n4926,n2887,n2792,n2818,n2844);
nand (n4927,n2749,n2792,n2890,n2888);
wire s0n4928,s1n4928,notn4928;
or (n4928,s0n4928,s1n4928);
not(notn4928,n4916);
and (s0n4928,notn4928,1'b0);
and (s1n4928,n4916,n4929);
xor (n4929,n4930,n4932);
xor (n4930,n4400,n4931);
and (n4931,n4402,n4840);
and (n4932,n2907,n4893);
wire s0n4933,s1n4933,notn4933;
or (n4933,s0n4933,s1n4933);
not(notn4933,n4916);
and (s0n4933,notn4933,1'b0);
and (s1n4933,n4916,n4934);
xor (n4934,n4935,n4937);
xor (n4935,n4400,n4936);
and (n4936,n2910,n4931);
and (n4937,n4930,n4932);
or (n4938,n4939,n2923);
or (n4939,n4940,n2922);
or (n4940,n2937,n2938);
or (n4941,1'b0,n4942,n4960,n4975,n4990);
and (n4942,n4943,n2710);
or (n4943,1'b0,n4944,n4951,n4957);
and (n4944,n4945,n4950);
or (n4945,1'b0,n4946,n4947,n4948,n4949);
and (n4946,n2920,n549);
and (n4947,n2946,n560);
and (n4948,n2954,n564);
and (n4949,n2963,n566);
not (n4950,n4927);
and (n4951,n4952,n2936);
or (n4952,1'b0,n4953,n4954,n4955,n4956);
and (n4953,n3017,n549);
and (n4954,n2703,n560);
and (n4955,n2705,n564);
and (n4956,n2707,n566);
and (n4957,n2701,n4958);
or (n4958,n2934,n4959);
not (n4959,n4926);
and (n4960,n4961,n2722);
or (n4961,1'b0,n4962,n4968,n4974);
and (n4962,n4963,n4950);
or (n4963,1'b0,n4964,n4965,n4966,n4967);
and (n4964,n2974,n549);
and (n4965,n2977,n560);
and (n4966,n2980,n564);
and (n4967,n2983,n566);
and (n4968,n4969,n2936);
or (n4969,1'b0,n4970,n4971,n4972,n4973);
and (n4970,n2709,n549);
and (n4971,n2715,n560);
and (n4972,n2717,n564);
and (n4973,n2719,n566);
and (n4974,n2713,n4958);
and (n4975,n4976,n2734);
or (n4976,1'b0,n4977,n4983,n4989);
and (n4977,n4978,n4950);
or (n4978,1'b0,n4979,n4980,n4981,n4982);
and (n4979,n2988,n549);
and (n4980,n2991,n560);
and (n4981,n2994,n564);
and (n4982,n2997,n566);
and (n4983,n4984,n2936);
or (n4984,1'b0,n4985,n4986,n4987,n4988);
and (n4985,n3032,n549);
and (n4986,n2727,n560);
and (n4987,n2729,n564);
and (n4988,n2731,n566);
and (n4989,n2725,n4958);
and (n4990,n4991,n2744);
or (n4991,1'b0,n4992,n4998,n5004);
and (n4992,n4993,n4950);
or (n4993,1'b0,n4994,n4995,n4996,n4997);
and (n4994,n3002,n549);
and (n4995,n3005,n560);
and (n4996,n3008,n564);
and (n4997,n3011,n566);
and (n4998,n4999,n2936);
or (n4999,1'b0,n5000,n5001,n5002,n5003);
and (n5000,n2733,n549);
and (n5001,n2739,n560);
and (n5002,n2741,n564);
and (n5003,n2164,n566);
and (n5004,n2737,n4958);
or (n5005,1'b0,n5006,n8043,n8045,n8048);
and (n5006,n5007,n2885);
wire s0n5007,s1n5007,notn5007;
or (n5007,s0n5007,s1n5007);
not(notn5007,n2883);
and (s0n5007,notn5007,1'b0);
and (s1n5007,n2883,n5008);
wire s0n5008,s1n5008,notn5008;
or (n5008,s0n5008,s1n5008);
not(notn5008,n8032);
and (s0n5008,notn5008,n5009);
and (s1n5008,n8032,1'b0);
wire s0n5009,s1n5009,notn5009;
or (n5009,s0n5009,s1n5009);
not(notn5009,n8017);
and (s0n5009,notn5009,n5010);
and (s1n5009,n8017,1'b1);
wire s0n5010,s1n5010,notn5010;
or (n5010,s0n5010,s1n5010);
not(notn5010,n5021);
and (s0n5010,notn5010,n5011);
and (s1n5010,n5021,n7777);
wire s0n5011,s1n5011,notn5011;
or (n5011,s0n5011,s1n5011);
not(notn5011,n5021);
and (s0n5011,notn5011,n5012);
and (s1n5011,n5021,n7774);
xor (n5012,n5013,n7751);
xor (n5013,n5014,n7694);
xor (n5014,n5015,n7625);
xor (n5015,n5016,n7615);
xor (n5016,n5017,n6069);
xor (n5017,n5018,n5031);
xor (n5018,n5019,n5029);
wire s0n5019,s1n5019,notn5019;
or (n5019,s0n5019,s1n5019);
not(notn5019,n5021);
and (s0n5019,notn5019,1'b0);
and (s1n5019,n5021,n5020);
or (n5021,n5022,n5028);
or (n5022,n5023,n5027);
and (n5023,n2942,n5024);
or (n5024,n5025,n549);
or (n5025,n5026,n560);
or (n5026,n566,n564);
and (n5027,n2885,n5024);
and (n5028,n2899,n2894);
wire s0n5029,s1n5029,notn5029;
or (n5029,s0n5029,s1n5029);
not(notn5029,n5021);
and (s0n5029,notn5029,1'b0);
and (s1n5029,n5021,n5030);
or (n5031,n5032,n5037,n6068);
and (n5032,n5033,n5035);
wire s0n5033,s1n5033,notn5033;
or (n5033,s0n5033,s1n5033);
not(notn5033,n5021);
and (s0n5033,notn5033,1'b0);
and (s1n5033,n5021,n5034);
wire s0n5035,s1n5035,notn5035;
or (n5035,s0n5035,s1n5035);
not(notn5035,n5021);
and (s0n5035,notn5035,1'b0);
and (s1n5035,n5021,n5036);
and (n5037,n5035,n5038);
or (n5038,n5039,n5044,n6067);
and (n5039,n5040,n5042);
wire s0n5040,s1n5040,notn5040;
or (n5040,s0n5040,s1n5040);
not(notn5040,n5021);
and (s0n5040,notn5040,1'b0);
and (s1n5040,n5021,n5041);
wire s0n5042,s1n5042,notn5042;
or (n5042,s0n5042,s1n5042);
not(notn5042,n5021);
and (s0n5042,notn5042,1'b0);
and (s1n5042,n5021,n5043);
and (n5044,n5042,n5045);
or (n5045,n5046,n5051,n6066);
and (n5046,n5047,n5049);
wire s0n5047,s1n5047,notn5047;
or (n5047,s0n5047,s1n5047);
not(notn5047,n5021);
and (s0n5047,notn5047,1'b0);
and (s1n5047,n5021,n5048);
wire s0n5049,s1n5049,notn5049;
or (n5049,s0n5049,s1n5049);
not(notn5049,n5021);
and (s0n5049,notn5049,1'b0);
and (s1n5049,n5021,n5050);
and (n5051,n5049,n5052);
or (n5052,n5053,n5058,n6065);
and (n5053,n5054,n5056);
wire s0n5054,s1n5054,notn5054;
or (n5054,s0n5054,s1n5054);
not(notn5054,n5021);
and (s0n5054,notn5054,1'b0);
and (s1n5054,n5021,n5055);
wire s0n5056,s1n5056,notn5056;
or (n5056,s0n5056,s1n5056);
not(notn5056,n5021);
and (s0n5056,notn5056,1'b0);
and (s1n5056,n5021,n5057);
and (n5058,n5056,n5059);
or (n5059,n5060,n5198,n6064);
and (n5060,n5061,n5137);
wire s0n5061,s1n5061,notn5061;
or (n5061,s0n5061,s1n5061);
not(notn5061,n5021);
and (s0n5061,notn5061,n5062);
and (s1n5061,n5021,n5136);
or (n5062,1'b0,n5063,n5095,n5109,n5124);
and (n5063,n5064,n2710);
or (n5064,1'b0,n5065,n5080,n5085,n5090);
and (n5065,n5066,n5071);
wire s0n5066,s1n5066,notn5066;
or (n5066,s0n5066,s1n5066);
not(notn5066,n5069);
and (s0n5066,notn5066,n5067);
and (s1n5066,n5069,n5068);
or (n5069,n5070,n2901);
or (n5070,n2938,n2923);
or (n5071,n5072,n2943);
and (n5072,n5073,n549);
or (n5073,n5074,n2923);
or (n5074,n5075,n2922);
or (n5075,n5076,n2938);
or (n5076,n5077,n2937);
or (n5077,n5078,n4950);
or (n5078,n5079,n4959);
nor (n5079,n2749,n2935,n2818,n2844);
and (n5080,n5081,n5083);
wire s0n5081,s1n5081,notn5081;
or (n5081,s0n5081,s1n5081);
not(notn5081,n5069);
and (s0n5081,notn5081,n5082);
and (s1n5081,n5069,n5067);
or (n5083,n5084,n2951);
and (n5084,n5073,n560);
and (n5085,n5086,n5088);
wire s0n5086,s1n5086,notn5086;
or (n5086,s0n5086,s1n5086);
not(notn5086,n5069);
and (s0n5086,notn5086,n5087);
and (s1n5086,n5069,n5082);
or (n5088,n5089,n2959);
and (n5089,n5073,n564);
and (n5090,n5091,n5093);
wire s0n5091,s1n5091,notn5091;
or (n5091,s0n5091,s1n5091);
not(notn5091,n5069);
and (s0n5091,notn5091,n5092);
and (s1n5091,n5069,n5087);
or (n5093,n5094,n2968);
and (n5094,n5073,n566);
and (n5095,n5096,n2722);
or (n5096,1'b0,n5097,n5100,n5103,n5106);
and (n5097,n5098,n5071);
wire s0n5098,s1n5098,notn5098;
or (n5098,s0n5098,s1n5098);
not(notn5098,n5069);
and (s0n5098,notn5098,n5099);
and (s1n5098,n5069,n5092);
and (n5100,n5101,n5083);
wire s0n5101,s1n5101,notn5101;
or (n5101,s0n5101,s1n5101);
not(notn5101,n5069);
and (s0n5101,notn5101,n5102);
and (s1n5101,n5069,n5099);
and (n5103,n5104,n5088);
wire s0n5104,s1n5104,notn5104;
or (n5104,s0n5104,s1n5104);
not(notn5104,n5069);
and (s0n5104,notn5104,n5105);
and (s1n5104,n5069,n5102);
and (n5106,n5107,n5093);
wire s0n5107,s1n5107,notn5107;
or (n5107,s0n5107,s1n5107);
not(notn5107,n5069);
and (s0n5107,notn5107,n5108);
and (s1n5107,n5069,n5105);
and (n5109,n5110,n2734);
or (n5110,1'b0,n5111,n5115,n5118,n5121);
and (n5111,n5112,n5071);
wire s0n5112,s1n5112,notn5112;
or (n5112,s0n5112,s1n5112);
not(notn5112,n5069);
and (s0n5112,notn5112,n5113);
and (s1n5112,n5069,n5114);
and (n5115,n5116,n5083);
wire s0n5116,s1n5116,notn5116;
or (n5116,s0n5116,s1n5116);
not(notn5116,n5069);
and (s0n5116,notn5116,n5117);
and (s1n5116,n5069,n5113);
and (n5118,n5119,n5088);
wire s0n5119,s1n5119,notn5119;
or (n5119,s0n5119,s1n5119);
not(notn5119,n5069);
and (s0n5119,notn5119,n5120);
and (s1n5119,n5069,n5117);
and (n5121,n5122,n5093);
wire s0n5122,s1n5122,notn5122;
or (n5122,s0n5122,s1n5122);
not(notn5122,n5069);
and (s0n5122,notn5122,n5123);
and (s1n5122,n5069,n5120);
and (n5124,n5125,n2744);
or (n5125,1'b0,n5126,n5129,n5132,n5134);
and (n5126,n5127,n5071);
wire s0n5127,s1n5127,notn5127;
or (n5127,s0n5127,s1n5127);
not(notn5127,n5069);
and (s0n5127,notn5127,n5128);
and (s1n5127,n5069,n5123);
and (n5129,n5130,n5083);
wire s0n5130,s1n5130,notn5130;
or (n5130,s0n5130,s1n5130);
not(notn5130,n5069);
and (s0n5130,notn5130,n5131);
and (s1n5130,n5069,n5128);
and (n5132,n5133,n5088);
wire s0n5133,s1n5133,notn5133;
or (n5133,s0n5133,s1n5133);
not(notn5133,n5069);
and (s0n5133,notn5133,n2168);
and (s1n5133,n5069,n5131);
and (n5134,n5135,n5093);
wire s0n5135,s1n5135,notn5135;
or (n5135,s0n5135,s1n5135);
not(notn5135,n5069);
and (s0n5135,notn5135,n1831);
and (s1n5135,n5069,n2168);
wire s0n5137,s1n5137,notn5137;
or (n5137,s0n5137,s1n5137);
not(notn5137,n5021);
and (s0n5137,notn5137,n5138);
and (s1n5137,n5021,n5197);
or (n5138,1'b0,n5139,n5154,n5168,n5183);
and (n5139,n5140,n2710);
or (n5140,1'b0,n5141,n5145,n5148,n5151);
and (n5141,n5142,n5071);
wire s0n5142,s1n5142,notn5142;
or (n5142,s0n5142,s1n5142);
not(notn5142,n5069);
and (s0n5142,notn5142,n5143);
and (s1n5142,n5069,n5144);
and (n5145,n5146,n5083);
wire s0n5146,s1n5146,notn5146;
or (n5146,s0n5146,s1n5146);
not(notn5146,n5069);
and (s0n5146,notn5146,n5147);
and (s1n5146,n5069,n5143);
and (n5148,n5149,n5088);
wire s0n5149,s1n5149,notn5149;
or (n5149,s0n5149,s1n5149);
not(notn5149,n5069);
and (s0n5149,notn5149,n5150);
and (s1n5149,n5069,n5147);
and (n5151,n5152,n5093);
wire s0n5152,s1n5152,notn5152;
or (n5152,s0n5152,s1n5152);
not(notn5152,n5069);
and (s0n5152,notn5152,n5153);
and (s1n5152,n5069,n5150);
and (n5154,n5155,n2722);
or (n5155,1'b0,n5156,n5159,n5162,n5165);
and (n5156,n5157,n5071);
wire s0n5157,s1n5157,notn5157;
or (n5157,s0n5157,s1n5157);
not(notn5157,n5069);
and (s0n5157,notn5157,n5158);
and (s1n5157,n5069,n5153);
and (n5159,n5160,n5083);
wire s0n5160,s1n5160,notn5160;
or (n5160,s0n5160,s1n5160);
not(notn5160,n5069);
and (s0n5160,notn5160,n5161);
and (s1n5160,n5069,n5158);
and (n5162,n5163,n5088);
wire s0n5163,s1n5163,notn5163;
or (n5163,s0n5163,s1n5163);
not(notn5163,n5069);
and (s0n5163,notn5163,n5164);
and (s1n5163,n5069,n5161);
and (n5165,n5166,n5093);
wire s0n5166,s1n5166,notn5166;
or (n5166,s0n5166,s1n5166);
not(notn5166,n5069);
and (s0n5166,notn5166,n5167);
and (s1n5166,n5069,n5164);
and (n5168,n5169,n2734);
or (n5169,1'b0,n5170,n5174,n5177,n5180);
and (n5170,n5171,n5071);
wire s0n5171,s1n5171,notn5171;
or (n5171,s0n5171,s1n5171);
not(notn5171,n5069);
and (s0n5171,notn5171,n5172);
and (s1n5171,n5069,n5173);
and (n5174,n5175,n5083);
wire s0n5175,s1n5175,notn5175;
or (n5175,s0n5175,s1n5175);
not(notn5175,n5069);
and (s0n5175,notn5175,n5176);
and (s1n5175,n5069,n5172);
and (n5177,n5178,n5088);
wire s0n5178,s1n5178,notn5178;
or (n5178,s0n5178,s1n5178);
not(notn5178,n5069);
and (s0n5178,notn5178,n5179);
and (s1n5178,n5069,n5176);
and (n5180,n5181,n5093);
wire s0n5181,s1n5181,notn5181;
or (n5181,s0n5181,s1n5181);
not(notn5181,n5069);
and (s0n5181,notn5181,n5182);
and (s1n5181,n5069,n5179);
and (n5183,n5184,n2744);
or (n5184,1'b0,n5185,n5188,n5191,n5194);
and (n5185,n5186,n5071);
wire s0n5186,s1n5186,notn5186;
or (n5186,s0n5186,s1n5186);
not(notn5186,n5069);
and (s0n5186,notn5186,n5187);
and (s1n5186,n5069,n5182);
and (n5188,n5189,n5083);
wire s0n5189,s1n5189,notn5189;
or (n5189,s0n5189,s1n5189);
not(notn5189,n5069);
and (s0n5189,notn5189,n5190);
and (s1n5189,n5069,n5187);
and (n5191,n5192,n5088);
wire s0n5192,s1n5192,notn5192;
or (n5192,s0n5192,s1n5192);
not(notn5192,n5069);
and (s0n5192,notn5192,n5193);
and (s1n5192,n5069,n5190);
and (n5194,n5195,n5093);
wire s0n5195,s1n5195,notn5195;
or (n5195,s0n5195,s1n5195);
not(notn5195,n5069);
and (s0n5195,notn5195,n5196);
and (s1n5195,n5069,n5193);
and (n5198,n5137,n5199);
or (n5199,n5200,n5321,n6063);
and (n5200,n5201,n5260);
wire s0n5201,s1n5201,notn5201;
or (n5201,s0n5201,s1n5201);
not(notn5201,n5021);
and (s0n5201,notn5201,n5202);
and (s1n5201,n5021,n5259);
or (n5202,1'b0,n5203,n5218,n5232,n5247);
and (n5203,n5204,n2710);
or (n5204,1'b0,n5205,n5209,n5212,n5215);
and (n5205,n5206,n5071);
wire s0n5206,s1n5206,notn5206;
or (n5206,s0n5206,s1n5206);
not(notn5206,n5069);
and (s0n5206,notn5206,n5207);
and (s1n5206,n5069,n5208);
and (n5209,n5210,n5083);
wire s0n5210,s1n5210,notn5210;
or (n5210,s0n5210,s1n5210);
not(notn5210,n5069);
and (s0n5210,notn5210,n5211);
and (s1n5210,n5069,n5207);
and (n5212,n5213,n5088);
wire s0n5213,s1n5213,notn5213;
or (n5213,s0n5213,s1n5213);
not(notn5213,n5069);
and (s0n5213,notn5213,n5214);
and (s1n5213,n5069,n5211);
and (n5215,n5216,n5093);
wire s0n5216,s1n5216,notn5216;
or (n5216,s0n5216,s1n5216);
not(notn5216,n5069);
and (s0n5216,notn5216,n5217);
and (s1n5216,n5069,n5214);
and (n5218,n5219,n2722);
or (n5219,1'b0,n5220,n5223,n5226,n5229);
and (n5220,n5221,n5071);
wire s0n5221,s1n5221,notn5221;
or (n5221,s0n5221,s1n5221);
not(notn5221,n5069);
and (s0n5221,notn5221,n5222);
and (s1n5221,n5069,n5217);
and (n5223,n5224,n5083);
wire s0n5224,s1n5224,notn5224;
or (n5224,s0n5224,s1n5224);
not(notn5224,n5069);
and (s0n5224,notn5224,n5225);
and (s1n5224,n5069,n5222);
and (n5226,n5227,n5088);
wire s0n5227,s1n5227,notn5227;
or (n5227,s0n5227,s1n5227);
not(notn5227,n5069);
and (s0n5227,notn5227,n5228);
and (s1n5227,n5069,n5225);
and (n5229,n5230,n5093);
wire s0n5230,s1n5230,notn5230;
or (n5230,s0n5230,s1n5230);
not(notn5230,n5069);
and (s0n5230,notn5230,n5231);
and (s1n5230,n5069,n5228);
and (n5232,n5233,n2734);
or (n5233,1'b0,n5234,n5238,n5241,n5244);
and (n5234,n5235,n5071);
wire s0n5235,s1n5235,notn5235;
or (n5235,s0n5235,s1n5235);
not(notn5235,n5069);
and (s0n5235,notn5235,n5236);
and (s1n5235,n5069,n5237);
and (n5238,n5239,n5083);
wire s0n5239,s1n5239,notn5239;
or (n5239,s0n5239,s1n5239);
not(notn5239,n5069);
and (s0n5239,notn5239,n5240);
and (s1n5239,n5069,n5236);
and (n5241,n5242,n5088);
wire s0n5242,s1n5242,notn5242;
or (n5242,s0n5242,s1n5242);
not(notn5242,n5069);
and (s0n5242,notn5242,n5243);
and (s1n5242,n5069,n5240);
and (n5244,n5245,n5093);
wire s0n5245,s1n5245,notn5245;
or (n5245,s0n5245,s1n5245);
not(notn5245,n5069);
and (s0n5245,notn5245,n5246);
and (s1n5245,n5069,n5243);
and (n5247,n5248,n2744);
or (n5248,1'b0,n5249,n5252,n5255,n5257);
and (n5249,n5250,n5071);
wire s0n5250,s1n5250,notn5250;
or (n5250,s0n5250,s1n5250);
not(notn5250,n5069);
and (s0n5250,notn5250,n5251);
and (s1n5250,n5069,n5246);
and (n5252,n5253,n5083);
wire s0n5253,s1n5253,notn5253;
or (n5253,s0n5253,s1n5253);
not(notn5253,n5069);
and (s0n5253,notn5253,n5254);
and (s1n5253,n5069,n5251);
and (n5255,n5256,n5088);
wire s0n5256,s1n5256,notn5256;
or (n5256,s0n5256,s1n5256);
not(notn5256,n5069);
and (s0n5256,notn5256,n2184);
and (s1n5256,n5069,n5254);
and (n5257,n5258,n5093);
wire s0n5258,s1n5258,notn5258;
or (n5258,s0n5258,s1n5258);
not(notn5258,n5069);
and (s0n5258,notn5258,n1848);
and (s1n5258,n5069,n2184);
wire s0n5260,s1n5260,notn5260;
or (n5260,s0n5260,s1n5260);
not(notn5260,n5021);
and (s0n5260,notn5260,n5261);
and (s1n5260,n5021,n5320);
or (n5261,1'b0,n5262,n5277,n5291,n5306);
and (n5262,n5263,n2710);
or (n5263,1'b0,n5264,n5268,n5271,n5274);
and (n5264,n5265,n5071);
wire s0n5265,s1n5265,notn5265;
or (n5265,s0n5265,s1n5265);
not(notn5265,n5069);
and (s0n5265,notn5265,n5266);
and (s1n5265,n5069,n5267);
and (n5268,n5269,n5083);
wire s0n5269,s1n5269,notn5269;
or (n5269,s0n5269,s1n5269);
not(notn5269,n5069);
and (s0n5269,notn5269,n5270);
and (s1n5269,n5069,n5266);
and (n5271,n5272,n5088);
wire s0n5272,s1n5272,notn5272;
or (n5272,s0n5272,s1n5272);
not(notn5272,n5069);
and (s0n5272,notn5272,n5273);
and (s1n5272,n5069,n5270);
and (n5274,n5275,n5093);
wire s0n5275,s1n5275,notn5275;
or (n5275,s0n5275,s1n5275);
not(notn5275,n5069);
and (s0n5275,notn5275,n5276);
and (s1n5275,n5069,n5273);
and (n5277,n5278,n2722);
or (n5278,1'b0,n5279,n5282,n5285,n5288);
and (n5279,n5280,n5071);
wire s0n5280,s1n5280,notn5280;
or (n5280,s0n5280,s1n5280);
not(notn5280,n5069);
and (s0n5280,notn5280,n5281);
and (s1n5280,n5069,n5276);
and (n5282,n5283,n5083);
wire s0n5283,s1n5283,notn5283;
or (n5283,s0n5283,s1n5283);
not(notn5283,n5069);
and (s0n5283,notn5283,n5284);
and (s1n5283,n5069,n5281);
and (n5285,n5286,n5088);
wire s0n5286,s1n5286,notn5286;
or (n5286,s0n5286,s1n5286);
not(notn5286,n5069);
and (s0n5286,notn5286,n5287);
and (s1n5286,n5069,n5284);
and (n5288,n5289,n5093);
wire s0n5289,s1n5289,notn5289;
or (n5289,s0n5289,s1n5289);
not(notn5289,n5069);
and (s0n5289,notn5289,n5290);
and (s1n5289,n5069,n5287);
and (n5291,n5292,n2734);
or (n5292,1'b0,n5293,n5297,n5300,n5303);
and (n5293,n5294,n5071);
wire s0n5294,s1n5294,notn5294;
or (n5294,s0n5294,s1n5294);
not(notn5294,n5069);
and (s0n5294,notn5294,n5295);
and (s1n5294,n5069,n5296);
and (n5297,n5298,n5083);
wire s0n5298,s1n5298,notn5298;
or (n5298,s0n5298,s1n5298);
not(notn5298,n5069);
and (s0n5298,notn5298,n5299);
and (s1n5298,n5069,n5295);
and (n5300,n5301,n5088);
wire s0n5301,s1n5301,notn5301;
or (n5301,s0n5301,s1n5301);
not(notn5301,n5069);
and (s0n5301,notn5301,n5302);
and (s1n5301,n5069,n5299);
and (n5303,n5304,n5093);
wire s0n5304,s1n5304,notn5304;
or (n5304,s0n5304,s1n5304);
not(notn5304,n5069);
and (s0n5304,notn5304,n5305);
and (s1n5304,n5069,n5302);
and (n5306,n5307,n2744);
or (n5307,1'b0,n5308,n5311,n5314,n5317);
and (n5308,n5309,n5071);
wire s0n5309,s1n5309,notn5309;
or (n5309,s0n5309,s1n5309);
not(notn5309,n5069);
and (s0n5309,notn5309,n5310);
and (s1n5309,n5069,n5305);
and (n5311,n5312,n5083);
wire s0n5312,s1n5312,notn5312;
or (n5312,s0n5312,s1n5312);
not(notn5312,n5069);
and (s0n5312,notn5312,n5313);
and (s1n5312,n5069,n5310);
and (n5314,n5315,n5088);
wire s0n5315,s1n5315,notn5315;
or (n5315,s0n5315,s1n5315);
not(notn5315,n5069);
and (s0n5315,notn5315,n5316);
and (s1n5315,n5069,n5313);
and (n5317,n5318,n5093);
wire s0n5318,s1n5318,notn5318;
or (n5318,s0n5318,s1n5318);
not(notn5318,n5069);
and (s0n5318,notn5318,n5319);
and (s1n5318,n5069,n5316);
and (n5321,n5260,n5322);
or (n5322,n5323,n5444,n6062);
and (n5323,n5324,n5383);
wire s0n5324,s1n5324,notn5324;
or (n5324,s0n5324,s1n5324);
not(notn5324,n5021);
and (s0n5324,notn5324,n5325);
and (s1n5324,n5021,n5382);
or (n5325,1'b0,n5326,n5341,n5355,n5370);
and (n5326,n5327,n2710);
or (n5327,1'b0,n5328,n5332,n5335,n5338);
and (n5328,n5329,n5071);
wire s0n5329,s1n5329,notn5329;
or (n5329,s0n5329,s1n5329);
not(notn5329,n5069);
and (s0n5329,notn5329,n5330);
and (s1n5329,n5069,n5331);
and (n5332,n5333,n5083);
wire s0n5333,s1n5333,notn5333;
or (n5333,s0n5333,s1n5333);
not(notn5333,n5069);
and (s0n5333,notn5333,n5334);
and (s1n5333,n5069,n5330);
and (n5335,n5336,n5088);
wire s0n5336,s1n5336,notn5336;
or (n5336,s0n5336,s1n5336);
not(notn5336,n5069);
and (s0n5336,notn5336,n5337);
and (s1n5336,n5069,n5334);
and (n5338,n5339,n5093);
wire s0n5339,s1n5339,notn5339;
or (n5339,s0n5339,s1n5339);
not(notn5339,n5069);
and (s0n5339,notn5339,n5340);
and (s1n5339,n5069,n5337);
and (n5341,n5342,n2722);
or (n5342,1'b0,n5343,n5346,n5349,n5352);
and (n5343,n5344,n5071);
wire s0n5344,s1n5344,notn5344;
or (n5344,s0n5344,s1n5344);
not(notn5344,n5069);
and (s0n5344,notn5344,n5345);
and (s1n5344,n5069,n5340);
and (n5346,n5347,n5083);
wire s0n5347,s1n5347,notn5347;
or (n5347,s0n5347,s1n5347);
not(notn5347,n5069);
and (s0n5347,notn5347,n5348);
and (s1n5347,n5069,n5345);
and (n5349,n5350,n5088);
wire s0n5350,s1n5350,notn5350;
or (n5350,s0n5350,s1n5350);
not(notn5350,n5069);
and (s0n5350,notn5350,n5351);
and (s1n5350,n5069,n5348);
and (n5352,n5353,n5093);
wire s0n5353,s1n5353,notn5353;
or (n5353,s0n5353,s1n5353);
not(notn5353,n5069);
and (s0n5353,notn5353,n5354);
and (s1n5353,n5069,n5351);
and (n5355,n5356,n2734);
or (n5356,1'b0,n5357,n5361,n5364,n5367);
and (n5357,n5358,n5071);
wire s0n5358,s1n5358,notn5358;
or (n5358,s0n5358,s1n5358);
not(notn5358,n5069);
and (s0n5358,notn5358,n5359);
and (s1n5358,n5069,n5360);
and (n5361,n5362,n5083);
wire s0n5362,s1n5362,notn5362;
or (n5362,s0n5362,s1n5362);
not(notn5362,n5069);
and (s0n5362,notn5362,n5363);
and (s1n5362,n5069,n5359);
and (n5364,n5365,n5088);
wire s0n5365,s1n5365,notn5365;
or (n5365,s0n5365,s1n5365);
not(notn5365,n5069);
and (s0n5365,notn5365,n5366);
and (s1n5365,n5069,n5363);
and (n5367,n5368,n5093);
wire s0n5368,s1n5368,notn5368;
or (n5368,s0n5368,s1n5368);
not(notn5368,n5069);
and (s0n5368,notn5368,n5369);
and (s1n5368,n5069,n5366);
and (n5370,n5371,n2744);
or (n5371,1'b0,n5372,n5375,n5378,n5380);
and (n5372,n5373,n5071);
wire s0n5373,s1n5373,notn5373;
or (n5373,s0n5373,s1n5373);
not(notn5373,n5069);
and (s0n5373,notn5373,n5374);
and (s1n5373,n5069,n5369);
and (n5375,n5376,n5083);
wire s0n5376,s1n5376,notn5376;
or (n5376,s0n5376,s1n5376);
not(notn5376,n5069);
and (s0n5376,notn5376,n5377);
and (s1n5376,n5069,n5374);
and (n5378,n5379,n5088);
wire s0n5379,s1n5379,notn5379;
or (n5379,s0n5379,s1n5379);
not(notn5379,n5069);
and (s0n5379,notn5379,n2200);
and (s1n5379,n5069,n5377);
and (n5380,n5381,n5093);
wire s0n5381,s1n5381,notn5381;
or (n5381,s0n5381,s1n5381);
not(notn5381,n5069);
and (s0n5381,notn5381,n1865);
and (s1n5381,n5069,n2200);
wire s0n5383,s1n5383,notn5383;
or (n5383,s0n5383,s1n5383);
not(notn5383,n5021);
and (s0n5383,notn5383,n5384);
and (s1n5383,n5021,n5443);
or (n5384,1'b0,n5385,n5400,n5414,n5429);
and (n5385,n5386,n2710);
or (n5386,1'b0,n5387,n5391,n5394,n5397);
and (n5387,n5388,n5071);
wire s0n5388,s1n5388,notn5388;
or (n5388,s0n5388,s1n5388);
not(notn5388,n5069);
and (s0n5388,notn5388,n5389);
and (s1n5388,n5069,n5390);
and (n5391,n5392,n5083);
wire s0n5392,s1n5392,notn5392;
or (n5392,s0n5392,s1n5392);
not(notn5392,n5069);
and (s0n5392,notn5392,n5393);
and (s1n5392,n5069,n5389);
and (n5394,n5395,n5088);
wire s0n5395,s1n5395,notn5395;
or (n5395,s0n5395,s1n5395);
not(notn5395,n5069);
and (s0n5395,notn5395,n5396);
and (s1n5395,n5069,n5393);
and (n5397,n5398,n5093);
wire s0n5398,s1n5398,notn5398;
or (n5398,s0n5398,s1n5398);
not(notn5398,n5069);
and (s0n5398,notn5398,n5399);
and (s1n5398,n5069,n5396);
and (n5400,n5401,n2722);
or (n5401,1'b0,n5402,n5405,n5408,n5411);
and (n5402,n5403,n5071);
wire s0n5403,s1n5403,notn5403;
or (n5403,s0n5403,s1n5403);
not(notn5403,n5069);
and (s0n5403,notn5403,n5404);
and (s1n5403,n5069,n5399);
and (n5405,n5406,n5083);
wire s0n5406,s1n5406,notn5406;
or (n5406,s0n5406,s1n5406);
not(notn5406,n5069);
and (s0n5406,notn5406,n5407);
and (s1n5406,n5069,n5404);
and (n5408,n5409,n5088);
wire s0n5409,s1n5409,notn5409;
or (n5409,s0n5409,s1n5409);
not(notn5409,n5069);
and (s0n5409,notn5409,n5410);
and (s1n5409,n5069,n5407);
and (n5411,n5412,n5093);
wire s0n5412,s1n5412,notn5412;
or (n5412,s0n5412,s1n5412);
not(notn5412,n5069);
and (s0n5412,notn5412,n5413);
and (s1n5412,n5069,n5410);
and (n5414,n5415,n2734);
or (n5415,1'b0,n5416,n5420,n5423,n5426);
and (n5416,n5417,n5071);
wire s0n5417,s1n5417,notn5417;
or (n5417,s0n5417,s1n5417);
not(notn5417,n5069);
and (s0n5417,notn5417,n5418);
and (s1n5417,n5069,n5419);
and (n5420,n5421,n5083);
wire s0n5421,s1n5421,notn5421;
or (n5421,s0n5421,s1n5421);
not(notn5421,n5069);
and (s0n5421,notn5421,n5422);
and (s1n5421,n5069,n5418);
and (n5423,n5424,n5088);
wire s0n5424,s1n5424,notn5424;
or (n5424,s0n5424,s1n5424);
not(notn5424,n5069);
and (s0n5424,notn5424,n5425);
and (s1n5424,n5069,n5422);
and (n5426,n5427,n5093);
wire s0n5427,s1n5427,notn5427;
or (n5427,s0n5427,s1n5427);
not(notn5427,n5069);
and (s0n5427,notn5427,n5428);
and (s1n5427,n5069,n5425);
and (n5429,n5430,n2744);
or (n5430,1'b0,n5431,n5434,n5437,n5440);
and (n5431,n5432,n5071);
wire s0n5432,s1n5432,notn5432;
or (n5432,s0n5432,s1n5432);
not(notn5432,n5069);
and (s0n5432,notn5432,n5433);
and (s1n5432,n5069,n5428);
and (n5434,n5435,n5083);
wire s0n5435,s1n5435,notn5435;
or (n5435,s0n5435,s1n5435);
not(notn5435,n5069);
and (s0n5435,notn5435,n5436);
and (s1n5435,n5069,n5433);
and (n5437,n5438,n5088);
wire s0n5438,s1n5438,notn5438;
or (n5438,s0n5438,s1n5438);
not(notn5438,n5069);
and (s0n5438,notn5438,n5439);
and (s1n5438,n5069,n5436);
and (n5440,n5441,n5093);
wire s0n5441,s1n5441,notn5441;
or (n5441,s0n5441,s1n5441);
not(notn5441,n5069);
and (s0n5441,notn5441,n5442);
and (s1n5441,n5069,n5439);
and (n5444,n5383,n5445);
or (n5445,n5446,n5567,n6061);
and (n5446,n5447,n5506);
wire s0n5447,s1n5447,notn5447;
or (n5447,s0n5447,s1n5447);
not(notn5447,n5021);
and (s0n5447,notn5447,n5448);
and (s1n5447,n5021,n5505);
or (n5448,1'b0,n5449,n5464,n5478,n5493);
and (n5449,n5450,n2710);
or (n5450,1'b0,n5451,n5455,n5458,n5461);
and (n5451,n5452,n5071);
wire s0n5452,s1n5452,notn5452;
or (n5452,s0n5452,s1n5452);
not(notn5452,n5069);
and (s0n5452,notn5452,n5453);
and (s1n5452,n5069,n5454);
and (n5455,n5456,n5083);
wire s0n5456,s1n5456,notn5456;
or (n5456,s0n5456,s1n5456);
not(notn5456,n5069);
and (s0n5456,notn5456,n5457);
and (s1n5456,n5069,n5453);
and (n5458,n5459,n5088);
wire s0n5459,s1n5459,notn5459;
or (n5459,s0n5459,s1n5459);
not(notn5459,n5069);
and (s0n5459,notn5459,n5460);
and (s1n5459,n5069,n5457);
and (n5461,n5462,n5093);
wire s0n5462,s1n5462,notn5462;
or (n5462,s0n5462,s1n5462);
not(notn5462,n5069);
and (s0n5462,notn5462,n5463);
and (s1n5462,n5069,n5460);
and (n5464,n5465,n2722);
or (n5465,1'b0,n5466,n5469,n5472,n5475);
and (n5466,n5467,n5071);
wire s0n5467,s1n5467,notn5467;
or (n5467,s0n5467,s1n5467);
not(notn5467,n5069);
and (s0n5467,notn5467,n5468);
and (s1n5467,n5069,n5463);
and (n5469,n5470,n5083);
wire s0n5470,s1n5470,notn5470;
or (n5470,s0n5470,s1n5470);
not(notn5470,n5069);
and (s0n5470,notn5470,n5471);
and (s1n5470,n5069,n5468);
and (n5472,n5473,n5088);
wire s0n5473,s1n5473,notn5473;
or (n5473,s0n5473,s1n5473);
not(notn5473,n5069);
and (s0n5473,notn5473,n5474);
and (s1n5473,n5069,n5471);
and (n5475,n5476,n5093);
wire s0n5476,s1n5476,notn5476;
or (n5476,s0n5476,s1n5476);
not(notn5476,n5069);
and (s0n5476,notn5476,n5477);
and (s1n5476,n5069,n5474);
and (n5478,n5479,n2734);
or (n5479,1'b0,n5480,n5484,n5487,n5490);
and (n5480,n5481,n5071);
wire s0n5481,s1n5481,notn5481;
or (n5481,s0n5481,s1n5481);
not(notn5481,n5069);
and (s0n5481,notn5481,n5482);
and (s1n5481,n5069,n5483);
and (n5484,n5485,n5083);
wire s0n5485,s1n5485,notn5485;
or (n5485,s0n5485,s1n5485);
not(notn5485,n5069);
and (s0n5485,notn5485,n5486);
and (s1n5485,n5069,n5482);
and (n5487,n5488,n5088);
wire s0n5488,s1n5488,notn5488;
or (n5488,s0n5488,s1n5488);
not(notn5488,n5069);
and (s0n5488,notn5488,n5489);
and (s1n5488,n5069,n5486);
and (n5490,n5491,n5093);
wire s0n5491,s1n5491,notn5491;
or (n5491,s0n5491,s1n5491);
not(notn5491,n5069);
and (s0n5491,notn5491,n5492);
and (s1n5491,n5069,n5489);
and (n5493,n5494,n2744);
or (n5494,1'b0,n5495,n5498,n5501,n5503);
and (n5495,n5496,n5071);
wire s0n5496,s1n5496,notn5496;
or (n5496,s0n5496,s1n5496);
not(notn5496,n5069);
and (s0n5496,notn5496,n5497);
and (s1n5496,n5069,n5492);
and (n5498,n5499,n5083);
wire s0n5499,s1n5499,notn5499;
or (n5499,s0n5499,s1n5499);
not(notn5499,n5069);
and (s0n5499,notn5499,n5500);
and (s1n5499,n5069,n5497);
and (n5501,n5502,n5088);
wire s0n5502,s1n5502,notn5502;
or (n5502,s0n5502,s1n5502);
not(notn5502,n5069);
and (s0n5502,notn5502,n2216);
and (s1n5502,n5069,n5500);
and (n5503,n5504,n5093);
wire s0n5504,s1n5504,notn5504;
or (n5504,s0n5504,s1n5504);
not(notn5504,n5069);
and (s0n5504,notn5504,n1890);
and (s1n5504,n5069,n2216);
wire s0n5506,s1n5506,notn5506;
or (n5506,s0n5506,s1n5506);
not(notn5506,n5021);
and (s0n5506,notn5506,n5507);
and (s1n5506,n5021,n5566);
or (n5507,1'b0,n5508,n5523,n5537,n5552);
and (n5508,n5509,n2710);
or (n5509,1'b0,n5510,n5514,n5517,n5520);
and (n5510,n5511,n5071);
wire s0n5511,s1n5511,notn5511;
or (n5511,s0n5511,s1n5511);
not(notn5511,n5069);
and (s0n5511,notn5511,n5512);
and (s1n5511,n5069,n5513);
and (n5514,n5515,n5083);
wire s0n5515,s1n5515,notn5515;
or (n5515,s0n5515,s1n5515);
not(notn5515,n5069);
and (s0n5515,notn5515,n5516);
and (s1n5515,n5069,n5512);
and (n5517,n5518,n5088);
wire s0n5518,s1n5518,notn5518;
or (n5518,s0n5518,s1n5518);
not(notn5518,n5069);
and (s0n5518,notn5518,n5519);
and (s1n5518,n5069,n5516);
and (n5520,n5521,n5093);
wire s0n5521,s1n5521,notn5521;
or (n5521,s0n5521,s1n5521);
not(notn5521,n5069);
and (s0n5521,notn5521,n5522);
and (s1n5521,n5069,n5519);
and (n5523,n5524,n2722);
or (n5524,1'b0,n5525,n5528,n5531,n5534);
and (n5525,n5526,n5071);
wire s0n5526,s1n5526,notn5526;
or (n5526,s0n5526,s1n5526);
not(notn5526,n5069);
and (s0n5526,notn5526,n5527);
and (s1n5526,n5069,n5522);
and (n5528,n5529,n5083);
wire s0n5529,s1n5529,notn5529;
or (n5529,s0n5529,s1n5529);
not(notn5529,n5069);
and (s0n5529,notn5529,n5530);
and (s1n5529,n5069,n5527);
and (n5531,n5532,n5088);
wire s0n5532,s1n5532,notn5532;
or (n5532,s0n5532,s1n5532);
not(notn5532,n5069);
and (s0n5532,notn5532,n5533);
and (s1n5532,n5069,n5530);
and (n5534,n5535,n5093);
wire s0n5535,s1n5535,notn5535;
or (n5535,s0n5535,s1n5535);
not(notn5535,n5069);
and (s0n5535,notn5535,n5536);
and (s1n5535,n5069,n5533);
and (n5537,n5538,n2734);
or (n5538,1'b0,n5539,n5543,n5546,n5549);
and (n5539,n5540,n5071);
wire s0n5540,s1n5540,notn5540;
or (n5540,s0n5540,s1n5540);
not(notn5540,n5069);
and (s0n5540,notn5540,n5541);
and (s1n5540,n5069,n5542);
and (n5543,n5544,n5083);
wire s0n5544,s1n5544,notn5544;
or (n5544,s0n5544,s1n5544);
not(notn5544,n5069);
and (s0n5544,notn5544,n5545);
and (s1n5544,n5069,n5541);
and (n5546,n5547,n5088);
wire s0n5547,s1n5547,notn5547;
or (n5547,s0n5547,s1n5547);
not(notn5547,n5069);
and (s0n5547,notn5547,n5548);
and (s1n5547,n5069,n5545);
and (n5549,n5550,n5093);
wire s0n5550,s1n5550,notn5550;
or (n5550,s0n5550,s1n5550);
not(notn5550,n5069);
and (s0n5550,notn5550,n5551);
and (s1n5550,n5069,n5548);
and (n5552,n5553,n2744);
or (n5553,1'b0,n5554,n5557,n5560,n5563);
and (n5554,n5555,n5071);
wire s0n5555,s1n5555,notn5555;
or (n5555,s0n5555,s1n5555);
not(notn5555,n5069);
and (s0n5555,notn5555,n5556);
and (s1n5555,n5069,n5551);
and (n5557,n5558,n5083);
wire s0n5558,s1n5558,notn5558;
or (n5558,s0n5558,s1n5558);
not(notn5558,n5069);
and (s0n5558,notn5558,n5559);
and (s1n5558,n5069,n5556);
and (n5560,n5561,n5088);
wire s0n5561,s1n5561,notn5561;
or (n5561,s0n5561,s1n5561);
not(notn5561,n5069);
and (s0n5561,notn5561,n5562);
and (s1n5561,n5069,n5559);
and (n5563,n5564,n5093);
wire s0n5564,s1n5564,notn5564;
or (n5564,s0n5564,s1n5564);
not(notn5564,n5069);
and (s0n5564,notn5564,n5565);
and (s1n5564,n5069,n5562);
and (n5567,n5506,n5568);
or (n5568,n5569,n5690,n6060);
and (n5569,n5570,n5629);
wire s0n5570,s1n5570,notn5570;
or (n5570,s0n5570,s1n5570);
not(notn5570,n5021);
and (s0n5570,notn5570,n5571);
and (s1n5570,n5021,n5628);
or (n5571,1'b0,n5572,n5587,n5601,n5616);
and (n5572,n5573,n2710);
or (n5573,1'b0,n5574,n5578,n5581,n5584);
and (n5574,n5575,n5071);
wire s0n5575,s1n5575,notn5575;
or (n5575,s0n5575,s1n5575);
not(notn5575,n5069);
and (s0n5575,notn5575,n5576);
and (s1n5575,n5069,n5577);
and (n5578,n5579,n5083);
wire s0n5579,s1n5579,notn5579;
or (n5579,s0n5579,s1n5579);
not(notn5579,n5069);
and (s0n5579,notn5579,n5580);
and (s1n5579,n5069,n5576);
and (n5581,n5582,n5088);
wire s0n5582,s1n5582,notn5582;
or (n5582,s0n5582,s1n5582);
not(notn5582,n5069);
and (s0n5582,notn5582,n5583);
and (s1n5582,n5069,n5580);
and (n5584,n5585,n5093);
wire s0n5585,s1n5585,notn5585;
or (n5585,s0n5585,s1n5585);
not(notn5585,n5069);
and (s0n5585,notn5585,n5586);
and (s1n5585,n5069,n5583);
and (n5587,n5588,n2722);
or (n5588,1'b0,n5589,n5592,n5595,n5598);
and (n5589,n5590,n5071);
wire s0n5590,s1n5590,notn5590;
or (n5590,s0n5590,s1n5590);
not(notn5590,n5069);
and (s0n5590,notn5590,n5591);
and (s1n5590,n5069,n5586);
and (n5592,n5593,n5083);
wire s0n5593,s1n5593,notn5593;
or (n5593,s0n5593,s1n5593);
not(notn5593,n5069);
and (s0n5593,notn5593,n5594);
and (s1n5593,n5069,n5591);
and (n5595,n5596,n5088);
wire s0n5596,s1n5596,notn5596;
or (n5596,s0n5596,s1n5596);
not(notn5596,n5069);
and (s0n5596,notn5596,n5597);
and (s1n5596,n5069,n5594);
and (n5598,n5599,n5093);
wire s0n5599,s1n5599,notn5599;
or (n5599,s0n5599,s1n5599);
not(notn5599,n5069);
and (s0n5599,notn5599,n5600);
and (s1n5599,n5069,n5597);
and (n5601,n5602,n2734);
or (n5602,1'b0,n5603,n5607,n5610,n5613);
and (n5603,n5604,n5071);
wire s0n5604,s1n5604,notn5604;
or (n5604,s0n5604,s1n5604);
not(notn5604,n5069);
and (s0n5604,notn5604,n5605);
and (s1n5604,n5069,n5606);
and (n5607,n5608,n5083);
wire s0n5608,s1n5608,notn5608;
or (n5608,s0n5608,s1n5608);
not(notn5608,n5069);
and (s0n5608,notn5608,n5609);
and (s1n5608,n5069,n5605);
and (n5610,n5611,n5088);
wire s0n5611,s1n5611,notn5611;
or (n5611,s0n5611,s1n5611);
not(notn5611,n5069);
and (s0n5611,notn5611,n5612);
and (s1n5611,n5069,n5609);
and (n5613,n5614,n5093);
wire s0n5614,s1n5614,notn5614;
or (n5614,s0n5614,s1n5614);
not(notn5614,n5069);
and (s0n5614,notn5614,n5615);
and (s1n5614,n5069,n5612);
and (n5616,n5617,n2744);
or (n5617,1'b0,n5618,n5621,n5624,n5626);
and (n5618,n5619,n5071);
wire s0n5619,s1n5619,notn5619;
or (n5619,s0n5619,s1n5619);
not(notn5619,n5069);
and (s0n5619,notn5619,n5620);
and (s1n5619,n5069,n5615);
and (n5621,n5622,n5083);
wire s0n5622,s1n5622,notn5622;
or (n5622,s0n5622,s1n5622);
not(notn5622,n5069);
and (s0n5622,notn5622,n5623);
and (s1n5622,n5069,n5620);
and (n5624,n5625,n5088);
wire s0n5625,s1n5625,notn5625;
or (n5625,s0n5625,s1n5625);
not(notn5625,n5069);
and (s0n5625,notn5625,n2232);
and (s1n5625,n5069,n5623);
and (n5626,n5627,n5093);
wire s0n5627,s1n5627,notn5627;
or (n5627,s0n5627,s1n5627);
not(notn5627,n5069);
and (s0n5627,notn5627,n1917);
and (s1n5627,n5069,n2232);
wire s0n5629,s1n5629,notn5629;
or (n5629,s0n5629,s1n5629);
not(notn5629,n5021);
and (s0n5629,notn5629,n5630);
and (s1n5629,n5021,n5689);
or (n5630,1'b0,n5631,n5646,n5660,n5675);
and (n5631,n5632,n2710);
or (n5632,1'b0,n5633,n5637,n5640,n5643);
and (n5633,n5634,n5071);
wire s0n5634,s1n5634,notn5634;
or (n5634,s0n5634,s1n5634);
not(notn5634,n5069);
and (s0n5634,notn5634,n5635);
and (s1n5634,n5069,n5636);
and (n5637,n5638,n5083);
wire s0n5638,s1n5638,notn5638;
or (n5638,s0n5638,s1n5638);
not(notn5638,n5069);
and (s0n5638,notn5638,n5639);
and (s1n5638,n5069,n5635);
and (n5640,n5641,n5088);
wire s0n5641,s1n5641,notn5641;
or (n5641,s0n5641,s1n5641);
not(notn5641,n5069);
and (s0n5641,notn5641,n5642);
and (s1n5641,n5069,n5639);
and (n5643,n5644,n5093);
wire s0n5644,s1n5644,notn5644;
or (n5644,s0n5644,s1n5644);
not(notn5644,n5069);
and (s0n5644,notn5644,n5645);
and (s1n5644,n5069,n5642);
and (n5646,n5647,n2722);
or (n5647,1'b0,n5648,n5651,n5654,n5657);
and (n5648,n5649,n5071);
wire s0n5649,s1n5649,notn5649;
or (n5649,s0n5649,s1n5649);
not(notn5649,n5069);
and (s0n5649,notn5649,n5650);
and (s1n5649,n5069,n5645);
and (n5651,n5652,n5083);
wire s0n5652,s1n5652,notn5652;
or (n5652,s0n5652,s1n5652);
not(notn5652,n5069);
and (s0n5652,notn5652,n5653);
and (s1n5652,n5069,n5650);
and (n5654,n5655,n5088);
wire s0n5655,s1n5655,notn5655;
or (n5655,s0n5655,s1n5655);
not(notn5655,n5069);
and (s0n5655,notn5655,n5656);
and (s1n5655,n5069,n5653);
and (n5657,n5658,n5093);
wire s0n5658,s1n5658,notn5658;
or (n5658,s0n5658,s1n5658);
not(notn5658,n5069);
and (s0n5658,notn5658,n5659);
and (s1n5658,n5069,n5656);
and (n5660,n5661,n2734);
or (n5661,1'b0,n5662,n5666,n5669,n5672);
and (n5662,n5663,n5071);
wire s0n5663,s1n5663,notn5663;
or (n5663,s0n5663,s1n5663);
not(notn5663,n5069);
and (s0n5663,notn5663,n5664);
and (s1n5663,n5069,n5665);
and (n5666,n5667,n5083);
wire s0n5667,s1n5667,notn5667;
or (n5667,s0n5667,s1n5667);
not(notn5667,n5069);
and (s0n5667,notn5667,n5668);
and (s1n5667,n5069,n5664);
and (n5669,n5670,n5088);
wire s0n5670,s1n5670,notn5670;
or (n5670,s0n5670,s1n5670);
not(notn5670,n5069);
and (s0n5670,notn5670,n5671);
and (s1n5670,n5069,n5668);
and (n5672,n5673,n5093);
wire s0n5673,s1n5673,notn5673;
or (n5673,s0n5673,s1n5673);
not(notn5673,n5069);
and (s0n5673,notn5673,n5674);
and (s1n5673,n5069,n5671);
and (n5675,n5676,n2744);
or (n5676,1'b0,n5677,n5680,n5683,n5686);
and (n5677,n5678,n5071);
wire s0n5678,s1n5678,notn5678;
or (n5678,s0n5678,s1n5678);
not(notn5678,n5069);
and (s0n5678,notn5678,n5679);
and (s1n5678,n5069,n5674);
and (n5680,n5681,n5083);
wire s0n5681,s1n5681,notn5681;
or (n5681,s0n5681,s1n5681);
not(notn5681,n5069);
and (s0n5681,notn5681,n5682);
and (s1n5681,n5069,n5679);
and (n5683,n5684,n5088);
wire s0n5684,s1n5684,notn5684;
or (n5684,s0n5684,s1n5684);
not(notn5684,n5069);
and (s0n5684,notn5684,n5685);
and (s1n5684,n5069,n5682);
and (n5686,n5687,n5093);
wire s0n5687,s1n5687,notn5687;
or (n5687,s0n5687,s1n5687);
not(notn5687,n5069);
and (s0n5687,notn5687,n5688);
and (s1n5687,n5069,n5685);
and (n5690,n5629,n5691);
or (n5691,n5692,n5813,n6059);
and (n5692,n5693,n5752);
wire s0n5693,s1n5693,notn5693;
or (n5693,s0n5693,s1n5693);
not(notn5693,n5021);
and (s0n5693,notn5693,n5694);
and (s1n5693,n5021,n5751);
or (n5694,1'b0,n5695,n5710,n5724,n5739);
and (n5695,n5696,n2710);
or (n5696,1'b0,n5697,n5701,n5704,n5707);
and (n5697,n5698,n5071);
wire s0n5698,s1n5698,notn5698;
or (n5698,s0n5698,s1n5698);
not(notn5698,n5069);
and (s0n5698,notn5698,n5699);
and (s1n5698,n5069,n5700);
and (n5701,n5702,n5083);
wire s0n5702,s1n5702,notn5702;
or (n5702,s0n5702,s1n5702);
not(notn5702,n5069);
and (s0n5702,notn5702,n5703);
and (s1n5702,n5069,n5699);
and (n5704,n5705,n5088);
wire s0n5705,s1n5705,notn5705;
or (n5705,s0n5705,s1n5705);
not(notn5705,n5069);
and (s0n5705,notn5705,n5706);
and (s1n5705,n5069,n5703);
and (n5707,n5708,n5093);
wire s0n5708,s1n5708,notn5708;
or (n5708,s0n5708,s1n5708);
not(notn5708,n5069);
and (s0n5708,notn5708,n5709);
and (s1n5708,n5069,n5706);
and (n5710,n5711,n2722);
or (n5711,1'b0,n5712,n5715,n5718,n5721);
and (n5712,n5713,n5071);
wire s0n5713,s1n5713,notn5713;
or (n5713,s0n5713,s1n5713);
not(notn5713,n5069);
and (s0n5713,notn5713,n5714);
and (s1n5713,n5069,n5709);
and (n5715,n5716,n5083);
wire s0n5716,s1n5716,notn5716;
or (n5716,s0n5716,s1n5716);
not(notn5716,n5069);
and (s0n5716,notn5716,n5717);
and (s1n5716,n5069,n5714);
and (n5718,n5719,n5088);
wire s0n5719,s1n5719,notn5719;
or (n5719,s0n5719,s1n5719);
not(notn5719,n5069);
and (s0n5719,notn5719,n5720);
and (s1n5719,n5069,n5717);
and (n5721,n5722,n5093);
wire s0n5722,s1n5722,notn5722;
or (n5722,s0n5722,s1n5722);
not(notn5722,n5069);
and (s0n5722,notn5722,n5723);
and (s1n5722,n5069,n5720);
and (n5724,n5725,n2734);
or (n5725,1'b0,n5726,n5730,n5733,n5736);
and (n5726,n5727,n5071);
wire s0n5727,s1n5727,notn5727;
or (n5727,s0n5727,s1n5727);
not(notn5727,n5069);
and (s0n5727,notn5727,n5728);
and (s1n5727,n5069,n5729);
and (n5730,n5731,n5083);
wire s0n5731,s1n5731,notn5731;
or (n5731,s0n5731,s1n5731);
not(notn5731,n5069);
and (s0n5731,notn5731,n5732);
and (s1n5731,n5069,n5728);
and (n5733,n5734,n5088);
wire s0n5734,s1n5734,notn5734;
or (n5734,s0n5734,s1n5734);
not(notn5734,n5069);
and (s0n5734,notn5734,n5735);
and (s1n5734,n5069,n5732);
and (n5736,n5737,n5093);
wire s0n5737,s1n5737,notn5737;
or (n5737,s0n5737,s1n5737);
not(notn5737,n5069);
and (s0n5737,notn5737,n5738);
and (s1n5737,n5069,n5735);
and (n5739,n5740,n2744);
or (n5740,1'b0,n5741,n5744,n5747,n5749);
and (n5741,n5742,n5071);
wire s0n5742,s1n5742,notn5742;
or (n5742,s0n5742,s1n5742);
not(notn5742,n5069);
and (s0n5742,notn5742,n5743);
and (s1n5742,n5069,n5738);
and (n5744,n5745,n5083);
wire s0n5745,s1n5745,notn5745;
or (n5745,s0n5745,s1n5745);
not(notn5745,n5069);
and (s0n5745,notn5745,n5746);
and (s1n5745,n5069,n5743);
and (n5747,n5748,n5088);
wire s0n5748,s1n5748,notn5748;
or (n5748,s0n5748,s1n5748);
not(notn5748,n5069);
and (s0n5748,notn5748,n2248);
and (s1n5748,n5069,n5746);
and (n5749,n5750,n5093);
wire s0n5750,s1n5750,notn5750;
or (n5750,s0n5750,s1n5750);
not(notn5750,n5069);
and (s0n5750,notn5750,n1943);
and (s1n5750,n5069,n2248);
wire s0n5752,s1n5752,notn5752;
or (n5752,s0n5752,s1n5752);
not(notn5752,n5021);
and (s0n5752,notn5752,n5753);
and (s1n5752,n5021,n5812);
or (n5753,1'b0,n5754,n5769,n5783,n5798);
and (n5754,n5755,n2710);
or (n5755,1'b0,n5756,n5760,n5763,n5766);
and (n5756,n5757,n5071);
wire s0n5757,s1n5757,notn5757;
or (n5757,s0n5757,s1n5757);
not(notn5757,n5069);
and (s0n5757,notn5757,n5758);
and (s1n5757,n5069,n5759);
and (n5760,n5761,n5083);
wire s0n5761,s1n5761,notn5761;
or (n5761,s0n5761,s1n5761);
not(notn5761,n5069);
and (s0n5761,notn5761,n5762);
and (s1n5761,n5069,n5758);
and (n5763,n5764,n5088);
wire s0n5764,s1n5764,notn5764;
or (n5764,s0n5764,s1n5764);
not(notn5764,n5069);
and (s0n5764,notn5764,n5765);
and (s1n5764,n5069,n5762);
and (n5766,n5767,n5093);
wire s0n5767,s1n5767,notn5767;
or (n5767,s0n5767,s1n5767);
not(notn5767,n5069);
and (s0n5767,notn5767,n5768);
and (s1n5767,n5069,n5765);
and (n5769,n5770,n2722);
or (n5770,1'b0,n5771,n5774,n5777,n5780);
and (n5771,n5772,n5071);
wire s0n5772,s1n5772,notn5772;
or (n5772,s0n5772,s1n5772);
not(notn5772,n5069);
and (s0n5772,notn5772,n5773);
and (s1n5772,n5069,n5768);
and (n5774,n5775,n5083);
wire s0n5775,s1n5775,notn5775;
or (n5775,s0n5775,s1n5775);
not(notn5775,n5069);
and (s0n5775,notn5775,n5776);
and (s1n5775,n5069,n5773);
and (n5777,n5778,n5088);
wire s0n5778,s1n5778,notn5778;
or (n5778,s0n5778,s1n5778);
not(notn5778,n5069);
and (s0n5778,notn5778,n5779);
and (s1n5778,n5069,n5776);
and (n5780,n5781,n5093);
wire s0n5781,s1n5781,notn5781;
or (n5781,s0n5781,s1n5781);
not(notn5781,n5069);
and (s0n5781,notn5781,n5782);
and (s1n5781,n5069,n5779);
and (n5783,n5784,n2734);
or (n5784,1'b0,n5785,n5789,n5792,n5795);
and (n5785,n5786,n5071);
wire s0n5786,s1n5786,notn5786;
or (n5786,s0n5786,s1n5786);
not(notn5786,n5069);
and (s0n5786,notn5786,n5787);
and (s1n5786,n5069,n5788);
and (n5789,n5790,n5083);
wire s0n5790,s1n5790,notn5790;
or (n5790,s0n5790,s1n5790);
not(notn5790,n5069);
and (s0n5790,notn5790,n5791);
and (s1n5790,n5069,n5787);
and (n5792,n5793,n5088);
wire s0n5793,s1n5793,notn5793;
or (n5793,s0n5793,s1n5793);
not(notn5793,n5069);
and (s0n5793,notn5793,n5794);
and (s1n5793,n5069,n5791);
and (n5795,n5796,n5093);
wire s0n5796,s1n5796,notn5796;
or (n5796,s0n5796,s1n5796);
not(notn5796,n5069);
and (s0n5796,notn5796,n5797);
and (s1n5796,n5069,n5794);
and (n5798,n5799,n2744);
or (n5799,1'b0,n5800,n5803,n5806,n5809);
and (n5800,n5801,n5071);
wire s0n5801,s1n5801,notn5801;
or (n5801,s0n5801,s1n5801);
not(notn5801,n5069);
and (s0n5801,notn5801,n5802);
and (s1n5801,n5069,n5797);
and (n5803,n5804,n5083);
wire s0n5804,s1n5804,notn5804;
or (n5804,s0n5804,s1n5804);
not(notn5804,n5069);
and (s0n5804,notn5804,n5805);
and (s1n5804,n5069,n5802);
and (n5806,n5807,n5088);
wire s0n5807,s1n5807,notn5807;
or (n5807,s0n5807,s1n5807);
not(notn5807,n5069);
and (s0n5807,notn5807,n5808);
and (s1n5807,n5069,n5805);
and (n5809,n5810,n5093);
wire s0n5810,s1n5810,notn5810;
or (n5810,s0n5810,s1n5810);
not(notn5810,n5069);
and (s0n5810,notn5810,n5811);
and (s1n5810,n5069,n5808);
and (n5813,n5752,n5814);
or (n5814,n5815,n5936,n6058);
and (n5815,n5816,n5875);
wire s0n5816,s1n5816,notn5816;
or (n5816,s0n5816,s1n5816);
not(notn5816,n5021);
and (s0n5816,notn5816,n5817);
and (s1n5816,n5021,n5874);
or (n5817,1'b0,n5818,n5833,n5847,n5862);
and (n5818,n5819,n2710);
or (n5819,1'b0,n5820,n5824,n5827,n5830);
and (n5820,n5821,n5071);
wire s0n5821,s1n5821,notn5821;
or (n5821,s0n5821,s1n5821);
not(notn5821,n5069);
and (s0n5821,notn5821,n5822);
and (s1n5821,n5069,n5823);
and (n5824,n5825,n5083);
wire s0n5825,s1n5825,notn5825;
or (n5825,s0n5825,s1n5825);
not(notn5825,n5069);
and (s0n5825,notn5825,n5826);
and (s1n5825,n5069,n5822);
and (n5827,n5828,n5088);
wire s0n5828,s1n5828,notn5828;
or (n5828,s0n5828,s1n5828);
not(notn5828,n5069);
and (s0n5828,notn5828,n5829);
and (s1n5828,n5069,n5826);
and (n5830,n5831,n5093);
wire s0n5831,s1n5831,notn5831;
or (n5831,s0n5831,s1n5831);
not(notn5831,n5069);
and (s0n5831,notn5831,n5832);
and (s1n5831,n5069,n5829);
and (n5833,n5834,n2722);
or (n5834,1'b0,n5835,n5838,n5841,n5844);
and (n5835,n5836,n5071);
wire s0n5836,s1n5836,notn5836;
or (n5836,s0n5836,s1n5836);
not(notn5836,n5069);
and (s0n5836,notn5836,n5837);
and (s1n5836,n5069,n5832);
and (n5838,n5839,n5083);
wire s0n5839,s1n5839,notn5839;
or (n5839,s0n5839,s1n5839);
not(notn5839,n5069);
and (s0n5839,notn5839,n5840);
and (s1n5839,n5069,n5837);
and (n5841,n5842,n5088);
wire s0n5842,s1n5842,notn5842;
or (n5842,s0n5842,s1n5842);
not(notn5842,n5069);
and (s0n5842,notn5842,n5843);
and (s1n5842,n5069,n5840);
and (n5844,n5845,n5093);
wire s0n5845,s1n5845,notn5845;
or (n5845,s0n5845,s1n5845);
not(notn5845,n5069);
and (s0n5845,notn5845,n5846);
and (s1n5845,n5069,n5843);
and (n5847,n5848,n2734);
or (n5848,1'b0,n5849,n5853,n5856,n5859);
and (n5849,n5850,n5071);
wire s0n5850,s1n5850,notn5850;
or (n5850,s0n5850,s1n5850);
not(notn5850,n5069);
and (s0n5850,notn5850,n5851);
and (s1n5850,n5069,n5852);
and (n5853,n5854,n5083);
wire s0n5854,s1n5854,notn5854;
or (n5854,s0n5854,s1n5854);
not(notn5854,n5069);
and (s0n5854,notn5854,n5855);
and (s1n5854,n5069,n5851);
and (n5856,n5857,n5088);
wire s0n5857,s1n5857,notn5857;
or (n5857,s0n5857,s1n5857);
not(notn5857,n5069);
and (s0n5857,notn5857,n5858);
and (s1n5857,n5069,n5855);
and (n5859,n5860,n5093);
wire s0n5860,s1n5860,notn5860;
or (n5860,s0n5860,s1n5860);
not(notn5860,n5069);
and (s0n5860,notn5860,n5861);
and (s1n5860,n5069,n5858);
and (n5862,n5863,n2744);
or (n5863,1'b0,n5864,n5867,n5870,n5872);
and (n5864,n5865,n5071);
wire s0n5865,s1n5865,notn5865;
or (n5865,s0n5865,s1n5865);
not(notn5865,n5069);
and (s0n5865,notn5865,n5866);
and (s1n5865,n5069,n5861);
and (n5867,n5868,n5083);
wire s0n5868,s1n5868,notn5868;
or (n5868,s0n5868,s1n5868);
not(notn5868,n5069);
and (s0n5868,notn5868,n5869);
and (s1n5868,n5069,n5866);
and (n5870,n5871,n5088);
wire s0n5871,s1n5871,notn5871;
or (n5871,s0n5871,s1n5871);
not(notn5871,n5069);
and (s0n5871,notn5871,n2264);
and (s1n5871,n5069,n5869);
and (n5872,n5873,n5093);
wire s0n5873,s1n5873,notn5873;
or (n5873,s0n5873,s1n5873);
not(notn5873,n5069);
and (s0n5873,notn5873,n1972);
and (s1n5873,n5069,n2264);
wire s0n5875,s1n5875,notn5875;
or (n5875,s0n5875,s1n5875);
not(notn5875,n5021);
and (s0n5875,notn5875,n5876);
and (s1n5875,n5021,n5935);
or (n5876,1'b0,n5877,n5892,n5906,n5921);
and (n5877,n5878,n2710);
or (n5878,1'b0,n5879,n5883,n5886,n5889);
and (n5879,n5880,n5071);
wire s0n5880,s1n5880,notn5880;
or (n5880,s0n5880,s1n5880);
not(notn5880,n5069);
and (s0n5880,notn5880,n5881);
and (s1n5880,n5069,n5882);
and (n5883,n5884,n5083);
wire s0n5884,s1n5884,notn5884;
or (n5884,s0n5884,s1n5884);
not(notn5884,n5069);
and (s0n5884,notn5884,n5885);
and (s1n5884,n5069,n5881);
and (n5886,n5887,n5088);
wire s0n5887,s1n5887,notn5887;
or (n5887,s0n5887,s1n5887);
not(notn5887,n5069);
and (s0n5887,notn5887,n5888);
and (s1n5887,n5069,n5885);
and (n5889,n5890,n5093);
wire s0n5890,s1n5890,notn5890;
or (n5890,s0n5890,s1n5890);
not(notn5890,n5069);
and (s0n5890,notn5890,n5891);
and (s1n5890,n5069,n5888);
and (n5892,n5893,n2722);
or (n5893,1'b0,n5894,n5897,n5900,n5903);
and (n5894,n5895,n5071);
wire s0n5895,s1n5895,notn5895;
or (n5895,s0n5895,s1n5895);
not(notn5895,n5069);
and (s0n5895,notn5895,n5896);
and (s1n5895,n5069,n5891);
and (n5897,n5898,n5083);
wire s0n5898,s1n5898,notn5898;
or (n5898,s0n5898,s1n5898);
not(notn5898,n5069);
and (s0n5898,notn5898,n5899);
and (s1n5898,n5069,n5896);
and (n5900,n5901,n5088);
wire s0n5901,s1n5901,notn5901;
or (n5901,s0n5901,s1n5901);
not(notn5901,n5069);
and (s0n5901,notn5901,n5902);
and (s1n5901,n5069,n5899);
and (n5903,n5904,n5093);
wire s0n5904,s1n5904,notn5904;
or (n5904,s0n5904,s1n5904);
not(notn5904,n5069);
and (s0n5904,notn5904,n5905);
and (s1n5904,n5069,n5902);
and (n5906,n5907,n2734);
or (n5907,1'b0,n5908,n5912,n5915,n5918);
and (n5908,n5909,n5071);
wire s0n5909,s1n5909,notn5909;
or (n5909,s0n5909,s1n5909);
not(notn5909,n5069);
and (s0n5909,notn5909,n5910);
and (s1n5909,n5069,n5911);
and (n5912,n5913,n5083);
wire s0n5913,s1n5913,notn5913;
or (n5913,s0n5913,s1n5913);
not(notn5913,n5069);
and (s0n5913,notn5913,n5914);
and (s1n5913,n5069,n5910);
and (n5915,n5916,n5088);
wire s0n5916,s1n5916,notn5916;
or (n5916,s0n5916,s1n5916);
not(notn5916,n5069);
and (s0n5916,notn5916,n5917);
and (s1n5916,n5069,n5914);
and (n5918,n5919,n5093);
wire s0n5919,s1n5919,notn5919;
or (n5919,s0n5919,s1n5919);
not(notn5919,n5069);
and (s0n5919,notn5919,n5920);
and (s1n5919,n5069,n5917);
and (n5921,n5922,n2744);
or (n5922,1'b0,n5923,n5926,n5929,n5932);
and (n5923,n5924,n5071);
wire s0n5924,s1n5924,notn5924;
or (n5924,s0n5924,s1n5924);
not(notn5924,n5069);
and (s0n5924,notn5924,n5925);
and (s1n5924,n5069,n5920);
and (n5926,n5927,n5083);
wire s0n5927,s1n5927,notn5927;
or (n5927,s0n5927,s1n5927);
not(notn5927,n5069);
and (s0n5927,notn5927,n5928);
and (s1n5927,n5069,n5925);
and (n5929,n5930,n5088);
wire s0n5930,s1n5930,notn5930;
or (n5930,s0n5930,s1n5930);
not(notn5930,n5069);
and (s0n5930,notn5930,n5931);
and (s1n5930,n5069,n5928);
and (n5932,n5933,n5093);
wire s0n5933,s1n5933,notn5933;
or (n5933,s0n5933,s1n5933);
not(notn5933,n5069);
and (s0n5933,notn5933,n5934);
and (s1n5933,n5069,n5931);
and (n5936,n5875,n5937);
and (n5937,n5938,n5997);
wire s0n5938,s1n5938,notn5938;
or (n5938,s0n5938,s1n5938);
not(notn5938,n5021);
and (s0n5938,notn5938,n5939);
and (s1n5938,n5021,n5996);
or (n5939,1'b0,n5940,n5955,n5969,n5984);
and (n5940,n5941,n2710);
or (n5941,1'b0,n5942,n5946,n5949,n5952);
and (n5942,n5943,n5071);
wire s0n5943,s1n5943,notn5943;
or (n5943,s0n5943,s1n5943);
not(notn5943,n5069);
and (s0n5943,notn5943,n5944);
and (s1n5943,n5069,n5945);
and (n5946,n5947,n5083);
wire s0n5947,s1n5947,notn5947;
or (n5947,s0n5947,s1n5947);
not(notn5947,n5069);
and (s0n5947,notn5947,n5948);
and (s1n5947,n5069,n5944);
and (n5949,n5950,n5088);
wire s0n5950,s1n5950,notn5950;
or (n5950,s0n5950,s1n5950);
not(notn5950,n5069);
and (s0n5950,notn5950,n5951);
and (s1n5950,n5069,n5948);
and (n5952,n5953,n5093);
wire s0n5953,s1n5953,notn5953;
or (n5953,s0n5953,s1n5953);
not(notn5953,n5069);
and (s0n5953,notn5953,n5954);
and (s1n5953,n5069,n5951);
and (n5955,n5956,n2722);
or (n5956,1'b0,n5957,n5960,n5963,n5966);
and (n5957,n5958,n5071);
wire s0n5958,s1n5958,notn5958;
or (n5958,s0n5958,s1n5958);
not(notn5958,n5069);
and (s0n5958,notn5958,n5959);
and (s1n5958,n5069,n5954);
and (n5960,n5961,n5083);
wire s0n5961,s1n5961,notn5961;
or (n5961,s0n5961,s1n5961);
not(notn5961,n5069);
and (s0n5961,notn5961,n5962);
and (s1n5961,n5069,n5959);
and (n5963,n5964,n5088);
wire s0n5964,s1n5964,notn5964;
or (n5964,s0n5964,s1n5964);
not(notn5964,n5069);
and (s0n5964,notn5964,n5965);
and (s1n5964,n5069,n5962);
and (n5966,n5967,n5093);
wire s0n5967,s1n5967,notn5967;
or (n5967,s0n5967,s1n5967);
not(notn5967,n5069);
and (s0n5967,notn5967,n5968);
and (s1n5967,n5069,n5965);
and (n5969,n5970,n2734);
or (n5970,1'b0,n5971,n5975,n5978,n5981);
and (n5971,n5972,n5071);
wire s0n5972,s1n5972,notn5972;
or (n5972,s0n5972,s1n5972);
not(notn5972,n5069);
and (s0n5972,notn5972,n5973);
and (s1n5972,n5069,n5974);
and (n5975,n5976,n5083);
wire s0n5976,s1n5976,notn5976;
or (n5976,s0n5976,s1n5976);
not(notn5976,n5069);
and (s0n5976,notn5976,n5977);
and (s1n5976,n5069,n5973);
and (n5978,n5979,n5088);
wire s0n5979,s1n5979,notn5979;
or (n5979,s0n5979,s1n5979);
not(notn5979,n5069);
and (s0n5979,notn5979,n5980);
and (s1n5979,n5069,n5977);
and (n5981,n5982,n5093);
wire s0n5982,s1n5982,notn5982;
or (n5982,s0n5982,s1n5982);
not(notn5982,n5069);
and (s0n5982,notn5982,n5983);
and (s1n5982,n5069,n5980);
and (n5984,n5985,n2744);
or (n5985,1'b0,n5986,n5989,n5992,n5994);
and (n5986,n5987,n5071);
wire s0n5987,s1n5987,notn5987;
or (n5987,s0n5987,s1n5987);
not(notn5987,n5069);
and (s0n5987,notn5987,n5988);
and (s1n5987,n5069,n5983);
and (n5989,n5990,n5083);
wire s0n5990,s1n5990,notn5990;
or (n5990,s0n5990,s1n5990);
not(notn5990,n5069);
and (s0n5990,notn5990,n5991);
and (s1n5990,n5069,n5988);
and (n5992,n5993,n5088);
wire s0n5993,s1n5993,notn5993;
or (n5993,s0n5993,s1n5993);
not(notn5993,n5069);
and (s0n5993,notn5993,n2279);
and (s1n5993,n5069,n5991);
and (n5994,n5995,n5093);
wire s0n5995,s1n5995,notn5995;
or (n5995,s0n5995,s1n5995);
not(notn5995,n5069);
and (s0n5995,notn5995,n1991);
and (s1n5995,n5069,n2279);
wire s0n5997,s1n5997,notn5997;
or (n5997,s0n5997,s1n5997);
not(notn5997,n5021);
and (s0n5997,notn5997,n5998);
and (s1n5997,n5021,n6057);
or (n5998,1'b0,n5999,n6014,n6028,n6043);
and (n5999,n6000,n2710);
or (n6000,1'b0,n6001,n6005,n6008,n6011);
and (n6001,n6002,n5071);
wire s0n6002,s1n6002,notn6002;
or (n6002,s0n6002,s1n6002);
not(notn6002,n5069);
and (s0n6002,notn6002,n6003);
and (s1n6002,n5069,n6004);
and (n6005,n6006,n5083);
wire s0n6006,s1n6006,notn6006;
or (n6006,s0n6006,s1n6006);
not(notn6006,n5069);
and (s0n6006,notn6006,n6007);
and (s1n6006,n5069,n6003);
and (n6008,n6009,n5088);
wire s0n6009,s1n6009,notn6009;
or (n6009,s0n6009,s1n6009);
not(notn6009,n5069);
and (s0n6009,notn6009,n6010);
and (s1n6009,n5069,n6007);
and (n6011,n6012,n5093);
wire s0n6012,s1n6012,notn6012;
or (n6012,s0n6012,s1n6012);
not(notn6012,n5069);
and (s0n6012,notn6012,n6013);
and (s1n6012,n5069,n6010);
and (n6014,n6015,n2722);
or (n6015,1'b0,n6016,n6019,n6022,n6025);
and (n6016,n6017,n5071);
wire s0n6017,s1n6017,notn6017;
or (n6017,s0n6017,s1n6017);
not(notn6017,n5069);
and (s0n6017,notn6017,n6018);
and (s1n6017,n5069,n6013);
and (n6019,n6020,n5083);
wire s0n6020,s1n6020,notn6020;
or (n6020,s0n6020,s1n6020);
not(notn6020,n5069);
and (s0n6020,notn6020,n6021);
and (s1n6020,n5069,n6018);
and (n6022,n6023,n5088);
wire s0n6023,s1n6023,notn6023;
or (n6023,s0n6023,s1n6023);
not(notn6023,n5069);
and (s0n6023,notn6023,n6024);
and (s1n6023,n5069,n6021);
and (n6025,n6026,n5093);
wire s0n6026,s1n6026,notn6026;
or (n6026,s0n6026,s1n6026);
not(notn6026,n5069);
and (s0n6026,notn6026,n6027);
and (s1n6026,n5069,n6024);
and (n6028,n6029,n2734);
or (n6029,1'b0,n6030,n6034,n6037,n6040);
and (n6030,n6031,n5071);
wire s0n6031,s1n6031,notn6031;
or (n6031,s0n6031,s1n6031);
not(notn6031,n5069);
and (s0n6031,notn6031,n6032);
and (s1n6031,n5069,n6033);
and (n6034,n6035,n5083);
wire s0n6035,s1n6035,notn6035;
or (n6035,s0n6035,s1n6035);
not(notn6035,n5069);
and (s0n6035,notn6035,n6036);
and (s1n6035,n5069,n6032);
and (n6037,n6038,n5088);
wire s0n6038,s1n6038,notn6038;
or (n6038,s0n6038,s1n6038);
not(notn6038,n5069);
and (s0n6038,notn6038,n6039);
and (s1n6038,n5069,n6036);
and (n6040,n6041,n5093);
wire s0n6041,s1n6041,notn6041;
or (n6041,s0n6041,s1n6041);
not(notn6041,n5069);
and (s0n6041,notn6041,n6042);
and (s1n6041,n5069,n6039);
and (n6043,n6044,n2744);
or (n6044,1'b0,n6045,n6048,n6051,n6054);
and (n6045,n6046,n5071);
wire s0n6046,s1n6046,notn6046;
or (n6046,s0n6046,s1n6046);
not(notn6046,n5069);
and (s0n6046,notn6046,n6047);
and (s1n6046,n5069,n6042);
and (n6048,n6049,n5083);
wire s0n6049,s1n6049,notn6049;
or (n6049,s0n6049,s1n6049);
not(notn6049,n5069);
and (s0n6049,notn6049,n6050);
and (s1n6049,n5069,n6047);
and (n6051,n6052,n5088);
wire s0n6052,s1n6052,notn6052;
or (n6052,s0n6052,s1n6052);
not(notn6052,n5069);
and (s0n6052,notn6052,n6053);
and (s1n6052,n5069,n6050);
and (n6054,n6055,n5093);
wire s0n6055,s1n6055,notn6055;
or (n6055,s0n6055,s1n6055);
not(notn6055,n5069);
and (s0n6055,notn6055,n6056);
and (s1n6055,n5069,n6053);
and (n6058,n5816,n5937);
and (n6059,n5693,n5814);
and (n6060,n5570,n5691);
and (n6061,n5447,n5568);
and (n6062,n5324,n5445);
and (n6063,n5201,n5322);
and (n6064,n5061,n5199);
and (n6065,n5054,n5059);
and (n6066,n5047,n5052);
and (n6067,n5040,n5045);
and (n6068,n5033,n5038);
xor (n6069,n6070,n7580);
xor (n6070,n6071,n7421);
xor (n6071,n6072,n6811);
xor (n6072,n6073,n6078);
xor (n6073,n6074,n6076);
wire s0n6074,s1n6074,notn6074;
or (n6074,s0n6074,s1n6074);
not(notn6074,n5021);
and (s0n6074,notn6074,1'b0);
and (s1n6074,n5021,n6075);
wire s0n6076,s1n6076,notn6076;
or (n6076,s0n6076,s1n6076);
not(notn6076,n5021);
and (s0n6076,notn6076,1'b0);
and (s1n6076,n5021,n6077);
or (n6078,n6079,n6084,n6810);
and (n6079,n6080,n6082);
wire s0n6080,s1n6080,notn6080;
or (n6080,s0n6080,s1n6080);
not(notn6080,n5021);
and (s0n6080,notn6080,1'b0);
and (s1n6080,n5021,n6081);
wire s0n6082,s1n6082,notn6082;
or (n6082,s0n6082,s1n6082);
not(notn6082,n5021);
and (s0n6082,notn6082,1'b0);
and (s1n6082,n5021,n6083);
and (n6084,n6082,n6085);
or (n6085,n6086,n6091,n6809);
and (n6086,n6087,n6089);
wire s0n6087,s1n6087,notn6087;
or (n6087,s0n6087,s1n6087);
not(notn6087,n5021);
and (s0n6087,notn6087,1'b0);
and (s1n6087,n5021,n6088);
wire s0n6089,s1n6089,notn6089;
or (n6089,s0n6089,s1n6089);
not(notn6089,n5021);
and (s0n6089,notn6089,1'b0);
and (s1n6089,n5021,n6090);
and (n6091,n6089,n6092);
or (n6092,n6093,n6180,n6808);
and (n6093,n6094,n6137);
wire s0n6094,s1n6094,notn6094;
or (n6094,s0n6094,s1n6094);
not(notn6094,n5021);
and (s0n6094,notn6094,n6095);
and (s1n6094,n5021,n6136);
or (n6095,1'b0,n6096,n6106,n6116,n6126);
and (n6096,n6097,n2710);
or (n6097,1'b0,n6098,n6100,n6102,n6104);
and (n6098,n6099,n5071);
wire s0n6099,s1n6099,notn6099;
or (n6099,s0n6099,s1n6099);
not(notn6099,n5069);
and (s0n6099,notn6099,n2703);
and (s1n6099,n5069,n3017);
and (n6100,n6101,n5083);
wire s0n6101,s1n6101,notn6101;
or (n6101,s0n6101,s1n6101);
not(notn6101,n5069);
and (s0n6101,notn6101,n2705);
and (s1n6101,n5069,n2703);
and (n6102,n6103,n5088);
wire s0n6103,s1n6103,notn6103;
or (n6103,s0n6103,s1n6103);
not(notn6103,n5069);
and (s0n6103,notn6103,n2707);
and (s1n6103,n5069,n2705);
and (n6104,n6105,n5093);
wire s0n6105,s1n6105,notn6105;
or (n6105,s0n6105,s1n6105);
not(notn6105,n5069);
and (s0n6105,notn6105,n2709);
and (s1n6105,n5069,n2707);
and (n6106,n6107,n2722);
or (n6107,1'b0,n6108,n6110,n6112,n6114);
and (n6108,n6109,n5071);
wire s0n6109,s1n6109,notn6109;
or (n6109,s0n6109,s1n6109);
not(notn6109,n5069);
and (s0n6109,notn6109,n2715);
and (s1n6109,n5069,n2709);
and (n6110,n6111,n5083);
wire s0n6111,s1n6111,notn6111;
or (n6111,s0n6111,s1n6111);
not(notn6111,n5069);
and (s0n6111,notn6111,n2717);
and (s1n6111,n5069,n2715);
and (n6112,n6113,n5088);
wire s0n6113,s1n6113,notn6113;
or (n6113,s0n6113,s1n6113);
not(notn6113,n5069);
and (s0n6113,notn6113,n2719);
and (s1n6113,n5069,n2717);
and (n6114,n6115,n5093);
wire s0n6115,s1n6115,notn6115;
or (n6115,s0n6115,s1n6115);
not(notn6115,n5069);
and (s0n6115,notn6115,n2721);
and (s1n6115,n5069,n2719);
and (n6116,n6117,n2734);
or (n6117,1'b0,n6118,n6120,n6122,n6124);
and (n6118,n6119,n5071);
wire s0n6119,s1n6119,notn6119;
or (n6119,s0n6119,s1n6119);
not(notn6119,n5069);
and (s0n6119,notn6119,n2727);
and (s1n6119,n5069,n3032);
and (n6120,n6121,n5083);
wire s0n6121,s1n6121,notn6121;
or (n6121,s0n6121,s1n6121);
not(notn6121,n5069);
and (s0n6121,notn6121,n2729);
and (s1n6121,n5069,n2727);
and (n6122,n6123,n5088);
wire s0n6123,s1n6123,notn6123;
or (n6123,s0n6123,s1n6123);
not(notn6123,n5069);
and (s0n6123,notn6123,n2731);
and (s1n6123,n5069,n2729);
and (n6124,n6125,n5093);
wire s0n6125,s1n6125,notn6125;
or (n6125,s0n6125,s1n6125);
not(notn6125,n5069);
and (s0n6125,notn6125,n2733);
and (s1n6125,n5069,n2731);
and (n6126,n6127,n2744);
or (n6127,1'b0,n6128,n6130,n6132,n6134);
and (n6128,n6129,n5071);
wire s0n6129,s1n6129,notn6129;
or (n6129,s0n6129,s1n6129);
not(notn6129,n5069);
and (s0n6129,notn6129,n2739);
and (s1n6129,n5069,n2733);
and (n6130,n6131,n5083);
wire s0n6131,s1n6131,notn6131;
or (n6131,s0n6131,s1n6131);
not(notn6131,n5069);
and (s0n6131,notn6131,n2741);
and (s1n6131,n5069,n2739);
and (n6132,n6133,n5088);
wire s0n6133,s1n6133,notn6133;
or (n6133,s0n6133,s1n6133);
not(notn6133,n5069);
and (s0n6133,notn6133,n2164);
and (s1n6133,n5069,n2741);
and (n6134,n6135,n5093);
wire s0n6135,s1n6135,notn6135;
or (n6135,s0n6135,s1n6135);
not(notn6135,n5069);
and (s0n6135,notn6135,n1827);
and (s1n6135,n5069,n2164);
wire s0n6137,s1n6137,notn6137;
or (n6137,s0n6137,s1n6137);
not(notn6137,n5021);
and (s0n6137,notn6137,n6138);
and (s1n6137,n5021,n6179);
or (n6138,1'b0,n6139,n6149,n6159,n6169);
and (n6139,n6140,n2710);
or (n6140,1'b0,n6141,n6143,n6145,n6147);
and (n6141,n6142,n5071);
wire s0n6142,s1n6142,notn6142;
or (n6142,s0n6142,s1n6142);
not(notn6142,n5069);
and (s0n6142,notn6142,n2920);
and (s1n6142,n5069,n3018);
and (n6143,n6144,n5083);
wire s0n6144,s1n6144,notn6144;
or (n6144,s0n6144,s1n6144);
not(notn6144,n5069);
and (s0n6144,notn6144,n2946);
and (s1n6144,n5069,n2920);
and (n6145,n6146,n5088);
wire s0n6146,s1n6146,notn6146;
or (n6146,s0n6146,s1n6146);
not(notn6146,n5069);
and (s0n6146,notn6146,n2954);
and (s1n6146,n5069,n2946);
and (n6147,n6148,n5093);
wire s0n6148,s1n6148,notn6148;
or (n6148,s0n6148,s1n6148);
not(notn6148,n5069);
and (s0n6148,notn6148,n2963);
and (s1n6148,n5069,n2954);
and (n6149,n6150,n2722);
or (n6150,1'b0,n6151,n6153,n6155,n6157);
and (n6151,n6152,n5071);
wire s0n6152,s1n6152,notn6152;
or (n6152,s0n6152,s1n6152);
not(notn6152,n5069);
and (s0n6152,notn6152,n2974);
and (s1n6152,n5069,n2963);
and (n6153,n6154,n5083);
wire s0n6154,s1n6154,notn6154;
or (n6154,s0n6154,s1n6154);
not(notn6154,n5069);
and (s0n6154,notn6154,n2977);
and (s1n6154,n5069,n2974);
and (n6155,n6156,n5088);
wire s0n6156,s1n6156,notn6156;
or (n6156,s0n6156,s1n6156);
not(notn6156,n5069);
and (s0n6156,notn6156,n2980);
and (s1n6156,n5069,n2977);
and (n6157,n6158,n5093);
wire s0n6158,s1n6158,notn6158;
or (n6158,s0n6158,s1n6158);
not(notn6158,n5069);
and (s0n6158,notn6158,n2983);
and (s1n6158,n5069,n2980);
and (n6159,n6160,n2734);
or (n6160,1'b0,n6161,n6163,n6165,n6167);
and (n6161,n6162,n5071);
wire s0n6162,s1n6162,notn6162;
or (n6162,s0n6162,s1n6162);
not(notn6162,n5069);
and (s0n6162,notn6162,n2988);
and (s1n6162,n5069,n3033);
and (n6163,n6164,n5083);
wire s0n6164,s1n6164,notn6164;
or (n6164,s0n6164,s1n6164);
not(notn6164,n5069);
and (s0n6164,notn6164,n2991);
and (s1n6164,n5069,n2988);
and (n6165,n6166,n5088);
wire s0n6166,s1n6166,notn6166;
or (n6166,s0n6166,s1n6166);
not(notn6166,n5069);
and (s0n6166,notn6166,n2994);
and (s1n6166,n5069,n2991);
and (n6167,n6168,n5093);
wire s0n6168,s1n6168,notn6168;
or (n6168,s0n6168,s1n6168);
not(notn6168,n5069);
and (s0n6168,notn6168,n2997);
and (s1n6168,n5069,n2994);
and (n6169,n6170,n2744);
or (n6170,1'b0,n6171,n6173,n6175,n6177);
and (n6171,n6172,n5071);
wire s0n6172,s1n6172,notn6172;
or (n6172,s0n6172,s1n6172);
not(notn6172,n5069);
and (s0n6172,notn6172,n3002);
and (s1n6172,n5069,n2997);
and (n6173,n6174,n5083);
wire s0n6174,s1n6174,notn6174;
or (n6174,s0n6174,s1n6174);
not(notn6174,n5069);
and (s0n6174,notn6174,n3005);
and (s1n6174,n5069,n3002);
and (n6175,n6176,n5088);
wire s0n6176,s1n6176,notn6176;
or (n6176,s0n6176,s1n6176);
not(notn6176,n5069);
and (s0n6176,notn6176,n3008);
and (s1n6176,n5069,n3005);
and (n6177,n6178,n5093);
wire s0n6178,s1n6178,notn6178;
or (n6178,s0n6178,s1n6178);
not(notn6178,n5069);
and (s0n6178,notn6178,n3011);
and (s1n6178,n5069,n3008);
and (n6180,n6137,n6181);
or (n6181,n6182,n6269,n6807);
and (n6182,n6183,n6226);
wire s0n6183,s1n6183,notn6183;
or (n6183,s0n6183,s1n6183);
not(notn6183,n5021);
and (s0n6183,notn6183,n6184);
and (s1n6183,n5021,n6225);
or (n6184,1'b0,n6185,n6195,n6205,n6215);
and (n6185,n6186,n2710);
or (n6186,1'b0,n6187,n6189,n6191,n6193);
and (n6187,n6188,n5071);
wire s0n6188,s1n6188,notn6188;
or (n6188,s0n6188,s1n6188);
not(notn6188,n5069);
and (s0n6188,notn6188,n3051);
and (s1n6188,n5069,n3122);
and (n6189,n6190,n5083);
wire s0n6190,s1n6190,notn6190;
or (n6190,s0n6190,s1n6190);
not(notn6190,n5069);
and (s0n6190,notn6190,n3055);
and (s1n6190,n5069,n3051);
and (n6191,n6192,n5088);
wire s0n6192,s1n6192,notn6192;
or (n6192,s0n6192,s1n6192);
not(notn6192,n5069);
and (s0n6192,notn6192,n3059);
and (s1n6192,n5069,n3055);
and (n6193,n6194,n5093);
wire s0n6194,s1n6194,notn6194;
or (n6194,s0n6194,s1n6194);
not(notn6194,n5069);
and (s0n6194,notn6194,n3063);
and (s1n6194,n5069,n3059);
and (n6195,n6196,n2722);
or (n6196,1'b0,n6197,n6199,n6201,n6203);
and (n6197,n6198,n5071);
wire s0n6198,s1n6198,notn6198;
or (n6198,s0n6198,s1n6198);
not(notn6198,n5069);
and (s0n6198,notn6198,n3069);
and (s1n6198,n5069,n3063);
and (n6199,n6200,n5083);
wire s0n6200,s1n6200,notn6200;
or (n6200,s0n6200,s1n6200);
not(notn6200,n5069);
and (s0n6200,notn6200,n3073);
and (s1n6200,n5069,n3069);
and (n6201,n6202,n5088);
wire s0n6202,s1n6202,notn6202;
or (n6202,s0n6202,s1n6202);
not(notn6202,n5069);
and (s0n6202,notn6202,n3077);
and (s1n6202,n5069,n3073);
and (n6203,n6204,n5093);
wire s0n6204,s1n6204,notn6204;
or (n6204,s0n6204,s1n6204);
not(notn6204,n5069);
and (s0n6204,notn6204,n3081);
and (s1n6204,n5069,n3077);
and (n6205,n6206,n2734);
or (n6206,1'b0,n6207,n6209,n6211,n6213);
and (n6207,n6208,n5071);
wire s0n6208,s1n6208,notn6208;
or (n6208,s0n6208,s1n6208);
not(notn6208,n5069);
and (s0n6208,notn6208,n3087);
and (s1n6208,n5069,n3137);
and (n6209,n6210,n5083);
wire s0n6210,s1n6210,notn6210;
or (n6210,s0n6210,s1n6210);
not(notn6210,n5069);
and (s0n6210,notn6210,n3091);
and (s1n6210,n5069,n3087);
and (n6211,n6212,n5088);
wire s0n6212,s1n6212,notn6212;
or (n6212,s0n6212,s1n6212);
not(notn6212,n5069);
and (s0n6212,notn6212,n3095);
and (s1n6212,n5069,n3091);
and (n6213,n6214,n5093);
wire s0n6214,s1n6214,notn6214;
or (n6214,s0n6214,s1n6214);
not(notn6214,n5069);
and (s0n6214,notn6214,n3099);
and (s1n6214,n5069,n3095);
and (n6215,n6216,n2744);
or (n6216,1'b0,n6217,n6219,n6221,n6223);
and (n6217,n6218,n5071);
wire s0n6218,s1n6218,notn6218;
or (n6218,s0n6218,s1n6218);
not(notn6218,n5069);
and (s0n6218,notn6218,n3105);
and (s1n6218,n5069,n3099);
and (n6219,n6220,n5083);
wire s0n6220,s1n6220,notn6220;
or (n6220,s0n6220,s1n6220);
not(notn6220,n5069);
and (s0n6220,notn6220,n3109);
and (s1n6220,n5069,n3105);
and (n6221,n6222,n5088);
wire s0n6222,s1n6222,notn6222;
or (n6222,s0n6222,s1n6222);
not(notn6222,n5069);
and (s0n6222,notn6222,n2180);
and (s1n6222,n5069,n3109);
and (n6223,n6224,n5093);
wire s0n6224,s1n6224,notn6224;
or (n6224,s0n6224,s1n6224);
not(notn6224,n5069);
and (s0n6224,notn6224,n1844);
and (s1n6224,n5069,n2180);
wire s0n6226,s1n6226,notn6226;
or (n6226,s0n6226,s1n6226);
not(notn6226,n5021);
and (s0n6226,notn6226,n6227);
and (s1n6226,n5021,n6268);
or (n6227,1'b0,n6228,n6238,n6248,n6258);
and (n6228,n6229,n2710);
or (n6229,1'b0,n6230,n6232,n6234,n6236);
and (n6230,n6231,n5071);
wire s0n6231,s1n6231,notn6231;
or (n6231,s0n6231,s1n6231);
not(notn6231,n5069);
and (s0n6231,notn6231,n3052);
and (s1n6231,n5069,n3123);
and (n6232,n6233,n5083);
wire s0n6233,s1n6233,notn6233;
or (n6233,s0n6233,s1n6233);
not(notn6233,n5069);
and (s0n6233,notn6233,n3056);
and (s1n6233,n5069,n3052);
and (n6234,n6235,n5088);
wire s0n6235,s1n6235,notn6235;
or (n6235,s0n6235,s1n6235);
not(notn6235,n5069);
and (s0n6235,notn6235,n3060);
and (s1n6235,n5069,n3056);
and (n6236,n6237,n5093);
wire s0n6237,s1n6237,notn6237;
or (n6237,s0n6237,s1n6237);
not(notn6237,n5069);
and (s0n6237,notn6237,n3064);
and (s1n6237,n5069,n3060);
and (n6238,n6239,n2722);
or (n6239,1'b0,n6240,n6242,n6244,n6246);
and (n6240,n6241,n5071);
wire s0n6241,s1n6241,notn6241;
or (n6241,s0n6241,s1n6241);
not(notn6241,n5069);
and (s0n6241,notn6241,n3070);
and (s1n6241,n5069,n3064);
and (n6242,n6243,n5083);
wire s0n6243,s1n6243,notn6243;
or (n6243,s0n6243,s1n6243);
not(notn6243,n5069);
and (s0n6243,notn6243,n3074);
and (s1n6243,n5069,n3070);
and (n6244,n6245,n5088);
wire s0n6245,s1n6245,notn6245;
or (n6245,s0n6245,s1n6245);
not(notn6245,n5069);
and (s0n6245,notn6245,n3078);
and (s1n6245,n5069,n3074);
and (n6246,n6247,n5093);
wire s0n6247,s1n6247,notn6247;
or (n6247,s0n6247,s1n6247);
not(notn6247,n5069);
and (s0n6247,notn6247,n3082);
and (s1n6247,n5069,n3078);
and (n6248,n6249,n2734);
or (n6249,1'b0,n6250,n6252,n6254,n6256);
and (n6250,n6251,n5071);
wire s0n6251,s1n6251,notn6251;
or (n6251,s0n6251,s1n6251);
not(notn6251,n5069);
and (s0n6251,notn6251,n3088);
and (s1n6251,n5069,n3138);
and (n6252,n6253,n5083);
wire s0n6253,s1n6253,notn6253;
or (n6253,s0n6253,s1n6253);
not(notn6253,n5069);
and (s0n6253,notn6253,n3092);
and (s1n6253,n5069,n3088);
and (n6254,n6255,n5088);
wire s0n6255,s1n6255,notn6255;
or (n6255,s0n6255,s1n6255);
not(notn6255,n5069);
and (s0n6255,notn6255,n3096);
and (s1n6255,n5069,n3092);
and (n6256,n6257,n5093);
wire s0n6257,s1n6257,notn6257;
or (n6257,s0n6257,s1n6257);
not(notn6257,n5069);
and (s0n6257,notn6257,n3100);
and (s1n6257,n5069,n3096);
and (n6258,n6259,n2744);
or (n6259,1'b0,n6260,n6262,n6264,n6266);
and (n6260,n6261,n5071);
wire s0n6261,s1n6261,notn6261;
or (n6261,s0n6261,s1n6261);
not(notn6261,n5069);
and (s0n6261,notn6261,n3106);
and (s1n6261,n5069,n3100);
and (n6262,n6263,n5083);
wire s0n6263,s1n6263,notn6263;
or (n6263,s0n6263,s1n6263);
not(notn6263,n5069);
and (s0n6263,notn6263,n3110);
and (s1n6263,n5069,n3106);
and (n6264,n6265,n5088);
wire s0n6265,s1n6265,notn6265;
or (n6265,s0n6265,s1n6265);
not(notn6265,n5069);
and (s0n6265,notn6265,n3113);
and (s1n6265,n5069,n3110);
and (n6266,n6267,n5093);
wire s0n6267,s1n6267,notn6267;
or (n6267,s0n6267,s1n6267);
not(notn6267,n5069);
and (s0n6267,notn6267,n3116);
and (s1n6267,n5069,n3113);
and (n6269,n6226,n6270);
or (n6270,n6271,n6358,n6806);
and (n6271,n6272,n6315);
wire s0n6272,s1n6272,notn6272;
or (n6272,s0n6272,s1n6272);
not(notn6272,n5021);
and (s0n6272,notn6272,n6273);
and (s1n6272,n5021,n6314);
or (n6273,1'b0,n6274,n6284,n6294,n6304);
and (n6274,n6275,n2710);
or (n6275,1'b0,n6276,n6278,n6280,n6282);
and (n6276,n6277,n5071);
wire s0n6277,s1n6277,notn6277;
or (n6277,s0n6277,s1n6277);
not(notn6277,n5069);
and (s0n6277,notn6277,n3156);
and (s1n6277,n5069,n3227);
and (n6278,n6279,n5083);
wire s0n6279,s1n6279,notn6279;
or (n6279,s0n6279,s1n6279);
not(notn6279,n5069);
and (s0n6279,notn6279,n3160);
and (s1n6279,n5069,n3156);
and (n6280,n6281,n5088);
wire s0n6281,s1n6281,notn6281;
or (n6281,s0n6281,s1n6281);
not(notn6281,n5069);
and (s0n6281,notn6281,n3164);
and (s1n6281,n5069,n3160);
and (n6282,n6283,n5093);
wire s0n6283,s1n6283,notn6283;
or (n6283,s0n6283,s1n6283);
not(notn6283,n5069);
and (s0n6283,notn6283,n3168);
and (s1n6283,n5069,n3164);
and (n6284,n6285,n2722);
or (n6285,1'b0,n6286,n6288,n6290,n6292);
and (n6286,n6287,n5071);
wire s0n6287,s1n6287,notn6287;
or (n6287,s0n6287,s1n6287);
not(notn6287,n5069);
and (s0n6287,notn6287,n3174);
and (s1n6287,n5069,n3168);
and (n6288,n6289,n5083);
wire s0n6289,s1n6289,notn6289;
or (n6289,s0n6289,s1n6289);
not(notn6289,n5069);
and (s0n6289,notn6289,n3178);
and (s1n6289,n5069,n3174);
and (n6290,n6291,n5088);
wire s0n6291,s1n6291,notn6291;
or (n6291,s0n6291,s1n6291);
not(notn6291,n5069);
and (s0n6291,notn6291,n3182);
and (s1n6291,n5069,n3178);
and (n6292,n6293,n5093);
wire s0n6293,s1n6293,notn6293;
or (n6293,s0n6293,s1n6293);
not(notn6293,n5069);
and (s0n6293,notn6293,n3186);
and (s1n6293,n5069,n3182);
and (n6294,n6295,n2734);
or (n6295,1'b0,n6296,n6298,n6300,n6302);
and (n6296,n6297,n5071);
wire s0n6297,s1n6297,notn6297;
or (n6297,s0n6297,s1n6297);
not(notn6297,n5069);
and (s0n6297,notn6297,n3192);
and (s1n6297,n5069,n3242);
and (n6298,n6299,n5083);
wire s0n6299,s1n6299,notn6299;
or (n6299,s0n6299,s1n6299);
not(notn6299,n5069);
and (s0n6299,notn6299,n3196);
and (s1n6299,n5069,n3192);
and (n6300,n6301,n5088);
wire s0n6301,s1n6301,notn6301;
or (n6301,s0n6301,s1n6301);
not(notn6301,n5069);
and (s0n6301,notn6301,n3200);
and (s1n6301,n5069,n3196);
and (n6302,n6303,n5093);
wire s0n6303,s1n6303,notn6303;
or (n6303,s0n6303,s1n6303);
not(notn6303,n5069);
and (s0n6303,notn6303,n3204);
and (s1n6303,n5069,n3200);
and (n6304,n6305,n2744);
or (n6305,1'b0,n6306,n6308,n6310,n6312);
and (n6306,n6307,n5071);
wire s0n6307,s1n6307,notn6307;
or (n6307,s0n6307,s1n6307);
not(notn6307,n5069);
and (s0n6307,notn6307,n3210);
and (s1n6307,n5069,n3204);
and (n6308,n6309,n5083);
wire s0n6309,s1n6309,notn6309;
or (n6309,s0n6309,s1n6309);
not(notn6309,n5069);
and (s0n6309,notn6309,n3214);
and (s1n6309,n5069,n3210);
and (n6310,n6311,n5088);
wire s0n6311,s1n6311,notn6311;
or (n6311,s0n6311,s1n6311);
not(notn6311,n5069);
and (s0n6311,notn6311,n2196);
and (s1n6311,n5069,n3214);
and (n6312,n6313,n5093);
wire s0n6313,s1n6313,notn6313;
or (n6313,s0n6313,s1n6313);
not(notn6313,n5069);
and (s0n6313,notn6313,n1861);
and (s1n6313,n5069,n2196);
wire s0n6315,s1n6315,notn6315;
or (n6315,s0n6315,s1n6315);
not(notn6315,n5021);
and (s0n6315,notn6315,n6316);
and (s1n6315,n5021,n6357);
or (n6316,1'b0,n6317,n6327,n6337,n6347);
and (n6317,n6318,n2710);
or (n6318,1'b0,n6319,n6321,n6323,n6325);
and (n6319,n6320,n5071);
wire s0n6320,s1n6320,notn6320;
or (n6320,s0n6320,s1n6320);
not(notn6320,n5069);
and (s0n6320,notn6320,n3157);
and (s1n6320,n5069,n3228);
and (n6321,n6322,n5083);
wire s0n6322,s1n6322,notn6322;
or (n6322,s0n6322,s1n6322);
not(notn6322,n5069);
and (s0n6322,notn6322,n3161);
and (s1n6322,n5069,n3157);
and (n6323,n6324,n5088);
wire s0n6324,s1n6324,notn6324;
or (n6324,s0n6324,s1n6324);
not(notn6324,n5069);
and (s0n6324,notn6324,n3165);
and (s1n6324,n5069,n3161);
and (n6325,n6326,n5093);
wire s0n6326,s1n6326,notn6326;
or (n6326,s0n6326,s1n6326);
not(notn6326,n5069);
and (s0n6326,notn6326,n3169);
and (s1n6326,n5069,n3165);
and (n6327,n6328,n2722);
or (n6328,1'b0,n6329,n6331,n6333,n6335);
and (n6329,n6330,n5071);
wire s0n6330,s1n6330,notn6330;
or (n6330,s0n6330,s1n6330);
not(notn6330,n5069);
and (s0n6330,notn6330,n3175);
and (s1n6330,n5069,n3169);
and (n6331,n6332,n5083);
wire s0n6332,s1n6332,notn6332;
or (n6332,s0n6332,s1n6332);
not(notn6332,n5069);
and (s0n6332,notn6332,n3179);
and (s1n6332,n5069,n3175);
and (n6333,n6334,n5088);
wire s0n6334,s1n6334,notn6334;
or (n6334,s0n6334,s1n6334);
not(notn6334,n5069);
and (s0n6334,notn6334,n3183);
and (s1n6334,n5069,n3179);
and (n6335,n6336,n5093);
wire s0n6336,s1n6336,notn6336;
or (n6336,s0n6336,s1n6336);
not(notn6336,n5069);
and (s0n6336,notn6336,n3187);
and (s1n6336,n5069,n3183);
and (n6337,n6338,n2734);
or (n6338,1'b0,n6339,n6341,n6343,n6345);
and (n6339,n6340,n5071);
wire s0n6340,s1n6340,notn6340;
or (n6340,s0n6340,s1n6340);
not(notn6340,n5069);
and (s0n6340,notn6340,n3193);
and (s1n6340,n5069,n3243);
and (n6341,n6342,n5083);
wire s0n6342,s1n6342,notn6342;
or (n6342,s0n6342,s1n6342);
not(notn6342,n5069);
and (s0n6342,notn6342,n3197);
and (s1n6342,n5069,n3193);
and (n6343,n6344,n5088);
wire s0n6344,s1n6344,notn6344;
or (n6344,s0n6344,s1n6344);
not(notn6344,n5069);
and (s0n6344,notn6344,n3201);
and (s1n6344,n5069,n3197);
and (n6345,n6346,n5093);
wire s0n6346,s1n6346,notn6346;
or (n6346,s0n6346,s1n6346);
not(notn6346,n5069);
and (s0n6346,notn6346,n3205);
and (s1n6346,n5069,n3201);
and (n6347,n6348,n2744);
or (n6348,1'b0,n6349,n6351,n6353,n6355);
and (n6349,n6350,n5071);
wire s0n6350,s1n6350,notn6350;
or (n6350,s0n6350,s1n6350);
not(notn6350,n5069);
and (s0n6350,notn6350,n3211);
and (s1n6350,n5069,n3205);
and (n6351,n6352,n5083);
wire s0n6352,s1n6352,notn6352;
or (n6352,s0n6352,s1n6352);
not(notn6352,n5069);
and (s0n6352,notn6352,n3215);
and (s1n6352,n5069,n3211);
and (n6353,n6354,n5088);
wire s0n6354,s1n6354,notn6354;
or (n6354,s0n6354,s1n6354);
not(notn6354,n5069);
and (s0n6354,notn6354,n3218);
and (s1n6354,n5069,n3215);
and (n6355,n6356,n5093);
wire s0n6356,s1n6356,notn6356;
or (n6356,s0n6356,s1n6356);
not(notn6356,n5069);
and (s0n6356,notn6356,n3221);
and (s1n6356,n5069,n3218);
and (n6358,n6315,n6359);
or (n6359,n6360,n6447,n6805);
and (n6360,n6361,n6404);
wire s0n6361,s1n6361,notn6361;
or (n6361,s0n6361,s1n6361);
not(notn6361,n5021);
and (s0n6361,notn6361,n6362);
and (s1n6361,n5021,n6403);
or (n6362,1'b0,n6363,n6373,n6383,n6393);
and (n6363,n6364,n2710);
or (n6364,1'b0,n6365,n6367,n6369,n6371);
and (n6365,n6366,n5071);
wire s0n6366,s1n6366,notn6366;
or (n6366,s0n6366,s1n6366);
not(notn6366,n5069);
and (s0n6366,notn6366,n3261);
and (s1n6366,n5069,n3332);
and (n6367,n6368,n5083);
wire s0n6368,s1n6368,notn6368;
or (n6368,s0n6368,s1n6368);
not(notn6368,n5069);
and (s0n6368,notn6368,n3265);
and (s1n6368,n5069,n3261);
and (n6369,n6370,n5088);
wire s0n6370,s1n6370,notn6370;
or (n6370,s0n6370,s1n6370);
not(notn6370,n5069);
and (s0n6370,notn6370,n3269);
and (s1n6370,n5069,n3265);
and (n6371,n6372,n5093);
wire s0n6372,s1n6372,notn6372;
or (n6372,s0n6372,s1n6372);
not(notn6372,n5069);
and (s0n6372,notn6372,n3273);
and (s1n6372,n5069,n3269);
and (n6373,n6374,n2722);
or (n6374,1'b0,n6375,n6377,n6379,n6381);
and (n6375,n6376,n5071);
wire s0n6376,s1n6376,notn6376;
or (n6376,s0n6376,s1n6376);
not(notn6376,n5069);
and (s0n6376,notn6376,n3279);
and (s1n6376,n5069,n3273);
and (n6377,n6378,n5083);
wire s0n6378,s1n6378,notn6378;
or (n6378,s0n6378,s1n6378);
not(notn6378,n5069);
and (s0n6378,notn6378,n3283);
and (s1n6378,n5069,n3279);
and (n6379,n6380,n5088);
wire s0n6380,s1n6380,notn6380;
or (n6380,s0n6380,s1n6380);
not(notn6380,n5069);
and (s0n6380,notn6380,n3287);
and (s1n6380,n5069,n3283);
and (n6381,n6382,n5093);
wire s0n6382,s1n6382,notn6382;
or (n6382,s0n6382,s1n6382);
not(notn6382,n5069);
and (s0n6382,notn6382,n3291);
and (s1n6382,n5069,n3287);
and (n6383,n6384,n2734);
or (n6384,1'b0,n6385,n6387,n6389,n6391);
and (n6385,n6386,n5071);
wire s0n6386,s1n6386,notn6386;
or (n6386,s0n6386,s1n6386);
not(notn6386,n5069);
and (s0n6386,notn6386,n3297);
and (s1n6386,n5069,n3347);
and (n6387,n6388,n5083);
wire s0n6388,s1n6388,notn6388;
or (n6388,s0n6388,s1n6388);
not(notn6388,n5069);
and (s0n6388,notn6388,n3301);
and (s1n6388,n5069,n3297);
and (n6389,n6390,n5088);
wire s0n6390,s1n6390,notn6390;
or (n6390,s0n6390,s1n6390);
not(notn6390,n5069);
and (s0n6390,notn6390,n3305);
and (s1n6390,n5069,n3301);
and (n6391,n6392,n5093);
wire s0n6392,s1n6392,notn6392;
or (n6392,s0n6392,s1n6392);
not(notn6392,n5069);
and (s0n6392,notn6392,n3309);
and (s1n6392,n5069,n3305);
and (n6393,n6394,n2744);
or (n6394,1'b0,n6395,n6397,n6399,n6401);
and (n6395,n6396,n5071);
wire s0n6396,s1n6396,notn6396;
or (n6396,s0n6396,s1n6396);
not(notn6396,n5069);
and (s0n6396,notn6396,n3315);
and (s1n6396,n5069,n3309);
and (n6397,n6398,n5083);
wire s0n6398,s1n6398,notn6398;
or (n6398,s0n6398,s1n6398);
not(notn6398,n5069);
and (s0n6398,notn6398,n3319);
and (s1n6398,n5069,n3315);
and (n6399,n6400,n5088);
wire s0n6400,s1n6400,notn6400;
or (n6400,s0n6400,s1n6400);
not(notn6400,n5069);
and (s0n6400,notn6400,n2212);
and (s1n6400,n5069,n3319);
and (n6401,n6402,n5093);
wire s0n6402,s1n6402,notn6402;
or (n6402,s0n6402,s1n6402);
not(notn6402,n5069);
and (s0n6402,notn6402,n1886);
and (s1n6402,n5069,n2212);
wire s0n6404,s1n6404,notn6404;
or (n6404,s0n6404,s1n6404);
not(notn6404,n5021);
and (s0n6404,notn6404,n6405);
and (s1n6404,n5021,n6446);
or (n6405,1'b0,n6406,n6416,n6426,n6436);
and (n6406,n6407,n2710);
or (n6407,1'b0,n6408,n6410,n6412,n6414);
and (n6408,n6409,n5071);
wire s0n6409,s1n6409,notn6409;
or (n6409,s0n6409,s1n6409);
not(notn6409,n5069);
and (s0n6409,notn6409,n3262);
and (s1n6409,n5069,n3333);
and (n6410,n6411,n5083);
wire s0n6411,s1n6411,notn6411;
or (n6411,s0n6411,s1n6411);
not(notn6411,n5069);
and (s0n6411,notn6411,n3266);
and (s1n6411,n5069,n3262);
and (n6412,n6413,n5088);
wire s0n6413,s1n6413,notn6413;
or (n6413,s0n6413,s1n6413);
not(notn6413,n5069);
and (s0n6413,notn6413,n3270);
and (s1n6413,n5069,n3266);
and (n6414,n6415,n5093);
wire s0n6415,s1n6415,notn6415;
or (n6415,s0n6415,s1n6415);
not(notn6415,n5069);
and (s0n6415,notn6415,n3274);
and (s1n6415,n5069,n3270);
and (n6416,n6417,n2722);
or (n6417,1'b0,n6418,n6420,n6422,n6424);
and (n6418,n6419,n5071);
wire s0n6419,s1n6419,notn6419;
or (n6419,s0n6419,s1n6419);
not(notn6419,n5069);
and (s0n6419,notn6419,n3280);
and (s1n6419,n5069,n3274);
and (n6420,n6421,n5083);
wire s0n6421,s1n6421,notn6421;
or (n6421,s0n6421,s1n6421);
not(notn6421,n5069);
and (s0n6421,notn6421,n3284);
and (s1n6421,n5069,n3280);
and (n6422,n6423,n5088);
wire s0n6423,s1n6423,notn6423;
or (n6423,s0n6423,s1n6423);
not(notn6423,n5069);
and (s0n6423,notn6423,n3288);
and (s1n6423,n5069,n3284);
and (n6424,n6425,n5093);
wire s0n6425,s1n6425,notn6425;
or (n6425,s0n6425,s1n6425);
not(notn6425,n5069);
and (s0n6425,notn6425,n3292);
and (s1n6425,n5069,n3288);
and (n6426,n6427,n2734);
or (n6427,1'b0,n6428,n6430,n6432,n6434);
and (n6428,n6429,n5071);
wire s0n6429,s1n6429,notn6429;
or (n6429,s0n6429,s1n6429);
not(notn6429,n5069);
and (s0n6429,notn6429,n3298);
and (s1n6429,n5069,n3348);
and (n6430,n6431,n5083);
wire s0n6431,s1n6431,notn6431;
or (n6431,s0n6431,s1n6431);
not(notn6431,n5069);
and (s0n6431,notn6431,n3302);
and (s1n6431,n5069,n3298);
and (n6432,n6433,n5088);
wire s0n6433,s1n6433,notn6433;
or (n6433,s0n6433,s1n6433);
not(notn6433,n5069);
and (s0n6433,notn6433,n3306);
and (s1n6433,n5069,n3302);
and (n6434,n6435,n5093);
wire s0n6435,s1n6435,notn6435;
or (n6435,s0n6435,s1n6435);
not(notn6435,n5069);
and (s0n6435,notn6435,n3310);
and (s1n6435,n5069,n3306);
and (n6436,n6437,n2744);
or (n6437,1'b0,n6438,n6440,n6442,n6444);
and (n6438,n6439,n5071);
wire s0n6439,s1n6439,notn6439;
or (n6439,s0n6439,s1n6439);
not(notn6439,n5069);
and (s0n6439,notn6439,n3316);
and (s1n6439,n5069,n3310);
and (n6440,n6441,n5083);
wire s0n6441,s1n6441,notn6441;
or (n6441,s0n6441,s1n6441);
not(notn6441,n5069);
and (s0n6441,notn6441,n3320);
and (s1n6441,n5069,n3316);
and (n6442,n6443,n5088);
wire s0n6443,s1n6443,notn6443;
or (n6443,s0n6443,s1n6443);
not(notn6443,n5069);
and (s0n6443,notn6443,n3323);
and (s1n6443,n5069,n3320);
and (n6444,n6445,n5093);
wire s0n6445,s1n6445,notn6445;
or (n6445,s0n6445,s1n6445);
not(notn6445,n5069);
and (s0n6445,notn6445,n3326);
and (s1n6445,n5069,n3323);
and (n6447,n6404,n6448);
or (n6448,n6449,n6536,n6804);
and (n6449,n6450,n6493);
wire s0n6450,s1n6450,notn6450;
or (n6450,s0n6450,s1n6450);
not(notn6450,n5021);
and (s0n6450,notn6450,n6451);
and (s1n6450,n5021,n6492);
or (n6451,1'b0,n6452,n6462,n6472,n6482);
and (n6452,n6453,n2710);
or (n6453,1'b0,n6454,n6456,n6458,n6460);
and (n6454,n6455,n5071);
wire s0n6455,s1n6455,notn6455;
or (n6455,s0n6455,s1n6455);
not(notn6455,n5069);
and (s0n6455,notn6455,n3366);
and (s1n6455,n5069,n3437);
and (n6456,n6457,n5083);
wire s0n6457,s1n6457,notn6457;
or (n6457,s0n6457,s1n6457);
not(notn6457,n5069);
and (s0n6457,notn6457,n3370);
and (s1n6457,n5069,n3366);
and (n6458,n6459,n5088);
wire s0n6459,s1n6459,notn6459;
or (n6459,s0n6459,s1n6459);
not(notn6459,n5069);
and (s0n6459,notn6459,n3374);
and (s1n6459,n5069,n3370);
and (n6460,n6461,n5093);
wire s0n6461,s1n6461,notn6461;
or (n6461,s0n6461,s1n6461);
not(notn6461,n5069);
and (s0n6461,notn6461,n3378);
and (s1n6461,n5069,n3374);
and (n6462,n6463,n2722);
or (n6463,1'b0,n6464,n6466,n6468,n6470);
and (n6464,n6465,n5071);
wire s0n6465,s1n6465,notn6465;
or (n6465,s0n6465,s1n6465);
not(notn6465,n5069);
and (s0n6465,notn6465,n3384);
and (s1n6465,n5069,n3378);
and (n6466,n6467,n5083);
wire s0n6467,s1n6467,notn6467;
or (n6467,s0n6467,s1n6467);
not(notn6467,n5069);
and (s0n6467,notn6467,n3388);
and (s1n6467,n5069,n3384);
and (n6468,n6469,n5088);
wire s0n6469,s1n6469,notn6469;
or (n6469,s0n6469,s1n6469);
not(notn6469,n5069);
and (s0n6469,notn6469,n3392);
and (s1n6469,n5069,n3388);
and (n6470,n6471,n5093);
wire s0n6471,s1n6471,notn6471;
or (n6471,s0n6471,s1n6471);
not(notn6471,n5069);
and (s0n6471,notn6471,n3396);
and (s1n6471,n5069,n3392);
and (n6472,n6473,n2734);
or (n6473,1'b0,n6474,n6476,n6478,n6480);
and (n6474,n6475,n5071);
wire s0n6475,s1n6475,notn6475;
or (n6475,s0n6475,s1n6475);
not(notn6475,n5069);
and (s0n6475,notn6475,n3402);
and (s1n6475,n5069,n3452);
and (n6476,n6477,n5083);
wire s0n6477,s1n6477,notn6477;
or (n6477,s0n6477,s1n6477);
not(notn6477,n5069);
and (s0n6477,notn6477,n3406);
and (s1n6477,n5069,n3402);
and (n6478,n6479,n5088);
wire s0n6479,s1n6479,notn6479;
or (n6479,s0n6479,s1n6479);
not(notn6479,n5069);
and (s0n6479,notn6479,n3410);
and (s1n6479,n5069,n3406);
and (n6480,n6481,n5093);
wire s0n6481,s1n6481,notn6481;
or (n6481,s0n6481,s1n6481);
not(notn6481,n5069);
and (s0n6481,notn6481,n3414);
and (s1n6481,n5069,n3410);
and (n6482,n6483,n2744);
or (n6483,1'b0,n6484,n6486,n6488,n6490);
and (n6484,n6485,n5071);
wire s0n6485,s1n6485,notn6485;
or (n6485,s0n6485,s1n6485);
not(notn6485,n5069);
and (s0n6485,notn6485,n3420);
and (s1n6485,n5069,n3414);
and (n6486,n6487,n5083);
wire s0n6487,s1n6487,notn6487;
or (n6487,s0n6487,s1n6487);
not(notn6487,n5069);
and (s0n6487,notn6487,n3424);
and (s1n6487,n5069,n3420);
and (n6488,n6489,n5088);
wire s0n6489,s1n6489,notn6489;
or (n6489,s0n6489,s1n6489);
not(notn6489,n5069);
and (s0n6489,notn6489,n2228);
and (s1n6489,n5069,n3424);
and (n6490,n6491,n5093);
wire s0n6491,s1n6491,notn6491;
or (n6491,s0n6491,s1n6491);
not(notn6491,n5069);
and (s0n6491,notn6491,n1913);
and (s1n6491,n5069,n2228);
wire s0n6493,s1n6493,notn6493;
or (n6493,s0n6493,s1n6493);
not(notn6493,n5021);
and (s0n6493,notn6493,n6494);
and (s1n6493,n5021,n6535);
or (n6494,1'b0,n6495,n6505,n6515,n6525);
and (n6495,n6496,n2710);
or (n6496,1'b0,n6497,n6499,n6501,n6503);
and (n6497,n6498,n5071);
wire s0n6498,s1n6498,notn6498;
or (n6498,s0n6498,s1n6498);
not(notn6498,n5069);
and (s0n6498,notn6498,n3367);
and (s1n6498,n5069,n3438);
and (n6499,n6500,n5083);
wire s0n6500,s1n6500,notn6500;
or (n6500,s0n6500,s1n6500);
not(notn6500,n5069);
and (s0n6500,notn6500,n3371);
and (s1n6500,n5069,n3367);
and (n6501,n6502,n5088);
wire s0n6502,s1n6502,notn6502;
or (n6502,s0n6502,s1n6502);
not(notn6502,n5069);
and (s0n6502,notn6502,n3375);
and (s1n6502,n5069,n3371);
and (n6503,n6504,n5093);
wire s0n6504,s1n6504,notn6504;
or (n6504,s0n6504,s1n6504);
not(notn6504,n5069);
and (s0n6504,notn6504,n3379);
and (s1n6504,n5069,n3375);
and (n6505,n6506,n2722);
or (n6506,1'b0,n6507,n6509,n6511,n6513);
and (n6507,n6508,n5071);
wire s0n6508,s1n6508,notn6508;
or (n6508,s0n6508,s1n6508);
not(notn6508,n5069);
and (s0n6508,notn6508,n3385);
and (s1n6508,n5069,n3379);
and (n6509,n6510,n5083);
wire s0n6510,s1n6510,notn6510;
or (n6510,s0n6510,s1n6510);
not(notn6510,n5069);
and (s0n6510,notn6510,n3389);
and (s1n6510,n5069,n3385);
and (n6511,n6512,n5088);
wire s0n6512,s1n6512,notn6512;
or (n6512,s0n6512,s1n6512);
not(notn6512,n5069);
and (s0n6512,notn6512,n3393);
and (s1n6512,n5069,n3389);
and (n6513,n6514,n5093);
wire s0n6514,s1n6514,notn6514;
or (n6514,s0n6514,s1n6514);
not(notn6514,n5069);
and (s0n6514,notn6514,n3397);
and (s1n6514,n5069,n3393);
and (n6515,n6516,n2734);
or (n6516,1'b0,n6517,n6519,n6521,n6523);
and (n6517,n6518,n5071);
wire s0n6518,s1n6518,notn6518;
or (n6518,s0n6518,s1n6518);
not(notn6518,n5069);
and (s0n6518,notn6518,n3403);
and (s1n6518,n5069,n3453);
and (n6519,n6520,n5083);
wire s0n6520,s1n6520,notn6520;
or (n6520,s0n6520,s1n6520);
not(notn6520,n5069);
and (s0n6520,notn6520,n3407);
and (s1n6520,n5069,n3403);
and (n6521,n6522,n5088);
wire s0n6522,s1n6522,notn6522;
or (n6522,s0n6522,s1n6522);
not(notn6522,n5069);
and (s0n6522,notn6522,n3411);
and (s1n6522,n5069,n3407);
and (n6523,n6524,n5093);
wire s0n6524,s1n6524,notn6524;
or (n6524,s0n6524,s1n6524);
not(notn6524,n5069);
and (s0n6524,notn6524,n3415);
and (s1n6524,n5069,n3411);
and (n6525,n6526,n2744);
or (n6526,1'b0,n6527,n6529,n6531,n6533);
and (n6527,n6528,n5071);
wire s0n6528,s1n6528,notn6528;
or (n6528,s0n6528,s1n6528);
not(notn6528,n5069);
and (s0n6528,notn6528,n3421);
and (s1n6528,n5069,n3415);
and (n6529,n6530,n5083);
wire s0n6530,s1n6530,notn6530;
or (n6530,s0n6530,s1n6530);
not(notn6530,n5069);
and (s0n6530,notn6530,n3425);
and (s1n6530,n5069,n3421);
and (n6531,n6532,n5088);
wire s0n6532,s1n6532,notn6532;
or (n6532,s0n6532,s1n6532);
not(notn6532,n5069);
and (s0n6532,notn6532,n3428);
and (s1n6532,n5069,n3425);
and (n6533,n6534,n5093);
wire s0n6534,s1n6534,notn6534;
or (n6534,s0n6534,s1n6534);
not(notn6534,n5069);
and (s0n6534,notn6534,n3431);
and (s1n6534,n5069,n3428);
and (n6536,n6493,n6537);
or (n6537,n6538,n6625,n6803);
and (n6538,n6539,n6582);
wire s0n6539,s1n6539,notn6539;
or (n6539,s0n6539,s1n6539);
not(notn6539,n5021);
and (s0n6539,notn6539,n6540);
and (s1n6539,n5021,n6581);
or (n6540,1'b0,n6541,n6551,n6561,n6571);
and (n6541,n6542,n2710);
or (n6542,1'b0,n6543,n6545,n6547,n6549);
and (n6543,n6544,n5071);
wire s0n6544,s1n6544,notn6544;
or (n6544,s0n6544,s1n6544);
not(notn6544,n5069);
and (s0n6544,notn6544,n3471);
and (s1n6544,n5069,n3542);
and (n6545,n6546,n5083);
wire s0n6546,s1n6546,notn6546;
or (n6546,s0n6546,s1n6546);
not(notn6546,n5069);
and (s0n6546,notn6546,n3475);
and (s1n6546,n5069,n3471);
and (n6547,n6548,n5088);
wire s0n6548,s1n6548,notn6548;
or (n6548,s0n6548,s1n6548);
not(notn6548,n5069);
and (s0n6548,notn6548,n3479);
and (s1n6548,n5069,n3475);
and (n6549,n6550,n5093);
wire s0n6550,s1n6550,notn6550;
or (n6550,s0n6550,s1n6550);
not(notn6550,n5069);
and (s0n6550,notn6550,n3483);
and (s1n6550,n5069,n3479);
and (n6551,n6552,n2722);
or (n6552,1'b0,n6553,n6555,n6557,n6559);
and (n6553,n6554,n5071);
wire s0n6554,s1n6554,notn6554;
or (n6554,s0n6554,s1n6554);
not(notn6554,n5069);
and (s0n6554,notn6554,n3489);
and (s1n6554,n5069,n3483);
and (n6555,n6556,n5083);
wire s0n6556,s1n6556,notn6556;
or (n6556,s0n6556,s1n6556);
not(notn6556,n5069);
and (s0n6556,notn6556,n3493);
and (s1n6556,n5069,n3489);
and (n6557,n6558,n5088);
wire s0n6558,s1n6558,notn6558;
or (n6558,s0n6558,s1n6558);
not(notn6558,n5069);
and (s0n6558,notn6558,n3497);
and (s1n6558,n5069,n3493);
and (n6559,n6560,n5093);
wire s0n6560,s1n6560,notn6560;
or (n6560,s0n6560,s1n6560);
not(notn6560,n5069);
and (s0n6560,notn6560,n3501);
and (s1n6560,n5069,n3497);
and (n6561,n6562,n2734);
or (n6562,1'b0,n6563,n6565,n6567,n6569);
and (n6563,n6564,n5071);
wire s0n6564,s1n6564,notn6564;
or (n6564,s0n6564,s1n6564);
not(notn6564,n5069);
and (s0n6564,notn6564,n3507);
and (s1n6564,n5069,n3557);
and (n6565,n6566,n5083);
wire s0n6566,s1n6566,notn6566;
or (n6566,s0n6566,s1n6566);
not(notn6566,n5069);
and (s0n6566,notn6566,n3511);
and (s1n6566,n5069,n3507);
and (n6567,n6568,n5088);
wire s0n6568,s1n6568,notn6568;
or (n6568,s0n6568,s1n6568);
not(notn6568,n5069);
and (s0n6568,notn6568,n3515);
and (s1n6568,n5069,n3511);
and (n6569,n6570,n5093);
wire s0n6570,s1n6570,notn6570;
or (n6570,s0n6570,s1n6570);
not(notn6570,n5069);
and (s0n6570,notn6570,n3519);
and (s1n6570,n5069,n3515);
and (n6571,n6572,n2744);
or (n6572,1'b0,n6573,n6575,n6577,n6579);
and (n6573,n6574,n5071);
wire s0n6574,s1n6574,notn6574;
or (n6574,s0n6574,s1n6574);
not(notn6574,n5069);
and (s0n6574,notn6574,n3525);
and (s1n6574,n5069,n3519);
and (n6575,n6576,n5083);
wire s0n6576,s1n6576,notn6576;
or (n6576,s0n6576,s1n6576);
not(notn6576,n5069);
and (s0n6576,notn6576,n3529);
and (s1n6576,n5069,n3525);
and (n6577,n6578,n5088);
wire s0n6578,s1n6578,notn6578;
or (n6578,s0n6578,s1n6578);
not(notn6578,n5069);
and (s0n6578,notn6578,n2244);
and (s1n6578,n5069,n3529);
and (n6579,n6580,n5093);
wire s0n6580,s1n6580,notn6580;
or (n6580,s0n6580,s1n6580);
not(notn6580,n5069);
and (s0n6580,notn6580,n1939);
and (s1n6580,n5069,n2244);
wire s0n6582,s1n6582,notn6582;
or (n6582,s0n6582,s1n6582);
not(notn6582,n5021);
and (s0n6582,notn6582,n6583);
and (s1n6582,n5021,n6624);
or (n6583,1'b0,n6584,n6594,n6604,n6614);
and (n6584,n6585,n2710);
or (n6585,1'b0,n6586,n6588,n6590,n6592);
and (n6586,n6587,n5071);
wire s0n6587,s1n6587,notn6587;
or (n6587,s0n6587,s1n6587);
not(notn6587,n5069);
and (s0n6587,notn6587,n3472);
and (s1n6587,n5069,n3543);
and (n6588,n6589,n5083);
wire s0n6589,s1n6589,notn6589;
or (n6589,s0n6589,s1n6589);
not(notn6589,n5069);
and (s0n6589,notn6589,n3476);
and (s1n6589,n5069,n3472);
and (n6590,n6591,n5088);
wire s0n6591,s1n6591,notn6591;
or (n6591,s0n6591,s1n6591);
not(notn6591,n5069);
and (s0n6591,notn6591,n3480);
and (s1n6591,n5069,n3476);
and (n6592,n6593,n5093);
wire s0n6593,s1n6593,notn6593;
or (n6593,s0n6593,s1n6593);
not(notn6593,n5069);
and (s0n6593,notn6593,n3484);
and (s1n6593,n5069,n3480);
and (n6594,n6595,n2722);
or (n6595,1'b0,n6596,n6598,n6600,n6602);
and (n6596,n6597,n5071);
wire s0n6597,s1n6597,notn6597;
or (n6597,s0n6597,s1n6597);
not(notn6597,n5069);
and (s0n6597,notn6597,n3490);
and (s1n6597,n5069,n3484);
and (n6598,n6599,n5083);
wire s0n6599,s1n6599,notn6599;
or (n6599,s0n6599,s1n6599);
not(notn6599,n5069);
and (s0n6599,notn6599,n3494);
and (s1n6599,n5069,n3490);
and (n6600,n6601,n5088);
wire s0n6601,s1n6601,notn6601;
or (n6601,s0n6601,s1n6601);
not(notn6601,n5069);
and (s0n6601,notn6601,n3498);
and (s1n6601,n5069,n3494);
and (n6602,n6603,n5093);
wire s0n6603,s1n6603,notn6603;
or (n6603,s0n6603,s1n6603);
not(notn6603,n5069);
and (s0n6603,notn6603,n3502);
and (s1n6603,n5069,n3498);
and (n6604,n6605,n2734);
or (n6605,1'b0,n6606,n6608,n6610,n6612);
and (n6606,n6607,n5071);
wire s0n6607,s1n6607,notn6607;
or (n6607,s0n6607,s1n6607);
not(notn6607,n5069);
and (s0n6607,notn6607,n3508);
and (s1n6607,n5069,n3558);
and (n6608,n6609,n5083);
wire s0n6609,s1n6609,notn6609;
or (n6609,s0n6609,s1n6609);
not(notn6609,n5069);
and (s0n6609,notn6609,n3512);
and (s1n6609,n5069,n3508);
and (n6610,n6611,n5088);
wire s0n6611,s1n6611,notn6611;
or (n6611,s0n6611,s1n6611);
not(notn6611,n5069);
and (s0n6611,notn6611,n3516);
and (s1n6611,n5069,n3512);
and (n6612,n6613,n5093);
wire s0n6613,s1n6613,notn6613;
or (n6613,s0n6613,s1n6613);
not(notn6613,n5069);
and (s0n6613,notn6613,n3520);
and (s1n6613,n5069,n3516);
and (n6614,n6615,n2744);
or (n6615,1'b0,n6616,n6618,n6620,n6622);
and (n6616,n6617,n5071);
wire s0n6617,s1n6617,notn6617;
or (n6617,s0n6617,s1n6617);
not(notn6617,n5069);
and (s0n6617,notn6617,n3526);
and (s1n6617,n5069,n3520);
and (n6618,n6619,n5083);
wire s0n6619,s1n6619,notn6619;
or (n6619,s0n6619,s1n6619);
not(notn6619,n5069);
and (s0n6619,notn6619,n3530);
and (s1n6619,n5069,n3526);
and (n6620,n6621,n5088);
wire s0n6621,s1n6621,notn6621;
or (n6621,s0n6621,s1n6621);
not(notn6621,n5069);
and (s0n6621,notn6621,n3533);
and (s1n6621,n5069,n3530);
and (n6622,n6623,n5093);
wire s0n6623,s1n6623,notn6623;
or (n6623,s0n6623,s1n6623);
not(notn6623,n5069);
and (s0n6623,notn6623,n3536);
and (s1n6623,n5069,n3533);
and (n6625,n6582,n6626);
or (n6626,n6627,n6714,n6802);
and (n6627,n6628,n6671);
wire s0n6628,s1n6628,notn6628;
or (n6628,s0n6628,s1n6628);
not(notn6628,n5021);
and (s0n6628,notn6628,n6629);
and (s1n6628,n5021,n6670);
or (n6629,1'b0,n6630,n6640,n6650,n6660);
and (n6630,n6631,n2710);
or (n6631,1'b0,n6632,n6634,n6636,n6638);
and (n6632,n6633,n5071);
wire s0n6633,s1n6633,notn6633;
or (n6633,s0n6633,s1n6633);
not(notn6633,n5069);
and (s0n6633,notn6633,n3576);
and (s1n6633,n5069,n3647);
and (n6634,n6635,n5083);
wire s0n6635,s1n6635,notn6635;
or (n6635,s0n6635,s1n6635);
not(notn6635,n5069);
and (s0n6635,notn6635,n3580);
and (s1n6635,n5069,n3576);
and (n6636,n6637,n5088);
wire s0n6637,s1n6637,notn6637;
or (n6637,s0n6637,s1n6637);
not(notn6637,n5069);
and (s0n6637,notn6637,n3584);
and (s1n6637,n5069,n3580);
and (n6638,n6639,n5093);
wire s0n6639,s1n6639,notn6639;
or (n6639,s0n6639,s1n6639);
not(notn6639,n5069);
and (s0n6639,notn6639,n3588);
and (s1n6639,n5069,n3584);
and (n6640,n6641,n2722);
or (n6641,1'b0,n6642,n6644,n6646,n6648);
and (n6642,n6643,n5071);
wire s0n6643,s1n6643,notn6643;
or (n6643,s0n6643,s1n6643);
not(notn6643,n5069);
and (s0n6643,notn6643,n3594);
and (s1n6643,n5069,n3588);
and (n6644,n6645,n5083);
wire s0n6645,s1n6645,notn6645;
or (n6645,s0n6645,s1n6645);
not(notn6645,n5069);
and (s0n6645,notn6645,n3598);
and (s1n6645,n5069,n3594);
and (n6646,n6647,n5088);
wire s0n6647,s1n6647,notn6647;
or (n6647,s0n6647,s1n6647);
not(notn6647,n5069);
and (s0n6647,notn6647,n3602);
and (s1n6647,n5069,n3598);
and (n6648,n6649,n5093);
wire s0n6649,s1n6649,notn6649;
or (n6649,s0n6649,s1n6649);
not(notn6649,n5069);
and (s0n6649,notn6649,n3606);
and (s1n6649,n5069,n3602);
and (n6650,n6651,n2734);
or (n6651,1'b0,n6652,n6654,n6656,n6658);
and (n6652,n6653,n5071);
wire s0n6653,s1n6653,notn6653;
or (n6653,s0n6653,s1n6653);
not(notn6653,n5069);
and (s0n6653,notn6653,n3612);
and (s1n6653,n5069,n3662);
and (n6654,n6655,n5083);
wire s0n6655,s1n6655,notn6655;
or (n6655,s0n6655,s1n6655);
not(notn6655,n5069);
and (s0n6655,notn6655,n3616);
and (s1n6655,n5069,n3612);
and (n6656,n6657,n5088);
wire s0n6657,s1n6657,notn6657;
or (n6657,s0n6657,s1n6657);
not(notn6657,n5069);
and (s0n6657,notn6657,n3620);
and (s1n6657,n5069,n3616);
and (n6658,n6659,n5093);
wire s0n6659,s1n6659,notn6659;
or (n6659,s0n6659,s1n6659);
not(notn6659,n5069);
and (s0n6659,notn6659,n3624);
and (s1n6659,n5069,n3620);
and (n6660,n6661,n2744);
or (n6661,1'b0,n6662,n6664,n6666,n6668);
and (n6662,n6663,n5071);
wire s0n6663,s1n6663,notn6663;
or (n6663,s0n6663,s1n6663);
not(notn6663,n5069);
and (s0n6663,notn6663,n3630);
and (s1n6663,n5069,n3624);
and (n6664,n6665,n5083);
wire s0n6665,s1n6665,notn6665;
or (n6665,s0n6665,s1n6665);
not(notn6665,n5069);
and (s0n6665,notn6665,n3634);
and (s1n6665,n5069,n3630);
and (n6666,n6667,n5088);
wire s0n6667,s1n6667,notn6667;
or (n6667,s0n6667,s1n6667);
not(notn6667,n5069);
and (s0n6667,notn6667,n2260);
and (s1n6667,n5069,n3634);
and (n6668,n6669,n5093);
wire s0n6669,s1n6669,notn6669;
or (n6669,s0n6669,s1n6669);
not(notn6669,n5069);
and (s0n6669,notn6669,n1968);
and (s1n6669,n5069,n2260);
wire s0n6671,s1n6671,notn6671;
or (n6671,s0n6671,s1n6671);
not(notn6671,n5021);
and (s0n6671,notn6671,n6672);
and (s1n6671,n5021,n6713);
or (n6672,1'b0,n6673,n6683,n6693,n6703);
and (n6673,n6674,n2710);
or (n6674,1'b0,n6675,n6677,n6679,n6681);
and (n6675,n6676,n5071);
wire s0n6676,s1n6676,notn6676;
or (n6676,s0n6676,s1n6676);
not(notn6676,n5069);
and (s0n6676,notn6676,n3577);
and (s1n6676,n5069,n3648);
and (n6677,n6678,n5083);
wire s0n6678,s1n6678,notn6678;
or (n6678,s0n6678,s1n6678);
not(notn6678,n5069);
and (s0n6678,notn6678,n3581);
and (s1n6678,n5069,n3577);
and (n6679,n6680,n5088);
wire s0n6680,s1n6680,notn6680;
or (n6680,s0n6680,s1n6680);
not(notn6680,n5069);
and (s0n6680,notn6680,n3585);
and (s1n6680,n5069,n3581);
and (n6681,n6682,n5093);
wire s0n6682,s1n6682,notn6682;
or (n6682,s0n6682,s1n6682);
not(notn6682,n5069);
and (s0n6682,notn6682,n3589);
and (s1n6682,n5069,n3585);
and (n6683,n6684,n2722);
or (n6684,1'b0,n6685,n6687,n6689,n6691);
and (n6685,n6686,n5071);
wire s0n6686,s1n6686,notn6686;
or (n6686,s0n6686,s1n6686);
not(notn6686,n5069);
and (s0n6686,notn6686,n3595);
and (s1n6686,n5069,n3589);
and (n6687,n6688,n5083);
wire s0n6688,s1n6688,notn6688;
or (n6688,s0n6688,s1n6688);
not(notn6688,n5069);
and (s0n6688,notn6688,n3599);
and (s1n6688,n5069,n3595);
and (n6689,n6690,n5088);
wire s0n6690,s1n6690,notn6690;
or (n6690,s0n6690,s1n6690);
not(notn6690,n5069);
and (s0n6690,notn6690,n3603);
and (s1n6690,n5069,n3599);
and (n6691,n6692,n5093);
wire s0n6692,s1n6692,notn6692;
or (n6692,s0n6692,s1n6692);
not(notn6692,n5069);
and (s0n6692,notn6692,n3607);
and (s1n6692,n5069,n3603);
and (n6693,n6694,n2734);
or (n6694,1'b0,n6695,n6697,n6699,n6701);
and (n6695,n6696,n5071);
wire s0n6696,s1n6696,notn6696;
or (n6696,s0n6696,s1n6696);
not(notn6696,n5069);
and (s0n6696,notn6696,n3613);
and (s1n6696,n5069,n3663);
and (n6697,n6698,n5083);
wire s0n6698,s1n6698,notn6698;
or (n6698,s0n6698,s1n6698);
not(notn6698,n5069);
and (s0n6698,notn6698,n3617);
and (s1n6698,n5069,n3613);
and (n6699,n6700,n5088);
wire s0n6700,s1n6700,notn6700;
or (n6700,s0n6700,s1n6700);
not(notn6700,n5069);
and (s0n6700,notn6700,n3621);
and (s1n6700,n5069,n3617);
and (n6701,n6702,n5093);
wire s0n6702,s1n6702,notn6702;
or (n6702,s0n6702,s1n6702);
not(notn6702,n5069);
and (s0n6702,notn6702,n3625);
and (s1n6702,n5069,n3621);
and (n6703,n6704,n2744);
or (n6704,1'b0,n6705,n6707,n6709,n6711);
and (n6705,n6706,n5071);
wire s0n6706,s1n6706,notn6706;
or (n6706,s0n6706,s1n6706);
not(notn6706,n5069);
and (s0n6706,notn6706,n3631);
and (s1n6706,n5069,n3625);
and (n6707,n6708,n5083);
wire s0n6708,s1n6708,notn6708;
or (n6708,s0n6708,s1n6708);
not(notn6708,n5069);
and (s0n6708,notn6708,n3635);
and (s1n6708,n5069,n3631);
and (n6709,n6710,n5088);
wire s0n6710,s1n6710,notn6710;
or (n6710,s0n6710,s1n6710);
not(notn6710,n5069);
and (s0n6710,notn6710,n3638);
and (s1n6710,n5069,n3635);
and (n6711,n6712,n5093);
wire s0n6712,s1n6712,notn6712;
or (n6712,s0n6712,s1n6712);
not(notn6712,n5069);
and (s0n6712,notn6712,n3641);
and (s1n6712,n5069,n3638);
and (n6714,n6671,n6715);
and (n6715,n6716,n6759);
wire s0n6716,s1n6716,notn6716;
or (n6716,s0n6716,s1n6716);
not(notn6716,n5021);
and (s0n6716,notn6716,n6717);
and (s1n6716,n5021,n6758);
or (n6717,1'b0,n6718,n6728,n6738,n6748);
and (n6718,n6719,n2710);
or (n6719,1'b0,n6720,n6722,n6724,n6726);
and (n6720,n6721,n5071);
wire s0n6721,s1n6721,notn6721;
or (n6721,s0n6721,s1n6721);
not(notn6721,n5069);
and (s0n6721,notn6721,n3680);
and (s1n6721,n5069,n3751);
and (n6722,n6723,n5083);
wire s0n6723,s1n6723,notn6723;
or (n6723,s0n6723,s1n6723);
not(notn6723,n5069);
and (s0n6723,notn6723,n3684);
and (s1n6723,n5069,n3680);
and (n6724,n6725,n5088);
wire s0n6725,s1n6725,notn6725;
or (n6725,s0n6725,s1n6725);
not(notn6725,n5069);
and (s0n6725,notn6725,n3688);
and (s1n6725,n5069,n3684);
and (n6726,n6727,n5093);
wire s0n6727,s1n6727,notn6727;
or (n6727,s0n6727,s1n6727);
not(notn6727,n5069);
and (s0n6727,notn6727,n3692);
and (s1n6727,n5069,n3688);
and (n6728,n6729,n2722);
or (n6729,1'b0,n6730,n6732,n6734,n6736);
and (n6730,n6731,n5071);
wire s0n6731,s1n6731,notn6731;
or (n6731,s0n6731,s1n6731);
not(notn6731,n5069);
and (s0n6731,notn6731,n3698);
and (s1n6731,n5069,n3692);
and (n6732,n6733,n5083);
wire s0n6733,s1n6733,notn6733;
or (n6733,s0n6733,s1n6733);
not(notn6733,n5069);
and (s0n6733,notn6733,n3702);
and (s1n6733,n5069,n3698);
and (n6734,n6735,n5088);
wire s0n6735,s1n6735,notn6735;
or (n6735,s0n6735,s1n6735);
not(notn6735,n5069);
and (s0n6735,notn6735,n3706);
and (s1n6735,n5069,n3702);
and (n6736,n6737,n5093);
wire s0n6737,s1n6737,notn6737;
or (n6737,s0n6737,s1n6737);
not(notn6737,n5069);
and (s0n6737,notn6737,n3710);
and (s1n6737,n5069,n3706);
and (n6738,n6739,n2734);
or (n6739,1'b0,n6740,n6742,n6744,n6746);
and (n6740,n6741,n5071);
wire s0n6741,s1n6741,notn6741;
or (n6741,s0n6741,s1n6741);
not(notn6741,n5069);
and (s0n6741,notn6741,n3716);
and (s1n6741,n5069,n3766);
and (n6742,n6743,n5083);
wire s0n6743,s1n6743,notn6743;
or (n6743,s0n6743,s1n6743);
not(notn6743,n5069);
and (s0n6743,notn6743,n3720);
and (s1n6743,n5069,n3716);
and (n6744,n6745,n5088);
wire s0n6745,s1n6745,notn6745;
or (n6745,s0n6745,s1n6745);
not(notn6745,n5069);
and (s0n6745,notn6745,n3724);
and (s1n6745,n5069,n3720);
and (n6746,n6747,n5093);
wire s0n6747,s1n6747,notn6747;
or (n6747,s0n6747,s1n6747);
not(notn6747,n5069);
and (s0n6747,notn6747,n3728);
and (s1n6747,n5069,n3724);
and (n6748,n6749,n2744);
or (n6749,1'b0,n6750,n6752,n6754,n6756);
and (n6750,n6751,n5071);
wire s0n6751,s1n6751,notn6751;
or (n6751,s0n6751,s1n6751);
not(notn6751,n5069);
and (s0n6751,notn6751,n3734);
and (s1n6751,n5069,n3728);
and (n6752,n6753,n5083);
wire s0n6753,s1n6753,notn6753;
or (n6753,s0n6753,s1n6753);
not(notn6753,n5069);
and (s0n6753,notn6753,n3738);
and (s1n6753,n5069,n3734);
and (n6754,n6755,n5088);
wire s0n6755,s1n6755,notn6755;
or (n6755,s0n6755,s1n6755);
not(notn6755,n5069);
and (s0n6755,notn6755,n2275);
and (s1n6755,n5069,n3738);
and (n6756,n6757,n5093);
wire s0n6757,s1n6757,notn6757;
or (n6757,s0n6757,s1n6757);
not(notn6757,n5069);
and (s0n6757,notn6757,n1987);
and (s1n6757,n5069,n2275);
wire s0n6759,s1n6759,notn6759;
or (n6759,s0n6759,s1n6759);
not(notn6759,n5021);
and (s0n6759,notn6759,n6760);
and (s1n6759,n5021,n6801);
or (n6760,1'b0,n6761,n6771,n6781,n6791);
and (n6761,n6762,n2710);
or (n6762,1'b0,n6763,n6765,n6767,n6769);
and (n6763,n6764,n5071);
wire s0n6764,s1n6764,notn6764;
or (n6764,s0n6764,s1n6764);
not(notn6764,n5069);
and (s0n6764,notn6764,n3681);
and (s1n6764,n5069,n3752);
and (n6765,n6766,n5083);
wire s0n6766,s1n6766,notn6766;
or (n6766,s0n6766,s1n6766);
not(notn6766,n5069);
and (s0n6766,notn6766,n3685);
and (s1n6766,n5069,n3681);
and (n6767,n6768,n5088);
wire s0n6768,s1n6768,notn6768;
or (n6768,s0n6768,s1n6768);
not(notn6768,n5069);
and (s0n6768,notn6768,n3689);
and (s1n6768,n5069,n3685);
and (n6769,n6770,n5093);
wire s0n6770,s1n6770,notn6770;
or (n6770,s0n6770,s1n6770);
not(notn6770,n5069);
and (s0n6770,notn6770,n3693);
and (s1n6770,n5069,n3689);
and (n6771,n6772,n2722);
or (n6772,1'b0,n6773,n6775,n6777,n6779);
and (n6773,n6774,n5071);
wire s0n6774,s1n6774,notn6774;
or (n6774,s0n6774,s1n6774);
not(notn6774,n5069);
and (s0n6774,notn6774,n3699);
and (s1n6774,n5069,n3693);
and (n6775,n6776,n5083);
wire s0n6776,s1n6776,notn6776;
or (n6776,s0n6776,s1n6776);
not(notn6776,n5069);
and (s0n6776,notn6776,n3703);
and (s1n6776,n5069,n3699);
and (n6777,n6778,n5088);
wire s0n6778,s1n6778,notn6778;
or (n6778,s0n6778,s1n6778);
not(notn6778,n5069);
and (s0n6778,notn6778,n3707);
and (s1n6778,n5069,n3703);
and (n6779,n6780,n5093);
wire s0n6780,s1n6780,notn6780;
or (n6780,s0n6780,s1n6780);
not(notn6780,n5069);
and (s0n6780,notn6780,n3711);
and (s1n6780,n5069,n3707);
and (n6781,n6782,n2734);
or (n6782,1'b0,n6783,n6785,n6787,n6789);
and (n6783,n6784,n5071);
wire s0n6784,s1n6784,notn6784;
or (n6784,s0n6784,s1n6784);
not(notn6784,n5069);
and (s0n6784,notn6784,n3717);
and (s1n6784,n5069,n3767);
and (n6785,n6786,n5083);
wire s0n6786,s1n6786,notn6786;
or (n6786,s0n6786,s1n6786);
not(notn6786,n5069);
and (s0n6786,notn6786,n3721);
and (s1n6786,n5069,n3717);
and (n6787,n6788,n5088);
wire s0n6788,s1n6788,notn6788;
or (n6788,s0n6788,s1n6788);
not(notn6788,n5069);
and (s0n6788,notn6788,n3725);
and (s1n6788,n5069,n3721);
and (n6789,n6790,n5093);
wire s0n6790,s1n6790,notn6790;
or (n6790,s0n6790,s1n6790);
not(notn6790,n5069);
and (s0n6790,notn6790,n3729);
and (s1n6790,n5069,n3725);
and (n6791,n6792,n2744);
or (n6792,1'b0,n6793,n6795,n6797,n6799);
and (n6793,n6794,n5071);
wire s0n6794,s1n6794,notn6794;
or (n6794,s0n6794,s1n6794);
not(notn6794,n5069);
and (s0n6794,notn6794,n3735);
and (s1n6794,n5069,n3729);
and (n6795,n6796,n5083);
wire s0n6796,s1n6796,notn6796;
or (n6796,s0n6796,s1n6796);
not(notn6796,n5069);
and (s0n6796,notn6796,n3739);
and (s1n6796,n5069,n3735);
and (n6797,n6798,n5088);
wire s0n6798,s1n6798,notn6798;
or (n6798,s0n6798,s1n6798);
not(notn6798,n5069);
and (s0n6798,notn6798,n3742);
and (s1n6798,n5069,n3739);
and (n6799,n6800,n5093);
wire s0n6800,s1n6800,notn6800;
or (n6800,s0n6800,s1n6800);
not(notn6800,n5069);
and (s0n6800,notn6800,n3745);
and (s1n6800,n5069,n3742);
and (n6802,n6628,n6715);
and (n6803,n6539,n6626);
and (n6804,n6450,n6537);
and (n6805,n6361,n6448);
and (n6806,n6272,n6359);
and (n6807,n6183,n6270);
and (n6808,n6094,n6181);
and (n6809,n6087,n6092);
and (n6810,n6080,n6085);
not (n6811,n6812);
nor (n6812,n6813,n7418);
and (n6813,n6814,n7413);
nand (n6814,n6815,n7397);
or (n6815,n6816,n6839);
nand (n6816,n6817,n6828);
and (n6817,n6818,n6823);
or (n6818,n6819,n6821);
wire s0n6819,s1n6819,notn6819;
or (n6819,s0n6819,s1n6819);
not(notn6819,n5021);
and (s0n6819,notn6819,1'b0);
and (s1n6819,n5021,n6820);
wire s0n6821,s1n6821,notn6821;
or (n6821,s0n6821,s1n6821);
not(notn6821,n5021);
and (s0n6821,notn6821,1'b0);
and (s1n6821,n5021,n6822);
or (n6823,n6824,n6826);
wire s0n6824,s1n6824,notn6824;
or (n6824,s0n6824,s1n6824);
not(notn6824,n5021);
and (s0n6824,notn6824,1'b0);
and (s1n6824,n5021,n6825);
wire s0n6826,s1n6826,notn6826;
or (n6826,s0n6826,s1n6826);
not(notn6826,n5021);
and (s0n6826,notn6826,1'b0);
and (s1n6826,n5021,n6827);
nor (n6828,n6829,n6834);
nor (n6829,n6830,n6832);
wire s0n6830,s1n6830,notn6830;
or (n6830,s0n6830,s1n6830);
not(notn6830,n5021);
and (s0n6830,notn6830,1'b0);
and (s1n6830,n5021,n6831);
wire s0n6832,s1n6832,notn6832;
or (n6832,s0n6832,s1n6832);
not(notn6832,n5021);
and (s0n6832,notn6832,1'b0);
and (s1n6832,n5021,n6833);
nor (n6834,n6835,n6837);
wire s0n6835,s1n6835,notn6835;
or (n6835,s0n6835,s1n6835);
not(notn6835,n5021);
and (s0n6835,notn6835,1'b0);
and (s1n6835,n5021,n6836);
wire s0n6837,s1n6837,notn6837;
or (n6837,s0n6837,s1n6837);
not(notn6837,n5021);
and (s0n6837,notn6837,1'b0);
and (s1n6837,n5021,n6838);
not (n6839,n6840);
or (n6840,n6841,n6908,n7396);
and (n6841,n6842,n6874);
wire s0n6842,s1n6842,notn6842;
or (n6842,s0n6842,s1n6842);
not(notn6842,n5021);
and (s0n6842,notn6842,n6843);
and (s1n6842,n5021,n6873);
or (n6843,1'b0,n6844,n6845,n6846,n6861);
and (n6844,n5169,n2710);
and (n6845,n5184,n2722);
and (n6846,n6847,n2734);
or (n6847,1'b0,n6848,n6852,n6855,n6858);
and (n6848,n6849,n5071);
wire s0n6849,s1n6849,notn6849;
or (n6849,s0n6849,s1n6849);
not(notn6849,n5069);
and (s0n6849,notn6849,n6850);
and (s1n6849,n5069,n6851);
and (n6852,n6853,n5083);
wire s0n6853,s1n6853,notn6853;
or (n6853,s0n6853,s1n6853);
not(notn6853,n5069);
and (s0n6853,notn6853,n6854);
and (s1n6853,n5069,n6850);
and (n6855,n6856,n5088);
wire s0n6856,s1n6856,notn6856;
or (n6856,s0n6856,s1n6856);
not(notn6856,n5069);
and (s0n6856,notn6856,n6857);
and (s1n6856,n5069,n6854);
and (n6858,n6859,n5093);
wire s0n6859,s1n6859,notn6859;
or (n6859,s0n6859,s1n6859);
not(notn6859,n5069);
and (s0n6859,notn6859,n6860);
and (s1n6859,n5069,n6857);
and (n6861,n6862,n2744);
or (n6862,1'b0,n6863,n6866,n6869,n6871);
and (n6863,n6864,n5071);
wire s0n6864,s1n6864,notn6864;
or (n6864,s0n6864,s1n6864);
not(notn6864,n5069);
and (s0n6864,notn6864,n6865);
and (s1n6864,n5069,n6860);
and (n6866,n6867,n5083);
wire s0n6867,s1n6867,notn6867;
or (n6867,s0n6867,s1n6867);
not(notn6867,n5069);
and (s0n6867,notn6867,n6868);
and (s1n6867,n5069,n6865);
and (n6869,n6870,n5088);
wire s0n6870,s1n6870,notn6870;
or (n6870,s0n6870,s1n6870);
not(notn6870,n5069);
and (s0n6870,notn6870,n1300);
and (s1n6870,n5069,n6868);
and (n6871,n6872,n5093);
wire s0n6872,s1n6872,notn6872;
or (n6872,s0n6872,s1n6872);
not(notn6872,n5069);
and (s0n6872,notn6872,n557);
and (s1n6872,n5069,n1300);
wire s0n6874,s1n6874,notn6874;
or (n6874,s0n6874,s1n6874);
not(notn6874,n5021);
and (s0n6874,notn6874,n6875);
and (s1n6874,n5021,n6907);
or (n6875,1'b0,n6876,n6891,n6905,n6906);
and (n6876,n6877,n2710);
or (n6877,1'b0,n6878,n6882,n6885,n6888);
and (n6878,n6879,n5071);
wire s0n6879,s1n6879,notn6879;
or (n6879,s0n6879,s1n6879);
not(notn6879,n5069);
and (s0n6879,notn6879,n6880);
and (s1n6879,n5069,n6881);
and (n6882,n6883,n5083);
wire s0n6883,s1n6883,notn6883;
or (n6883,s0n6883,s1n6883);
not(notn6883,n5069);
and (s0n6883,notn6883,n6884);
and (s1n6883,n5069,n6880);
and (n6885,n6886,n5088);
wire s0n6886,s1n6886,notn6886;
or (n6886,s0n6886,s1n6886);
not(notn6886,n5069);
and (s0n6886,notn6886,n6887);
and (s1n6886,n5069,n6884);
and (n6888,n6889,n5093);
wire s0n6889,s1n6889,notn6889;
or (n6889,s0n6889,s1n6889);
not(notn6889,n5069);
and (s0n6889,notn6889,n6890);
and (s1n6889,n5069,n6887);
and (n6891,n6892,n2722);
or (n6892,1'b0,n6893,n6896,n6899,n6902);
and (n6893,n6894,n5071);
wire s0n6894,s1n6894,notn6894;
or (n6894,s0n6894,s1n6894);
not(notn6894,n5069);
and (s0n6894,notn6894,n6895);
and (s1n6894,n5069,n6890);
and (n6896,n6897,n5083);
wire s0n6897,s1n6897,notn6897;
or (n6897,s0n6897,s1n6897);
not(notn6897,n5069);
and (s0n6897,notn6897,n6898);
and (s1n6897,n5069,n6895);
and (n6899,n6900,n5088);
wire s0n6900,s1n6900,notn6900;
or (n6900,s0n6900,s1n6900);
not(notn6900,n5069);
and (s0n6900,notn6900,n6901);
and (s1n6900,n5069,n6898);
and (n6902,n6903,n5093);
wire s0n6903,s1n6903,notn6903;
or (n6903,s0n6903,s1n6903);
not(notn6903,n5069);
and (s0n6903,notn6903,n6904);
and (s1n6903,n5069,n6901);
and (n6905,n5064,n2734);
and (n6906,n5096,n2744);
and (n6908,n6874,n6909);
or (n6909,n6910,n6977,n7395);
and (n6910,n6911,n6943);
wire s0n6911,s1n6911,notn6911;
or (n6911,s0n6911,s1n6911);
not(notn6911,n5021);
and (s0n6911,notn6911,n6912);
and (s1n6911,n5021,n6942);
or (n6912,1'b0,n6913,n6914,n6915,n6930);
and (n6913,n5292,n2710);
and (n6914,n5307,n2722);
and (n6915,n6916,n2734);
or (n6916,1'b0,n6917,n6921,n6924,n6927);
and (n6917,n6918,n5071);
wire s0n6918,s1n6918,notn6918;
or (n6918,s0n6918,s1n6918);
not(notn6918,n5069);
and (s0n6918,notn6918,n6919);
and (s1n6918,n5069,n6920);
and (n6921,n6922,n5083);
wire s0n6922,s1n6922,notn6922;
or (n6922,s0n6922,s1n6922);
not(notn6922,n5069);
and (s0n6922,notn6922,n6923);
and (s1n6922,n5069,n6919);
and (n6924,n6925,n5088);
wire s0n6925,s1n6925,notn6925;
or (n6925,s0n6925,s1n6925);
not(notn6925,n5069);
and (s0n6925,notn6925,n6926);
and (s1n6925,n5069,n6923);
and (n6927,n6928,n5093);
wire s0n6928,s1n6928,notn6928;
or (n6928,s0n6928,s1n6928);
not(notn6928,n5069);
and (s0n6928,notn6928,n6929);
and (s1n6928,n5069,n6926);
and (n6930,n6931,n2744);
or (n6931,1'b0,n6932,n6935,n6938,n6940);
and (n6932,n6933,n5071);
wire s0n6933,s1n6933,notn6933;
or (n6933,s0n6933,s1n6933);
not(notn6933,n5069);
and (s0n6933,notn6933,n6934);
and (s1n6933,n5069,n6929);
and (n6935,n6936,n5083);
wire s0n6936,s1n6936,notn6936;
or (n6936,s0n6936,s1n6936);
not(notn6936,n5069);
and (s0n6936,notn6936,n6937);
and (s1n6936,n5069,n6934);
and (n6938,n6939,n5088);
wire s0n6939,s1n6939,notn6939;
or (n6939,s0n6939,s1n6939);
not(notn6939,n5069);
and (s0n6939,notn6939,n1316);
and (s1n6939,n5069,n6937);
and (n6940,n6941,n5093);
wire s0n6941,s1n6941,notn6941;
or (n6941,s0n6941,s1n6941);
not(notn6941,n5069);
and (s0n6941,notn6941,n749);
and (s1n6941,n5069,n1316);
wire s0n6943,s1n6943,notn6943;
or (n6943,s0n6943,s1n6943);
not(notn6943,n5021);
and (s0n6943,notn6943,n6944);
and (s1n6943,n5021,n6976);
or (n6944,1'b0,n6945,n6960,n6974,n6975);
and (n6945,n6946,n2710);
or (n6946,1'b0,n6947,n6951,n6954,n6957);
and (n6947,n6948,n5071);
wire s0n6948,s1n6948,notn6948;
or (n6948,s0n6948,s1n6948);
not(notn6948,n5069);
and (s0n6948,notn6948,n6949);
and (s1n6948,n5069,n6950);
and (n6951,n6952,n5083);
wire s0n6952,s1n6952,notn6952;
or (n6952,s0n6952,s1n6952);
not(notn6952,n5069);
and (s0n6952,notn6952,n6953);
and (s1n6952,n5069,n6949);
and (n6954,n6955,n5088);
wire s0n6955,s1n6955,notn6955;
or (n6955,s0n6955,s1n6955);
not(notn6955,n5069);
and (s0n6955,notn6955,n6956);
and (s1n6955,n5069,n6953);
and (n6957,n6958,n5093);
wire s0n6958,s1n6958,notn6958;
or (n6958,s0n6958,s1n6958);
not(notn6958,n5069);
and (s0n6958,notn6958,n6959);
and (s1n6958,n5069,n6956);
and (n6960,n6961,n2722);
or (n6961,1'b0,n6962,n6965,n6968,n6971);
and (n6962,n6963,n5071);
wire s0n6963,s1n6963,notn6963;
or (n6963,s0n6963,s1n6963);
not(notn6963,n5069);
and (s0n6963,notn6963,n6964);
and (s1n6963,n5069,n6959);
and (n6965,n6966,n5083);
wire s0n6966,s1n6966,notn6966;
or (n6966,s0n6966,s1n6966);
not(notn6966,n5069);
and (s0n6966,notn6966,n6967);
and (s1n6966,n5069,n6964);
and (n6968,n6969,n5088);
wire s0n6969,s1n6969,notn6969;
or (n6969,s0n6969,s1n6969);
not(notn6969,n5069);
and (s0n6969,notn6969,n6970);
and (s1n6969,n5069,n6967);
and (n6971,n6972,n5093);
wire s0n6972,s1n6972,notn6972;
or (n6972,s0n6972,s1n6972);
not(notn6972,n5069);
and (s0n6972,notn6972,n6973);
and (s1n6972,n5069,n6970);
and (n6974,n5204,n2734);
and (n6975,n5219,n2744);
and (n6977,n6943,n6978);
or (n6978,n6979,n7046,n7394);
and (n6979,n6980,n7012);
wire s0n6980,s1n6980,notn6980;
or (n6980,s0n6980,s1n6980);
not(notn6980,n5021);
and (s0n6980,notn6980,n6981);
and (s1n6980,n5021,n7011);
or (n6981,1'b0,n6982,n6983,n6984,n6999);
and (n6982,n5415,n2710);
and (n6983,n5430,n2722);
and (n6984,n6985,n2734);
or (n6985,1'b0,n6986,n6990,n6993,n6996);
and (n6986,n6987,n5071);
wire s0n6987,s1n6987,notn6987;
or (n6987,s0n6987,s1n6987);
not(notn6987,n5069);
and (s0n6987,notn6987,n6988);
and (s1n6987,n5069,n6989);
and (n6990,n6991,n5083);
wire s0n6991,s1n6991,notn6991;
or (n6991,s0n6991,s1n6991);
not(notn6991,n5069);
and (s0n6991,notn6991,n6992);
and (s1n6991,n5069,n6988);
and (n6993,n6994,n5088);
wire s0n6994,s1n6994,notn6994;
or (n6994,s0n6994,s1n6994);
not(notn6994,n5069);
and (s0n6994,notn6994,n6995);
and (s1n6994,n5069,n6992);
and (n6996,n6997,n5093);
wire s0n6997,s1n6997,notn6997;
or (n6997,s0n6997,s1n6997);
not(notn6997,n5069);
and (s0n6997,notn6997,n6998);
and (s1n6997,n5069,n6995);
and (n6999,n7000,n2744);
or (n7000,1'b0,n7001,n7004,n7007,n7009);
and (n7001,n7002,n5071);
wire s0n7002,s1n7002,notn7002;
or (n7002,s0n7002,s1n7002);
not(notn7002,n5069);
and (s0n7002,notn7002,n7003);
and (s1n7002,n5069,n6998);
and (n7004,n7005,n5083);
wire s0n7005,s1n7005,notn7005;
or (n7005,s0n7005,s1n7005);
not(notn7005,n5069);
and (s0n7005,notn7005,n7006);
and (s1n7005,n5069,n7003);
and (n7007,n7008,n5088);
wire s0n7008,s1n7008,notn7008;
or (n7008,s0n7008,s1n7008);
not(notn7008,n5069);
and (s0n7008,notn7008,n1332);
and (s1n7008,n5069,n7006);
and (n7009,n7010,n5093);
wire s0n7010,s1n7010,notn7010;
or (n7010,s0n7010,s1n7010);
not(notn7010,n5069);
and (s0n7010,notn7010,n770);
and (s1n7010,n5069,n1332);
wire s0n7012,s1n7012,notn7012;
or (n7012,s0n7012,s1n7012);
not(notn7012,n5021);
and (s0n7012,notn7012,n7013);
and (s1n7012,n5021,n7045);
or (n7013,1'b0,n7014,n7029,n7043,n7044);
and (n7014,n7015,n2710);
or (n7015,1'b0,n7016,n7020,n7023,n7026);
and (n7016,n7017,n5071);
wire s0n7017,s1n7017,notn7017;
or (n7017,s0n7017,s1n7017);
not(notn7017,n5069);
and (s0n7017,notn7017,n7018);
and (s1n7017,n5069,n7019);
and (n7020,n7021,n5083);
wire s0n7021,s1n7021,notn7021;
or (n7021,s0n7021,s1n7021);
not(notn7021,n5069);
and (s0n7021,notn7021,n7022);
and (s1n7021,n5069,n7018);
and (n7023,n7024,n5088);
wire s0n7024,s1n7024,notn7024;
or (n7024,s0n7024,s1n7024);
not(notn7024,n5069);
and (s0n7024,notn7024,n7025);
and (s1n7024,n5069,n7022);
and (n7026,n7027,n5093);
wire s0n7027,s1n7027,notn7027;
or (n7027,s0n7027,s1n7027);
not(notn7027,n5069);
and (s0n7027,notn7027,n7028);
and (s1n7027,n5069,n7025);
and (n7029,n7030,n2722);
or (n7030,1'b0,n7031,n7034,n7037,n7040);
and (n7031,n7032,n5071);
wire s0n7032,s1n7032,notn7032;
or (n7032,s0n7032,s1n7032);
not(notn7032,n5069);
and (s0n7032,notn7032,n7033);
and (s1n7032,n5069,n7028);
and (n7034,n7035,n5083);
wire s0n7035,s1n7035,notn7035;
or (n7035,s0n7035,s1n7035);
not(notn7035,n5069);
and (s0n7035,notn7035,n7036);
and (s1n7035,n5069,n7033);
and (n7037,n7038,n5088);
wire s0n7038,s1n7038,notn7038;
or (n7038,s0n7038,s1n7038);
not(notn7038,n5069);
and (s0n7038,notn7038,n7039);
and (s1n7038,n5069,n7036);
and (n7040,n7041,n5093);
wire s0n7041,s1n7041,notn7041;
or (n7041,s0n7041,s1n7041);
not(notn7041,n5069);
and (s0n7041,notn7041,n7042);
and (s1n7041,n5069,n7039);
and (n7043,n5327,n2734);
and (n7044,n5342,n2744);
and (n7046,n7012,n7047);
or (n7047,n7048,n7115,n7393);
and (n7048,n7049,n7081);
wire s0n7049,s1n7049,notn7049;
or (n7049,s0n7049,s1n7049);
not(notn7049,n5021);
and (s0n7049,notn7049,n7050);
and (s1n7049,n5021,n7080);
or (n7050,1'b0,n7051,n7052,n7053,n7068);
and (n7051,n5538,n2710);
and (n7052,n5553,n2722);
and (n7053,n7054,n2734);
or (n7054,1'b0,n7055,n7059,n7062,n7065);
and (n7055,n7056,n5071);
wire s0n7056,s1n7056,notn7056;
or (n7056,s0n7056,s1n7056);
not(notn7056,n5069);
and (s0n7056,notn7056,n7057);
and (s1n7056,n5069,n7058);
and (n7059,n7060,n5083);
wire s0n7060,s1n7060,notn7060;
or (n7060,s0n7060,s1n7060);
not(notn7060,n5069);
and (s0n7060,notn7060,n7061);
and (s1n7060,n5069,n7057);
and (n7062,n7063,n5088);
wire s0n7063,s1n7063,notn7063;
or (n7063,s0n7063,s1n7063);
not(notn7063,n5069);
and (s0n7063,notn7063,n7064);
and (s1n7063,n5069,n7061);
and (n7065,n7066,n5093);
wire s0n7066,s1n7066,notn7066;
or (n7066,s0n7066,s1n7066);
not(notn7066,n5069);
and (s0n7066,notn7066,n7067);
and (s1n7066,n5069,n7064);
and (n7068,n7069,n2744);
or (n7069,1'b0,n7070,n7073,n7076,n7078);
and (n7070,n7071,n5071);
wire s0n7071,s1n7071,notn7071;
or (n7071,s0n7071,s1n7071);
not(notn7071,n5069);
and (s0n7071,notn7071,n7072);
and (s1n7071,n5069,n7067);
and (n7073,n7074,n5083);
wire s0n7074,s1n7074,notn7074;
or (n7074,s0n7074,s1n7074);
not(notn7074,n5069);
and (s0n7074,notn7074,n7075);
and (s1n7074,n5069,n7072);
and (n7076,n7077,n5088);
wire s0n7077,s1n7077,notn7077;
or (n7077,s0n7077,s1n7077);
not(notn7077,n5069);
and (s0n7077,notn7077,n1348);
and (s1n7077,n5069,n7075);
and (n7078,n7079,n5093);
wire s0n7079,s1n7079,notn7079;
or (n7079,s0n7079,s1n7079);
not(notn7079,n5069);
and (s0n7079,notn7079,n796);
and (s1n7079,n5069,n1348);
wire s0n7081,s1n7081,notn7081;
or (n7081,s0n7081,s1n7081);
not(notn7081,n5021);
and (s0n7081,notn7081,n7082);
and (s1n7081,n5021,n7114);
or (n7082,1'b0,n7083,n7098,n7112,n7113);
and (n7083,n7084,n2710);
or (n7084,1'b0,n7085,n7089,n7092,n7095);
and (n7085,n7086,n5071);
wire s0n7086,s1n7086,notn7086;
or (n7086,s0n7086,s1n7086);
not(notn7086,n5069);
and (s0n7086,notn7086,n7087);
and (s1n7086,n5069,n7088);
and (n7089,n7090,n5083);
wire s0n7090,s1n7090,notn7090;
or (n7090,s0n7090,s1n7090);
not(notn7090,n5069);
and (s0n7090,notn7090,n7091);
and (s1n7090,n5069,n7087);
and (n7092,n7093,n5088);
wire s0n7093,s1n7093,notn7093;
or (n7093,s0n7093,s1n7093);
not(notn7093,n5069);
and (s0n7093,notn7093,n7094);
and (s1n7093,n5069,n7091);
and (n7095,n7096,n5093);
wire s0n7096,s1n7096,notn7096;
or (n7096,s0n7096,s1n7096);
not(notn7096,n5069);
and (s0n7096,notn7096,n7097);
and (s1n7096,n5069,n7094);
and (n7098,n7099,n2722);
or (n7099,1'b0,n7100,n7103,n7106,n7109);
and (n7100,n7101,n5071);
wire s0n7101,s1n7101,notn7101;
or (n7101,s0n7101,s1n7101);
not(notn7101,n5069);
and (s0n7101,notn7101,n7102);
and (s1n7101,n5069,n7097);
and (n7103,n7104,n5083);
wire s0n7104,s1n7104,notn7104;
or (n7104,s0n7104,s1n7104);
not(notn7104,n5069);
and (s0n7104,notn7104,n7105);
and (s1n7104,n5069,n7102);
and (n7106,n7107,n5088);
wire s0n7107,s1n7107,notn7107;
or (n7107,s0n7107,s1n7107);
not(notn7107,n5069);
and (s0n7107,notn7107,n7108);
and (s1n7107,n5069,n7105);
and (n7109,n7110,n5093);
wire s0n7110,s1n7110,notn7110;
or (n7110,s0n7110,s1n7110);
not(notn7110,n5069);
and (s0n7110,notn7110,n7111);
and (s1n7110,n5069,n7108);
and (n7112,n5450,n2734);
and (n7113,n5465,n2744);
and (n7115,n7081,n7116);
or (n7116,n7117,n7184,n7392);
and (n7117,n7118,n7150);
wire s0n7118,s1n7118,notn7118;
or (n7118,s0n7118,s1n7118);
not(notn7118,n5021);
and (s0n7118,notn7118,n7119);
and (s1n7118,n5021,n7149);
or (n7119,1'b0,n7120,n7121,n7122,n7137);
and (n7120,n5661,n2710);
and (n7121,n5676,n2722);
and (n7122,n7123,n2734);
or (n7123,1'b0,n7124,n7128,n7131,n7134);
and (n7124,n7125,n5071);
wire s0n7125,s1n7125,notn7125;
or (n7125,s0n7125,s1n7125);
not(notn7125,n5069);
and (s0n7125,notn7125,n7126);
and (s1n7125,n5069,n7127);
and (n7128,n7129,n5083);
wire s0n7129,s1n7129,notn7129;
or (n7129,s0n7129,s1n7129);
not(notn7129,n5069);
and (s0n7129,notn7129,n7130);
and (s1n7129,n5069,n7126);
and (n7131,n7132,n5088);
wire s0n7132,s1n7132,notn7132;
or (n7132,s0n7132,s1n7132);
not(notn7132,n5069);
and (s0n7132,notn7132,n7133);
and (s1n7132,n5069,n7130);
and (n7134,n7135,n5093);
wire s0n7135,s1n7135,notn7135;
or (n7135,s0n7135,s1n7135);
not(notn7135,n5069);
and (s0n7135,notn7135,n7136);
and (s1n7135,n5069,n7133);
and (n7137,n7138,n2744);
or (n7138,1'b0,n7139,n7142,n7145,n7147);
and (n7139,n7140,n5071);
wire s0n7140,s1n7140,notn7140;
or (n7140,s0n7140,s1n7140);
not(notn7140,n5069);
and (s0n7140,notn7140,n7141);
and (s1n7140,n5069,n7136);
and (n7142,n7143,n5083);
wire s0n7143,s1n7143,notn7143;
or (n7143,s0n7143,s1n7143);
not(notn7143,n5069);
and (s0n7143,notn7143,n7144);
and (s1n7143,n5069,n7141);
and (n7145,n7146,n5088);
wire s0n7146,s1n7146,notn7146;
or (n7146,s0n7146,s1n7146);
not(notn7146,n5069);
and (s0n7146,notn7146,n1364);
and (s1n7146,n5069,n7144);
and (n7147,n7148,n5093);
wire s0n7148,s1n7148,notn7148;
or (n7148,s0n7148,s1n7148);
not(notn7148,n5069);
and (s0n7148,notn7148,n812);
and (s1n7148,n5069,n1364);
wire s0n7150,s1n7150,notn7150;
or (n7150,s0n7150,s1n7150);
not(notn7150,n5021);
and (s0n7150,notn7150,n7151);
and (s1n7150,n5021,n7183);
or (n7151,1'b0,n7152,n7167,n7181,n7182);
and (n7152,n7153,n2710);
or (n7153,1'b0,n7154,n7158,n7161,n7164);
and (n7154,n7155,n5071);
wire s0n7155,s1n7155,notn7155;
or (n7155,s0n7155,s1n7155);
not(notn7155,n5069);
and (s0n7155,notn7155,n7156);
and (s1n7155,n5069,n7157);
and (n7158,n7159,n5083);
wire s0n7159,s1n7159,notn7159;
or (n7159,s0n7159,s1n7159);
not(notn7159,n5069);
and (s0n7159,notn7159,n7160);
and (s1n7159,n5069,n7156);
and (n7161,n7162,n5088);
wire s0n7162,s1n7162,notn7162;
or (n7162,s0n7162,s1n7162);
not(notn7162,n5069);
and (s0n7162,notn7162,n7163);
and (s1n7162,n5069,n7160);
and (n7164,n7165,n5093);
wire s0n7165,s1n7165,notn7165;
or (n7165,s0n7165,s1n7165);
not(notn7165,n5069);
and (s0n7165,notn7165,n7166);
and (s1n7165,n5069,n7163);
and (n7167,n7168,n2722);
or (n7168,1'b0,n7169,n7172,n7175,n7178);
and (n7169,n7170,n5071);
wire s0n7170,s1n7170,notn7170;
or (n7170,s0n7170,s1n7170);
not(notn7170,n5069);
and (s0n7170,notn7170,n7171);
and (s1n7170,n5069,n7166);
and (n7172,n7173,n5083);
wire s0n7173,s1n7173,notn7173;
or (n7173,s0n7173,s1n7173);
not(notn7173,n5069);
and (s0n7173,notn7173,n7174);
and (s1n7173,n5069,n7171);
and (n7175,n7176,n5088);
wire s0n7176,s1n7176,notn7176;
or (n7176,s0n7176,s1n7176);
not(notn7176,n5069);
and (s0n7176,notn7176,n7177);
and (s1n7176,n5069,n7174);
and (n7178,n7179,n5093);
wire s0n7179,s1n7179,notn7179;
or (n7179,s0n7179,s1n7179);
not(notn7179,n5069);
and (s0n7179,notn7179,n7180);
and (s1n7179,n5069,n7177);
and (n7181,n5573,n2734);
and (n7182,n5588,n2744);
and (n7184,n7150,n7185);
or (n7185,n7186,n7253,n7391);
and (n7186,n7187,n7219);
wire s0n7187,s1n7187,notn7187;
or (n7187,s0n7187,s1n7187);
not(notn7187,n5021);
and (s0n7187,notn7187,n7188);
and (s1n7187,n5021,n7218);
or (n7188,1'b0,n7189,n7190,n7191,n7206);
and (n7189,n5784,n2710);
and (n7190,n5799,n2722);
and (n7191,n7192,n2734);
or (n7192,1'b0,n7193,n7197,n7200,n7203);
and (n7193,n7194,n5071);
wire s0n7194,s1n7194,notn7194;
or (n7194,s0n7194,s1n7194);
not(notn7194,n5069);
and (s0n7194,notn7194,n7195);
and (s1n7194,n5069,n7196);
and (n7197,n7198,n5083);
wire s0n7198,s1n7198,notn7198;
or (n7198,s0n7198,s1n7198);
not(notn7198,n5069);
and (s0n7198,notn7198,n7199);
and (s1n7198,n5069,n7195);
and (n7200,n7201,n5088);
wire s0n7201,s1n7201,notn7201;
or (n7201,s0n7201,s1n7201);
not(notn7201,n5069);
and (s0n7201,notn7201,n7202);
and (s1n7201,n5069,n7199);
and (n7203,n7204,n5093);
wire s0n7204,s1n7204,notn7204;
or (n7204,s0n7204,s1n7204);
not(notn7204,n5069);
and (s0n7204,notn7204,n7205);
and (s1n7204,n5069,n7202);
and (n7206,n7207,n2744);
or (n7207,1'b0,n7208,n7211,n7214,n7216);
and (n7208,n7209,n5071);
wire s0n7209,s1n7209,notn7209;
or (n7209,s0n7209,s1n7209);
not(notn7209,n5069);
and (s0n7209,notn7209,n7210);
and (s1n7209,n5069,n7205);
and (n7211,n7212,n5083);
wire s0n7212,s1n7212,notn7212;
or (n7212,s0n7212,s1n7212);
not(notn7212,n5069);
and (s0n7212,notn7212,n7213);
and (s1n7212,n5069,n7210);
and (n7214,n7215,n5088);
wire s0n7215,s1n7215,notn7215;
or (n7215,s0n7215,s1n7215);
not(notn7215,n5069);
and (s0n7215,notn7215,n1380);
and (s1n7215,n5069,n7213);
and (n7216,n7217,n5093);
wire s0n7217,s1n7217,notn7217;
or (n7217,s0n7217,s1n7217);
not(notn7217,n5069);
and (s0n7217,notn7217,n833);
and (s1n7217,n5069,n1380);
wire s0n7219,s1n7219,notn7219;
or (n7219,s0n7219,s1n7219);
not(notn7219,n5021);
and (s0n7219,notn7219,n7220);
and (s1n7219,n5021,n7252);
or (n7220,1'b0,n7221,n7236,n7250,n7251);
and (n7221,n7222,n2710);
or (n7222,1'b0,n7223,n7227,n7230,n7233);
and (n7223,n7224,n5071);
wire s0n7224,s1n7224,notn7224;
or (n7224,s0n7224,s1n7224);
not(notn7224,n5069);
and (s0n7224,notn7224,n7225);
and (s1n7224,n5069,n7226);
and (n7227,n7228,n5083);
wire s0n7228,s1n7228,notn7228;
or (n7228,s0n7228,s1n7228);
not(notn7228,n5069);
and (s0n7228,notn7228,n7229);
and (s1n7228,n5069,n7225);
and (n7230,n7231,n5088);
wire s0n7231,s1n7231,notn7231;
or (n7231,s0n7231,s1n7231);
not(notn7231,n5069);
and (s0n7231,notn7231,n7232);
and (s1n7231,n5069,n7229);
and (n7233,n7234,n5093);
wire s0n7234,s1n7234,notn7234;
or (n7234,s0n7234,s1n7234);
not(notn7234,n5069);
and (s0n7234,notn7234,n7235);
and (s1n7234,n5069,n7232);
and (n7236,n7237,n2722);
or (n7237,1'b0,n7238,n7241,n7244,n7247);
and (n7238,n7239,n5071);
wire s0n7239,s1n7239,notn7239;
or (n7239,s0n7239,s1n7239);
not(notn7239,n5069);
and (s0n7239,notn7239,n7240);
and (s1n7239,n5069,n7235);
and (n7241,n7242,n5083);
wire s0n7242,s1n7242,notn7242;
or (n7242,s0n7242,s1n7242);
not(notn7242,n5069);
and (s0n7242,notn7242,n7243);
and (s1n7242,n5069,n7240);
and (n7244,n7245,n5088);
wire s0n7245,s1n7245,notn7245;
or (n7245,s0n7245,s1n7245);
not(notn7245,n5069);
and (s0n7245,notn7245,n7246);
and (s1n7245,n5069,n7243);
and (n7247,n7248,n5093);
wire s0n7248,s1n7248,notn7248;
or (n7248,s0n7248,s1n7248);
not(notn7248,n5069);
and (s0n7248,notn7248,n7249);
and (s1n7248,n5069,n7246);
and (n7250,n5696,n2734);
and (n7251,n5711,n2744);
and (n7253,n7219,n7254);
or (n7254,n7255,n7322,n7390);
and (n7255,n7256,n7288);
wire s0n7256,s1n7256,notn7256;
or (n7256,s0n7256,s1n7256);
not(notn7256,n5021);
and (s0n7256,notn7256,n7257);
and (s1n7256,n5021,n7287);
or (n7257,1'b0,n7258,n7259,n7260,n7275);
and (n7258,n5907,n2710);
and (n7259,n5922,n2722);
and (n7260,n7261,n2734);
or (n7261,1'b0,n7262,n7266,n7269,n7272);
and (n7262,n7263,n5071);
wire s0n7263,s1n7263,notn7263;
or (n7263,s0n7263,s1n7263);
not(notn7263,n5069);
and (s0n7263,notn7263,n7264);
and (s1n7263,n5069,n7265);
and (n7266,n7267,n5083);
wire s0n7267,s1n7267,notn7267;
or (n7267,s0n7267,s1n7267);
not(notn7267,n5069);
and (s0n7267,notn7267,n7268);
and (s1n7267,n5069,n7264);
and (n7269,n7270,n5088);
wire s0n7270,s1n7270,notn7270;
or (n7270,s0n7270,s1n7270);
not(notn7270,n5069);
and (s0n7270,notn7270,n7271);
and (s1n7270,n5069,n7268);
and (n7272,n7273,n5093);
wire s0n7273,s1n7273,notn7273;
or (n7273,s0n7273,s1n7273);
not(notn7273,n5069);
and (s0n7273,notn7273,n7274);
and (s1n7273,n5069,n7271);
and (n7275,n7276,n2744);
or (n7276,1'b0,n7277,n7280,n7283,n7285);
and (n7277,n7278,n5071);
wire s0n7278,s1n7278,notn7278;
or (n7278,s0n7278,s1n7278);
not(notn7278,n5069);
and (s0n7278,notn7278,n7279);
and (s1n7278,n5069,n7274);
and (n7280,n7281,n5083);
wire s0n7281,s1n7281,notn7281;
or (n7281,s0n7281,s1n7281);
not(notn7281,n5069);
and (s0n7281,notn7281,n7282);
and (s1n7281,n5069,n7279);
and (n7283,n7284,n5088);
wire s0n7284,s1n7284,notn7284;
or (n7284,s0n7284,s1n7284);
not(notn7284,n5069);
and (s0n7284,notn7284,n1397);
and (s1n7284,n5069,n7282);
and (n7285,n7286,n5093);
wire s0n7286,s1n7286,notn7286;
or (n7286,s0n7286,s1n7286);
not(notn7286,n5069);
and (s0n7286,notn7286,n863);
and (s1n7286,n5069,n1397);
wire s0n7288,s1n7288,notn7288;
or (n7288,s0n7288,s1n7288);
not(notn7288,n5021);
and (s0n7288,notn7288,n7289);
and (s1n7288,n5021,n7321);
or (n7289,1'b0,n7290,n7305,n7319,n7320);
and (n7290,n7291,n2710);
or (n7291,1'b0,n7292,n7296,n7299,n7302);
and (n7292,n7293,n5071);
wire s0n7293,s1n7293,notn7293;
or (n7293,s0n7293,s1n7293);
not(notn7293,n5069);
and (s0n7293,notn7293,n7294);
and (s1n7293,n5069,n7295);
and (n7296,n7297,n5083);
wire s0n7297,s1n7297,notn7297;
or (n7297,s0n7297,s1n7297);
not(notn7297,n5069);
and (s0n7297,notn7297,n7298);
and (s1n7297,n5069,n7294);
and (n7299,n7300,n5088);
wire s0n7300,s1n7300,notn7300;
or (n7300,s0n7300,s1n7300);
not(notn7300,n5069);
and (s0n7300,notn7300,n7301);
and (s1n7300,n5069,n7298);
and (n7302,n7303,n5093);
wire s0n7303,s1n7303,notn7303;
or (n7303,s0n7303,s1n7303);
not(notn7303,n5069);
and (s0n7303,notn7303,n7304);
and (s1n7303,n5069,n7301);
and (n7305,n7306,n2722);
or (n7306,1'b0,n7307,n7310,n7313,n7316);
and (n7307,n7308,n5071);
wire s0n7308,s1n7308,notn7308;
or (n7308,s0n7308,s1n7308);
not(notn7308,n5069);
and (s0n7308,notn7308,n7309);
and (s1n7308,n5069,n7304);
and (n7310,n7311,n5083);
wire s0n7311,s1n7311,notn7311;
or (n7311,s0n7311,s1n7311);
not(notn7311,n5069);
and (s0n7311,notn7311,n7312);
and (s1n7311,n5069,n7309);
and (n7313,n7314,n5088);
wire s0n7314,s1n7314,notn7314;
or (n7314,s0n7314,s1n7314);
not(notn7314,n5069);
and (s0n7314,notn7314,n7315);
and (s1n7314,n5069,n7312);
and (n7316,n7317,n5093);
wire s0n7317,s1n7317,notn7317;
or (n7317,s0n7317,s1n7317);
not(notn7317,n5069);
and (s0n7317,notn7317,n7318);
and (s1n7317,n5069,n7315);
and (n7319,n5819,n2734);
and (n7320,n5834,n2744);
and (n7322,n7288,n7323);
and (n7323,n7324,n7356);
wire s0n7324,s1n7324,notn7324;
or (n7324,s0n7324,s1n7324);
not(notn7324,n5021);
and (s0n7324,notn7324,n7325);
and (s1n7324,n5021,n7355);
or (n7325,1'b0,n7326,n7327,n7328,n7343);
and (n7326,n6029,n2710);
and (n7327,n6044,n2722);
and (n7328,n7329,n2734);
or (n7329,1'b0,n7330,n7334,n7337,n7340);
and (n7330,n7331,n5071);
wire s0n7331,s1n7331,notn7331;
or (n7331,s0n7331,s1n7331);
not(notn7331,n5069);
and (s0n7331,notn7331,n7332);
and (s1n7331,n5069,n7333);
and (n7334,n7335,n5083);
wire s0n7335,s1n7335,notn7335;
or (n7335,s0n7335,s1n7335);
not(notn7335,n5069);
and (s0n7335,notn7335,n7336);
and (s1n7335,n5069,n7332);
and (n7337,n7338,n5088);
wire s0n7338,s1n7338,notn7338;
or (n7338,s0n7338,s1n7338);
not(notn7338,n5069);
and (s0n7338,notn7338,n7339);
and (s1n7338,n5069,n7336);
and (n7340,n7341,n5093);
wire s0n7341,s1n7341,notn7341;
or (n7341,s0n7341,s1n7341);
not(notn7341,n5069);
and (s0n7341,notn7341,n7342);
and (s1n7341,n5069,n7339);
and (n7343,n7344,n2744);
or (n7344,1'b0,n7345,n7348,n7351,n7353);
and (n7345,n7346,n5071);
wire s0n7346,s1n7346,notn7346;
or (n7346,s0n7346,s1n7346);
not(notn7346,n5069);
and (s0n7346,notn7346,n7347);
and (s1n7346,n5069,n7342);
and (n7348,n7349,n5083);
wire s0n7349,s1n7349,notn7349;
or (n7349,s0n7349,s1n7349);
not(notn7349,n5069);
and (s0n7349,notn7349,n7350);
and (s1n7349,n5069,n7347);
and (n7351,n7352,n5088);
wire s0n7352,s1n7352,notn7352;
or (n7352,s0n7352,s1n7352);
not(notn7352,n5069);
and (s0n7352,notn7352,n1412);
and (s1n7352,n5069,n7350);
and (n7353,n7354,n5093);
wire s0n7354,s1n7354,notn7354;
or (n7354,s0n7354,s1n7354);
not(notn7354,n5069);
and (s0n7354,notn7354,n886);
and (s1n7354,n5069,n1412);
wire s0n7356,s1n7356,notn7356;
or (n7356,s0n7356,s1n7356);
not(notn7356,n5021);
and (s0n7356,notn7356,n7357);
and (s1n7356,n5021,n7389);
or (n7357,1'b0,n7358,n7373,n7387,n7388);
and (n7358,n7359,n2710);
or (n7359,1'b0,n7360,n7364,n7367,n7370);
and (n7360,n7361,n5071);
wire s0n7361,s1n7361,notn7361;
or (n7361,s0n7361,s1n7361);
not(notn7361,n5069);
and (s0n7361,notn7361,n7362);
and (s1n7361,n5069,n7363);
and (n7364,n7365,n5083);
wire s0n7365,s1n7365,notn7365;
or (n7365,s0n7365,s1n7365);
not(notn7365,n5069);
and (s0n7365,notn7365,n7366);
and (s1n7365,n5069,n7362);
and (n7367,n7368,n5088);
wire s0n7368,s1n7368,notn7368;
or (n7368,s0n7368,s1n7368);
not(notn7368,n5069);
and (s0n7368,notn7368,n7369);
and (s1n7368,n5069,n7366);
and (n7370,n7371,n5093);
wire s0n7371,s1n7371,notn7371;
or (n7371,s0n7371,s1n7371);
not(notn7371,n5069);
and (s0n7371,notn7371,n7372);
and (s1n7371,n5069,n7369);
and (n7373,n7374,n2722);
or (n7374,1'b0,n7375,n7378,n7381,n7384);
and (n7375,n7376,n5071);
wire s0n7376,s1n7376,notn7376;
or (n7376,s0n7376,s1n7376);
not(notn7376,n5069);
and (s0n7376,notn7376,n7377);
and (s1n7376,n5069,n7372);
and (n7378,n7379,n5083);
wire s0n7379,s1n7379,notn7379;
or (n7379,s0n7379,s1n7379);
not(notn7379,n5069);
and (s0n7379,notn7379,n7380);
and (s1n7379,n5069,n7377);
and (n7381,n7382,n5088);
wire s0n7382,s1n7382,notn7382;
or (n7382,s0n7382,s1n7382);
not(notn7382,n5069);
and (s0n7382,notn7382,n7383);
and (s1n7382,n5069,n7380);
and (n7384,n7385,n5093);
wire s0n7385,s1n7385,notn7385;
or (n7385,s0n7385,s1n7385);
not(notn7385,n5069);
and (s0n7385,notn7385,n7386);
and (s1n7385,n5069,n7383);
and (n7387,n5941,n2734);
and (n7388,n5956,n2744);
and (n7390,n7256,n7323);
and (n7391,n7187,n7254);
and (n7392,n7118,n7185);
and (n7393,n7049,n7116);
and (n7394,n6980,n7047);
and (n7395,n6911,n6978);
and (n7396,n6842,n6909);
not (n7397,n7398);
nand (n7398,n7399,n7408);
or (n7399,n7400,n7401);
not (n7400,n6828);
not (n7401,n7402);
nand (n7402,n7403,n7407);
or (n7403,n7404,n7405);
not (n7404,n6823);
not (n7405,n7406);
and (n7406,n6819,n6821);
nand (n7407,n6824,n6826);
nor (n7408,n7409,n7412);
and (n7409,n7410,n7411);
not (n7410,n6829);
and (n7411,n6835,n6837);
and (n7412,n6830,n6832);
xor (n7413,n7414,n7416);
wire s0n7414,s1n7414,notn7414;
or (n7414,s0n7414,s1n7414);
not(notn7414,n5021);
and (s0n7414,notn7414,1'b0);
and (s1n7414,n5021,n7415);
wire s0n7416,s1n7416,notn7416;
or (n7416,s0n7416,s1n7416);
not(notn7416,n5021);
and (s0n7416,notn7416,1'b0);
and (s1n7416,n5021,n7417);
and (n7418,n7419,n7420);
not (n7419,n6814);
not (n7420,n7413);
or (n7421,n7422,n7439,n7579);
and (n7422,n7423,n7425);
xor (n7423,n7424,n6085);
xor (n7424,n6080,n6082);
not (n7425,n7426);
nand (n7426,n7427,n7438);
or (n7427,n7428,n7430);
not (n7428,n7429);
xor (n7429,n6830,n6832);
nand (n7430,n7431,n7435);
or (n7431,n7432,n6839);
not (n7432,n7433);
nor (n7433,n7434,n6834);
not (n7434,n6817);
nor (n7435,n7436,n7411);
and (n7436,n7402,n7437);
not (n7437,n6834);
nand (n7438,n7430,n7428);
and (n7439,n7425,n7440);
or (n7440,n7441,n7506,n7578);
and (n7441,n7442,n7444);
xor (n7442,n7443,n6092);
xor (n7443,n6087,n6089);
not (n7444,n7445);
xor (n7445,n7446,n7447);
xor (n7446,n6835,n6837);
nand (n7447,n7448,n7491);
or (n7448,n7449,n7470);
not (n7449,n7450);
and (n7450,n7451,n7463);
nor (n7451,n7452,n7459);
nand (n7452,n7453,n7456);
nand (n7453,n7454,n7455);
not (n7454,n7049);
not (n7455,n7081);
nand (n7456,n7457,n7458);
not (n7457,n7118);
not (n7458,n7150);
not (n7459,n7460);
nand (n7460,n7461,n7462);
not (n7461,n6842);
not (n7462,n6874);
not (n7463,n7464);
nor (n7464,n7465,n7467);
not (n7465,n7466);
not (n7466,n7117);
nand (n7467,n7468,n7469);
not (n7468,n7219);
not (n7469,n7187);
not (n7470,n7471);
nor (n7471,n7472,n7481);
nand (n7472,n7473,n6817);
not (n7473,n7474);
nand (n7474,n7475,n7478);
nand (n7475,n7476,n7477);
not (n7476,n6980);
not (n7477,n7012);
nand (n7478,n7479,n7480);
not (n7479,n6911);
not (n7480,n6943);
not (n7481,n7482);
nand (n7482,n7483,n7485,n7490);
and (n7483,n7484,n7466);
not (n7484,n7255);
nand (n7485,n7486,n7488);
not (n7486,n7487);
nor (n7487,n7256,n7288);
not (n7488,n7489);
not (n7489,n7323);
not (n7490,n7186);
nor (n7491,n7492,n7499);
and (n7492,n7493,n7494,n6817);
and (n7493,n7460,n7478);
not (n7494,n7495);
nand (n7495,n7496,n7475);
nand (n7496,n7497,n7498);
not (n7497,n7048);
not (n7498,n6979);
nand (n7499,n7500,n7401);
or (n7500,n7434,n7501);
not (n7501,n7502);
nand (n7502,n7503,n7505);
or (n7503,n7504,n7459);
not (n7504,n6910);
not (n7505,n6841);
and (n7506,n7444,n7507);
or (n7507,n7508,n7517,n7577);
and (n7508,n7509,n7511);
xor (n7509,n7510,n6181);
xor (n7510,n6094,n6137);
not (n7511,n7512);
xor (n7512,n7513,n7514);
xor (n7513,n6824,n6826);
or (n7514,n7406,n7515,n7516);
and (n7515,n6821,n6840);
and (n7516,n6819,n6840);
and (n7517,n7511,n7518);
or (n7518,n7519,n7525,n7576);
and (n7519,n7520,n7522);
xor (n7520,n7521,n6270);
xor (n7521,n6183,n6226);
not (n7522,n7523);
xor (n7523,n7524,n6840);
xor (n7524,n6819,n6821);
and (n7525,n7522,n7526);
or (n7526,n7527,n7533,n7575);
and (n7527,n7528,n7530);
xor (n7528,n7529,n6359);
xor (n7529,n6272,n6315);
not (n7530,n7531);
xor (n7531,n7532,n6909);
xor (n7532,n6842,n6874);
and (n7533,n7530,n7534);
or (n7534,n7535,n7541,n7574);
and (n7535,n7536,n7538);
xor (n7536,n7537,n6448);
xor (n7537,n6361,n6404);
not (n7538,n7539);
xor (n7539,n7540,n6978);
xor (n7540,n6911,n6943);
and (n7541,n7538,n7542);
or (n7542,n7543,n7549,n7573);
and (n7543,n7544,n7546);
xor (n7544,n7545,n6537);
xor (n7545,n6450,n6493);
not (n7546,n7547);
xor (n7547,n7548,n7047);
xor (n7548,n6980,n7012);
and (n7549,n7546,n7550);
or (n7550,n7551,n7557,n7572);
and (n7551,n7552,n7554);
xor (n7552,n7553,n6626);
xor (n7553,n6539,n6582);
not (n7554,n7555);
xor (n7555,n7556,n7116);
xor (n7556,n7049,n7081);
and (n7557,n7554,n7558);
or (n7558,n7559,n7565,n7571);
and (n7559,n7560,n7562);
xor (n7560,n7561,n6715);
xor (n7561,n6628,n6671);
not (n7562,n7563);
xor (n7563,n7564,n7185);
xor (n7564,n7118,n7150);
and (n7565,n7562,n7566);
and (n7566,n7567,n7568);
xor (n7567,n6716,n6759);
not (n7568,n7569);
xor (n7569,n7570,n7254);
xor (n7570,n7187,n7219);
and (n7571,n7560,n7566);
and (n7572,n7552,n7558);
and (n7573,n7544,n7550);
and (n7574,n7536,n7542);
and (n7575,n7528,n7534);
and (n7576,n7520,n7526);
and (n7577,n7509,n7518);
and (n7578,n7442,n7507);
and (n7579,n7423,n7440);
and (n7580,n7581,n7583);
xor (n7581,n7582,n7440);
xor (n7582,n7423,n7425);
and (n7583,n7584,n7586);
xor (n7584,n7585,n7507);
xor (n7585,n7442,n7444);
and (n7586,n7587,n7589);
xor (n7587,n7588,n7518);
xor (n7588,n7509,n7511);
and (n7589,n7590,n7592);
xor (n7590,n7591,n7526);
xor (n7591,n7520,n7522);
and (n7592,n7593,n7595);
xor (n7593,n7594,n7534);
xor (n7594,n7528,n7530);
and (n7595,n7596,n7598);
xor (n7596,n7597,n7542);
xor (n7597,n7536,n7538);
and (n7598,n7599,n7601);
xor (n7599,n7600,n7550);
xor (n7600,n7544,n7546);
and (n7601,n7602,n7604);
xor (n7602,n7603,n7558);
xor (n7603,n7552,n7554);
and (n7604,n7605,n7607);
xor (n7605,n7606,n7566);
xor (n7606,n7560,n7562);
and (n7607,n7608,n7609);
xor (n7608,n7567,n7568);
and (n7609,n7610,n7613);
not (n7610,n7611);
xor (n7611,n7612,n7323);
xor (n7612,n7256,n7288);
not (n7613,n7614);
xor (n7614,n7324,n7356);
or (n7615,n7616,n7620,n7693);
and (n7616,n7617,n7619);
xor (n7617,n7618,n5038);
xor (n7618,n5033,n5035);
xor (n7619,n7581,n7583);
and (n7620,n7619,n7621);
or (n7621,n7622,n7626,n7692);
and (n7622,n7623,n7625);
xor (n7623,n7624,n5045);
xor (n7624,n5040,n5042);
xor (n7625,n7584,n7586);
and (n7626,n7625,n7627);
or (n7627,n7628,n7632,n7691);
and (n7628,n7629,n7631);
xor (n7629,n7630,n5052);
xor (n7630,n5047,n5049);
xor (n7631,n7587,n7589);
and (n7632,n7631,n7633);
or (n7633,n7634,n7638,n7690);
and (n7634,n7635,n7637);
xor (n7635,n7636,n5059);
xor (n7636,n5054,n5056);
xor (n7637,n7590,n7592);
and (n7638,n7637,n7639);
or (n7639,n7640,n7644,n7689);
and (n7640,n7641,n7643);
xor (n7641,n7642,n5199);
xor (n7642,n5061,n5137);
xor (n7643,n7593,n7595);
and (n7644,n7643,n7645);
or (n7645,n7646,n7650,n7688);
and (n7646,n7647,n7649);
xor (n7647,n7648,n5322);
xor (n7648,n5201,n5260);
xor (n7649,n7596,n7598);
and (n7650,n7649,n7651);
or (n7651,n7652,n7656,n7687);
and (n7652,n7653,n7655);
xor (n7653,n7654,n5445);
xor (n7654,n5324,n5383);
xor (n7655,n7599,n7601);
and (n7656,n7655,n7657);
or (n7657,n7658,n7662,n7686);
and (n7658,n7659,n7661);
xor (n7659,n7660,n5568);
xor (n7660,n5447,n5506);
xor (n7661,n7602,n7604);
and (n7662,n7661,n7663);
or (n7663,n7664,n7668,n7685);
and (n7664,n7665,n7667);
xor (n7665,n7666,n5691);
xor (n7666,n5570,n5629);
xor (n7667,n7605,n7607);
and (n7668,n7667,n7669);
or (n7669,n7670,n7674,n7684);
and (n7670,n7671,n7673);
xor (n7671,n7672,n5814);
xor (n7672,n5693,n5752);
xor (n7673,n7608,n7609);
and (n7674,n7673,n7675);
or (n7675,n7676,n7680,n7683);
and (n7676,n7677,n7679);
xor (n7677,n7678,n5937);
xor (n7678,n5816,n5875);
xor (n7679,n7610,n7613);
and (n7680,n7679,n7681);
and (n7681,n7682,n7614);
xor (n7682,n5938,n5997);
and (n7683,n7677,n7681);
and (n7684,n7671,n7675);
and (n7685,n7665,n7669);
and (n7686,n7659,n7663);
and (n7687,n7653,n7657);
and (n7688,n7647,n7651);
and (n7689,n7641,n7645);
and (n7690,n7635,n7639);
and (n7691,n7629,n7633);
and (n7692,n7623,n7627);
and (n7693,n7617,n7621);
or (n7694,n7695,n7698,n7750);
and (n7695,n7696,n7631);
xor (n7696,n7697,n7621);
xor (n7697,n7617,n7619);
and (n7698,n7631,n7699);
or (n7699,n7700,n7703,n7749);
and (n7700,n7701,n7637);
xor (n7701,n7702,n7627);
xor (n7702,n7623,n7625);
and (n7703,n7637,n7704);
or (n7704,n7705,n7708,n7748);
and (n7705,n7706,n7643);
xor (n7706,n7707,n7633);
xor (n7707,n7629,n7631);
and (n7708,n7643,n7709);
or (n7709,n7710,n7713,n7747);
and (n7710,n7711,n7649);
xor (n7711,n7712,n7639);
xor (n7712,n7635,n7637);
and (n7713,n7649,n7714);
or (n7714,n7715,n7718,n7746);
and (n7715,n7716,n7655);
xor (n7716,n7717,n7645);
xor (n7717,n7641,n7643);
and (n7718,n7655,n7719);
or (n7719,n7720,n7723,n7745);
and (n7720,n7721,n7661);
xor (n7721,n7722,n7651);
xor (n7722,n7647,n7649);
and (n7723,n7661,n7724);
or (n7724,n7725,n7728,n7744);
and (n7725,n7726,n7667);
xor (n7726,n7727,n7657);
xor (n7727,n7653,n7655);
and (n7728,n7667,n7729);
or (n7729,n7730,n7733,n7743);
and (n7730,n7731,n7673);
xor (n7731,n7732,n7663);
xor (n7732,n7659,n7661);
and (n7733,n7673,n7734);
or (n7734,n7735,n7738,n7742);
and (n7735,n7736,n7679);
xor (n7736,n7737,n7669);
xor (n7737,n7665,n7667);
and (n7738,n7679,n7739);
and (n7739,n7740,n7614);
xor (n7740,n7741,n7675);
xor (n7741,n7671,n7673);
and (n7742,n7736,n7739);
and (n7743,n7731,n7734);
and (n7744,n7726,n7729);
and (n7745,n7721,n7724);
and (n7746,n7716,n7719);
and (n7747,n7711,n7714);
and (n7748,n7706,n7709);
and (n7749,n7701,n7704);
and (n7750,n7696,n7699);
and (n7751,n7752,n7754);
xor (n7752,n7753,n7699);
xor (n7753,n7696,n7631);
and (n7754,n7755,n7757);
xor (n7755,n7756,n7704);
xor (n7756,n7701,n7637);
and (n7757,n7758,n7760);
xor (n7758,n7759,n7709);
xor (n7759,n7706,n7643);
and (n7760,n7761,n7763);
xor (n7761,n7762,n7714);
xor (n7762,n7711,n7649);
and (n7763,n7764,n7766);
xor (n7764,n7765,n7719);
xor (n7765,n7716,n7655);
and (n7766,n7767,n7769);
xor (n7767,n7768,n7724);
xor (n7768,n7721,n7661);
and (n7769,n7770,n7772);
xor (n7770,n7771,n7729);
xor (n7771,n7726,n7667);
xor (n7772,n7773,n7734);
xor (n7773,n7731,n7673);
xor (n7774,n5013,n7775);
and (n7775,n7752,n7776);
and (n7776,n7755,n7758);
wire s0n7777,s1n7777,notn7777;
or (n7777,s0n7777,s1n7777);
not(notn7777,n5021);
and (s0n7777,notn7777,n7778);
and (s1n7777,n5021,n8011);
xor (n7778,n7779,n7998);
xor (n7779,n7780,n7970);
xor (n7780,n7781,n7949);
xor (n7781,n7782,n7943);
xor (n7782,n7783,n7805);
xor (n7783,n7784,n7789);
xor (n7784,n7785,n7787);
wire s0n7785,s1n7785,notn7785;
or (n7785,s0n7785,s1n7785);
not(notn7785,n5021);
and (s0n7785,notn7785,1'b0);
and (s1n7785,n5021,n7786);
wire s0n7787,s1n7787,notn7787;
or (n7787,s0n7787,s1n7787);
not(notn7787,n5021);
and (s0n7787,notn7787,1'b0);
and (s1n7787,n5021,n7788);
or (n7789,n7790,n7791,n7804);
and (n7790,n7785,n7787);
and (n7791,n7787,n7792);
or (n7792,n7793,n7798,n7803);
and (n7793,n7794,n7796);
wire s0n7794,s1n7794,notn7794;
or (n7794,s0n7794,s1n7794);
not(notn7794,n5021);
and (s0n7794,notn7794,1'b0);
and (s1n7794,n5021,n7795);
wire s0n7796,s1n7796,notn7796;
or (n7796,s0n7796,s1n7796);
not(notn7796,n5021);
and (s0n7796,notn7796,1'b0);
and (s1n7796,n5021,n7797);
and (n7798,n7796,n7799);
or (n7799,n7800,n7801,n7802);
and (n7800,n5019,n5029);
and (n7801,n5029,n5031);
and (n7802,n5019,n5031);
and (n7803,n7794,n7799);
and (n7804,n7785,n7792);
xor (n7805,n7806,n7930);
xor (n7806,n7807,n7875);
xor (n7807,n7808,n7846);
xor (n7808,n7809,n7814);
xor (n7809,n7810,n7812);
wire s0n7810,s1n7810,notn7810;
or (n7810,s0n7810,s1n7810);
not(notn7810,n5021);
and (s0n7810,notn7810,1'b0);
and (s1n7810,n5021,n7811);
wire s0n7812,s1n7812,notn7812;
or (n7812,s0n7812,s1n7812);
not(notn7812,n5021);
and (s0n7812,notn7812,1'b0);
and (s1n7812,n5021,n7813);
or (n7814,n7815,n7816,n7845);
and (n7815,n7810,n7812);
and (n7816,n7812,n7817);
or (n7817,n7818,n7823,n7844);
and (n7818,n7819,n7821);
wire s0n7819,s1n7819,notn7819;
or (n7819,s0n7819,s1n7819);
not(notn7819,n5021);
and (s0n7819,notn7819,1'b0);
and (s1n7819,n5021,n7820);
wire s0n7821,s1n7821,notn7821;
or (n7821,s0n7821,s1n7821);
not(notn7821,n5021);
and (s0n7821,notn7821,1'b0);
and (s1n7821,n5021,n7822);
and (n7823,n7821,n7824);
or (n7824,n7825,n7830,n7843);
and (n7825,n7826,n7828);
wire s0n7826,s1n7826,notn7826;
or (n7826,s0n7826,s1n7826);
not(notn7826,n5021);
and (s0n7826,notn7826,1'b0);
and (s1n7826,n5021,n7827);
wire s0n7828,s1n7828,notn7828;
or (n7828,s0n7828,s1n7828);
not(notn7828,n5021);
and (s0n7828,notn7828,1'b0);
and (s1n7828,n5021,n7829);
and (n7830,n7828,n7831);
or (n7831,n7832,n7837,n7842);
and (n7832,n7833,n7835);
wire s0n7833,s1n7833,notn7833;
or (n7833,s0n7833,s1n7833);
not(notn7833,n5021);
and (s0n7833,notn7833,1'b0);
and (s1n7833,n5021,n7834);
wire s0n7835,s1n7835,notn7835;
or (n7835,s0n7835,s1n7835);
not(notn7835,n5021);
and (s0n7835,notn7835,1'b0);
and (s1n7835,n5021,n7836);
and (n7837,n7835,n7838);
or (n7838,n7839,n7840,n7841);
and (n7839,n6074,n6076);
and (n7840,n6076,n6078);
and (n7841,n6074,n6078);
and (n7842,n7833,n7838);
and (n7843,n7826,n7831);
and (n7844,n7819,n7824);
and (n7845,n7810,n7817);
not (n7846,n7847);
nor (n7847,n7848,n7864);
and (n7848,n6840,n7849);
nor (n7849,n7850,n6816);
not (n7850,n7851);
nor (n7851,n7852,n7859);
nand (n7852,n7853,n7854);
or (n7853,n7414,n7416);
or (n7854,n7855,n7857);
wire s0n7855,s1n7855,notn7855;
or (n7855,s0n7855,s1n7855);
not(notn7855,n5021);
and (s0n7855,notn7855,1'b0);
and (s1n7855,n5021,n7856);
wire s0n7857,s1n7857,notn7857;
or (n7857,s0n7857,s1n7857);
not(notn7857,n5021);
and (s0n7857,notn7857,1'b0);
and (s1n7857,n5021,n7858);
and (n7859,n7860,n7862);
wire s0n7860,s1n7860,notn7860;
or (n7860,s0n7860,s1n7860);
not(notn7860,n5021);
and (s0n7860,notn7860,1'b0);
and (s1n7860,n5021,n7861);
wire s0n7862,s1n7862,notn7862;
or (n7862,s0n7862,s1n7862);
not(notn7862,n5021);
and (s0n7862,notn7862,1'b0);
and (s1n7862,n5021,n7863);
nand (n7864,n7865,n7866);
or (n7865,n7397,n7850);
nor (n7866,n7867,n7874);
and (n7867,n7868,n7873);
nand (n7868,n7869,n7872);
or (n7869,n7870,n7871);
nand (n7870,n7414,n7416);
not (n7871,n7854);
nand (n7872,n7855,n7857);
not (n7873,n7859);
nor (n7874,n7860,n7862);
or (n7875,n7876,n7878,n7929);
and (n7876,n7877,n7846);
xor (n7877,n7809,n7817);
and (n7878,n7846,n7879);
or (n7879,n7880,n7883,n7928);
and (n7880,n7881,n7846);
xor (n7881,n7882,n7824);
xor (n7882,n7819,n7821);
and (n7883,n7846,n7884);
or (n7884,n7885,n7901,n7927);
and (n7885,n7886,n7888);
xor (n7886,n7887,n7831);
xor (n7887,n7826,n7828);
not (n7888,n7889);
nand (n7889,n7890,n7900);
or (n7890,n7891,n7893);
not (n7891,n7892);
xor (n7892,n7860,n7862);
nand (n7893,n7894,n7897);
or (n7894,n7895,n6839);
not (n7895,n7896);
nor (n7896,n6816,n7852);
nor (n7897,n7898,n7868);
and (n7898,n7398,n7899);
not (n7899,n7852);
nand (n7900,n7893,n7891);
and (n7901,n7888,n7902);
or (n7902,n7903,n7921,n7926);
and (n7903,n7904,n7906);
xor (n7904,n7905,n7838);
xor (n7905,n7833,n7835);
not (n7906,n7907);
nor (n7907,n7908,n7918);
and (n7908,n7909,n7917);
nand (n7909,n7910,n7914);
or (n7910,n7911,n6839);
not (n7911,n7912);
nor (n7912,n7913,n6816);
not (n7913,n7853);
nor (n7914,n7915,n7916);
and (n7915,n7398,n7853);
not (n7916,n7870);
xor (n7917,n7855,n7857);
and (n7918,n7919,n7920);
not (n7919,n7909);
not (n7920,n7917);
and (n7921,n7906,n7922);
or (n7922,n7923,n7924,n7925);
and (n7923,n6072,n6811);
and (n7924,n6811,n7421);
and (n7925,n6072,n7421);
and (n7926,n7904,n7922);
and (n7927,n7886,n7902);
and (n7928,n7881,n7884);
and (n7929,n7877,n7879);
and (n7930,n7931,n7933);
xor (n7931,n7932,n7879);
xor (n7932,n7877,n7846);
and (n7933,n7934,n7936);
xor (n7934,n7935,n7884);
xor (n7935,n7881,n7846);
and (n7936,n7937,n7939);
xor (n7937,n7938,n7902);
xor (n7938,n7886,n7888);
and (n7939,n7940,n7942);
xor (n7940,n7941,n7922);
xor (n7941,n7904,n7906);
and (n7942,n6070,n7580);
or (n7943,n7944,n7946,n7969);
and (n7944,n7783,n7945);
xor (n7945,n7931,n7933);
and (n7946,n7945,n7947);
or (n7947,n7948,n7950,n7968);
and (n7948,n7783,n7949);
xor (n7949,n7934,n7936);
and (n7950,n7949,n7951);
or (n7951,n7952,n7955,n7967);
and (n7952,n7953,n7954);
xor (n7953,n7784,n7792);
xor (n7954,n7937,n7939);
and (n7955,n7954,n7956);
or (n7956,n7957,n7961,n7966);
and (n7957,n7958,n7960);
xor (n7958,n7959,n7799);
xor (n7959,n7794,n7796);
xor (n7960,n7940,n7942);
and (n7961,n7960,n7962);
or (n7962,n7963,n7964,n7965);
and (n7963,n5017,n6069);
and (n7964,n6069,n7615);
and (n7965,n5017,n7615);
and (n7966,n7958,n7962);
and (n7967,n7953,n7956);
and (n7968,n7783,n7951);
and (n7969,n7783,n7947);
or (n7970,n7971,n7974,n7997);
and (n7971,n7972,n7954);
xor (n7972,n7973,n7947);
xor (n7973,n7783,n7945);
and (n7974,n7954,n7975);
or (n7975,n7976,n7979,n7996);
and (n7976,n7977,n7960);
xor (n7977,n7978,n7951);
xor (n7978,n7783,n7949);
and (n7979,n7960,n7980);
or (n7980,n7981,n7984,n7995);
and (n7981,n7982,n6069);
xor (n7982,n7983,n7956);
xor (n7983,n7953,n7954);
and (n7984,n6069,n7985);
or (n7985,n7986,n7989,n7994);
and (n7986,n7987,n7619);
xor (n7987,n7988,n7962);
xor (n7988,n7958,n7960);
and (n7989,n7619,n7990);
or (n7990,n7991,n7992,n7993);
and (n7991,n5015,n7625);
and (n7992,n7625,n7694);
and (n7993,n5015,n7694);
and (n7994,n7987,n7990);
and (n7995,n7982,n7985);
and (n7996,n7977,n7980);
and (n7997,n7972,n7975);
and (n7998,n7999,n8001);
xor (n7999,n8000,n7975);
xor (n8000,n7972,n7954);
and (n8001,n8002,n8004);
xor (n8002,n8003,n7980);
xor (n8003,n7977,n7960);
and (n8004,n8005,n8007);
xor (n8005,n8006,n7985);
xor (n8006,n7982,n6069);
and (n8007,n8008,n8010);
xor (n8008,n8009,n7990);
xor (n8009,n7987,n7619);
and (n8010,n5013,n7751);
xor (n8011,n7779,n8012);
and (n8012,n7999,n8013);
and (n8013,n8002,n8014);
and (n8014,n8005,n8015);
and (n8015,n8008,n8016);
and (n8016,n5013,n7775);
wire s0n8017,s1n8017,notn8017;
or (n8017,s0n8017,s1n8017);
not(notn8017,n5021);
and (s0n8017,notn8017,n8018);
and (s1n8017,n5021,n8021);
wire s0n8018,s1n8018,notn8018;
or (n8018,s0n8018,s1n8018);
not(notn8018,n5021);
and (s0n8018,notn8018,n8019);
and (s1n8018,n5021,n8020);
xor (n8019,n8008,n8010);
xor (n8020,n8008,n8016);
wire s0n8021,s1n8021,notn8021;
or (n8021,s0n8021,s1n8021);
not(notn8021,n5021);
and (s0n8021,notn8021,n8022);
and (s1n8021,n5021,n8030);
xor (n8022,n8023,n8029);
xor (n8023,n8024,n8025);
xor (n8024,n7781,n7945);
or (n8025,n8026,n8027,n8028);
and (n8026,n7781,n7949);
and (n8027,n7949,n7970);
and (n8028,n7781,n7970);
and (n8029,n7779,n7998);
xor (n8030,n8023,n8031);
and (n8031,n7779,n8012);
wire s0n8032,s1n8032,notn8032;
or (n8032,s0n8032,s1n8032);
not(notn8032,n5021);
and (s0n8032,notn8032,n8033);
and (s1n8032,n5021,n8041);
xor (n8033,n8034,n8040);
xor (n8034,n8035,n8036);
xor (n8035,n7781,n7805);
or (n8036,n8037,n8038,n8039);
and (n8037,n7781,n7945);
and (n8038,n7945,n8025);
and (n8039,n7781,n8025);
and (n8040,n8023,n8029);
xor (n8041,n8034,n8042);
and (n8042,n8023,n8031);
and (n8043,n8044,n2899);
wire s0n8044,s1n8044,notn8044;
or (n8044,s0n8044,s1n8044);
not(notn8044,n2894);
and (s0n8044,notn8044,1'b0);
and (s1n8044,n2894,n5008);
and (n8045,n5008,n8046);
or (n8046,n8047,n4938);
or (n8047,n4959,n4950);
and (n8048,n2903,n8049);
or (n8049,n2934,n2936);
and (n8050,n5005,n8051);
or (n8051,n8052,n8162,n8822);
and (n8052,n8053,n8146);
or (n8053,1'b0,n8054,n8057,n8060,n8065);
and (n8054,n8055,n2885);
wire s0n8055,s1n8055,notn8055;
or (n8055,s0n8055,s1n8055);
not(notn8055,n2883);
and (s0n8055,notn8055,1'b0);
and (s1n8055,n2883,n8056);
and (n8057,n8058,n2899);
wire s0n8058,s1n8058,notn8058;
or (n8058,s0n8058,s1n8058);
not(notn8058,n2894);
and (s0n8058,notn8058,1'b0);
and (s1n8058,n2894,n8059);
and (n8060,n8061,n4938);
wire s0n8061,s1n8061,notn8061;
or (n8061,s0n8061,s1n8061);
not(notn8061,n4933);
and (s0n8061,notn8061,n8062);
and (s1n8061,n4933,1'b0);
wire s0n8062,s1n8062,notn8062;
or (n8062,s0n8062,s1n8062);
not(notn8062,n4928);
and (s0n8062,notn8062,n8063);
and (s1n8062,n4928,1'b1);
wire s0n8063,s1n8063,notn8063;
or (n8063,s0n8063,s1n8063);
not(notn8063,n4916);
and (s0n8063,notn8063,1'b0);
and (s1n8063,n4916,n8064);
xor (n8064,n4894,n4896);
or (n8065,1'b0,n8066,n8086,n8106,n8126);
and (n8066,n8067,n2710);
or (n8067,1'b0,n8068,n8074,n8080);
and (n8068,n8069,n4950);
or (n8069,1'b0,n8070,n8071,n8072,n8073);
and (n8070,n3052,n549);
and (n8071,n3056,n560);
and (n8072,n3060,n564);
and (n8073,n3064,n566);
and (n8074,n8075,n2936);
or (n8075,1'b0,n8076,n8077,n8078,n8079);
and (n8076,n3122,n549);
and (n8077,n3051,n560);
and (n8078,n3055,n564);
and (n8079,n3059,n566);
and (n8080,n8081,n4958);
or (n8081,1'b0,n8082,n8083,n8084,n8085);
and (n8082,n3051,n549);
and (n8083,n3055,n560);
and (n8084,n3059,n564);
and (n8085,n3063,n566);
and (n8086,n8087,n2722);
or (n8087,1'b0,n8088,n8094,n8100);
and (n8088,n8089,n4950);
or (n8089,1'b0,n8090,n8091,n8092,n8093);
and (n8090,n3070,n549);
and (n8091,n3074,n560);
and (n8092,n3078,n564);
and (n8093,n3082,n566);
and (n8094,n8095,n2936);
or (n8095,1'b0,n8096,n8097,n8098,n8099);
and (n8096,n3063,n549);
and (n8097,n3069,n560);
and (n8098,n3073,n564);
and (n8099,n3077,n566);
and (n8100,n8101,n4958);
or (n8101,1'b0,n8102,n8103,n8104,n8105);
and (n8102,n3069,n549);
and (n8103,n3073,n560);
and (n8104,n3077,n564);
and (n8105,n3081,n566);
and (n8106,n8107,n2734);
or (n8107,1'b0,n8108,n8114,n8120);
and (n8108,n8109,n4950);
or (n8109,1'b0,n8110,n8111,n8112,n8113);
and (n8110,n3088,n549);
and (n8111,n3092,n560);
and (n8112,n3096,n564);
and (n8113,n3100,n566);
and (n8114,n8115,n2936);
or (n8115,1'b0,n8116,n8117,n8118,n8119);
and (n8116,n3137,n549);
and (n8117,n3087,n560);
and (n8118,n3091,n564);
and (n8119,n3095,n566);
and (n8120,n8121,n4958);
or (n8121,1'b0,n8122,n8123,n8124,n8125);
and (n8122,n3087,n549);
and (n8123,n3091,n560);
and (n8124,n3095,n564);
and (n8125,n3099,n566);
and (n8126,n8127,n2744);
or (n8127,1'b0,n8128,n8134,n8140);
and (n8128,n8129,n4950);
or (n8129,1'b0,n8130,n8131,n8132,n8133);
and (n8130,n3106,n549);
and (n8131,n3110,n560);
and (n8132,n3113,n564);
and (n8133,n3116,n566);
and (n8134,n8135,n2936);
or (n8135,1'b0,n8136,n8137,n8138,n8139);
and (n8136,n3099,n549);
and (n8137,n3105,n560);
and (n8138,n3109,n564);
and (n8139,n2180,n566);
and (n8140,n8141,n4958);
or (n8141,1'b0,n8142,n8143,n8144,n8145);
and (n8142,n3105,n549);
and (n8143,n3109,n560);
and (n8144,n2180,n564);
and (n8145,n1844,n566);
or (n8146,1'b0,n8147,n8158,n8160,n8161);
and (n8147,n8148,n2885);
wire s0n8148,s1n8148,notn8148;
or (n8148,s0n8148,s1n8148);
not(notn8148,n2883);
and (s0n8148,notn8148,1'b0);
and (s1n8148,n2883,n8149);
wire s0n8149,s1n8149,notn8149;
or (n8149,s0n8149,s1n8149);
not(notn8149,n8032);
and (s0n8149,notn8149,n8150);
and (s1n8149,n8032,1'b0);
wire s0n8150,s1n8150,notn8150;
or (n8150,s0n8150,s1n8150);
not(notn8150,n8017);
and (s0n8150,notn8150,n8151);
and (s1n8150,n8017,1'b1);
wire s0n8151,s1n8151,notn8151;
or (n8151,s0n8151,s1n8151);
not(notn8151,n5021);
and (s0n8151,notn8151,n8152);
and (s1n8151,n5021,n8155);
wire s0n8152,s1n8152,notn8152;
or (n8152,s0n8152,s1n8152);
not(notn8152,n5021);
and (s0n8152,notn8152,n8153);
and (s1n8152,n5021,n8154);
xor (n8153,n7752,n7754);
xor (n8154,n7752,n7776);
wire s0n8155,s1n8155,notn8155;
or (n8155,s0n8155,s1n8155);
not(notn8155,n5021);
and (s0n8155,notn8155,n8156);
and (s1n8155,n5021,n8157);
xor (n8156,n7999,n8001);
xor (n8157,n7999,n8013);
and (n8158,n8159,n2899);
wire s0n8159,s1n8159,notn8159;
or (n8159,s0n8159,s1n8159);
not(notn8159,n2894);
and (s0n8159,notn8159,1'b0);
and (s1n8159,n2894,n8149);
and (n8160,n8149,n8046);
and (n8161,n8061,n8049);
and (n8162,n8146,n8163);
or (n8163,n8164,n8274,n8821);
and (n8164,n8165,n8258);
or (n8165,1'b0,n8166,n8169,n8172,n8177);
and (n8166,n8167,n2885);
wire s0n8167,s1n8167,notn8167;
or (n8167,s0n8167,s1n8167);
not(notn8167,n2883);
and (s0n8167,notn8167,1'b0);
and (s1n8167,n2883,n8168);
and (n8169,n8170,n2899);
wire s0n8170,s1n8170,notn8170;
or (n8170,s0n8170,s1n8170);
not(notn8170,n2894);
and (s0n8170,notn8170,1'b0);
and (s1n8170,n2894,n8171);
and (n8172,n8173,n4938);
wire s0n8173,s1n8173,notn8173;
or (n8173,s0n8173,s1n8173);
not(notn8173,n4933);
and (s0n8173,notn8173,n8174);
and (s1n8173,n4933,1'b0);
wire s0n8174,s1n8174,notn8174;
or (n8174,s0n8174,s1n8174);
not(notn8174,n4928);
and (s0n8174,notn8174,n8175);
and (s1n8174,n4928,1'b1);
wire s0n8175,s1n8175,notn8175;
or (n8175,s0n8175,s1n8175);
not(notn8175,n4916);
and (s0n8175,notn8175,1'b0);
and (s1n8175,n4916,n8176);
xor (n8176,n4897,n4899);
or (n8177,1'b0,n8178,n8198,n8218,n8238);
and (n8178,n8179,n2710);
or (n8179,1'b0,n8180,n8186,n8192);
and (n8180,n8181,n4950);
or (n8181,1'b0,n8182,n8183,n8184,n8185);
and (n8182,n3157,n549);
and (n8183,n3161,n560);
and (n8184,n3165,n564);
and (n8185,n3169,n566);
and (n8186,n8187,n2936);
or (n8187,1'b0,n8188,n8189,n8190,n8191);
and (n8188,n3227,n549);
and (n8189,n3156,n560);
and (n8190,n3160,n564);
and (n8191,n3164,n566);
and (n8192,n8193,n4958);
or (n8193,1'b0,n8194,n8195,n8196,n8197);
and (n8194,n3156,n549);
and (n8195,n3160,n560);
and (n8196,n3164,n564);
and (n8197,n3168,n566);
and (n8198,n8199,n2722);
or (n8199,1'b0,n8200,n8206,n8212);
and (n8200,n8201,n4950);
or (n8201,1'b0,n8202,n8203,n8204,n8205);
and (n8202,n3175,n549);
and (n8203,n3179,n560);
and (n8204,n3183,n564);
and (n8205,n3187,n566);
and (n8206,n8207,n2936);
or (n8207,1'b0,n8208,n8209,n8210,n8211);
and (n8208,n3168,n549);
and (n8209,n3174,n560);
and (n8210,n3178,n564);
and (n8211,n3182,n566);
and (n8212,n8213,n4958);
or (n8213,1'b0,n8214,n8215,n8216,n8217);
and (n8214,n3174,n549);
and (n8215,n3178,n560);
and (n8216,n3182,n564);
and (n8217,n3186,n566);
and (n8218,n8219,n2734);
or (n8219,1'b0,n8220,n8226,n8232);
and (n8220,n8221,n4950);
or (n8221,1'b0,n8222,n8223,n8224,n8225);
and (n8222,n3193,n549);
and (n8223,n3197,n560);
and (n8224,n3201,n564);
and (n8225,n3205,n566);
and (n8226,n8227,n2936);
or (n8227,1'b0,n8228,n8229,n8230,n8231);
and (n8228,n3242,n549);
and (n8229,n3192,n560);
and (n8230,n3196,n564);
and (n8231,n3200,n566);
and (n8232,n8233,n4958);
or (n8233,1'b0,n8234,n8235,n8236,n8237);
and (n8234,n3192,n549);
and (n8235,n3196,n560);
and (n8236,n3200,n564);
and (n8237,n3204,n566);
and (n8238,n8239,n2744);
or (n8239,1'b0,n8240,n8246,n8252);
and (n8240,n8241,n4950);
or (n8241,1'b0,n8242,n8243,n8244,n8245);
and (n8242,n3211,n549);
and (n8243,n3215,n560);
and (n8244,n3218,n564);
and (n8245,n3221,n566);
and (n8246,n8247,n2936);
or (n8247,1'b0,n8248,n8249,n8250,n8251);
and (n8248,n3204,n549);
and (n8249,n3210,n560);
and (n8250,n3214,n564);
and (n8251,n2196,n566);
and (n8252,n8253,n4958);
or (n8253,1'b0,n8254,n8255,n8256,n8257);
and (n8254,n3210,n549);
and (n8255,n3214,n560);
and (n8256,n2196,n564);
and (n8257,n1861,n566);
or (n8258,1'b0,n8259,n8270,n8272,n8273);
and (n8259,n8260,n2885);
wire s0n8260,s1n8260,notn8260;
or (n8260,s0n8260,s1n8260);
not(notn8260,n2883);
and (s0n8260,notn8260,1'b0);
and (s1n8260,n2883,n8261);
wire s0n8261,s1n8261,notn8261;
or (n8261,s0n8261,s1n8261);
not(notn8261,n8032);
and (s0n8261,notn8261,n8262);
and (s1n8261,n8032,1'b0);
wire s0n8262,s1n8262,notn8262;
or (n8262,s0n8262,s1n8262);
not(notn8262,n8017);
and (s0n8262,notn8262,n8263);
and (s1n8262,n8017,1'b1);
wire s0n8263,s1n8263,notn8263;
or (n8263,s0n8263,s1n8263);
not(notn8263,n5021);
and (s0n8263,notn8263,n8264);
and (s1n8263,n5021,n8267);
wire s0n8264,s1n8264,notn8264;
or (n8264,s0n8264,s1n8264);
not(notn8264,n5021);
and (s0n8264,notn8264,n8265);
and (s1n8264,n5021,n8266);
xor (n8265,n7755,n7757);
xor (n8266,n7755,n7758);
wire s0n8267,s1n8267,notn8267;
or (n8267,s0n8267,s1n8267);
not(notn8267,n5021);
and (s0n8267,notn8267,n8268);
and (s1n8267,n5021,n8269);
xor (n8268,n8002,n8004);
xor (n8269,n8002,n8014);
and (n8270,n8271,n2899);
wire s0n8271,s1n8271,notn8271;
or (n8271,s0n8271,s1n8271);
not(notn8271,n2894);
and (s0n8271,notn8271,1'b0);
and (s1n8271,n2894,n8261);
and (n8272,n8261,n8046);
and (n8273,n8173,n8049);
and (n8274,n8258,n8275);
or (n8275,n8276,n8386,n8820);
and (n8276,n8277,n8370);
or (n8277,1'b0,n8278,n8281,n8284,n8289);
and (n8278,n8279,n2885);
wire s0n8279,s1n8279,notn8279;
or (n8279,s0n8279,s1n8279);
not(notn8279,n2883);
and (s0n8279,notn8279,1'b0);
and (s1n8279,n2883,n8280);
and (n8281,n8282,n2899);
wire s0n8282,s1n8282,notn8282;
or (n8282,s0n8282,s1n8282);
not(notn8282,n2894);
and (s0n8282,notn8282,1'b0);
and (s1n8282,n2894,n8283);
and (n8284,n8285,n4938);
wire s0n8285,s1n8285,notn8285;
or (n8285,s0n8285,s1n8285);
not(notn8285,n4933);
and (s0n8285,notn8285,n8286);
and (s1n8285,n4933,1'b0);
wire s0n8286,s1n8286,notn8286;
or (n8286,s0n8286,s1n8286);
not(notn8286,n4928);
and (s0n8286,notn8286,n8287);
and (s1n8286,n4928,1'b1);
wire s0n8287,s1n8287,notn8287;
or (n8287,s0n8287,s1n8287);
not(notn8287,n4916);
and (s0n8287,notn8287,1'b0);
and (s1n8287,n4916,n8288);
xor (n8288,n4900,n4902);
or (n8289,1'b0,n8290,n8310,n8330,n8350);
and (n8290,n8291,n2710);
or (n8291,1'b0,n8292,n8298,n8304);
and (n8292,n8293,n4950);
or (n8293,1'b0,n8294,n8295,n8296,n8297);
and (n8294,n3262,n549);
and (n8295,n3266,n560);
and (n8296,n3270,n564);
and (n8297,n3274,n566);
and (n8298,n8299,n2936);
or (n8299,1'b0,n8300,n8301,n8302,n8303);
and (n8300,n3332,n549);
and (n8301,n3261,n560);
and (n8302,n3265,n564);
and (n8303,n3269,n566);
and (n8304,n8305,n4958);
or (n8305,1'b0,n8306,n8307,n8308,n8309);
and (n8306,n3261,n549);
and (n8307,n3265,n560);
and (n8308,n3269,n564);
and (n8309,n3273,n566);
and (n8310,n8311,n2722);
or (n8311,1'b0,n8312,n8318,n8324);
and (n8312,n8313,n4950);
or (n8313,1'b0,n8314,n8315,n8316,n8317);
and (n8314,n3280,n549);
and (n8315,n3284,n560);
and (n8316,n3288,n564);
and (n8317,n3292,n566);
and (n8318,n8319,n2936);
or (n8319,1'b0,n8320,n8321,n8322,n8323);
and (n8320,n3273,n549);
and (n8321,n3279,n560);
and (n8322,n3283,n564);
and (n8323,n3287,n566);
and (n8324,n8325,n4958);
or (n8325,1'b0,n8326,n8327,n8328,n8329);
and (n8326,n3279,n549);
and (n8327,n3283,n560);
and (n8328,n3287,n564);
and (n8329,n3291,n566);
and (n8330,n8331,n2734);
or (n8331,1'b0,n8332,n8338,n8344);
and (n8332,n8333,n4950);
or (n8333,1'b0,n8334,n8335,n8336,n8337);
and (n8334,n3298,n549);
and (n8335,n3302,n560);
and (n8336,n3306,n564);
and (n8337,n3310,n566);
and (n8338,n8339,n2936);
or (n8339,1'b0,n8340,n8341,n8342,n8343);
and (n8340,n3347,n549);
and (n8341,n3297,n560);
and (n8342,n3301,n564);
and (n8343,n3305,n566);
and (n8344,n8345,n4958);
or (n8345,1'b0,n8346,n8347,n8348,n8349);
and (n8346,n3297,n549);
and (n8347,n3301,n560);
and (n8348,n3305,n564);
and (n8349,n3309,n566);
and (n8350,n8351,n2744);
or (n8351,1'b0,n8352,n8358,n8364);
and (n8352,n8353,n4950);
or (n8353,1'b0,n8354,n8355,n8356,n8357);
and (n8354,n3316,n549);
and (n8355,n3320,n560);
and (n8356,n3323,n564);
and (n8357,n3326,n566);
and (n8358,n8359,n2936);
or (n8359,1'b0,n8360,n8361,n8362,n8363);
and (n8360,n3309,n549);
and (n8361,n3315,n560);
and (n8362,n3319,n564);
and (n8363,n2212,n566);
and (n8364,n8365,n4958);
or (n8365,1'b0,n8366,n8367,n8368,n8369);
and (n8366,n3315,n549);
and (n8367,n3319,n560);
and (n8368,n2212,n564);
and (n8369,n1886,n566);
or (n8370,1'b0,n8371,n8382,n8384,n8385);
and (n8371,n8372,n2885);
wire s0n8372,s1n8372,notn8372;
or (n8372,s0n8372,s1n8372);
not(notn8372,n2883);
and (s0n8372,notn8372,1'b0);
and (s1n8372,n2883,n8373);
wire s0n8373,s1n8373,notn8373;
or (n8373,s0n8373,s1n8373);
not(notn8373,n8032);
and (s0n8373,notn8373,n8374);
and (s1n8373,n8032,1'b0);
wire s0n8374,s1n8374,notn8374;
or (n8374,s0n8374,s1n8374);
not(notn8374,n8017);
and (s0n8374,notn8374,n8375);
and (s1n8374,n8017,1'b1);
wire s0n8375,s1n8375,notn8375;
or (n8375,s0n8375,s1n8375);
not(notn8375,n5021);
and (s0n8375,notn8375,n8376);
and (s1n8375,n5021,n8379);
wire s0n8376,s1n8376,notn8376;
or (n8376,s0n8376,s1n8376);
not(notn8376,n5021);
and (s0n8376,notn8376,n8377);
and (s1n8376,n5021,n8378);
xor (n8377,n7758,n7760);
not (n8378,n7758);
wire s0n8379,s1n8379,notn8379;
or (n8379,s0n8379,s1n8379);
not(notn8379,n5021);
and (s0n8379,notn8379,n8380);
and (s1n8379,n5021,n8381);
xor (n8380,n8005,n8007);
xor (n8381,n8005,n8015);
and (n8382,n8383,n2899);
wire s0n8383,s1n8383,notn8383;
or (n8383,s0n8383,s1n8383);
not(notn8383,n2894);
and (s0n8383,notn8383,1'b0);
and (s1n8383,n2894,n8373);
and (n8384,n8373,n8046);
and (n8385,n8285,n8049);
and (n8386,n8370,n8387);
or (n8387,n8388,n8494,n8819);
and (n8388,n8389,n8482);
or (n8389,1'b0,n8390,n8393,n8396,n8401);
and (n8390,n8391,n2885);
wire s0n8391,s1n8391,notn8391;
or (n8391,s0n8391,s1n8391);
not(notn8391,n2883);
and (s0n8391,notn8391,1'b0);
and (s1n8391,n2883,n8392);
and (n8393,n8394,n2899);
wire s0n8394,s1n8394,notn8394;
or (n8394,s0n8394,s1n8394);
not(notn8394,n2894);
and (s0n8394,notn8394,1'b0);
and (s1n8394,n2894,n8395);
and (n8396,n8397,n4938);
wire s0n8397,s1n8397,notn8397;
or (n8397,s0n8397,s1n8397);
not(notn8397,n4933);
and (s0n8397,notn8397,n8398);
and (s1n8397,n4933,1'b0);
wire s0n8398,s1n8398,notn8398;
or (n8398,s0n8398,s1n8398);
not(notn8398,n4928);
and (s0n8398,notn8398,n8399);
and (s1n8398,n4928,1'b1);
wire s0n8399,s1n8399,notn8399;
or (n8399,s0n8399,s1n8399);
not(notn8399,n4916);
and (s0n8399,notn8399,1'b0);
and (s1n8399,n4916,n8400);
xor (n8400,n4903,n4905);
or (n8401,1'b0,n8402,n8422,n8442,n8462);
and (n8402,n8403,n2710);
or (n8403,1'b0,n8404,n8410,n8416);
and (n8404,n8405,n4950);
or (n8405,1'b0,n8406,n8407,n8408,n8409);
and (n8406,n3367,n549);
and (n8407,n3371,n560);
and (n8408,n3375,n564);
and (n8409,n3379,n566);
and (n8410,n8411,n2936);
or (n8411,1'b0,n8412,n8413,n8414,n8415);
and (n8412,n3437,n549);
and (n8413,n3366,n560);
and (n8414,n3370,n564);
and (n8415,n3374,n566);
and (n8416,n8417,n4958);
or (n8417,1'b0,n8418,n8419,n8420,n8421);
and (n8418,n3366,n549);
and (n8419,n3370,n560);
and (n8420,n3374,n564);
and (n8421,n3378,n566);
and (n8422,n8423,n2722);
or (n8423,1'b0,n8424,n8430,n8436);
and (n8424,n8425,n4950);
or (n8425,1'b0,n8426,n8427,n8428,n8429);
and (n8426,n3385,n549);
and (n8427,n3389,n560);
and (n8428,n3393,n564);
and (n8429,n3397,n566);
and (n8430,n8431,n2936);
or (n8431,1'b0,n8432,n8433,n8434,n8435);
and (n8432,n3378,n549);
and (n8433,n3384,n560);
and (n8434,n3388,n564);
and (n8435,n3392,n566);
and (n8436,n8437,n4958);
or (n8437,1'b0,n8438,n8439,n8440,n8441);
and (n8438,n3384,n549);
and (n8439,n3388,n560);
and (n8440,n3392,n564);
and (n8441,n3396,n566);
and (n8442,n8443,n2734);
or (n8443,1'b0,n8444,n8450,n8456);
and (n8444,n8445,n4950);
or (n8445,1'b0,n8446,n8447,n8448,n8449);
and (n8446,n3403,n549);
and (n8447,n3407,n560);
and (n8448,n3411,n564);
and (n8449,n3415,n566);
and (n8450,n8451,n2936);
or (n8451,1'b0,n8452,n8453,n8454,n8455);
and (n8452,n3452,n549);
and (n8453,n3402,n560);
and (n8454,n3406,n564);
and (n8455,n3410,n566);
and (n8456,n8457,n4958);
or (n8457,1'b0,n8458,n8459,n8460,n8461);
and (n8458,n3402,n549);
and (n8459,n3406,n560);
and (n8460,n3410,n564);
and (n8461,n3414,n566);
and (n8462,n8463,n2744);
or (n8463,1'b0,n8464,n8470,n8476);
and (n8464,n8465,n4950);
or (n8465,1'b0,n8466,n8467,n8468,n8469);
and (n8466,n3421,n549);
and (n8467,n3425,n560);
and (n8468,n3428,n564);
and (n8469,n3431,n566);
and (n8470,n8471,n2936);
or (n8471,1'b0,n8472,n8473,n8474,n8475);
and (n8472,n3414,n549);
and (n8473,n3420,n560);
and (n8474,n3424,n564);
and (n8475,n2228,n566);
and (n8476,n8477,n4958);
or (n8477,1'b0,n8478,n8479,n8480,n8481);
and (n8478,n3420,n549);
and (n8479,n3424,n560);
and (n8480,n2228,n564);
and (n8481,n1913,n566);
or (n8482,1'b0,n8483,n8490,n8492,n8493);
and (n8483,n8484,n2885);
wire s0n8484,s1n8484,notn8484;
or (n8484,s0n8484,s1n8484);
not(notn8484,n2883);
and (s0n8484,notn8484,1'b0);
and (s1n8484,n2883,n8485);
wire s0n8485,s1n8485,notn8485;
or (n8485,s0n8485,s1n8485);
not(notn8485,n8032);
and (s0n8485,notn8485,n8486);
and (s1n8485,n8032,1'b0);
wire s0n8486,s1n8486,notn8486;
or (n8486,s0n8486,s1n8486);
not(notn8486,n8017);
and (s0n8486,notn8486,n8487);
and (s1n8486,n8017,1'b1);
wire s0n8487,s1n8487,notn8487;
or (n8487,s0n8487,s1n8487);
not(notn8487,n5021);
and (s0n8487,notn8487,n8488);
and (s1n8487,n5021,n8018);
wire s0n8488,s1n8488,notn8488;
or (n8488,s0n8488,s1n8488);
not(notn8488,n5021);
and (s0n8488,notn8488,n8489);
and (s1n8488,n5021,n7761);
xor (n8489,n7761,n7763);
and (n8490,n8491,n2899);
wire s0n8491,s1n8491,notn8491;
or (n8491,s0n8491,s1n8491);
not(notn8491,n2894);
and (s0n8491,notn8491,1'b0);
and (s1n8491,n2894,n8485);
and (n8492,n8485,n8046);
and (n8493,n8397,n8049);
and (n8494,n8482,n8495);
or (n8495,n8496,n8602,n8818);
and (n8496,n8497,n8590);
or (n8497,1'b0,n8498,n8501,n8504,n8509);
and (n8498,n8499,n2885);
wire s0n8499,s1n8499,notn8499;
or (n8499,s0n8499,s1n8499);
not(notn8499,n2883);
and (s0n8499,notn8499,1'b0);
and (s1n8499,n2883,n8500);
and (n8501,n8502,n2899);
wire s0n8502,s1n8502,notn8502;
or (n8502,s0n8502,s1n8502);
not(notn8502,n2894);
and (s0n8502,notn8502,1'b0);
and (s1n8502,n2894,n8503);
and (n8504,n8505,n4938);
wire s0n8505,s1n8505,notn8505;
or (n8505,s0n8505,s1n8505);
not(notn8505,n4933);
and (s0n8505,notn8505,n8506);
and (s1n8505,n4933,1'b0);
wire s0n8506,s1n8506,notn8506;
or (n8506,s0n8506,s1n8506);
not(notn8506,n4928);
and (s0n8506,notn8506,n8507);
and (s1n8506,n4928,1'b1);
wire s0n8507,s1n8507,notn8507;
or (n8507,s0n8507,s1n8507);
not(notn8507,n4916);
and (s0n8507,notn8507,1'b0);
and (s1n8507,n4916,n8508);
xor (n8508,n4906,n4908);
or (n8509,1'b0,n8510,n8530,n8550,n8570);
and (n8510,n8511,n2710);
or (n8511,1'b0,n8512,n8518,n8524);
and (n8512,n8513,n4950);
or (n8513,1'b0,n8514,n8515,n8516,n8517);
and (n8514,n3472,n549);
and (n8515,n3476,n560);
and (n8516,n3480,n564);
and (n8517,n3484,n566);
and (n8518,n8519,n2936);
or (n8519,1'b0,n8520,n8521,n8522,n8523);
and (n8520,n3542,n549);
and (n8521,n3471,n560);
and (n8522,n3475,n564);
and (n8523,n3479,n566);
and (n8524,n8525,n4958);
or (n8525,1'b0,n8526,n8527,n8528,n8529);
and (n8526,n3471,n549);
and (n8527,n3475,n560);
and (n8528,n3479,n564);
and (n8529,n3483,n566);
and (n8530,n8531,n2722);
or (n8531,1'b0,n8532,n8538,n8544);
and (n8532,n8533,n4950);
or (n8533,1'b0,n8534,n8535,n8536,n8537);
and (n8534,n3490,n549);
and (n8535,n3494,n560);
and (n8536,n3498,n564);
and (n8537,n3502,n566);
and (n8538,n8539,n2936);
or (n8539,1'b0,n8540,n8541,n8542,n8543);
and (n8540,n3483,n549);
and (n8541,n3489,n560);
and (n8542,n3493,n564);
and (n8543,n3497,n566);
and (n8544,n8545,n4958);
or (n8545,1'b0,n8546,n8547,n8548,n8549);
and (n8546,n3489,n549);
and (n8547,n3493,n560);
and (n8548,n3497,n564);
and (n8549,n3501,n566);
and (n8550,n8551,n2734);
or (n8551,1'b0,n8552,n8558,n8564);
and (n8552,n8553,n4950);
or (n8553,1'b0,n8554,n8555,n8556,n8557);
and (n8554,n3508,n549);
and (n8555,n3512,n560);
and (n8556,n3516,n564);
and (n8557,n3520,n566);
and (n8558,n8559,n2936);
or (n8559,1'b0,n8560,n8561,n8562,n8563);
and (n8560,n3557,n549);
and (n8561,n3507,n560);
and (n8562,n3511,n564);
and (n8563,n3515,n566);
and (n8564,n8565,n4958);
or (n8565,1'b0,n8566,n8567,n8568,n8569);
and (n8566,n3507,n549);
and (n8567,n3511,n560);
and (n8568,n3515,n564);
and (n8569,n3519,n566);
and (n8570,n8571,n2744);
or (n8571,1'b0,n8572,n8578,n8584);
and (n8572,n8573,n4950);
or (n8573,1'b0,n8574,n8575,n8576,n8577);
and (n8574,n3526,n549);
and (n8575,n3530,n560);
and (n8576,n3533,n564);
and (n8577,n3536,n566);
and (n8578,n8579,n2936);
or (n8579,1'b0,n8580,n8581,n8582,n8583);
and (n8580,n3519,n549);
and (n8581,n3525,n560);
and (n8582,n3529,n564);
and (n8583,n2244,n566);
and (n8584,n8585,n4958);
or (n8585,1'b0,n8586,n8587,n8588,n8589);
and (n8586,n3525,n549);
and (n8587,n3529,n560);
and (n8588,n2244,n564);
and (n8589,n1939,n566);
or (n8590,1'b0,n8591,n8598,n8600,n8601);
and (n8591,n8592,n2885);
wire s0n8592,s1n8592,notn8592;
or (n8592,s0n8592,s1n8592);
not(notn8592,n2883);
and (s0n8592,notn8592,1'b0);
and (s1n8592,n2883,n8593);
wire s0n8593,s1n8593,notn8593;
or (n8593,s0n8593,s1n8593);
not(notn8593,n8032);
and (s0n8593,notn8593,n8594);
and (s1n8593,n8032,1'b0);
wire s0n8594,s1n8594,notn8594;
or (n8594,s0n8594,s1n8594);
not(notn8594,n8017);
and (s0n8594,notn8594,n8595);
and (s1n8594,n8017,1'b1);
wire s0n8595,s1n8595,notn8595;
or (n8595,s0n8595,s1n8595);
not(notn8595,n5021);
and (s0n8595,notn8595,n8596);
and (s1n8595,n5021,n5011);
wire s0n8596,s1n8596,notn8596;
or (n8596,s0n8596,s1n8596);
not(notn8596,n5021);
and (s0n8596,notn8596,n8597);
and (s1n8596,n5021,n7764);
xor (n8597,n7764,n7766);
and (n8598,n8599,n2899);
wire s0n8599,s1n8599,notn8599;
or (n8599,s0n8599,s1n8599);
not(notn8599,n2894);
and (s0n8599,notn8599,1'b0);
and (s1n8599,n2894,n8593);
and (n8600,n8593,n8046);
and (n8601,n8505,n8049);
and (n8602,n8590,n8603);
or (n8603,n8604,n8710,n8817);
and (n8604,n8605,n8698);
or (n8605,1'b0,n8606,n8609,n8612,n8617);
and (n8606,n8607,n2885);
wire s0n8607,s1n8607,notn8607;
or (n8607,s0n8607,s1n8607);
not(notn8607,n2883);
and (s0n8607,notn8607,1'b0);
and (s1n8607,n2883,n8608);
and (n8609,n8610,n2899);
wire s0n8610,s1n8610,notn8610;
or (n8610,s0n8610,s1n8610);
not(notn8610,n2894);
and (s0n8610,notn8610,1'b0);
and (s1n8610,n2894,n8611);
and (n8612,n8613,n4938);
wire s0n8613,s1n8613,notn8613;
or (n8613,s0n8613,s1n8613);
not(notn8613,n4933);
and (s0n8613,notn8613,n8614);
and (s1n8613,n4933,1'b0);
wire s0n8614,s1n8614,notn8614;
or (n8614,s0n8614,s1n8614);
not(notn8614,n4928);
and (s0n8614,notn8614,n8615);
and (s1n8614,n4928,1'b1);
wire s0n8615,s1n8615,notn8615;
or (n8615,s0n8615,s1n8615);
not(notn8615,n4916);
and (s0n8615,notn8615,1'b0);
and (s1n8615,n4916,n8616);
xor (n8616,n4909,n4911);
or (n8617,1'b0,n8618,n8638,n8658,n8678);
and (n8618,n8619,n2710);
or (n8619,1'b0,n8620,n8626,n8632);
and (n8620,n8621,n4950);
or (n8621,1'b0,n8622,n8623,n8624,n8625);
and (n8622,n3577,n549);
and (n8623,n3581,n560);
and (n8624,n3585,n564);
and (n8625,n3589,n566);
and (n8626,n8627,n2936);
or (n8627,1'b0,n8628,n8629,n8630,n8631);
and (n8628,n3647,n549);
and (n8629,n3576,n560);
and (n8630,n3580,n564);
and (n8631,n3584,n566);
and (n8632,n8633,n4958);
or (n8633,1'b0,n8634,n8635,n8636,n8637);
and (n8634,n3576,n549);
and (n8635,n3580,n560);
and (n8636,n3584,n564);
and (n8637,n3588,n566);
and (n8638,n8639,n2722);
or (n8639,1'b0,n8640,n8646,n8652);
and (n8640,n8641,n4950);
or (n8641,1'b0,n8642,n8643,n8644,n8645);
and (n8642,n3595,n549);
and (n8643,n3599,n560);
and (n8644,n3603,n564);
and (n8645,n3607,n566);
and (n8646,n8647,n2936);
or (n8647,1'b0,n8648,n8649,n8650,n8651);
and (n8648,n3588,n549);
and (n8649,n3594,n560);
and (n8650,n3598,n564);
and (n8651,n3602,n566);
and (n8652,n8653,n4958);
or (n8653,1'b0,n8654,n8655,n8656,n8657);
and (n8654,n3594,n549);
and (n8655,n3598,n560);
and (n8656,n3602,n564);
and (n8657,n3606,n566);
and (n8658,n8659,n2734);
or (n8659,1'b0,n8660,n8666,n8672);
and (n8660,n8661,n4950);
or (n8661,1'b0,n8662,n8663,n8664,n8665);
and (n8662,n3613,n549);
and (n8663,n3617,n560);
and (n8664,n3621,n564);
and (n8665,n3625,n566);
and (n8666,n8667,n2936);
or (n8667,1'b0,n8668,n8669,n8670,n8671);
and (n8668,n3662,n549);
and (n8669,n3612,n560);
and (n8670,n3616,n564);
and (n8671,n3620,n566);
and (n8672,n8673,n4958);
or (n8673,1'b0,n8674,n8675,n8676,n8677);
and (n8674,n3612,n549);
and (n8675,n3616,n560);
and (n8676,n3620,n564);
and (n8677,n3624,n566);
and (n8678,n8679,n2744);
or (n8679,1'b0,n8680,n8686,n8692);
and (n8680,n8681,n4950);
or (n8681,1'b0,n8682,n8683,n8684,n8685);
and (n8682,n3631,n549);
and (n8683,n3635,n560);
and (n8684,n3638,n564);
and (n8685,n3641,n566);
and (n8686,n8687,n2936);
or (n8687,1'b0,n8688,n8689,n8690,n8691);
and (n8688,n3624,n549);
and (n8689,n3630,n560);
and (n8690,n3634,n564);
and (n8691,n2260,n566);
and (n8692,n8693,n4958);
or (n8693,1'b0,n8694,n8695,n8696,n8697);
and (n8694,n3630,n549);
and (n8695,n3634,n560);
and (n8696,n2260,n564);
and (n8697,n1968,n566);
or (n8698,1'b0,n8699,n8706,n8708,n8709);
and (n8699,n8700,n2885);
wire s0n8700,s1n8700,notn8700;
or (n8700,s0n8700,s1n8700);
not(notn8700,n2883);
and (s0n8700,notn8700,1'b0);
and (s1n8700,n2883,n8701);
wire s0n8701,s1n8701,notn8701;
or (n8701,s0n8701,s1n8701);
not(notn8701,n8032);
and (s0n8701,notn8701,n8702);
and (s1n8701,n8032,1'b0);
wire s0n8702,s1n8702,notn8702;
or (n8702,s0n8702,s1n8702);
not(notn8702,n8017);
and (s0n8702,notn8702,n8703);
and (s1n8702,n8017,1'b1);
wire s0n8703,s1n8703,notn8703;
or (n8703,s0n8703,s1n8703);
not(notn8703,n5021);
and (s0n8703,notn8703,n8704);
and (s1n8703,n5021,n8152);
wire s0n8704,s1n8704,notn8704;
or (n8704,s0n8704,s1n8704);
not(notn8704,n5021);
and (s0n8704,notn8704,n8705);
and (s1n8704,n5021,n7767);
xor (n8705,n7767,n7769);
and (n8706,n8707,n2899);
wire s0n8707,s1n8707,notn8707;
or (n8707,s0n8707,s1n8707);
not(notn8707,n2894);
and (s0n8707,notn8707,1'b0);
and (s1n8707,n2894,n8701);
and (n8708,n8701,n8046);
and (n8709,n8613,n8049);
and (n8710,n8698,n8711);
and (n8711,n8712,n8805);
or (n8712,1'b0,n8713,n8716,n8719,n8724);
and (n8713,n8714,n2885);
wire s0n8714,s1n8714,notn8714;
or (n8714,s0n8714,s1n8714);
not(notn8714,n2883);
and (s0n8714,notn8714,1'b0);
and (s1n8714,n2883,n8715);
and (n8716,n8717,n2899);
wire s0n8717,s1n8717,notn8717;
or (n8717,s0n8717,s1n8717);
not(notn8717,n2894);
and (s0n8717,notn8717,1'b0);
and (s1n8717,n2894,n8718);
and (n8719,n8720,n4938);
wire s0n8720,s1n8720,notn8720;
or (n8720,s0n8720,s1n8720);
not(notn8720,n4933);
and (s0n8720,notn8720,n8721);
and (s1n8720,n4933,1'b0);
wire s0n8721,s1n8721,notn8721;
or (n8721,s0n8721,s1n8721);
not(notn8721,n4928);
and (s0n8721,notn8721,n8722);
and (s1n8721,n4928,1'b1);
wire s0n8722,s1n8722,notn8722;
or (n8722,s0n8722,s1n8722);
not(notn8722,n4916);
and (s0n8722,notn8722,1'b0);
and (s1n8722,n4916,n8723);
xor (n8723,n4912,n4914);
or (n8724,1'b0,n8725,n8745,n8765,n8785);
and (n8725,n8726,n2710);
or (n8726,1'b0,n8727,n8733,n8739);
and (n8727,n8728,n4950);
or (n8728,1'b0,n8729,n8730,n8731,n8732);
and (n8729,n3681,n549);
and (n8730,n3685,n560);
and (n8731,n3689,n564);
and (n8732,n3693,n566);
and (n8733,n8734,n2936);
or (n8734,1'b0,n8735,n8736,n8737,n8738);
and (n8735,n3751,n549);
and (n8736,n3680,n560);
and (n8737,n3684,n564);
and (n8738,n3688,n566);
and (n8739,n8740,n4958);
or (n8740,1'b0,n8741,n8742,n8743,n8744);
and (n8741,n3680,n549);
and (n8742,n3684,n560);
and (n8743,n3688,n564);
and (n8744,n3692,n566);
and (n8745,n8746,n2722);
or (n8746,1'b0,n8747,n8753,n8759);
and (n8747,n8748,n4950);
or (n8748,1'b0,n8749,n8750,n8751,n8752);
and (n8749,n3699,n549);
and (n8750,n3703,n560);
and (n8751,n3707,n564);
and (n8752,n3711,n566);
and (n8753,n8754,n2936);
or (n8754,1'b0,n8755,n8756,n8757,n8758);
and (n8755,n3692,n549);
and (n8756,n3698,n560);
and (n8757,n3702,n564);
and (n8758,n3706,n566);
and (n8759,n8760,n4958);
or (n8760,1'b0,n8761,n8762,n8763,n8764);
and (n8761,n3698,n549);
and (n8762,n3702,n560);
and (n8763,n3706,n564);
and (n8764,n3710,n566);
and (n8765,n8766,n2734);
or (n8766,1'b0,n8767,n8773,n8779);
and (n8767,n8768,n4950);
or (n8768,1'b0,n8769,n8770,n8771,n8772);
and (n8769,n3717,n549);
and (n8770,n3721,n560);
and (n8771,n3725,n564);
and (n8772,n3729,n566);
and (n8773,n8774,n2936);
or (n8774,1'b0,n8775,n8776,n8777,n8778);
and (n8775,n3766,n549);
and (n8776,n3716,n560);
and (n8777,n3720,n564);
and (n8778,n3724,n566);
and (n8779,n8780,n4958);
or (n8780,1'b0,n8781,n8782,n8783,n8784);
and (n8781,n3716,n549);
and (n8782,n3720,n560);
and (n8783,n3724,n564);
and (n8784,n3728,n566);
and (n8785,n8786,n2744);
or (n8786,1'b0,n8787,n8793,n8799);
and (n8787,n8788,n4950);
or (n8788,1'b0,n8789,n8790,n8791,n8792);
and (n8789,n3735,n549);
and (n8790,n3739,n560);
and (n8791,n3742,n564);
and (n8792,n3745,n566);
and (n8793,n8794,n2936);
or (n8794,1'b0,n8795,n8796,n8797,n8798);
and (n8795,n3728,n549);
and (n8796,n3734,n560);
and (n8797,n3738,n564);
and (n8798,n2275,n566);
and (n8799,n8800,n4958);
or (n8800,1'b0,n8801,n8802,n8803,n8804);
and (n8801,n3734,n549);
and (n8802,n3738,n560);
and (n8803,n2275,n564);
and (n8804,n1987,n566);
or (n8805,1'b0,n8806,n8813,n8815,n8816);
and (n8806,n8807,n2885);
wire s0n8807,s1n8807,notn8807;
or (n8807,s0n8807,s1n8807);
not(notn8807,n2883);
and (s0n8807,notn8807,1'b0);
and (s1n8807,n2883,n8808);
wire s0n8808,s1n8808,notn8808;
or (n8808,s0n8808,s1n8808);
not(notn8808,n8032);
and (s0n8808,notn8808,n8809);
and (s1n8808,n8032,1'b0);
wire s0n8809,s1n8809,notn8809;
or (n8809,s0n8809,s1n8809);
not(notn8809,n8017);
and (s0n8809,notn8809,n8810);
and (s1n8809,n8017,1'b1);
wire s0n8810,s1n8810,notn8810;
or (n8810,s0n8810,s1n8810);
not(notn8810,n5021);
and (s0n8810,notn8810,n8811);
and (s1n8810,n5021,n8264);
wire s0n8811,s1n8811,notn8811;
or (n8811,s0n8811,s1n8811);
not(notn8811,n5021);
and (s0n8811,notn8811,n8812);
and (s1n8811,n5021,n7770);
xor (n8812,n7770,n7772);
and (n8813,n8814,n2899);
wire s0n8814,s1n8814,notn8814;
or (n8814,s0n8814,s1n8814);
not(notn8814,n2894);
and (s0n8814,notn8814,1'b0);
and (s1n8814,n2894,n8808);
and (n8815,n8808,n8046);
and (n8816,n8720,n8049);
and (n8817,n8605,n8711);
and (n8818,n8497,n8603);
and (n8819,n8389,n8495);
and (n8820,n8277,n8387);
and (n8821,n8165,n8275);
and (n8822,n8053,n8163);
and (n8823,n2879,n8051);
and (n8824,n8825,n8827);
xor (n8825,n8826,n8051);
xor (n8826,n2879,n5005);
and (n8827,n8828,n8830);
xor (n8828,n8829,n8163);
xor (n8829,n8053,n8146);
and (n8830,n8831,n8833);
xor (n8831,n8832,n8275);
xor (n8832,n8165,n8258);
and (n8833,n8834,n8836);
xor (n8834,n8835,n8387);
xor (n8835,n8277,n8370);
and (n8836,n8837,n8839);
xor (n8837,n8838,n8495);
xor (n8838,n8389,n8482);
and (n8839,n8840,n8842);
xor (n8840,n8841,n8603);
xor (n8841,n8497,n8590);
and (n8842,n8843,n8845);
xor (n8843,n8844,n8711);
xor (n8844,n8605,n8698);
xor (n8845,n8712,n8805);
and (n8846,n8847,n8848);
wire s0n8847,s1n8847,notn8847;
or (n8847,s0n8847,s1n8847);
not(notn8847,n5024);
and (s0n8847,notn8847,1'b0);
and (s1n8847,n5024,n2876);
or (n8848,n8849,n2889);
or (n8849,n8850,n2886);
or (n8850,n8851,n2923);
or (n8851,n8852,n2922);
or (n8852,n8853,n4950);
or (n8853,n8854,n2938);
or (n8854,n8855,n2937);
or (n8855,n8049,n4959);
and (n8856,n5007,n2942);
and (n8857,n5008,n5079);
and (n8858,n2903,n2933);
nor (n8859,n2748,n2900,n2901);
and (n8860,n583,n2696);
nand (n8861,n8862,n8863);
not (n8862,n2873);
nor (n8863,n2692,n8864);
and (n8864,n8865,n9686);
nand (n8865,n8866,n9661);
not (n8866,n8867);
or (n8867,n8868,n9660);
and (n8868,n8869,n9261);
xor (n8869,n8870,n9203);
xor (n8870,n8871,n9152);
xor (n8871,n8872,n9127);
or (n8872,n8873,n9126);
and (n8873,n8874,n8996);
xor (n8874,n8875,n8971);
xor (n8875,n8876,n8920);
xor (n8876,n8877,n8879);
xor (n8877,n8878,n1209);
xor (n8878,n1082,n2088);
xor (n8879,n8880,n2334);
xor (n8880,n8881,n8918);
or (n8881,n8882,n8917);
and (n8882,n8883,n2415);
xor (n8883,n8884,n1645);
and (n8884,n8885,n1653);
xor (n8885,n1652,n8886);
xor (n8886,n8887,n8897);
xor (n8887,n8888,n8894);
xor (n8888,n8889,n8893);
xor (n8889,n8890,n8892);
nor (n8890,n8891,n1026);
not (n8891,n2158);
and (n8892,n1294,n1027);
and (n8893,n8892,n1310);
and (n8894,n8890,n8895);
not (n8895,n8896);
not (n8896,n2174);
or (n8897,n8898,n8916);
and (n8898,n8899,n8908);
xor (n8899,n8900,n8901);
nor (n8900,n1505,n1026);
and (n8901,n8902,n1027);
nand (n8902,n8903,n8907);
or (n8903,n8904,n8905);
not (n8904,n2171);
not (n8905,n8906);
not (n8906,n2289);
or (n8907,n8906,n2171);
and (n8908,n8909,n1027);
or (n8909,n8910,n8914);
nor (n8910,n8911,n8896);
and (n8911,n8912,n8913);
not (n8912,n2294);
not (n8913,n2186);
nor (n8914,n8915,n8891);
not (n8915,n2218);
and (n8916,n8900,n8901);
and (n8917,n8884,n1645);
xor (n8918,n8919,n1638);
xor (n8919,n1485,n1637);
or (n8920,n8921,n8970);
and (n8921,n8922,n8928);
xor (n8922,n8923,n8927);
or (n8923,n8924,n8926);
and (n8924,n8925,n1224);
xor (n8925,n2099,n2028);
and (n8926,n2099,n2028);
xor (n8927,n8883,n2415);
and (n8928,n8929,n1091);
xor (n8929,n1223,n8930);
or (n8930,n8931,n8969);
and (n8931,n8932,n8954);
xor (n8932,n2427,n8933);
and (n8933,n8934,n8948);
or (n8934,n8935,n8947);
and (n8935,n8936,n8946);
xor (n8936,n8937,n8945);
and (n8937,n8938,n1027);
nand (n8938,n8939,n8941,n8944);
or (n8939,n8940,n8912);
not (n8940,n2250);
or (n8941,n8942,n8943);
not (n8942,n2300);
not (n8943,n2222);
not (n8944,n2205);
and (n8945,n1529,n1027);
nor (n8946,n1526,n1026);
and (n8947,n8937,n8945);
and (n8948,n8949,n1027);
nor (n8949,n8950,n8952);
and (n8950,n8951,n8895);
xor (n8951,n8912,n8913);
and (n8952,n8953,n8896);
not (n8953,n8951);
or (n8954,n8955,n8968);
and (n8955,n8956,n2433);
xor (n8956,n1669,n8957);
xor (n8957,n8958,n8967);
xor (n8958,n8959,n8960);
and (n8959,n1516,n1027);
and (n8960,n8961,n1027);
nand (n8961,n8962,n8966);
or (n8962,n8963,n8942);
and (n8963,n8964,n8965);
not (n8964,n2190);
not (n8965,n2202);
not (n8966,n2189);
and (n8967,n1511,n1027);
and (n8968,n1669,n8957);
and (n8969,n2427,n8933);
and (n8970,n8923,n8927);
xor (n8971,n8972,n8992);
xor (n8972,n8973,n8982);
xor (n8973,n8974,n2410);
xor (n8974,n1208,n8975);
and (n8975,n8976,n8979);
or (n8976,n8977,n8978);
and (n8977,n8887,n8897);
and (n8978,n8888,n8894);
or (n8979,n8980,n8981);
and (n8980,n8889,n8893);
and (n8981,n8890,n8892);
or (n8982,n8983,n8991);
and (n8983,n8984,n1216);
xor (n8984,n8985,n2093);
or (n8985,n8986,n8990);
and (n8986,n8987,n2344);
xor (n8987,n8988,n8989);
xor (n8988,n8885,n1653);
and (n8989,n1659,n1581);
and (n8990,n8988,n8989);
and (n8991,n8985,n2093);
or (n8992,n8993,n8995);
and (n8993,n8994,n1086);
xor (n8994,n1087,n2024);
and (n8995,n1087,n2024);
or (n8996,n8997,n9125);
and (n8997,n8998,n9023);
xor (n8998,n8999,n9000);
xor (n8999,n8922,n8928);
or (n9000,n9001,n9022);
and (n9001,n9002,n9009);
xor (n9002,n9003,n9008);
or (n9003,n9004,n9007);
and (n9004,n9005,n2036);
xor (n9005,n1232,n9006);
xor (n9006,n8932,n8954);
and (n9007,n1232,n9006);
xor (n9008,n8929,n1091);
or (n9009,n9010,n9021);
and (n9010,n9011,n1148);
xor (n9011,n2034,n9012);
or (n9012,n9013,n9020);
and (n9013,n9014,n1239);
xor (n9014,n9015,n9017);
xor (n9015,n9016,n1668);
xor (n9016,n8934,n8948);
and (n9017,n9018,n2439);
xor (n9018,n9019,n1676);
xor (n9019,n8936,n8946);
and (n9020,n9015,n9017);
and (n9021,n2034,n9012);
and (n9022,n9003,n9008);
or (n9023,n9024,n9124);
and (n9024,n9025,n9111);
xor (n9025,n9026,n9110);
or (n9026,n9027,n9109);
and (n9027,n9028,n1152);
xor (n9028,n9029,n9085);
or (n9029,n9030,n9084);
and (n9030,n9031,n1240);
xor (n9031,n9032,n9052);
xor (n9032,n9033,n2358);
xor (n9033,n1587,n9034);
or (n9034,n9035,n9051);
and (n9035,n9036,n1677);
xor (n9036,n9037,n9049);
or (n9037,n9038,n9039);
and (n9038,n1540,n1027);
and (n9039,n9040,n1027);
nand (n9040,n9041,n9042);
not (n9041,n2221);
nand (n9042,n9043,n9047);
or (n9043,n9044,n9045);
not (n9044,n8943);
not (n9045,n9046);
not (n9046,n2234);
not (n9047,n9048);
not (n9048,n2312);
nor (n9049,n1026,n9050);
xor (n9050,n2302,n8942);
and (n9051,n9037,n9049);
and (n9052,n9053,n9083);
xor (n9053,n9054,n9081);
or (n9054,n9055,n9080);
and (n9055,n9056,n2445);
xor (n9056,n9057,n9065);
and (n9057,n9058,n9061);
xor (n9058,n9059,n1692);
and (n9059,n9060,n1027);
xnor (n9060,n9048,n2314);
and (n9061,n9062,n9063);
and (n9062,n2557,n9047);
nor (n9063,n9064,n1559);
not (n9064,n1801);
or (n9065,n9066,n9079);
and (n9066,n9067,n9078);
xor (n9067,n9068,n9077);
and (n9068,n9069,n1027);
not (n9069,n9070);
nor (n9070,n9071,n9072);
and (n9071,n9047,n2254);
and (n9072,n9073,n9076);
nand (n9073,n9074,n9075);
not (n9074,n2318);
not (n9075,n2238);
not (n9076,n8940);
and (n9077,n1552,n1027);
and (n9078,n1558,n1027);
and (n9079,n9068,n9077);
and (n9080,n9057,n9065);
and (n9081,n9082,n1600);
xor (n9082,n2372,n1684);
xor (n9083,n9018,n2439);
and (n9084,n9032,n9052);
or (n9085,n9086,n9108);
and (n9086,n9087,n2111);
xor (n9087,n9088,n9089);
xor (n9088,n8956,n2433);
or (n9089,n9090,n9107);
and (n9090,n9091,n2365);
xor (n9091,n1594,n9092);
or (n9092,n9093,n9106);
and (n9093,n9094,n1685);
xor (n9094,n9095,n9105);
and (n9095,n9096,n1027);
not (n9096,n9097);
nor (n9097,n9098,n9104);
and (n9098,n9099,n9102);
not (n9099,n9100);
xor (n9100,n8915,n9101);
not (n9101,n2306);
not (n9102,n9103);
not (n9103,n2206);
and (n9104,n9100,n9103);
and (n9105,n1546,n1027);
and (n9106,n9095,n9105);
and (n9107,n1594,n9092);
and (n9108,n9088,n9089);
and (n9109,n9029,n9085);
xor (n9110,n8925,n1224);
xor (n9111,n9112,n1144);
xor (n9112,n2030,n9113);
xor (n9113,n9114,n2421);
xor (n9114,n1493,n9115);
or (n9115,n9116,n9123);
and (n9116,n9117,n9120);
xor (n9117,n9118,n9119);
xor (n9118,n8899,n8908);
and (n9119,n1496,n1027);
or (n9120,n9121,n9122);
and (n9121,n8958,n8967);
and (n9122,n8959,n8960);
and (n9123,n9118,n9119);
and (n9124,n9026,n9110);
and (n9125,n8999,n9000);
and (n9126,n8875,n8971);
xor (n9127,n9128,n9149);
xor (n9128,n9129,n9136);
xor (n9129,n9130,n9133);
xor (n9130,n9131,n9132);
and (n9131,n8974,n2410);
and (n9132,n8919,n1638);
or (n9133,n9134,n9135);
and (n9134,n8878,n1209);
and (n9135,n1082,n2088);
and (n9136,n9137,n9144);
xor (n9137,n9138,n2019);
or (n9138,n9139,n9143);
and (n9139,n9140,n2022);
xor (n9140,n1488,n9141);
xor (n9141,n9142,n1644);
xor (n9142,n8976,n8979);
and (n9143,n1488,n9141);
and (n9144,n9145,n2337);
xor (n9145,n1215,n9146);
or (n9146,n9147,n9148);
and (n9147,n9114,n2421);
and (n9148,n1493,n9115);
or (n9149,n9150,n9151);
and (n9150,n8972,n8992);
and (n9151,n8973,n8982);
xor (n9152,n9153,n9165);
xor (n9153,n9154,n9157);
or (n9154,n9155,n9156);
and (n9155,n8876,n8920);
and (n9156,n8877,n8879);
xor (n9157,n9158,n9163);
xor (n9158,n9159,n9162);
or (n9159,n9160,n9161);
and (n9160,n8880,n2334);
and (n9161,n8881,n8918);
xor (n9162,n1479,n1077);
xor (n9163,n9164,n1079);
xor (n9164,n1818,n2155);
or (n9165,n9166,n9202);
and (n9166,n9167,n9178);
xor (n9167,n9168,n9177);
or (n9168,n9169,n9176);
and (n9169,n9170,n9175);
xor (n9170,n9171,n9174);
or (n9171,n9172,n9173);
and (n9172,n9112,n1144);
and (n9173,n2030,n9113);
xor (n9174,n9140,n2022);
xor (n9175,n8984,n1216);
and (n9176,n9171,n9174);
xor (n9177,n9137,n9144);
or (n9178,n9179,n9201);
and (n9179,n9180,n9200);
xor (n9180,n9181,n9182);
xor (n9181,n9145,n2337);
or (n9182,n9183,n9199);
and (n9183,n9184,n9194);
xor (n9184,n9185,n9186);
xor (n9185,n8987,n2344);
or (n9186,n9187,n9193);
and (n9187,n9188,n2351);
xor (n9188,n9189,n9192);
or (n9189,n9190,n9191);
and (n9190,n9033,n2358);
and (n9191,n1587,n9034);
xor (n9192,n9117,n9120);
and (n9193,n9189,n9192);
or (n9194,n9195,n9198);
and (n9195,n9196,n2105);
xor (n9196,n1231,n9197);
xor (n9197,n1659,n1581);
and (n9198,n1231,n9197);
and (n9199,n9185,n9186);
xor (n9200,n8994,n1086);
and (n9201,n9181,n9182);
and (n9202,n9168,n9177);
or (n9203,n9204,n9260);
and (n9204,n9205,n9259);
xor (n9205,n9206,n9258);
or (n9206,n9207,n9257);
and (n9207,n9208,n9211);
xor (n9208,n9209,n9210);
xor (n9209,n9180,n9200);
xor (n9210,n9170,n9175);
or (n9211,n9212,n9256);
and (n9212,n9213,n9246);
xor (n9213,n9214,n9245);
or (n9214,n9215,n9244);
and (n9215,n9216,n9219);
xor (n9216,n9217,n9218);
xor (n9217,n9196,n2105);
xor (n9218,n9188,n2351);
or (n9219,n9220,n9243);
and (n9220,n9221,n2042);
xor (n9221,n9222,n9225);
and (n9222,n9223,n2117);
xor (n9223,n1247,n9224);
xor (n9224,n9036,n1677);
or (n9225,n9226,n9242);
and (n9226,n9227,n1248);
xor (n9227,n9228,n9229);
xor (n9228,n9091,n2365);
or (n9229,n9230,n9241);
and (n9230,n9231,n9237);
xor (n9231,n9232,n9233);
xor (n9232,n9094,n1685);
nand (n9233,n9234,n9037);
or (n9234,n9235,n9236);
not (n9235,n9039);
not (n9236,n9038);
or (n9237,n9238,n9240);
and (n9238,n9239,n1606);
xor (n9239,n1693,n2451);
and (n9240,n1693,n2451);
and (n9241,n9232,n9233);
and (n9242,n9228,n9229);
and (n9243,n9222,n9225);
and (n9244,n9217,n9218);
xor (n9245,n9184,n9194);
or (n9246,n9247,n9255);
and (n9247,n9248,n9254);
xor (n9248,n9249,n9250);
xor (n9249,n9005,n2036);
or (n9250,n9251,n9253);
and (n9251,n9252,n1159);
xor (n9252,n1156,n2040);
and (n9253,n1156,n2040);
xor (n9254,n9011,n1148);
and (n9255,n9249,n9250);
and (n9256,n9214,n9245);
and (n9257,n9209,n9210);
xor (n9258,n9167,n9178);
xor (n9259,n8874,n8996);
and (n9260,n9206,n9258);
or (n9261,n9262,n9659);
and (n9262,n9263,n9334);
xor (n9263,n9264,n9265);
xor (n9264,n9205,n9259);
or (n9265,n9266,n9333);
and (n9266,n9267,n9332);
xor (n9267,n9268,n9331);
or (n9268,n9269,n9330);
and (n9269,n9270,n9329);
xor (n9270,n9271,n9272);
xor (n9271,n9002,n9009);
or (n9272,n9273,n9328);
and (n9273,n9274,n9305);
xor (n9274,n9275,n9276);
xor (n9275,n9028,n1152);
or (n9276,n9277,n9304);
and (n9277,n9278,n9281);
xor (n9278,n9279,n9280);
xor (n9279,n9014,n1239);
xor (n9280,n9087,n2111);
or (n9281,n9282,n9303);
and (n9282,n9283,n2046);
xor (n9283,n9284,n1163);
and (n9284,n9285,n9302);
and (n9285,n9286,n9291);
or (n9286,n9287,n9290);
and (n9287,n9288,n2386);
xor (n9288,n1701,n9289);
xor (n9289,n9062,n9063);
and (n9290,n1701,n9289);
and (n9291,n9292,n9301);
xor (n9292,n9293,n1271);
and (n9293,n9294,n1027);
nand (n9294,n9295,n9300);
or (n9295,n9075,n9296);
nand (n9296,n9297,n9299);
or (n9297,n9298,n8940);
not (n9298,n9074);
nand (n9299,n9298,n8940);
nand (n9300,n9296,n9075);
and (n9301,n1564,n1027);
xor (n9302,n9056,n2445);
and (n9303,n9284,n1163);
and (n9304,n9279,n9280);
or (n9305,n9306,n9327);
and (n9306,n9307,n9326);
xor (n9307,n9308,n9325);
or (n9308,n9309,n9324);
and (n9309,n9310,n1166);
xor (n9310,n9311,n9323);
or (n9311,n9312,n9322);
and (n9312,n9313,n1256);
xor (n9313,n9314,n9315);
xor (n9314,n9082,n1600);
or (n9315,n9316,n9321);
and (n9316,n9317,n2379);
xor (n9317,n9318,n9319);
xor (n9318,n9067,n9078);
and (n9319,n2457,n9320);
and (n9320,n2462,n2140);
and (n9321,n9318,n9319);
and (n9322,n9314,n9315);
xor (n9323,n9053,n9083);
and (n9324,n9311,n9323);
xor (n9325,n9031,n1240);
xor (n9326,n9252,n1159);
and (n9327,n9308,n9325);
and (n9328,n9275,n9276);
xor (n9329,n9025,n9111);
and (n9330,n9271,n9272);
xor (n9331,n8998,n9023);
xor (n9332,n9208,n9211);
and (n9333,n9268,n9331);
or (n9334,n9335,n9658);
and (n9335,n9336,n9427);
xor (n9336,n9337,n9338);
xor (n9337,n9267,n9332);
or (n9338,n9339,n9426);
and (n9339,n9340,n9425);
xor (n9340,n9341,n9342);
xor (n9341,n9213,n9246);
or (n9342,n9343,n9424);
and (n9343,n9344,n9423);
xor (n9344,n9345,n9346);
xor (n9345,n9216,n9219);
or (n9346,n9347,n9422);
and (n9347,n9348,n9364);
xor (n9348,n9349,n9363);
or (n9349,n9350,n9362);
and (n9350,n9351,n9353);
xor (n9351,n2048,n9352);
xor (n9352,n9223,n2117);
or (n9353,n9354,n9361);
and (n9354,n9355,n1170);
xor (n9355,n9356,n2123);
or (n9356,n9357,n9360);
and (n9357,n9358,n1264);
xor (n9358,n2129,n9359);
xor (n9359,n9058,n9061);
and (n9360,n2129,n9359);
and (n9361,n9356,n2123);
and (n9362,n2048,n9352);
xor (n9363,n9221,n2042);
or (n9364,n9365,n9421);
and (n9365,n9366,n9420);
xor (n9366,n9367,n9368);
xor (n9367,n9227,n1248);
or (n9368,n9369,n9419);
and (n9369,n9370,n2054);
xor (n9370,n2052,n9371);
or (n9371,n9372,n9418);
and (n9372,n9373,n9396);
xor (n9373,n9374,n9375);
xor (n9374,n9239,n1606);
or (n9375,n9376,n9395);
and (n9376,n9377,n1612);
xor (n9377,n9378,n9385);
or (n9378,n9379,n9384);
and (n9379,n9380,n9382);
xor (n9380,n9381,n2392);
xor (n9381,n2462,n2140);
and (n9382,n9383,n1027);
not (n9383,n1570);
and (n9384,n9381,n2392);
or (n9385,n9386,n9394);
and (n9386,n9387,n9390);
xor (n9387,n9388,n9389);
and (n9388,n1390,n1027);
and (n9389,n2254,n1027);
and (n9390,n9391,n1027);
xor (n9391,n9392,n9393);
not (n9392,n2266);
not (n9393,n2323);
and (n9394,n9388,n9389);
and (n9395,n9378,n9385);
or (n9396,n9397,n9417);
and (n9397,n9398,n2135);
xor (n9398,n9399,n9415);
or (n9399,n9400,n9414);
and (n9400,n9401,n1277);
xor (n9401,n9402,n9409);
or (n9402,n9403,n9408);
and (n9403,n9404,n9406);
xor (n9404,n9405,n2397);
nor (n9405,n1556,n1026);
nor (n9406,n9407,n1026);
not (n9407,n2281);
and (n9408,n9405,n2397);
and (n9409,n9410,n9412);
nor (n9410,n9411,n1026);
not (n9411,n1406);
nor (n9412,n9413,n1026);
not (n9413,n2269);
and (n9414,n9402,n9409);
xor (n9415,n9416,n1700);
xor (n9416,n2457,n9320);
and (n9417,n9399,n9415);
and (n9418,n9374,n9375);
and (n9419,n2052,n9371);
xor (n9420,n9283,n2046);
and (n9421,n9367,n9368);
and (n9422,n9349,n9363);
xor (n9423,n9248,n9254);
and (n9424,n9345,n9346);
xor (n9425,n9270,n9329);
and (n9426,n9341,n9342);
or (n9427,n9428,n9657);
and (n9428,n9429,n9481);
xor (n9429,n9430,n9480);
or (n9430,n9431,n9479);
and (n9431,n9432,n9478);
xor (n9432,n9433,n9477);
or (n9433,n9434,n9476);
and (n9434,n9435,n9475);
xor (n9435,n9436,n9474);
or (n9436,n9437,n9473);
and (n9437,n9438,n9472);
xor (n9438,n9439,n9466);
or (n9439,n9440,n9465);
and (n9440,n9441,n9460);
xor (n9441,n9442,n9444);
xor (n9442,n9443,n1255);
xor (n9443,n9285,n9302);
or (n9444,n9445,n9459);
and (n9445,n9446,n1177);
xor (n9446,n9447,n9457);
or (n9447,n9448,n9456);
and (n9448,n9449,n9455);
xor (n9449,n1272,n9450);
or (n9450,n9451,n9454);
and (n9451,n9452,n1706);
xor (n9452,n9453,n1618);
xor (n9453,n9387,n9390);
and (n9454,n9453,n1618);
xor (n9455,n9288,n2386);
and (n9456,n1272,n9450);
xor (n9457,n9458,n1263);
xor (n9458,n9286,n9291);
and (n9459,n9447,n9457);
or (n9460,n9461,n9464);
and (n9461,n9462,n1179);
xor (n9462,n2058,n9463);
xor (n9463,n9317,n2379);
and (n9464,n2058,n9463);
and (n9465,n9442,n9444);
or (n9466,n9467,n9471);
and (n9467,n9468,n1173);
xor (n9468,n9469,n9470);
xor (n9469,n9231,n9237);
xor (n9470,n9313,n1256);
and (n9471,n9469,n9470);
xor (n9472,n9310,n1166);
and (n9473,n9439,n9466);
xor (n9474,n9278,n9281);
xor (n9475,n9307,n9326);
and (n9476,n9436,n9474);
xor (n9477,n9274,n9305);
xor (n9478,n9344,n9423);
and (n9479,n9433,n9477);
xor (n9480,n9340,n9425);
or (n9481,n9482,n9656);
and (n9482,n9483,n9548);
xor (n9483,n9484,n9547);
or (n9484,n9485,n9546);
and (n9485,n9486,n9545);
xor (n9486,n9487,n9488);
xor (n9487,n9348,n9364);
or (n9488,n9489,n9544);
and (n9489,n9490,n9543);
xor (n9490,n9491,n9492);
xor (n9491,n9351,n9353);
or (n9492,n9493,n9542);
and (n9493,n9494,n9506);
xor (n9494,n9495,n9496);
xor (n9495,n9355,n1170);
or (n9496,n9497,n9505);
and (n9497,n9498,n2060);
xor (n9498,n9499,n9500);
xor (n9499,n9358,n1264);
or (n9500,n9501,n9504);
and (n9501,n9502,n1183);
xor (n9502,n2064,n9503);
xor (n9503,n9292,n9301);
and (n9504,n2064,n9503);
and (n9505,n9499,n9500);
or (n9506,n9507,n9541);
and (n9507,n9508,n9526);
xor (n9508,n9509,n9510);
xor (n9509,n9373,n9396);
or (n9510,n9511,n9525);
and (n9511,n9512,n2066);
xor (n9512,n9513,n9524);
or (n9513,n9514,n9523);
and (n9514,n9515,n1189);
xor (n9515,n9516,n9517);
xor (n9516,n9380,n9382);
or (n9517,n9518,n9522);
and (n9518,n9519,n9521);
xor (n9519,n9520,n2075);
and (n9520,n1801,n2556);
xor (n9521,n9410,n9412);
and (n9522,n9520,n2075);
and (n9523,n9516,n9517);
xor (n9524,n9377,n1612);
and (n9525,n9513,n9524);
or (n9526,n9527,n9540);
and (n9527,n9528,n1185);
xor (n9528,n9529,n9530);
xor (n9529,n9398,n2135);
or (n9530,n9531,n9539);
and (n9531,n9532,n2070);
xor (n9532,n9533,n9534);
xor (n9533,n9452,n1706);
or (n9534,n9535,n9538);
and (n9535,n9536,n1623);
xor (n9536,n1194,n9537);
xor (n9537,n9404,n9406);
and (n9538,n1194,n9537);
and (n9539,n9533,n9534);
and (n9540,n9529,n9530);
and (n9541,n9509,n9510);
and (n9542,n9495,n9496);
xor (n9543,n9366,n9420);
and (n9544,n9491,n9492);
xor (n9545,n9435,n9475);
and (n9546,n9487,n9488);
xor (n9547,n9432,n9478);
nand (n9548,n9549,n9655);
or (n9549,n9550,n9565);
nor (n9550,n9551,n9552);
xor (n9551,n9486,n9545);
or (n9552,n9553,n9564);
and (n9553,n9554,n9563);
xor (n9554,n9555,n9556);
xor (n9555,n9438,n9472);
or (n9556,n9557,n9562);
and (n9557,n9558,n9561);
xor (n9558,n9559,n9560);
xor (n9559,n9370,n2054);
xor (n9560,n9468,n1173);
xor (n9561,n9441,n9460);
and (n9562,n9559,n9560);
xor (n9563,n9490,n9543);
and (n9564,n9555,n9556);
and (n9565,n9566,n9654);
nand (n9566,n9567,n9582);
or (n9567,n9568,n9569);
xor (n9568,n9554,n9563);
or (n9569,n9570,n9581);
and (n9570,n9571,n9580);
xor (n9571,n9572,n9579);
or (n9572,n9573,n9578);
and (n9573,n9574,n9577);
xor (n9574,n9575,n9576);
xor (n9575,n9462,n1179);
xor (n9576,n9446,n1177);
xor (n9577,n9498,n2060);
and (n9578,n9575,n9576);
xor (n9579,n9494,n9506);
xor (n9580,n9558,n9561);
and (n9581,n9572,n9579);
nand (n9582,n9583,n9647);
nand (n9583,n9584,n9619,n9622);
or (n9584,n9585,n9618);
or (n9585,n9586,n9617);
and (n9586,n9587,n9616);
xor (n9587,n9588,n9605);
or (n9588,n9589,n9604);
and (n9589,n9590,n9603);
xor (n9590,n9591,n9592);
xor (n9591,n9512,n2066);
or (n9592,n9593,n9602);
and (n9593,n9594,n9601);
xor (n9594,n9595,n9596);
xor (n9595,n9515,n1189);
or (n9596,n9597,n9600);
and (n9597,n9598,n2077);
xor (n9598,n9599,n1196);
xor (n9599,n9519,n9521);
and (n9600,n9599,n1196);
xor (n9601,n9532,n2070);
and (n9602,n9595,n9596);
xor (n9603,n9528,n1185);
and (n9604,n9591,n9592);
or (n9605,n9606,n9615);
and (n9606,n9607,n9614);
xor (n9607,n9608,n9613);
or (n9608,n9609,n9612);
and (n9609,n9610,n1191);
xor (n9610,n2072,n9611);
xor (n9611,n9401,n1277);
and (n9612,n2072,n9611);
xor (n9613,n9449,n9455);
xor (n9614,n9502,n1183);
and (n9615,n9608,n9613);
xor (n9616,n9508,n9526);
and (n9617,n9588,n9605);
xor (n9618,n9571,n9580);
or (n9619,n9620,n9621);
xor (n9620,n9587,n9616);
xor (n9621,n9574,n9577);
nand (n9622,n9623,n9643);
or (n9623,n9624,n9627);
nor (n9624,n9625,n9626);
xor (n9625,n9590,n9603);
xor (n9626,n9607,n9614);
nand (n9627,n9628,n9631,n9634);
or (n9628,n9629,n9630);
xor (n9629,n9610,n1191);
xor (n9630,n9594,n9601);
or (n9631,n9632,n9633);
xor (n9632,n9536,n1623);
xor (n9633,n9598,n2077);
nand (n9634,n9635,n9638);
or (n9635,n9636,n9637);
not (n9636,n9632);
not (n9637,n9633);
nor (n9638,n9639,n9642);
and (n9639,n9640,n9641);
xor (n9640,n1801,n2556);
or (n9641,n1800,n2557);
and (n9642,n1800,n2557);
nor (n9643,n9644,n9646);
and (n9644,n9645,n9629,n9630);
not (n9645,n9624);
and (n9646,n9625,n9626);
nor (n9647,n9648,n9652);
and (n9648,n9618,n9649);
nand (n9649,n9650,n9651);
not (n9650,n9585);
nand (n9651,n9620,n9621);
and (n9652,n9653,n9585);
not (n9653,n9651);
nand (n9654,n9568,n9569);
nand (n9655,n9551,n9552);
and (n9656,n9484,n9547);
and (n9657,n9430,n9480);
and (n9658,n9337,n9338);
and (n9659,n9264,n9265);
and (n9660,n8870,n9203);
not (n9661,n9662);
or (n9662,n9663,n9666);
or (n9663,n9664,n9665);
and (n9664,n8871,n9152);
and (n9665,n8872,n9127);
nand (n9666,n9667,n9671);
not (n9667,n9668);
or (n9668,n9669,n9670);
and (n9669,n9153,n9165);
and (n9670,n9154,n9157);
nor (n9671,n9672,n9685);
not (n9672,n9673);
nor (n9673,n9674,n9682);
not (n9674,n9675);
nor (n9675,n9676,n9677);
and (n9676,n9164,n1079);
not (n9677,n9678);
nor (n9678,n9679,n9680);
and (n9679,n1479,n1077);
not (n9680,n9681);
xnor (n9681,n8,n1291);
or (n9682,n9683,n9684);
and (n9683,n9158,n9163);
and (n9684,n9159,n9162);
and (n9685,n9128,n9149);
nor (n9686,n9687,n2697);
not (n9687,n9688);
and (n9688,n33,n2696);
endmodule
