module top (out,n13,n14,n16,n17,n20,n21,n25,n26,n28
        ,n29,n43,n48,n103,n131,n184,n294,n296,n299,n303
        ,n305,n322,n401,n453);
output out;
input n13;
input n14;
input n16;
input n17;
input n20;
input n21;
input n25;
input n26;
input n28;
input n29;
input n43;
input n48;
input n103;
input n131;
input n184;
input n294;
input n296;
input n299;
input n303;
input n305;
input n322;
input n401;
input n453;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n15;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n295;
wire n297;
wire n298;
wire n300;
wire n301;
wire n302;
wire n304;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
xor (out,n0,n613);
xor (n0,n1,n552);
xor (n1,n2,n283);
xor (n2,n3,n120);
xor (n3,n4,n80);
xor (n4,n5,n63);
xor (n5,n6,n60);
or (n6,n7,n50,n59);
and (n7,n8,n37);
or (n8,n9,n30,n36);
and (n9,n10,n23);
or (n10,n11,n18,n22);
and (n11,n12,n15);
and (n12,n13,n14);
and (n15,n16,n17);
and (n18,n15,n19);
and (n19,n20,n21);
and (n22,n12,n19);
and (n23,n24,n27);
and (n24,n25,n26);
and (n27,n28,n29);
and (n30,n23,n31);
xor (n31,n32,n35);
xor (n32,n33,n34);
and (n33,n13,n29);
and (n34,n16,n14);
and (n35,n20,n17);
and (n36,n10,n31);
xor (n37,n38,n45);
xor (n38,n39,n44);
nor (n39,n40,n41);
not (n40,n28);
and (n41,n42,n28);
not (n42,n43);
and (n44,n13,n26);
nor (n45,n46,n49);
and (n46,n47,n17);
not (n47,n48);
not (n49,n17);
and (n50,n37,n51);
xor (n51,n52,n58);
xor (n52,n53,n57);
or (n53,n54,n55,n56);
and (n54,n33,n34);
and (n55,n34,n35);
and (n56,n33,n35);
and (n57,n16,n29);
and (n58,n20,n14);
and (n59,n8,n51);
nor (n60,n61,n62);
and (n61,n47,n14);
not (n62,n14);
xor (n63,n64,n73);
xor (n64,n65,n69);
or (n65,n66,n67,n68);
and (n66,n39,n44);
and (n67,n44,n45);
and (n68,n39,n45);
or (n69,n70,n71,n72);
and (n70,n53,n57);
and (n71,n57,n58);
and (n72,n53,n58);
xor (n73,n74,n79);
xor (n74,n75,n78);
nor (n75,n76,n77);
not (n76,n13);
and (n77,n42,n13);
and (n78,n16,n26);
and (n79,n20,n29);
or (n80,n81,n116,n119);
and (n81,n82,n93);
or (n82,n83,n88,n92);
and (n83,n84,n87);
nor (n84,n85,n86);
not (n85,n25);
and (n86,n42,n25);
and (n87,n28,n26);
and (n88,n87,n89);
nor (n89,n90,n91);
and (n90,n47,n21);
not (n91,n21);
and (n92,n84,n89);
or (n93,n94,n112,n115);
and (n94,n95,n110);
or (n95,n96,n107,n109);
and (n96,n97,n105);
or (n97,n98,n101,n104);
and (n98,n99,n100);
and (n99,n13,n17);
and (n100,n16,n21);
and (n101,n100,n102);
and (n102,n20,n103);
and (n104,n99,n102);
xor (n105,n106,n19);
xor (n106,n12,n15);
and (n107,n105,n108);
xor (n108,n24,n27);
and (n109,n97,n108);
xor (n110,n111,n89);
xor (n111,n84,n87);
and (n112,n110,n113);
xor (n113,n114,n31);
xor (n114,n10,n23);
and (n115,n95,n113);
and (n116,n93,n117);
xor (n117,n118,n51);
xor (n118,n8,n37);
and (n119,n82,n117);
or (n120,n121,n167);
and (n121,n122,n124);
xor (n122,n123,n117);
xor (n123,n82,n93);
or (n124,n125,n163,n166);
and (n125,n126,n144);
or (n126,n127,n139,n143);
and (n127,n128,n136);
or (n128,n129,n133,n135);
and (n129,n130,n132);
and (n130,n131,n26);
and (n132,n25,n29);
and (n133,n132,n134);
and (n134,n28,n14);
and (n135,n130,n134);
nor (n136,n137,n138);
not (n137,n131);
and (n138,n42,n131);
and (n139,n136,n140);
nor (n140,n141,n142);
and (n141,n47,n103);
not (n142,n103);
and (n143,n128,n140);
or (n144,n145,n159,n162);
and (n145,n146,n157);
or (n146,n147,n153,n156);
and (n147,n148,n151);
and (n148,n149,n150);
and (n149,n13,n21);
and (n150,n16,n103);
xor (n151,n152,n134);
xor (n152,n130,n132);
and (n153,n151,n154);
xor (n154,n155,n102);
xor (n155,n99,n100);
and (n156,n148,n154);
xor (n157,n158,n140);
xor (n158,n128,n136);
and (n159,n157,n160);
xor (n160,n161,n108);
xor (n161,n97,n105);
and (n162,n146,n160);
and (n163,n144,n164);
xor (n164,n165,n113);
xor (n165,n95,n110);
and (n166,n126,n164);
and (n167,n168,n169);
xor (n168,n122,n124);
or (n169,n170,n189);
and (n170,n171,n173);
xor (n171,n172,n164);
xor (n172,n126,n144);
and (n173,n174,n187);
or (n174,n175,n181,n186);
and (n175,n176,n179);
and (n176,n177,n178);
and (n177,n28,n17);
xor (n178,n149,n150);
xor (n179,n180,n154);
xor (n180,n148,n151);
and (n181,n179,n182);
nor (n182,n183,n185);
not (n183,n184);
and (n185,n42,n184);
and (n186,n176,n182);
xor (n187,n188,n160);
xor (n188,n146,n157);
and (n189,n190,n191);
xor (n190,n171,n173);
or (n191,n192,n222);
and (n192,n193,n194);
xor (n193,n174,n187);
or (n194,n195,n218,n221);
and (n195,n196,n203);
or (n196,n197,n200,n202);
and (n197,n198,n199);
and (n198,n184,n26);
and (n199,n131,n29);
and (n200,n199,n201);
and (n201,n25,n14);
and (n202,n198,n201);
or (n203,n204,n215,n217);
and (n204,n205,n213);
or (n205,n206,n209,n212);
and (n206,n207,n208);
and (n207,n25,n21);
and (n208,n28,n103);
and (n209,n210,n211);
and (n210,n28,n21);
and (n211,n13,n103);
and (n212,n206,n211);
xor (n213,n214,n201);
xor (n214,n198,n199);
and (n215,n213,n216);
xor (n216,n177,n178);
and (n217,n205,n216);
and (n218,n203,n219);
xor (n219,n220,n182);
xor (n220,n176,n179);
and (n221,n196,n219);
and (n222,n223,n224);
xor (n223,n193,n194);
or (n224,n225,n253);
and (n225,n226,n228);
xor (n226,n227,n219);
xor (n227,n196,n203);
or (n228,n229,n249,n252);
and (n229,n230,n233);
and (n230,n231,n232);
and (n231,n131,n14);
and (n232,n25,n17);
or (n233,n234,n245,n248);
and (n234,n235,n244);
or (n235,n236,n241,n243);
and (n236,n237,n240);
and (n237,n238,n239);
and (n238,n131,n21);
and (n239,n25,n103);
and (n240,n131,n17);
and (n241,n240,n242);
xor (n242,n207,n208);
and (n243,n237,n242);
xor (n244,n231,n232);
and (n245,n244,n246);
xor (n246,n247,n211);
xor (n247,n206,n210);
and (n248,n235,n246);
and (n249,n233,n250);
xor (n250,n251,n216);
xor (n251,n205,n213);
and (n252,n230,n250);
and (n253,n254,n255);
xor (n254,n226,n228);
or (n255,n256,n278);
and (n256,n257,n259);
xor (n257,n258,n250);
xor (n258,n230,n233);
and (n259,n260,n276);
or (n260,n261,n272,n275);
and (n261,n262,n271);
or (n262,n263,n268,n270);
and (n263,n264,n267);
and (n264,n265,n266);
and (n265,n184,n21);
and (n266,n131,n103);
and (n267,n184,n17);
and (n268,n267,n269);
xor (n269,n238,n239);
and (n270,n264,n269);
and (n271,n184,n14);
and (n272,n271,n273);
xor (n273,n274,n242);
xor (n274,n237,n240);
and (n275,n262,n273);
xor (n276,n277,n246);
xor (n277,n235,n244);
and (n278,n279,n280);
xor (n279,n257,n259);
and (n280,n281,n282);
and (n281,n184,n29);
xor (n282,n260,n276);
xor (n283,n284,n390);
xor (n284,n285,n352);
xor (n285,n286,n335);
xor (n286,n287,n333);
or (n287,n288,n323,n332);
and (n288,n289,n313);
or (n289,n290,n306,n312);
and (n290,n291,n301);
or (n291,n292,n297,n300);
and (n292,n293,n295);
and (n293,n294,n14);
and (n295,n296,n17);
and (n297,n295,n298);
and (n298,n299,n21);
and (n300,n293,n298);
and (n301,n302,n304);
and (n302,n303,n26);
and (n304,n305,n29);
and (n306,n301,n307);
xor (n307,n308,n311);
xor (n308,n309,n310);
and (n309,n294,n29);
and (n310,n296,n14);
and (n311,n299,n17);
and (n312,n291,n307);
xor (n313,n314,n319);
xor (n314,n315,n318);
nor (n315,n316,n317);
not (n316,n305);
and (n317,n42,n305);
and (n318,n294,n26);
nor (n319,n320,n49);
and (n320,n321,n17);
not (n321,n322);
and (n323,n313,n324);
xor (n324,n325,n331);
xor (n325,n326,n330);
or (n326,n327,n328,n329);
and (n327,n309,n310);
and (n328,n310,n311);
and (n329,n309,n311);
and (n330,n296,n29);
and (n331,n299,n14);
and (n332,n289,n324);
nor (n333,n334,n62);
and (n334,n321,n14);
xor (n335,n336,n345);
xor (n336,n337,n341);
or (n337,n338,n339,n340);
and (n338,n315,n318);
and (n339,n318,n319);
and (n340,n315,n319);
or (n341,n342,n343,n344);
and (n342,n326,n330);
and (n343,n330,n331);
and (n344,n326,n331);
xor (n345,n346,n351);
xor (n346,n347,n350);
nor (n347,n348,n349);
not (n348,n294);
and (n349,n42,n294);
and (n350,n296,n26);
and (n351,n299,n29);
or (n352,n353,n386,n389);
and (n353,n354,n364);
or (n354,n355,n360,n363);
and (n355,n356,n359);
nor (n356,n357,n358);
not (n357,n303);
and (n358,n42,n303);
and (n359,n305,n26);
and (n360,n359,n361);
nor (n361,n362,n91);
and (n362,n321,n21);
and (n363,n356,n361);
or (n364,n365,n382,n385);
and (n365,n366,n380);
or (n366,n367,n377,n379);
and (n367,n368,n375);
or (n368,n369,n372,n374);
and (n369,n370,n371);
and (n370,n294,n17);
and (n371,n296,n21);
and (n372,n371,n373);
and (n373,n299,n103);
and (n374,n370,n373);
xor (n375,n376,n298);
xor (n376,n293,n295);
and (n377,n375,n378);
xor (n378,n302,n304);
and (n379,n368,n378);
xor (n380,n381,n361);
xor (n381,n356,n359);
and (n382,n380,n383);
xor (n383,n384,n307);
xor (n384,n291,n301);
and (n385,n366,n383);
and (n386,n364,n387);
xor (n387,n388,n324);
xor (n388,n289,n313);
and (n389,n354,n387);
or (n390,n391,n436);
and (n391,n392,n394);
xor (n392,n393,n387);
xor (n393,n354,n364);
or (n394,n395,n432,n435);
and (n395,n396,n413);
or (n396,n397,n409,n412);
and (n397,n398,n406);
or (n398,n399,n403,n405);
and (n399,n400,n402);
and (n400,n401,n26);
and (n402,n303,n29);
and (n403,n402,n404);
and (n404,n305,n14);
and (n405,n400,n404);
nor (n406,n407,n408);
not (n407,n401);
and (n408,n42,n401);
and (n409,n406,n410);
nor (n410,n411,n142);
and (n411,n321,n103);
and (n412,n398,n410);
or (n413,n414,n428,n431);
and (n414,n415,n426);
or (n415,n416,n422,n425);
and (n416,n417,n420);
and (n417,n418,n419);
and (n418,n294,n21);
and (n419,n296,n103);
xor (n420,n421,n404);
xor (n421,n400,n402);
and (n422,n420,n423);
xor (n423,n424,n373);
xor (n424,n370,n371);
and (n425,n417,n423);
xor (n426,n427,n410);
xor (n427,n398,n406);
and (n428,n426,n429);
xor (n429,n430,n378);
xor (n430,n368,n375);
and (n431,n415,n429);
and (n432,n413,n433);
xor (n433,n434,n383);
xor (n434,n366,n380);
and (n435,n396,n433);
and (n436,n437,n438);
xor (n437,n392,n394);
or (n438,n439,n458);
and (n439,n440,n442);
xor (n440,n441,n433);
xor (n441,n396,n413);
and (n442,n443,n456);
or (n443,n444,n450,n455);
and (n444,n445,n448);
and (n445,n446,n447);
and (n446,n305,n17);
xor (n447,n418,n419);
xor (n448,n449,n423);
xor (n449,n417,n420);
and (n450,n448,n451);
nor (n451,n452,n454);
not (n452,n453);
and (n454,n42,n453);
and (n455,n445,n451);
xor (n456,n457,n429);
xor (n457,n415,n426);
and (n458,n459,n460);
xor (n459,n440,n442);
or (n460,n461,n491);
and (n461,n462,n463);
xor (n462,n443,n456);
or (n463,n464,n487,n490);
and (n464,n465,n472);
or (n465,n466,n469,n471);
and (n466,n467,n468);
and (n467,n453,n26);
and (n468,n401,n29);
and (n469,n468,n470);
and (n470,n303,n14);
and (n471,n467,n470);
or (n472,n473,n484,n486);
and (n473,n474,n482);
or (n474,n475,n478,n481);
and (n475,n476,n477);
and (n476,n303,n21);
and (n477,n305,n103);
and (n478,n479,n480);
and (n479,n305,n21);
and (n480,n294,n103);
and (n481,n475,n480);
xor (n482,n483,n470);
xor (n483,n467,n468);
and (n484,n482,n485);
xor (n485,n446,n447);
and (n486,n474,n485);
and (n487,n472,n488);
xor (n488,n489,n451);
xor (n489,n445,n448);
and (n490,n465,n488);
and (n491,n492,n493);
xor (n492,n462,n463);
or (n493,n494,n522);
and (n494,n495,n497);
xor (n495,n496,n488);
xor (n496,n465,n472);
or (n497,n498,n518,n521);
and (n498,n499,n502);
and (n499,n500,n501);
and (n500,n401,n14);
and (n501,n303,n17);
or (n502,n503,n514,n517);
and (n503,n504,n513);
or (n504,n505,n510,n512);
and (n505,n506,n509);
and (n506,n507,n508);
and (n507,n401,n21);
and (n508,n303,n103);
and (n509,n401,n17);
and (n510,n509,n511);
xor (n511,n476,n477);
and (n512,n506,n511);
xor (n513,n500,n501);
and (n514,n513,n515);
xor (n515,n516,n480);
xor (n516,n475,n479);
and (n517,n504,n515);
and (n518,n502,n519);
xor (n519,n520,n485);
xor (n520,n474,n482);
and (n521,n499,n519);
and (n522,n523,n524);
xor (n523,n495,n497);
or (n524,n525,n547);
and (n525,n526,n528);
xor (n526,n527,n519);
xor (n527,n499,n502);
and (n528,n529,n545);
or (n529,n530,n541,n544);
and (n530,n531,n540);
or (n531,n532,n537,n539);
and (n532,n533,n536);
and (n533,n534,n535);
and (n534,n453,n21);
and (n535,n401,n103);
and (n536,n453,n17);
and (n537,n536,n538);
xor (n538,n507,n508);
and (n539,n533,n538);
and (n540,n453,n14);
and (n541,n540,n542);
xor (n542,n543,n511);
xor (n543,n506,n509);
and (n544,n531,n542);
xor (n545,n546,n515);
xor (n546,n504,n513);
and (n547,n548,n549);
xor (n548,n526,n528);
and (n549,n550,n551);
and (n550,n453,n29);
xor (n551,n529,n545);
or (n552,n553,n556,n612);
and (n553,n554,n555);
xor (n554,n168,n169);
xor (n555,n437,n438);
and (n556,n555,n557);
or (n557,n558,n561,n611);
and (n558,n559,n560);
xor (n559,n190,n191);
xor (n560,n459,n460);
and (n561,n560,n562);
or (n562,n563,n566,n610);
and (n563,n564,n565);
xor (n564,n223,n224);
xor (n565,n492,n493);
and (n566,n565,n567);
or (n567,n568,n571,n609);
and (n568,n569,n570);
xor (n569,n254,n255);
xor (n570,n523,n524);
and (n571,n570,n572);
or (n572,n573,n576,n608);
and (n573,n574,n575);
xor (n574,n279,n280);
xor (n575,n548,n549);
and (n576,n575,n577);
or (n577,n578,n581,n607);
and (n578,n579,n580);
xor (n579,n281,n282);
xor (n580,n550,n551);
and (n581,n580,n582);
or (n582,n583,n588,n606);
and (n583,n584,n586);
xor (n584,n585,n273);
xor (n585,n262,n271);
xor (n586,n587,n542);
xor (n587,n531,n540);
and (n588,n586,n589);
or (n589,n590,n595,n605);
and (n590,n591,n593);
xor (n591,n592,n269);
xor (n592,n264,n267);
xor (n593,n594,n538);
xor (n594,n533,n536);
and (n595,n593,n596);
or (n596,n597,n600,n604);
and (n597,n598,n599);
xor (n598,n265,n266);
xor (n599,n534,n535);
and (n600,n599,n601);
and (n601,n602,n603);
and (n602,n184,n103);
and (n603,n453,n103);
and (n604,n598,n601);
and (n605,n591,n596);
and (n606,n584,n589);
and (n607,n579,n582);
and (n608,n574,n577);
and (n609,n569,n572);
and (n610,n564,n567);
and (n611,n559,n562);
and (n612,n554,n557);
xor (n613,n614,n771);
xor (n614,n615,n735);
xor (n615,n616,n713);
xor (n616,n617,n661);
or (n617,n618,n640,n660);
and (n618,n619,n633);
nor (n619,n620,n632);
not (n620,n621);
xor (n621,n622,n623);
xor (n622,n28,n305);
or (n623,n624,n625,n631);
and (n624,n25,n303);
and (n625,n303,n626);
or (n626,n627,n628,n630);
and (n627,n131,n401);
and (n628,n401,n629);
and (n629,n184,n453);
and (n630,n131,n629);
and (n631,n25,n626);
and (n632,n42,n621);
and (n633,n634,n26);
xor (n634,n635,n636);
xor (n635,n13,n294);
or (n636,n637,n638,n639);
and (n637,n28,n305);
and (n638,n305,n623);
and (n639,n28,n623);
and (n640,n633,n641);
nor (n641,n642,n91);
and (n642,n643,n21);
not (n643,n644);
or (n644,n645,n646,n659);
and (n645,n48,n322);
and (n646,n322,n647);
or (n647,n648,n649,n658);
and (n648,n20,n299);
and (n649,n299,n650);
or (n650,n651,n652,n657);
and (n651,n16,n296);
and (n652,n296,n653);
or (n653,n654,n655,n656);
and (n654,n13,n294);
and (n655,n294,n636);
and (n656,n13,n636);
and (n657,n16,n653);
and (n658,n20,n650);
and (n659,n48,n647);
and (n660,n619,n641);
or (n661,n662,n696,n712);
and (n662,n663,n694);
or (n663,n664,n683,n693);
and (n664,n665,n678);
or (n665,n666,n673,n677);
and (n666,n667,n670);
and (n667,n668,n17);
xor (n668,n669,n653);
xor (n669,n16,n296);
and (n670,n671,n21);
xor (n671,n672,n650);
xor (n672,n20,n299);
and (n673,n670,n674);
and (n674,n675,n103);
xor (n675,n676,n647);
xor (n676,n48,n322);
and (n677,n667,n674);
xor (n678,n679,n682);
xor (n679,n680,n681);
and (n680,n668,n14);
and (n681,n671,n17);
and (n682,n675,n21);
and (n683,n678,n684);
xor (n684,n685,n692);
xor (n685,n686,n691);
nor (n686,n687,n690);
not (n687,n688);
xor (n688,n689,n626);
xor (n689,n25,n303);
and (n690,n42,n688);
and (n691,n621,n26);
and (n692,n634,n29);
and (n693,n665,n684);
xor (n694,n695,n641);
xor (n695,n619,n633);
and (n696,n694,n697);
xor (n697,n698,n707);
xor (n698,n699,n703);
or (n699,n700,n701,n702);
and (n700,n680,n681);
and (n701,n681,n682);
and (n702,n680,n682);
or (n703,n704,n705,n706);
and (n704,n686,n691);
and (n705,n691,n692);
and (n706,n686,n692);
xor (n707,n708,n711);
xor (n708,n709,n710);
and (n709,n668,n29);
and (n710,n671,n14);
and (n711,n675,n17);
and (n712,n663,n697);
xor (n713,n714,n727);
xor (n714,n715,n719);
or (n715,n716,n717,n718);
and (n716,n699,n703);
and (n717,n703,n707);
and (n718,n699,n707);
xor (n719,n720,n725);
xor (n720,n721,n724);
nor (n721,n722,n723);
not (n722,n634);
and (n723,n42,n634);
and (n724,n668,n26);
nor (n725,n726,n49);
and (n726,n643,n17);
xor (n727,n728,n734);
xor (n728,n729,n733);
or (n729,n730,n731,n732);
and (n730,n709,n710);
and (n731,n710,n711);
and (n732,n709,n711);
and (n733,n671,n29);
and (n734,n675,n14);
or (n735,n736,n767,n770);
and (n736,n737,n747);
and (n737,n738,n745);
or (n738,n739,n742,n744);
and (n739,n740,n741);
and (n740,n688,n26);
and (n741,n621,n29);
and (n742,n741,n743);
and (n743,n634,n14);
and (n744,n740,n743);
nor (n745,n746,n142);
and (n746,n643,n103);
or (n747,n748,n764,n766);
and (n748,n749,n762);
or (n749,n750,n758,n761);
and (n750,n751,n756);
nor (n751,n752,n755);
not (n752,n753);
xor (n753,n754,n629);
xor (n754,n131,n401);
and (n755,n42,n753);
xor (n756,n757,n674);
xor (n757,n667,n670);
and (n758,n756,n759);
xor (n759,n760,n743);
xor (n760,n740,n741);
and (n761,n751,n759);
xor (n762,n763,n684);
xor (n763,n665,n678);
and (n764,n762,n765);
xor (n765,n738,n745);
and (n766,n749,n765);
and (n767,n747,n768);
xor (n768,n769,n697);
xor (n769,n663,n694);
and (n770,n737,n768);
or (n771,n772,n809);
and (n772,n773,n775);
xor (n773,n774,n768);
xor (n774,n737,n747);
or (n775,n776,n805,n808);
and (n776,n777,n788);
and (n777,n778,n785);
or (n778,n779,n782,n784);
and (n779,n780,n781);
and (n780,n688,n29);
and (n781,n621,n14);
and (n782,n781,n783);
and (n783,n634,n17);
and (n784,n780,n783);
and (n785,n786,n787);
and (n786,n668,n21);
and (n787,n671,n103);
or (n788,n789,n801,n804);
and (n789,n790,n800);
or (n790,n791,n797,n799);
and (n791,n792,n795);
and (n792,n793,n794);
and (n793,n634,n21);
and (n794,n668,n103);
xor (n795,n796,n783);
xor (n796,n780,n781);
and (n797,n795,n798);
xor (n798,n786,n787);
and (n799,n792,n798);
xor (n800,n778,n785);
and (n801,n800,n802);
xor (n802,n803,n759);
xor (n803,n751,n756);
and (n804,n790,n802);
and (n805,n788,n806);
xor (n806,n807,n765);
xor (n807,n749,n762);
and (n808,n777,n806);
and (n809,n810,n811);
xor (n810,n773,n775);
or (n811,n812,n837);
and (n812,n813,n815);
xor (n813,n814,n806);
xor (n814,n777,n788);
or (n815,n816,n833,n836);
and (n816,n817,n823);
and (n817,n818,n822);
nor (n818,n819,n821);
not (n819,n820);
xor (n820,n184,n453);
and (n821,n42,n820);
and (n822,n753,n26);
or (n823,n824,n830,n832);
and (n824,n825,n828);
and (n825,n826,n827);
and (n826,n621,n17);
xor (n827,n793,n794);
xor (n828,n829,n798);
xor (n829,n792,n795);
and (n830,n828,n831);
xor (n831,n818,n822);
and (n832,n825,n831);
and (n833,n823,n834);
xor (n834,n835,n802);
xor (n835,n790,n800);
and (n836,n817,n834);
and (n837,n838,n839);
xor (n838,n813,n815);
or (n839,n840,n871);
and (n840,n841,n843);
xor (n841,n842,n834);
xor (n842,n817,n823);
or (n843,n844,n867,n870);
and (n844,n845,n852);
or (n845,n846,n849,n851);
and (n846,n847,n848);
and (n847,n820,n26);
and (n848,n753,n29);
and (n849,n848,n850);
and (n850,n688,n14);
and (n851,n847,n850);
or (n852,n853,n864,n866);
and (n853,n854,n862);
or (n854,n855,n858,n861);
and (n855,n856,n857);
and (n856,n688,n21);
and (n857,n621,n103);
and (n858,n859,n860);
and (n859,n621,n21);
and (n860,n634,n103);
and (n861,n855,n860);
xor (n862,n863,n850);
xor (n863,n847,n848);
and (n864,n862,n865);
xor (n865,n826,n827);
and (n866,n854,n865);
and (n867,n852,n868);
xor (n868,n869,n831);
xor (n869,n825,n828);
and (n870,n845,n868);
and (n871,n872,n873);
xor (n872,n841,n843);
or (n873,n874,n902);
and (n874,n875,n877);
xor (n875,n876,n868);
xor (n876,n845,n852);
or (n877,n878,n898,n901);
and (n878,n879,n882);
and (n879,n880,n881);
and (n880,n753,n14);
and (n881,n688,n17);
or (n882,n883,n894,n897);
and (n883,n884,n893);
or (n884,n885,n890,n892);
and (n885,n886,n889);
and (n886,n887,n888);
and (n887,n753,n21);
and (n888,n688,n103);
and (n889,n753,n17);
and (n890,n889,n891);
xor (n891,n856,n857);
and (n892,n886,n891);
xor (n893,n880,n881);
and (n894,n893,n895);
xor (n895,n896,n860);
xor (n896,n855,n859);
and (n897,n884,n895);
and (n898,n882,n899);
xor (n899,n900,n865);
xor (n900,n854,n862);
and (n901,n879,n899);
and (n902,n903,n904);
xor (n903,n875,n877);
or (n904,n905,n927);
and (n905,n906,n908);
xor (n906,n907,n899);
xor (n907,n879,n882);
and (n908,n909,n925);
or (n909,n910,n921,n924);
and (n910,n911,n920);
or (n911,n912,n917,n919);
and (n912,n913,n916);
and (n913,n914,n915);
and (n914,n820,n21);
and (n915,n753,n103);
and (n916,n820,n17);
and (n917,n916,n918);
xor (n918,n887,n888);
and (n919,n913,n918);
and (n920,n820,n14);
and (n921,n920,n922);
xor (n922,n923,n891);
xor (n923,n886,n889);
and (n924,n911,n922);
xor (n925,n926,n895);
xor (n926,n884,n893);
and (n927,n928,n929);
xor (n928,n906,n908);
and (n929,n930,n931);
and (n930,n820,n29);
xor (n931,n909,n925);
endmodule
