module top (out,n4,n21,n23,n24,n33,n34,n36,n37,n47
        ,n57,n61,n71,n72,n74,n75,n82,n88,n100,n101
        ,n103,n104,n107,n113,n125,n126,n135,n141,n171,n211
        ,n242,n273,n597,n603,n613,n950);
output out;
input n4;
input n21;
input n23;
input n24;
input n33;
input n34;
input n36;
input n37;
input n47;
input n57;
input n61;
input n71;
input n72;
input n74;
input n75;
input n82;
input n88;
input n100;
input n101;
input n103;
input n104;
input n107;
input n113;
input n125;
input n126;
input n135;
input n141;
input n171;
input n211;
input n242;
input n273;
input n597;
input n603;
input n613;
input n950;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n35;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n102;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
xnor (out,n0,n951);
nand (n0,n1,n950);
nand (n1,n2,n554);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
nand (n6,n7,n553);
or (n7,n8,n253);
not (n8,n9);
nand (n9,n10,n252);
nand (n10,n11,n221);
not (n11,n12);
xor (n12,n13,n180);
xor (n13,n14,n91);
xor (n14,n15,n63);
xor (n15,n16,n51);
nand (n16,n17,n43);
or (n17,n18,n28);
not (n18,n19);
nor (n19,n20,n25);
and (n20,n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n4);
and (s0n22,notn22,n23);
and (s1n22,n4,n24);
and (n25,n26,n27);
not (n26,n21);
not (n27,n22);
nand (n28,n29,n40);
nor (n29,n30,n38);
and (n30,n31,n35);
not (n31,n32);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n4);
and (s0n32,notn32,n33);
and (s1n32,n4,n34);
wire s0n35,s1n35,notn35;
or (n35,s0n35,s1n35);
not(notn35,n4);
and (s0n35,notn35,n36);
and (s1n35,n4,n37);
and (n38,n32,n39);
not (n39,n35);
nand (n40,n41,n42);
or (n41,n31,n22);
nand (n42,n22,n31);
nand (n43,n44,n50);
not (n44,n45);
nor (n45,n46,n48);
and (n46,n27,n47);
and (n48,n22,n49);
not (n49,n47);
not (n50,n29);
nor (n51,n52,n58);
nand (n52,n22,n53);
not (n53,n54);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n4);
and (s0n54,notn54,1'b0);
and (s1n54,n4,n56);
and (n56,n57,n24);
nor (n58,n59,n62);
and (n59,n54,n60);
not (n60,n61);
and (n62,n53,n61);
nand (n63,n64,n85);
or (n64,n65,n80);
nand (n65,n66,n77);
not (n66,n67);
nand (n67,n68,n76);
or (n68,n69,n73);
not (n69,n70);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n4);
and (s0n70,notn70,n71);
and (s1n70,n4,n72);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n4);
and (s0n73,notn73,n74);
and (s1n73,n4,n75);
nand (n76,n73,n69);
nand (n77,n78,n79);
or (n78,n69,n35);
nand (n79,n35,n69);
nor (n80,n81,n83);
and (n81,n39,n82);
and (n83,n35,n84);
not (n84,n82);
or (n85,n66,n86);
nor (n86,n87,n89);
and (n87,n39,n88);
and (n89,n35,n90);
not (n90,n88);
xor (n91,n92,n157);
xor (n92,n93,n144);
xor (n93,n94,n117);
nand (n94,n95,n110);
or (n95,n96,n105);
not (n96,n97);
nor (n97,n98,n102);
not (n98,n99);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n4);
and (s0n99,notn99,n100);
and (s1n99,n4,n101);
wire s0n102,s1n102,notn102;
or (n102,s0n102,s1n102);
not(notn102,n4);
and (s0n102,notn102,n103);
and (s1n102,n4,n104);
nor (n105,n106,n108);
and (n106,n98,n107);
and (n108,n99,n109);
not (n109,n107);
or (n110,n111,n116);
nor (n111,n112,n114);
and (n112,n98,n113);
and (n114,n99,n115);
not (n115,n113);
not (n116,n102);
nand (n117,n118,n138);
or (n118,n119,n132);
not (n119,n120);
and (n120,n121,n128);
nand (n121,n122,n127);
or (n122,n123,n73);
not (n123,n124);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n4);
and (s0n124,notn124,n125);
and (s1n124,n4,n126);
nand (n127,n73,n123);
not (n128,n129);
nand (n129,n130,n131);
or (n130,n123,n99);
nand (n131,n99,n123);
nor (n132,n133,n136);
and (n133,n134,n135);
not (n134,n73);
and (n136,n73,n137);
not (n137,n135);
or (n138,n139,n128);
nor (n139,n140,n142);
and (n140,n134,n141);
and (n142,n73,n143);
not (n143,n141);
and (n144,n145,n151);
nand (n145,n146,n150);
or (n146,n96,n147);
nor (n147,n148,n149);
and (n148,n98,n141);
and (n149,n99,n143);
or (n150,n105,n116);
nand (n151,n152,n156);
or (n152,n119,n153);
nor (n153,n154,n155);
and (n154,n134,n88);
and (n155,n73,n90);
or (n156,n128,n132);
or (n157,n158,n179);
and (n158,n159,n173);
xor (n159,n160,n167);
nand (n160,n161,n166);
or (n161,n162,n28);
not (n162,n163);
nor (n163,n164,n165);
and (n164,n61,n22);
and (n165,n60,n27);
nand (n166,n50,n19);
nor (n167,n52,n168);
nor (n168,n169,n172);
and (n169,n54,n170);
not (n170,n171);
and (n172,n53,n171);
nand (n173,n174,n178);
or (n174,n65,n175);
nor (n175,n176,n177);
and (n176,n39,n47);
and (n177,n35,n49);
or (n178,n66,n80);
and (n179,n160,n167);
or (n180,n181,n220);
and (n181,n182,n197);
xor (n182,n183,n184);
xor (n183,n145,n151);
and (n184,n185,n191);
nand (n185,n186,n190);
or (n186,n96,n187);
nor (n187,n188,n189);
and (n188,n98,n135);
and (n189,n99,n137);
or (n190,n147,n116);
nand (n191,n192,n196);
or (n192,n119,n193);
nor (n193,n194,n195);
and (n194,n134,n82);
and (n195,n73,n84);
or (n196,n153,n128);
or (n197,n198,n219);
and (n198,n199,n213);
xor (n199,n200,n207);
nand (n200,n201,n206);
or (n201,n202,n28);
not (n202,n203);
nor (n203,n204,n205);
and (n204,n171,n22);
and (n205,n170,n27);
nand (n206,n50,n163);
nor (n207,n52,n208);
nor (n208,n209,n212);
and (n209,n54,n210);
not (n210,n211);
and (n212,n53,n211);
nand (n213,n214,n218);
or (n214,n65,n215);
nor (n215,n216,n217);
and (n216,n39,n21);
and (n217,n35,n26);
or (n218,n66,n175);
and (n219,n200,n207);
and (n220,n183,n184);
not (n221,n222);
or (n222,n223,n251);
and (n223,n224,n227);
xor (n224,n225,n226);
xor (n225,n159,n173);
xor (n226,n182,n197);
and (n227,n228,n229);
xor (n228,n185,n191);
or (n229,n230,n250);
and (n230,n231,n244);
xor (n231,n232,n238);
nand (n232,n233,n237);
or (n233,n234,n28);
nor (n234,n235,n236);
and (n235,n211,n27);
and (n236,n210,n22);
nand (n237,n203,n50);
nor (n238,n52,n239);
nor (n239,n240,n243);
and (n240,n54,n241);
not (n241,n242);
and (n243,n53,n242);
nand (n244,n245,n249);
or (n245,n96,n246);
nor (n246,n247,n248);
and (n247,n98,n88);
and (n248,n99,n90);
or (n249,n187,n116);
and (n250,n232,n238);
and (n251,n225,n226);
nand (n252,n12,n222);
not (n253,n254);
nand (n254,n255,n408,n552);
nand (n255,n256,n401);
nand (n256,n257,n400);
or (n257,n258,n389);
nor (n258,n259,n388);
and (n259,n260,n360);
not (n260,n261);
nor (n261,n262,n343);
or (n262,n263,n342);
and (n263,n264,n313);
xor (n264,n265,n300);
or (n265,n266,n299);
and (n266,n267,n290);
xor (n267,n268,n280);
nand (n268,n269,n276);
or (n269,n270,n28);
not (n270,n271);
nand (n271,n272,n274);
or (n272,n27,n273);
or (n274,n22,n275);
not (n275,n273);
or (n276,n29,n277);
nor (n277,n278,n279);
and (n278,n242,n27);
and (n279,n241,n22);
nand (n280,n281,n286);
or (n281,n282,n119);
not (n282,n283);
nand (n283,n284,n285);
or (n284,n73,n60);
or (n285,n134,n61);
nand (n286,n129,n287);
nor (n287,n288,n289);
and (n288,n21,n73);
and (n289,n26,n134);
nand (n290,n291,n295);
or (n291,n65,n292);
nor (n292,n293,n294);
and (n293,n39,n211);
and (n294,n35,n210);
or (n295,n66,n296);
nor (n296,n297,n298);
and (n297,n39,n171);
and (n298,n35,n170);
and (n299,n268,n280);
xor (n300,n301,n310);
xor (n301,n302,n304);
and (n302,n303,n273);
not (n303,n52);
nand (n304,n305,n309);
or (n305,n96,n306);
nor (n306,n307,n308);
and (n307,n84,n99);
and (n308,n82,n98);
or (n309,n246,n116);
nand (n310,n311,n312);
or (n311,n28,n277);
or (n312,n29,n234);
xor (n313,n314,n328);
xor (n314,n315,n322);
nand (n315,n316,n318);
or (n316,n119,n317);
not (n317,n287);
or (n318,n128,n319);
nor (n319,n320,n321);
and (n320,n134,n47);
and (n321,n73,n49);
nand (n322,n323,n324);
or (n323,n65,n296);
or (n324,n66,n325);
nor (n325,n326,n327);
and (n326,n39,n61);
and (n327,n35,n60);
and (n328,n329,n334);
nor (n329,n330,n27);
nor (n330,n331,n333);
and (n331,n39,n332);
nand (n332,n32,n273);
and (n333,n31,n275);
nand (n334,n335,n340);
or (n335,n336,n96);
not (n336,n337);
nor (n337,n338,n339);
and (n338,n47,n99);
and (n339,n49,n98);
nand (n340,n341,n102);
not (n341,n306);
and (n342,n265,n300);
xor (n343,n344,n349);
xor (n344,n345,n346);
xor (n345,n231,n244);
or (n346,n347,n348);
and (n347,n314,n328);
and (n348,n315,n322);
xor (n349,n350,n357);
xor (n350,n351,n354);
nand (n351,n352,n353);
or (n352,n65,n325);
or (n353,n66,n215);
nand (n354,n355,n356);
or (n355,n119,n319);
or (n356,n193,n128);
or (n357,n358,n359);
and (n358,n301,n310);
and (n359,n302,n304);
not (n360,n361);
nand (n361,n362,n363);
xor (n362,n264,n313);
or (n363,n364,n387);
and (n364,n365,n386);
xor (n365,n366,n367);
xor (n366,n329,n334);
or (n367,n368,n385);
and (n368,n369,n378);
xor (n369,n370,n371);
and (n370,n50,n273);
nand (n371,n372,n373);
or (n372,n116,n336);
nand (n373,n374,n97);
not (n374,n375);
nor (n375,n376,n377);
and (n376,n21,n98);
and (n377,n26,n99);
nand (n378,n379,n384);
or (n379,n380,n119);
not (n380,n381);
nor (n381,n382,n383);
and (n382,n171,n73);
and (n383,n134,n170);
nand (n384,n129,n283);
and (n385,n370,n371);
xor (n386,n267,n290);
and (n387,n366,n367);
and (n388,n262,n343);
nor (n389,n390,n397);
xor (n390,n391,n394);
xor (n391,n392,n393);
xor (n392,n199,n213);
xor (n393,n228,n229);
or (n394,n395,n396);
and (n395,n350,n357);
and (n396,n351,n354);
or (n397,n398,n399);
and (n398,n344,n349);
and (n399,n345,n346);
nand (n400,n390,n397);
nand (n401,n402,n404);
not (n402,n403);
xor (n403,n224,n227);
not (n404,n405);
or (n405,n406,n407);
and (n406,n391,n394);
and (n407,n392,n393);
nand (n408,n401,n409,n551);
nor (n409,n410,n548);
nor (n410,n411,n546);
and (n411,n412,n541);
or (n412,n413,n540);
and (n413,n414,n456);
xor (n414,n415,n449);
or (n415,n416,n448);
and (n416,n417,n436);
xor (n417,n418,n425);
nand (n418,n419,n424);
or (n419,n420,n119);
not (n420,n421);
nor (n421,n422,n423);
and (n422,n210,n134);
and (n423,n211,n73);
nand (n424,n129,n381);
nand (n425,n426,n431);
or (n426,n427,n66);
not (n427,n428);
nor (n428,n429,n430);
and (n429,n242,n35);
and (n430,n241,n39);
nand (n431,n432,n433);
not (n432,n65);
nand (n433,n434,n435);
or (n434,n39,n273);
or (n435,n35,n275);
xor (n436,n437,n442);
and (n437,n438,n35);
nand (n438,n439,n441);
or (n439,n73,n440);
and (n440,n273,n70);
or (n441,n70,n273);
nand (n442,n443,n447);
or (n443,n96,n444);
nor (n444,n445,n446);
and (n445,n98,n61);
and (n446,n99,n60);
or (n447,n375,n116);
and (n448,n418,n425);
xor (n449,n450,n455);
xor (n450,n451,n454);
nand (n451,n452,n453);
or (n452,n427,n65);
or (n453,n66,n292);
and (n454,n437,n442);
xor (n455,n369,n378);
or (n456,n457,n539);
and (n457,n458,n479);
xor (n458,n459,n478);
or (n459,n460,n477);
and (n460,n461,n470);
xor (n461,n462,n463);
and (n462,n67,n273);
nand (n463,n464,n469);
or (n464,n465,n119);
not (n465,n466);
nor (n466,n467,n468);
and (n467,n242,n73);
and (n468,n241,n134);
nand (n469,n421,n129);
nand (n470,n471,n476);
or (n471,n96,n472);
not (n472,n473);
nor (n473,n474,n475);
and (n474,n170,n98);
and (n475,n171,n99);
or (n476,n444,n116);
and (n477,n462,n463);
xor (n478,n417,n436);
or (n479,n480,n538);
and (n480,n481,n537);
xor (n481,n482,n496);
nor (n482,n483,n491);
not (n483,n484);
nand (n484,n485,n490);
or (n485,n486,n96);
not (n486,n487);
nand (n487,n488,n489);
or (n488,n210,n99);
nand (n489,n99,n210);
nand (n490,n473,n102);
nand (n491,n492,n73);
nand (n492,n493,n495);
or (n493,n99,n494);
and (n494,n273,n124);
or (n495,n124,n273);
nand (n496,n497,n535);
or (n497,n498,n521);
not (n498,n499);
nand (n499,n500,n520);
or (n500,n501,n510);
nor (n501,n502,n509);
nand (n502,n503,n508);
or (n503,n504,n96);
not (n504,n505);
nand (n505,n506,n507);
or (n506,n241,n99);
nand (n507,n99,n241);
nand (n508,n487,n102);
nor (n509,n128,n275);
nand (n510,n511,n518);
nand (n511,n512,n517);
or (n512,n513,n96);
not (n513,n514);
nand (n514,n515,n516);
or (n515,n98,n273);
or (n516,n99,n275);
nand (n517,n505,n102);
nor (n518,n519,n98);
and (n519,n273,n102);
nand (n520,n502,n509);
not (n521,n522);
nand (n522,n523,n531);
not (n523,n524);
nand (n524,n525,n530);
or (n525,n526,n119);
not (n526,n527);
nand (n527,n528,n529);
or (n528,n134,n273);
or (n529,n73,n275);
nand (n530,n129,n466);
nor (n531,n532,n534);
and (n532,n483,n533);
not (n533,n491);
and (n534,n484,n491);
nand (n535,n536,n524);
not (n536,n531);
xor (n537,n461,n470);
and (n538,n482,n496);
and (n539,n459,n478);
and (n540,n415,n449);
or (n541,n542,n543);
xor (n542,n365,n386);
or (n543,n544,n545);
and (n544,n450,n455);
and (n545,n451,n454);
not (n546,n547);
nand (n547,n542,n543);
nand (n548,n549,n260);
not (n549,n550);
nor (n550,n362,n363);
not (n551,n389);
nand (n552,n403,n405);
or (n553,n254,n9);
nand (n554,n555,n3);
xnor (n555,n556,n916);
nand (n556,n557,n903);
or (n557,n558,n849);
not (n558,n559);
and (n559,n560,n771,n843);
nor (n560,n561,n720);
nor (n561,n562,n675);
or (n562,n563,n674);
and (n563,n564,n648);
xor (n564,n565,n590);
xor (n565,n566,n581);
xor (n566,n567,n577);
nand (n567,n568,n573);
or (n568,n569,n28);
not (n569,n570);
nor (n570,n571,n572);
and (n571,n88,n22);
and (n572,n90,n27);
nand (n573,n50,n574);
nor (n574,n575,n576);
and (n575,n135,n22);
and (n576,n137,n27);
nor (n577,n52,n578);
nor (n578,n579,n580);
and (n579,n54,n84);
and (n580,n53,n82);
nand (n581,n582,n586);
or (n582,n65,n583);
nor (n583,n584,n585);
and (n584,n39,n141);
and (n585,n35,n143);
or (n586,n66,n587);
nor (n587,n588,n589);
and (n588,n39,n107);
and (n589,n35,n109);
xor (n590,n591,n628);
xor (n591,n592,n614);
xor (n592,n593,n606);
nand (n593,n594,n600);
or (n594,n96,n595);
nor (n595,n596,n598);
and (n596,n98,n597);
and (n598,n99,n599);
not (n599,n597);
or (n600,n601,n116);
nor (n601,n602,n604);
and (n602,n98,n603);
and (n604,n99,n605);
not (n605,n603);
nand (n606,n607,n611);
or (n607,n119,n608);
nor (n608,n609,n610);
and (n609,n134,n113);
and (n610,n73,n115);
or (n611,n612,n128);
xor (n612,n613,n134);
and (n614,n615,n622);
nand (n615,n616,n621);
or (n616,n96,n617);
nor (n617,n618,n619);
and (n618,n98,n613);
and (n619,n99,n620);
not (n620,n613);
or (n621,n595,n116);
nand (n622,n623,n627);
or (n623,n119,n624);
nor (n624,n625,n626);
and (n625,n134,n107);
and (n626,n73,n109);
or (n627,n128,n608);
or (n628,n629,n647);
and (n629,n630,n641);
xor (n630,n631,n637);
nand (n631,n632,n636);
or (n632,n633,n28);
nor (n633,n634,n635);
and (n634,n82,n27);
and (n635,n84,n22);
nand (n636,n50,n570);
nor (n637,n52,n638);
nor (n638,n639,n640);
and (n639,n54,n49);
and (n640,n53,n47);
nand (n641,n642,n646);
or (n642,n65,n643);
nor (n643,n644,n645);
and (n644,n39,n135);
and (n645,n35,n137);
or (n646,n66,n583);
and (n647,n631,n637);
or (n648,n649,n673);
and (n649,n650,n659);
xor (n650,n651,n652);
xor (n651,n615,n622);
and (n652,n653,n656);
nand (n653,n654,n655);
or (n654,n96,n111);
or (n655,n617,n116);
nand (n656,n657,n658);
or (n657,n119,n139);
or (n658,n624,n128);
or (n659,n660,n672);
and (n660,n661,n669);
xor (n661,n662,n665);
nand (n662,n663,n664);
or (n663,n28,n45);
or (n664,n29,n633);
nor (n665,n52,n666);
nor (n666,n667,n668);
and (n667,n54,n26);
and (n668,n53,n21);
nand (n669,n670,n671);
or (n670,n643,n66);
or (n671,n65,n86);
and (n672,n662,n665);
and (n673,n651,n652);
and (n674,n565,n590);
xor (n675,n676,n717);
xor (n676,n677,n696);
xor (n677,n678,n690);
xor (n678,n679,n686);
nand (n679,n680,n682);
or (n680,n681,n28);
not (n681,n574);
or (n682,n29,n683);
nor (n683,n684,n685);
and (n684,n27,n141);
and (n685,n22,n143);
nor (n686,n52,n687);
nor (n687,n688,n689);
and (n688,n54,n90);
and (n689,n53,n88);
nand (n690,n691,n692);
or (n691,n65,n587);
or (n692,n66,n693);
nor (n693,n694,n695);
and (n694,n39,n113);
and (n695,n35,n115);
xor (n696,n697,n714);
xor (n697,n698,n713);
xor (n698,n699,n707);
nand (n699,n700,n701);
or (n700,n96,n601);
or (n701,n702,n116);
nor (n702,n703,n705);
and (n703,n98,n704);
and (n704,n57,n603);
and (n705,n99,n706);
not (n706,n704);
nand (n707,n708,n709);
or (n708,n612,n119);
nand (n709,n129,n710);
nand (n710,n711,n712);
or (n711,n73,n599);
or (n712,n134,n597);
and (n713,n593,n606);
or (n714,n715,n716);
and (n715,n566,n581);
and (n716,n567,n577);
or (n717,n718,n719);
and (n718,n591,n628);
and (n719,n592,n614);
not (n720,n721);
nand (n721,n722,n767);
not (n722,n723);
xor (n723,n724,n743);
xor (n724,n725,n740);
xor (n725,n726,n734);
xor (n726,n727,n731);
nor (n727,n52,n728);
nor (n728,n729,n730);
and (n729,n54,n137);
and (n730,n53,n135);
nand (n731,n732,n733);
or (n732,n102,n97);
not (n733,n702);
nand (n734,n735,n739);
or (n735,n736,n66);
nor (n736,n737,n738);
and (n737,n613,n39);
and (n738,n620,n35);
or (n739,n65,n693);
or (n740,n741,n742);
and (n741,n697,n714);
and (n742,n698,n713);
xor (n743,n744,n749);
xor (n744,n745,n746);
and (n745,n699,n707);
or (n746,n747,n748);
and (n747,n678,n690);
and (n748,n679,n686);
nand (n749,n750,n766);
or (n750,n751,n759);
not (n751,n752);
nand (n752,n753,n755);
or (n753,n119,n754);
not (n754,n710);
or (n755,n128,n756);
nor (n756,n757,n758);
and (n757,n134,n603);
and (n758,n73,n605);
not (n759,n760);
nand (n760,n761,n762);
or (n761,n28,n683);
or (n762,n29,n763);
nor (n763,n764,n765);
and (n764,n27,n107);
and (n765,n22,n109);
or (n766,n760,n752);
not (n767,n768);
or (n768,n769,n770);
and (n769,n676,n717);
and (n770,n677,n696);
nand (n771,n772,n833);
not (n772,n773);
xor (n773,n774,n825);
xor (n774,n775,n795);
xor (n775,n776,n791);
xor (n776,n777,n782);
nand (n777,n778,n779);
or (n778,n120,n129);
nand (n779,n780,n781);
or (n780,n73,n706);
or (n781,n134,n704);
nand (n782,n783,n787);
or (n783,n65,n784);
nor (n784,n785,n786);
and (n785,n39,n597);
and (n786,n35,n599);
or (n787,n66,n788);
nor (n788,n789,n790);
and (n789,n39,n603);
and (n790,n35,n605);
nor (n791,n52,n792);
nor (n792,n793,n794);
and (n793,n54,n109);
and (n794,n53,n107);
xor (n795,n796,n811);
xor (n796,n797,n806);
nand (n797,n798,n802);
or (n798,n28,n799);
nor (n799,n800,n801);
and (n800,n27,n113);
and (n801,n22,n115);
or (n802,n29,n803);
nor (n803,n804,n805);
and (n804,n27,n613);
and (n805,n22,n620);
nand (n806,n807,n809);
or (n807,n808,n128);
not (n808,n779);
nand (n809,n810,n120);
not (n810,n756);
or (n811,n812,n824);
and (n812,n813,n821);
xor (n813,n814,n818);
nor (n814,n52,n815);
nor (n815,n816,n817);
and (n816,n54,n143);
and (n817,n53,n141);
nand (n818,n819,n820);
or (n819,n65,n736);
or (n820,n66,n784);
nand (n821,n822,n823);
or (n822,n28,n763);
or (n823,n29,n799);
and (n824,n814,n818);
or (n825,n826,n832);
and (n826,n827,n829);
xor (n827,n828,n766);
not (n828,n806);
or (n829,n830,n831);
and (n830,n726,n734);
and (n831,n727,n731);
and (n832,n828,n766);
not (n833,n834);
or (n834,n835,n842);
and (n835,n836,n839);
xor (n836,n837,n838);
xor (n837,n813,n821);
xor (n838,n827,n829);
or (n839,n840,n841);
and (n840,n744,n749);
and (n841,n745,n746);
and (n842,n837,n838);
not (n843,n844);
nor (n844,n845,n846);
xor (n845,n836,n839);
or (n846,n847,n848);
and (n847,n724,n743);
and (n848,n725,n740);
not (n849,n850);
nand (n850,n851,n893,n902);
nand (n851,n254,n852);
nor (n852,n853,n872);
nand (n853,n854,n10);
not (n854,n855);
nor (n855,n856,n869);
xor (n856,n857,n866);
xor (n857,n858,n859);
xor (n858,n661,n669);
xor (n859,n860,n863);
xor (n860,n861,n862);
xor (n861,n653,n656);
and (n862,n94,n117);
or (n863,n864,n865);
and (n864,n15,n63);
and (n865,n16,n51);
or (n866,n867,n868);
and (n867,n92,n157);
and (n868,n93,n144);
or (n869,n870,n871);
and (n870,n13,n180);
and (n871,n14,n91);
nand (n872,n873,n886);
nand (n873,n874,n882);
not (n874,n875);
xor (n875,n876,n879);
xor (n876,n877,n878);
xor (n877,n630,n641);
xor (n878,n650,n659);
or (n879,n880,n881);
and (n880,n860,n863);
and (n881,n861,n862);
not (n882,n883);
or (n883,n884,n885);
and (n884,n857,n866);
and (n885,n858,n859);
nand (n886,n887,n889);
not (n887,n888);
xor (n888,n564,n648);
not (n889,n890);
or (n890,n891,n892);
and (n891,n876,n879);
and (n892,n877,n878);
nand (n893,n894,n886);
nand (n894,n895,n901);
or (n895,n896,n897);
not (n896,n873);
not (n897,n898);
nand (n898,n899,n900);
or (n899,n855,n252);
nand (n900,n856,n869);
nand (n901,n875,n883);
nand (n902,n890,n888);
not (n903,n904);
nand (n904,n905,n915);
or (n905,n906,n907);
not (n906,n771);
not (n907,n908);
nand (n908,n909,n914);
or (n909,n910,n844);
nor (n910,n911,n913);
and (n911,n912,n721);
and (n912,n562,n675);
nor (n913,n722,n767);
nand (n914,n845,n846);
or (n915,n772,n833);
nand (n916,n917,n949);
not (n917,n918);
nor (n918,n919,n922);
or (n919,n920,n921);
and (n920,n774,n825);
and (n921,n775,n795);
xor (n922,n923,n946);
xor (n923,n924,n927);
or (n924,n925,n926);
and (n925,n776,n791);
and (n926,n777,n782);
xor (n927,n928,n939);
xor (n928,n929,n935);
nand (n929,n930,n931);
or (n930,n28,n803);
or (n931,n29,n932);
nor (n932,n933,n934);
and (n933,n27,n597);
and (n934,n22,n599);
nor (n935,n52,n936);
nor (n936,n937,n938);
and (n937,n54,n115);
and (n938,n53,n113);
nor (n939,n940,n942);
and (n940,n432,n941);
not (n941,n788);
and (n942,n67,n943);
nand (n943,n944,n945);
or (n944,n35,n706);
or (n945,n39,n704);
or (n946,n947,n948);
and (n947,n796,n811);
and (n948,n797,n806);
nand (n949,n919,n922);
and (n951,n950,n952);
wire s0n952,s1n952,notn952;
or (n952,s0n952,s1n952);
not(notn952,n4);
and (s0n952,notn952,n953);
and (s1n952,n4,n1971);
xor (n953,n954,n1673);
xor (n954,n955,n1969);
xor (n955,n956,n1668);
xor (n956,n957,n1962);
xor (n957,n958,n1662);
xor (n958,n959,n1950);
xor (n959,n960,n1656);
xor (n960,n961,n1933);
xor (n961,n962,n1650);
xor (n962,n963,n1911);
xor (n963,n964,n1644);
xor (n964,n965,n1884);
xor (n965,n966,n1638);
xor (n966,n967,n1852);
xor (n967,n968,n1632);
xor (n968,n969,n1815);
xor (n969,n970,n1626);
xor (n970,n971,n1773);
xor (n971,n972,n1620);
xor (n972,n973,n1726);
xor (n973,n974,n1614);
xor (n974,n975,n1674);
xor (n975,n976,n1608);
xor (n976,n977,n1605);
xor (n977,n978,n1604);
xor (n978,n979,n1534);
xor (n979,n980,n1533);
xor (n980,n981,n1452);
xor (n981,n982,n1451);
xor (n982,n983,n1365);
xor (n983,n984,n1364);
xor (n984,n985,n1272);
xor (n985,n986,n1271);
xor (n986,n987,n998);
xor (n987,n988,n997);
xor (n988,n989,n996);
xor (n989,n990,n995);
xor (n990,n991,n994);
xor (n991,n992,n993);
and (n992,n704,n102);
and (n993,n704,n99);
and (n994,n992,n993);
and (n995,n704,n124);
and (n996,n990,n995);
and (n997,n704,n73);
or (n998,n999,n1000);
and (n999,n988,n997);
and (n1000,n987,n1001);
or (n1001,n1002,n1186);
and (n1002,n1003,n1185);
xor (n1003,n989,n1004);
or (n1004,n1005,n1097);
and (n1005,n1006,n1096);
xor (n1006,n991,n1007);
or (n1007,n994,n1008);
and (n1008,n1009,n1011);
xor (n1009,n992,n1010);
and (n1010,n603,n99);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
and (n1013,n603,n102);
and (n1014,n597,n99);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
and (n1019,n597,n102);
and (n1020,n613,n99);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
or (n1023,n1024,n1027);
and (n1024,n1025,n1026);
and (n1025,n613,n102);
and (n1026,n113,n99);
and (n1027,n1028,n1029);
xor (n1028,n1025,n1026);
or (n1029,n1030,n1033);
and (n1030,n1031,n1032);
and (n1031,n113,n102);
and (n1032,n107,n99);
and (n1033,n1034,n1035);
xor (n1034,n1031,n1032);
or (n1035,n1036,n1039);
and (n1036,n1037,n1038);
and (n1037,n107,n102);
and (n1038,n141,n99);
and (n1039,n1040,n1041);
xor (n1040,n1037,n1038);
or (n1041,n1042,n1045);
and (n1042,n1043,n1044);
and (n1043,n141,n102);
and (n1044,n135,n99);
and (n1045,n1046,n1047);
xor (n1046,n1043,n1044);
or (n1047,n1048,n1051);
and (n1048,n1049,n1050);
and (n1049,n135,n102);
and (n1050,n88,n99);
and (n1051,n1052,n1053);
xor (n1052,n1049,n1050);
or (n1053,n1054,n1057);
and (n1054,n1055,n1056);
and (n1055,n88,n102);
and (n1056,n82,n99);
and (n1057,n1058,n1059);
xor (n1058,n1055,n1056);
or (n1059,n1060,n1062);
and (n1060,n1061,n338);
and (n1061,n82,n102);
and (n1062,n1063,n1064);
xor (n1063,n1061,n338);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
and (n1066,n47,n102);
and (n1067,n21,n99);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1074);
and (n1071,n1072,n1073);
and (n1072,n21,n102);
and (n1073,n61,n99);
and (n1074,n1075,n1076);
xor (n1075,n1072,n1073);
or (n1076,n1077,n1079);
and (n1077,n1078,n475);
and (n1078,n61,n102);
and (n1079,n1080,n1081);
xor (n1080,n1078,n475);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
and (n1083,n171,n102);
and (n1084,n211,n99);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
and (n1089,n211,n102);
and (n1090,n242,n99);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
and (n1093,n1094,n1095);
and (n1094,n242,n102);
and (n1095,n273,n99);
and (n1096,n603,n124);
and (n1097,n1098,n1099);
xor (n1098,n1006,n1096);
or (n1099,n1100,n1103);
and (n1100,n1101,n1102);
xor (n1101,n1009,n1011);
and (n1102,n597,n124);
and (n1103,n1104,n1105);
xor (n1104,n1101,n1102);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
xor (n1107,n1016,n1017);
and (n1108,n613,n124);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
xor (n1113,n1022,n1023);
and (n1114,n113,n124);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
xor (n1119,n1028,n1029);
and (n1120,n107,n124);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
xor (n1125,n1034,n1035);
and (n1126,n141,n124);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
xor (n1131,n1040,n1041);
and (n1132,n135,n124);
and (n1133,n1134,n1135);
xor (n1134,n1131,n1132);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
xor (n1137,n1046,n1047);
and (n1138,n88,n124);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
xor (n1143,n1052,n1053);
and (n1144,n82,n124);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
xor (n1149,n1058,n1059);
and (n1150,n47,n124);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
xor (n1155,n1063,n1064);
and (n1156,n21,n124);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1163);
and (n1160,n1161,n1162);
xor (n1161,n1069,n1070);
and (n1162,n61,n124);
and (n1163,n1164,n1165);
xor (n1164,n1161,n1162);
or (n1165,n1166,n1169);
and (n1166,n1167,n1168);
xor (n1167,n1075,n1076);
and (n1168,n171,n124);
and (n1169,n1170,n1171);
xor (n1170,n1167,n1168);
or (n1171,n1172,n1175);
and (n1172,n1173,n1174);
xor (n1173,n1080,n1081);
and (n1174,n211,n124);
and (n1175,n1176,n1177);
xor (n1176,n1173,n1174);
or (n1177,n1178,n1181);
and (n1178,n1179,n1180);
xor (n1179,n1086,n1087);
and (n1180,n242,n124);
and (n1181,n1182,n1183);
xor (n1182,n1179,n1180);
and (n1183,n1184,n494);
xor (n1184,n1092,n1093);
and (n1185,n603,n73);
and (n1186,n1187,n1188);
xor (n1187,n1003,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1098,n1099);
and (n1191,n597,n73);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1104,n1105);
and (n1197,n613,n73);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1110,n1111);
and (n1203,n113,n73);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1116,n1117);
and (n1209,n107,n73);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1122,n1123);
and (n1215,n141,n73);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1128,n1129);
and (n1221,n135,n73);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1134,n1135);
and (n1227,n88,n73);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1140,n1141);
and (n1233,n82,n73);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1146,n1147);
and (n1239,n47,n73);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1245);
and (n1243,n1244,n288);
xor (n1244,n1152,n1153);
and (n1245,n1246,n1247);
xor (n1246,n1244,n288);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1158,n1159);
and (n1250,n61,n73);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1256);
and (n1254,n1255,n382);
xor (n1255,n1164,n1165);
and (n1256,n1257,n1258);
xor (n1257,n1255,n382);
or (n1258,n1259,n1261);
and (n1259,n1260,n423);
xor (n1260,n1170,n1171);
and (n1261,n1262,n1263);
xor (n1262,n1260,n423);
or (n1263,n1264,n1266);
and (n1264,n1265,n467);
xor (n1265,n1176,n1177);
and (n1266,n1267,n1268);
xor (n1267,n1265,n467);
and (n1268,n1269,n1270);
xor (n1269,n1182,n1183);
and (n1270,n273,n73);
and (n1271,n704,n70);
or (n1272,n1273,n1276);
and (n1273,n1274,n1275);
xor (n1274,n987,n1001);
and (n1275,n603,n70);
and (n1276,n1277,n1278);
xor (n1277,n1274,n1275);
or (n1278,n1279,n1282);
and (n1279,n1280,n1281);
xor (n1280,n1187,n1188);
and (n1281,n597,n70);
and (n1282,n1283,n1284);
xor (n1283,n1280,n1281);
or (n1284,n1285,n1288);
and (n1285,n1286,n1287);
xor (n1286,n1193,n1194);
and (n1287,n613,n70);
and (n1288,n1289,n1290);
xor (n1289,n1286,n1287);
or (n1290,n1291,n1294);
and (n1291,n1292,n1293);
xor (n1292,n1199,n1200);
and (n1293,n113,n70);
and (n1294,n1295,n1296);
xor (n1295,n1292,n1293);
or (n1296,n1297,n1300);
and (n1297,n1298,n1299);
xor (n1298,n1205,n1206);
and (n1299,n107,n70);
and (n1300,n1301,n1302);
xor (n1301,n1298,n1299);
or (n1302,n1303,n1306);
and (n1303,n1304,n1305);
xor (n1304,n1211,n1212);
and (n1305,n141,n70);
and (n1306,n1307,n1308);
xor (n1307,n1304,n1305);
or (n1308,n1309,n1312);
and (n1309,n1310,n1311);
xor (n1310,n1217,n1218);
and (n1311,n135,n70);
and (n1312,n1313,n1314);
xor (n1313,n1310,n1311);
or (n1314,n1315,n1318);
and (n1315,n1316,n1317);
xor (n1316,n1223,n1224);
and (n1317,n88,n70);
and (n1318,n1319,n1320);
xor (n1319,n1316,n1317);
or (n1320,n1321,n1324);
and (n1321,n1322,n1323);
xor (n1322,n1229,n1230);
and (n1323,n82,n70);
and (n1324,n1325,n1326);
xor (n1325,n1322,n1323);
or (n1326,n1327,n1330);
and (n1327,n1328,n1329);
xor (n1328,n1235,n1236);
and (n1329,n47,n70);
and (n1330,n1331,n1332);
xor (n1331,n1328,n1329);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1241,n1242);
and (n1335,n21,n70);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1246,n1247);
and (n1341,n61,n70);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1252,n1253);
and (n1347,n171,n70);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1257,n1258);
and (n1353,n211,n70);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1262,n1263);
and (n1359,n242,n70);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
and (n1362,n1363,n440);
xor (n1363,n1267,n1268);
and (n1364,n603,n35);
or (n1365,n1366,n1369);
and (n1366,n1367,n1368);
xor (n1367,n1277,n1278);
and (n1368,n597,n35);
and (n1369,n1370,n1371);
xor (n1370,n1367,n1368);
or (n1371,n1372,n1375);
and (n1372,n1373,n1374);
xor (n1373,n1283,n1284);
and (n1374,n613,n35);
and (n1375,n1376,n1377);
xor (n1376,n1373,n1374);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1289,n1290);
and (n1380,n113,n35);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1295,n1296);
and (n1386,n107,n35);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1301,n1302);
and (n1392,n141,n35);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1307,n1308);
and (n1398,n135,n35);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
or (n1401,n1402,n1405);
and (n1402,n1403,n1404);
xor (n1403,n1313,n1314);
and (n1404,n88,n35);
and (n1405,n1406,n1407);
xor (n1406,n1403,n1404);
or (n1407,n1408,n1411);
and (n1408,n1409,n1410);
xor (n1409,n1319,n1320);
and (n1410,n82,n35);
and (n1411,n1412,n1413);
xor (n1412,n1409,n1410);
or (n1413,n1414,n1417);
and (n1414,n1415,n1416);
xor (n1415,n1325,n1326);
and (n1416,n47,n35);
and (n1417,n1418,n1419);
xor (n1418,n1415,n1416);
or (n1419,n1420,n1423);
and (n1420,n1421,n1422);
xor (n1421,n1331,n1332);
and (n1422,n21,n35);
and (n1423,n1424,n1425);
xor (n1424,n1421,n1422);
or (n1425,n1426,n1429);
and (n1426,n1427,n1428);
xor (n1427,n1337,n1338);
and (n1428,n61,n35);
and (n1429,n1430,n1431);
xor (n1430,n1427,n1428);
or (n1431,n1432,n1435);
and (n1432,n1433,n1434);
xor (n1433,n1343,n1344);
and (n1434,n171,n35);
and (n1435,n1436,n1437);
xor (n1436,n1433,n1434);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1349,n1350);
and (n1440,n211,n35);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
or (n1443,n1444,n1446);
and (n1444,n1445,n429);
xor (n1445,n1355,n1356);
and (n1446,n1447,n1448);
xor (n1447,n1445,n429);
and (n1448,n1449,n1450);
xor (n1449,n1361,n1362);
and (n1450,n273,n35);
and (n1451,n597,n32);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1370,n1371);
and (n1455,n613,n32);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1376,n1377);
and (n1461,n113,n32);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1382,n1383);
and (n1467,n107,n32);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
or (n1470,n1471,n1474);
and (n1471,n1472,n1473);
xor (n1472,n1388,n1389);
and (n1473,n141,n32);
and (n1474,n1475,n1476);
xor (n1475,n1472,n1473);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1394,n1395);
and (n1479,n135,n32);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1400,n1401);
and (n1485,n88,n32);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1406,n1407);
and (n1491,n82,n32);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1412,n1413);
and (n1497,n47,n32);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1418,n1419);
and (n1503,n21,n32);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1424,n1425);
and (n1509,n61,n32);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1430,n1431);
and (n1515,n171,n32);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1436,n1437);
and (n1521,n211,n32);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1442,n1443);
and (n1527,n242,n32);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
and (n1530,n1531,n1532);
xor (n1531,n1447,n1448);
not (n1532,n332);
and (n1533,n613,n22);
or (n1534,n1535,n1538);
and (n1535,n1536,n1537);
xor (n1536,n1457,n1458);
and (n1537,n113,n22);
and (n1538,n1539,n1540);
xor (n1539,n1536,n1537);
or (n1540,n1541,n1544);
and (n1541,n1542,n1543);
xor (n1542,n1463,n1464);
and (n1543,n107,n22);
and (n1544,n1545,n1546);
xor (n1545,n1542,n1543);
or (n1546,n1547,n1550);
and (n1547,n1548,n1549);
xor (n1548,n1469,n1470);
and (n1549,n141,n22);
and (n1550,n1551,n1552);
xor (n1551,n1548,n1549);
or (n1552,n1553,n1555);
and (n1553,n1554,n575);
xor (n1554,n1475,n1476);
and (n1555,n1556,n1557);
xor (n1556,n1554,n575);
or (n1557,n1558,n1560);
and (n1558,n1559,n571);
xor (n1559,n1481,n1482);
and (n1560,n1561,n1562);
xor (n1561,n1559,n571);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
xor (n1564,n1487,n1488);
and (n1565,n82,n22);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
or (n1568,n1569,n1572);
and (n1569,n1570,n1571);
xor (n1570,n1493,n1494);
and (n1571,n47,n22);
and (n1572,n1573,n1574);
xor (n1573,n1570,n1571);
or (n1574,n1575,n1577);
and (n1575,n1576,n20);
xor (n1576,n1499,n1500);
and (n1577,n1578,n1579);
xor (n1578,n1576,n20);
or (n1579,n1580,n1582);
and (n1580,n1581,n164);
xor (n1581,n1505,n1506);
and (n1582,n1583,n1584);
xor (n1583,n1581,n164);
or (n1584,n1585,n1587);
and (n1585,n1586,n204);
xor (n1586,n1511,n1512);
and (n1587,n1588,n1589);
xor (n1588,n1586,n204);
or (n1589,n1590,n1593);
and (n1590,n1591,n1592);
xor (n1591,n1517,n1518);
and (n1592,n211,n22);
and (n1593,n1594,n1595);
xor (n1594,n1591,n1592);
or (n1595,n1596,n1599);
and (n1596,n1597,n1598);
xor (n1597,n1523,n1524);
and (n1598,n242,n22);
and (n1599,n1600,n1601);
xor (n1600,n1597,n1598);
and (n1601,n1602,n1603);
xor (n1602,n1529,n1530);
and (n1603,n273,n22);
and (n1604,n113,n54);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1539,n1540);
and (n1608,n107,n54);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1545,n1546);
and (n1614,n141,n54);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1551,n1552);
and (n1620,n135,n54);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1556,n1557);
and (n1626,n88,n54);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1633);
and (n1630,n1631,n1632);
xor (n1631,n1561,n1562);
and (n1632,n82,n54);
and (n1633,n1634,n1635);
xor (n1634,n1631,n1632);
or (n1635,n1636,n1639);
and (n1636,n1637,n1638);
xor (n1637,n1567,n1568);
and (n1638,n47,n54);
and (n1639,n1640,n1641);
xor (n1640,n1637,n1638);
or (n1641,n1642,n1645);
and (n1642,n1643,n1644);
xor (n1643,n1573,n1574);
and (n1644,n21,n54);
and (n1645,n1646,n1647);
xor (n1646,n1643,n1644);
or (n1647,n1648,n1651);
and (n1648,n1649,n1650);
xor (n1649,n1578,n1579);
and (n1650,n61,n54);
and (n1651,n1652,n1653);
xor (n1652,n1649,n1650);
or (n1653,n1654,n1657);
and (n1654,n1655,n1656);
xor (n1655,n1583,n1584);
and (n1656,n171,n54);
and (n1657,n1658,n1659);
xor (n1658,n1655,n1656);
or (n1659,n1660,n1663);
and (n1660,n1661,n1662);
xor (n1661,n1588,n1589);
and (n1662,n211,n54);
and (n1663,n1664,n1665);
xor (n1664,n1661,n1662);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n1594,n1595);
and (n1668,n242,n54);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
and (n1671,n1672,n1673);
xor (n1672,n1600,n1601);
and (n1673,n273,n54);
or (n1674,n1675,n1677);
and (n1675,n1676,n1614);
xor (n1676,n1610,n1611);
and (n1677,n1678,n1679);
xor (n1678,n1676,n1614);
or (n1679,n1680,n1682);
and (n1680,n1681,n1620);
xor (n1681,n1616,n1617);
and (n1682,n1683,n1684);
xor (n1683,n1681,n1620);
or (n1684,n1685,n1687);
and (n1685,n1686,n1626);
xor (n1686,n1622,n1623);
and (n1687,n1688,n1689);
xor (n1688,n1686,n1626);
or (n1689,n1690,n1692);
and (n1690,n1691,n1632);
xor (n1691,n1628,n1629);
and (n1692,n1693,n1694);
xor (n1693,n1691,n1632);
or (n1694,n1695,n1697);
and (n1695,n1696,n1638);
xor (n1696,n1634,n1635);
and (n1697,n1698,n1699);
xor (n1698,n1696,n1638);
or (n1699,n1700,n1702);
and (n1700,n1701,n1644);
xor (n1701,n1640,n1641);
and (n1702,n1703,n1704);
xor (n1703,n1701,n1644);
or (n1704,n1705,n1707);
and (n1705,n1706,n1650);
xor (n1706,n1646,n1647);
and (n1707,n1708,n1709);
xor (n1708,n1706,n1650);
or (n1709,n1710,n1712);
and (n1710,n1711,n1656);
xor (n1711,n1652,n1653);
and (n1712,n1713,n1714);
xor (n1713,n1711,n1656);
or (n1714,n1715,n1717);
and (n1715,n1716,n1662);
xor (n1716,n1658,n1659);
and (n1717,n1718,n1719);
xor (n1718,n1716,n1662);
or (n1719,n1720,n1722);
and (n1720,n1721,n1668);
xor (n1721,n1664,n1665);
and (n1722,n1723,n1724);
xor (n1723,n1721,n1668);
and (n1724,n1725,n1673);
xor (n1725,n1670,n1671);
or (n1726,n1727,n1729);
and (n1727,n1728,n1620);
xor (n1728,n1678,n1679);
and (n1729,n1730,n1731);
xor (n1730,n1728,n1620);
or (n1731,n1732,n1734);
and (n1732,n1733,n1626);
xor (n1733,n1683,n1684);
and (n1734,n1735,n1736);
xor (n1735,n1733,n1626);
or (n1736,n1737,n1739);
and (n1737,n1738,n1632);
xor (n1738,n1688,n1689);
and (n1739,n1740,n1741);
xor (n1740,n1738,n1632);
or (n1741,n1742,n1744);
and (n1742,n1743,n1638);
xor (n1743,n1693,n1694);
and (n1744,n1745,n1746);
xor (n1745,n1743,n1638);
or (n1746,n1747,n1749);
and (n1747,n1748,n1644);
xor (n1748,n1698,n1699);
and (n1749,n1750,n1751);
xor (n1750,n1748,n1644);
or (n1751,n1752,n1754);
and (n1752,n1753,n1650);
xor (n1753,n1703,n1704);
and (n1754,n1755,n1756);
xor (n1755,n1753,n1650);
or (n1756,n1757,n1759);
and (n1757,n1758,n1656);
xor (n1758,n1708,n1709);
and (n1759,n1760,n1761);
xor (n1760,n1758,n1656);
or (n1761,n1762,n1764);
and (n1762,n1763,n1662);
xor (n1763,n1713,n1714);
and (n1764,n1765,n1766);
xor (n1765,n1763,n1662);
or (n1766,n1767,n1769);
and (n1767,n1768,n1668);
xor (n1768,n1718,n1719);
and (n1769,n1770,n1771);
xor (n1770,n1768,n1668);
and (n1771,n1772,n1673);
xor (n1772,n1723,n1724);
or (n1773,n1774,n1776);
and (n1774,n1775,n1626);
xor (n1775,n1730,n1731);
and (n1776,n1777,n1778);
xor (n1777,n1775,n1626);
or (n1778,n1779,n1781);
and (n1779,n1780,n1632);
xor (n1780,n1735,n1736);
and (n1781,n1782,n1783);
xor (n1782,n1780,n1632);
or (n1783,n1784,n1786);
and (n1784,n1785,n1638);
xor (n1785,n1740,n1741);
and (n1786,n1787,n1788);
xor (n1787,n1785,n1638);
or (n1788,n1789,n1791);
and (n1789,n1790,n1644);
xor (n1790,n1745,n1746);
and (n1791,n1792,n1793);
xor (n1792,n1790,n1644);
or (n1793,n1794,n1796);
and (n1794,n1795,n1650);
xor (n1795,n1750,n1751);
and (n1796,n1797,n1798);
xor (n1797,n1795,n1650);
or (n1798,n1799,n1801);
and (n1799,n1800,n1656);
xor (n1800,n1755,n1756);
and (n1801,n1802,n1803);
xor (n1802,n1800,n1656);
or (n1803,n1804,n1806);
and (n1804,n1805,n1662);
xor (n1805,n1760,n1761);
and (n1806,n1807,n1808);
xor (n1807,n1805,n1662);
or (n1808,n1809,n1811);
and (n1809,n1810,n1668);
xor (n1810,n1765,n1766);
and (n1811,n1812,n1813);
xor (n1812,n1810,n1668);
and (n1813,n1814,n1673);
xor (n1814,n1770,n1771);
or (n1815,n1816,n1818);
and (n1816,n1817,n1632);
xor (n1817,n1777,n1778);
and (n1818,n1819,n1820);
xor (n1819,n1817,n1632);
or (n1820,n1821,n1823);
and (n1821,n1822,n1638);
xor (n1822,n1782,n1783);
and (n1823,n1824,n1825);
xor (n1824,n1822,n1638);
or (n1825,n1826,n1828);
and (n1826,n1827,n1644);
xor (n1827,n1787,n1788);
and (n1828,n1829,n1830);
xor (n1829,n1827,n1644);
or (n1830,n1831,n1833);
and (n1831,n1832,n1650);
xor (n1832,n1792,n1793);
and (n1833,n1834,n1835);
xor (n1834,n1832,n1650);
or (n1835,n1836,n1838);
and (n1836,n1837,n1656);
xor (n1837,n1797,n1798);
and (n1838,n1839,n1840);
xor (n1839,n1837,n1656);
or (n1840,n1841,n1843);
and (n1841,n1842,n1662);
xor (n1842,n1802,n1803);
and (n1843,n1844,n1845);
xor (n1844,n1842,n1662);
or (n1845,n1846,n1848);
and (n1846,n1847,n1668);
xor (n1847,n1807,n1808);
and (n1848,n1849,n1850);
xor (n1849,n1847,n1668);
and (n1850,n1851,n1673);
xor (n1851,n1812,n1813);
or (n1852,n1853,n1855);
and (n1853,n1854,n1638);
xor (n1854,n1819,n1820);
and (n1855,n1856,n1857);
xor (n1856,n1854,n1638);
or (n1857,n1858,n1860);
and (n1858,n1859,n1644);
xor (n1859,n1824,n1825);
and (n1860,n1861,n1862);
xor (n1861,n1859,n1644);
or (n1862,n1863,n1865);
and (n1863,n1864,n1650);
xor (n1864,n1829,n1830);
and (n1865,n1866,n1867);
xor (n1866,n1864,n1650);
or (n1867,n1868,n1870);
and (n1868,n1869,n1656);
xor (n1869,n1834,n1835);
and (n1870,n1871,n1872);
xor (n1871,n1869,n1656);
or (n1872,n1873,n1875);
and (n1873,n1874,n1662);
xor (n1874,n1839,n1840);
and (n1875,n1876,n1877);
xor (n1876,n1874,n1662);
or (n1877,n1878,n1880);
and (n1878,n1879,n1668);
xor (n1879,n1844,n1845);
and (n1880,n1881,n1882);
xor (n1881,n1879,n1668);
and (n1882,n1883,n1673);
xor (n1883,n1849,n1850);
or (n1884,n1885,n1887);
and (n1885,n1886,n1644);
xor (n1886,n1856,n1857);
and (n1887,n1888,n1889);
xor (n1888,n1886,n1644);
or (n1889,n1890,n1892);
and (n1890,n1891,n1650);
xor (n1891,n1861,n1862);
and (n1892,n1893,n1894);
xor (n1893,n1891,n1650);
or (n1894,n1895,n1897);
and (n1895,n1896,n1656);
xor (n1896,n1866,n1867);
and (n1897,n1898,n1899);
xor (n1898,n1896,n1656);
or (n1899,n1900,n1902);
and (n1900,n1901,n1662);
xor (n1901,n1871,n1872);
and (n1902,n1903,n1904);
xor (n1903,n1901,n1662);
or (n1904,n1905,n1907);
and (n1905,n1906,n1668);
xor (n1906,n1876,n1877);
and (n1907,n1908,n1909);
xor (n1908,n1906,n1668);
and (n1909,n1910,n1673);
xor (n1910,n1881,n1882);
or (n1911,n1912,n1914);
and (n1912,n1913,n1650);
xor (n1913,n1888,n1889);
and (n1914,n1915,n1916);
xor (n1915,n1913,n1650);
or (n1916,n1917,n1919);
and (n1917,n1918,n1656);
xor (n1918,n1893,n1894);
and (n1919,n1920,n1921);
xor (n1920,n1918,n1656);
or (n1921,n1922,n1924);
and (n1922,n1923,n1662);
xor (n1923,n1898,n1899);
and (n1924,n1925,n1926);
xor (n1925,n1923,n1662);
or (n1926,n1927,n1929);
and (n1927,n1928,n1668);
xor (n1928,n1903,n1904);
and (n1929,n1930,n1931);
xor (n1930,n1928,n1668);
and (n1931,n1932,n1673);
xor (n1932,n1908,n1909);
or (n1933,n1934,n1936);
and (n1934,n1935,n1656);
xor (n1935,n1915,n1916);
and (n1936,n1937,n1938);
xor (n1937,n1935,n1656);
or (n1938,n1939,n1941);
and (n1939,n1940,n1662);
xor (n1940,n1920,n1921);
and (n1941,n1942,n1943);
xor (n1942,n1940,n1662);
or (n1943,n1944,n1946);
and (n1944,n1945,n1668);
xor (n1945,n1925,n1926);
and (n1946,n1947,n1948);
xor (n1947,n1945,n1668);
and (n1948,n1949,n1673);
xor (n1949,n1930,n1931);
or (n1950,n1951,n1953);
and (n1951,n1952,n1662);
xor (n1952,n1937,n1938);
and (n1953,n1954,n1955);
xor (n1954,n1952,n1662);
or (n1955,n1956,n1958);
and (n1956,n1957,n1668);
xor (n1957,n1942,n1943);
and (n1958,n1959,n1960);
xor (n1959,n1957,n1668);
and (n1960,n1961,n1673);
xor (n1961,n1947,n1948);
or (n1962,n1963,n1965);
and (n1963,n1964,n1668);
xor (n1964,n1954,n1955);
and (n1965,n1966,n1967);
xor (n1966,n1964,n1668);
and (n1967,n1968,n1673);
xor (n1968,n1959,n1960);
and (n1969,n1970,n1673);
xor (n1970,n1966,n1967);
xor (n1971,n1851,n1673);
endmodule
