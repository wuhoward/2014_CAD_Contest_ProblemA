module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n434,n493,n546,n593,n634,n690,n691,n695,n697,n704
        ,n711,n718,n725,n732,n739,n746,n753,n760,n766,n768
        ,n835,n902,n969,n1036,n1101,n1160,n1213,n1260,n1301,n1335);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n434;
input n493;
input n546;
input n593;
input n634;
input n690;
input n691;
input n695;
input n697;
input n704;
input n711;
input n718;
input n725;
input n732;
input n739;
input n746;
input n753;
input n760;
input n766;
input n768;
input n835;
input n902;
input n969;
input n1036;
input n1101;
input n1160;
input n1213;
input n1260;
input n1301;
input n1335;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n692;
wire n693;
wire n694;
wire n696;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n767;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
xor (out,n0,n1336);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1335);
and (s0n0,notn0,n1);
and (s1n0,n1335,n668);
xor (n1,n2,n635);
xor (n2,n3,n633);
xor (n3,n4,n594);
xor (n4,n5,n592);
xor (n5,n6,n547);
xor (n6,n7,n545);
xor (n7,n8,n494);
xor (n8,n9,n492);
xor (n9,n10,n435);
xor (n10,n11,n433);
xor (n11,n12,n370);
xor (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
or (n370,n371,n374);
and (n371,n372,n373);
xor (n372,n304,n305);
and (n373,n30,n369);
and (n374,n375,n376);
xor (n375,n372,n373);
or (n376,n377,n380);
and (n377,n378,n379);
xor (n378,n310,n311);
and (n379,n37,n369);
and (n380,n381,n382);
xor (n381,n378,n379);
or (n382,n383,n386);
and (n383,n384,n385);
xor (n384,n316,n317);
and (n385,n44,n369);
and (n386,n387,n388);
xor (n387,n384,n385);
or (n388,n389,n392);
and (n389,n390,n391);
xor (n390,n322,n323);
and (n391,n51,n369);
and (n392,n393,n394);
xor (n393,n390,n391);
or (n394,n395,n398);
and (n395,n396,n397);
xor (n396,n328,n329);
and (n397,n58,n369);
and (n398,n399,n400);
xor (n399,n396,n397);
or (n400,n401,n404);
and (n401,n402,n403);
xor (n402,n334,n335);
and (n403,n65,n369);
and (n404,n405,n406);
xor (n405,n402,n403);
or (n406,n407,n410);
and (n407,n408,n409);
xor (n408,n340,n341);
and (n409,n72,n369);
and (n410,n411,n412);
xor (n411,n408,n409);
or (n412,n413,n416);
and (n413,n414,n415);
xor (n414,n346,n347);
and (n415,n79,n369);
and (n416,n417,n418);
xor (n417,n414,n415);
or (n418,n419,n422);
and (n419,n420,n421);
xor (n420,n352,n353);
and (n421,n86,n369);
and (n422,n423,n424);
xor (n423,n420,n421);
or (n424,n425,n428);
and (n425,n426,n427);
xor (n426,n358,n359);
and (n427,n93,n369);
and (n428,n429,n430);
xor (n429,n426,n427);
and (n430,n431,n432);
xor (n431,n364,n365);
and (n432,n99,n369);
and (n433,n30,n434);
or (n435,n436,n439);
and (n436,n437,n438);
xor (n437,n375,n376);
and (n438,n37,n434);
and (n439,n440,n441);
xor (n440,n437,n438);
or (n441,n442,n445);
and (n442,n443,n444);
xor (n443,n381,n382);
and (n444,n44,n434);
and (n445,n446,n447);
xor (n446,n443,n444);
or (n447,n448,n451);
and (n448,n449,n450);
xor (n449,n387,n388);
and (n450,n51,n434);
and (n451,n452,n453);
xor (n452,n449,n450);
or (n453,n454,n457);
and (n454,n455,n456);
xor (n455,n393,n394);
and (n456,n58,n434);
and (n457,n458,n459);
xor (n458,n455,n456);
or (n459,n460,n463);
and (n460,n461,n462);
xor (n461,n399,n400);
and (n462,n65,n434);
and (n463,n464,n465);
xor (n464,n461,n462);
or (n465,n466,n469);
and (n466,n467,n468);
xor (n467,n405,n406);
and (n468,n72,n434);
and (n469,n470,n471);
xor (n470,n467,n468);
or (n471,n472,n475);
and (n472,n473,n474);
xor (n473,n411,n412);
and (n474,n79,n434);
and (n475,n476,n477);
xor (n476,n473,n474);
or (n477,n478,n481);
and (n478,n479,n480);
xor (n479,n417,n418);
and (n480,n86,n434);
and (n481,n482,n483);
xor (n482,n479,n480);
or (n483,n484,n487);
and (n484,n485,n486);
xor (n485,n423,n424);
and (n486,n93,n434);
and (n487,n488,n489);
xor (n488,n485,n486);
and (n489,n490,n491);
xor (n490,n429,n430);
and (n491,n99,n434);
and (n492,n37,n493);
or (n494,n495,n498);
and (n495,n496,n497);
xor (n496,n440,n441);
and (n497,n44,n493);
and (n498,n499,n500);
xor (n499,n496,n497);
or (n500,n501,n504);
and (n501,n502,n503);
xor (n502,n446,n447);
and (n503,n51,n493);
and (n504,n505,n506);
xor (n505,n502,n503);
or (n506,n507,n510);
and (n507,n508,n509);
xor (n508,n452,n453);
and (n509,n58,n493);
and (n510,n511,n512);
xor (n511,n508,n509);
or (n512,n513,n516);
and (n513,n514,n515);
xor (n514,n458,n459);
and (n515,n65,n493);
and (n516,n517,n518);
xor (n517,n514,n515);
or (n518,n519,n522);
and (n519,n520,n521);
xor (n520,n464,n465);
and (n521,n72,n493);
and (n522,n523,n524);
xor (n523,n520,n521);
or (n524,n525,n528);
and (n525,n526,n527);
xor (n526,n470,n471);
and (n527,n79,n493);
and (n528,n529,n530);
xor (n529,n526,n527);
or (n530,n531,n534);
and (n531,n532,n533);
xor (n532,n476,n477);
and (n533,n86,n493);
and (n534,n535,n536);
xor (n535,n532,n533);
or (n536,n537,n540);
and (n537,n538,n539);
xor (n538,n482,n483);
and (n539,n93,n493);
and (n540,n541,n542);
xor (n541,n538,n539);
and (n542,n543,n544);
xor (n543,n488,n489);
and (n544,n99,n493);
and (n545,n44,n546);
or (n547,n548,n551);
and (n548,n549,n550);
xor (n549,n499,n500);
and (n550,n51,n546);
and (n551,n552,n553);
xor (n552,n549,n550);
or (n553,n554,n557);
and (n554,n555,n556);
xor (n555,n505,n506);
and (n556,n58,n546);
and (n557,n558,n559);
xor (n558,n555,n556);
or (n559,n560,n563);
and (n560,n561,n562);
xor (n561,n511,n512);
and (n562,n65,n546);
and (n563,n564,n565);
xor (n564,n561,n562);
or (n565,n566,n569);
and (n566,n567,n568);
xor (n567,n517,n518);
and (n568,n72,n546);
and (n569,n570,n571);
xor (n570,n567,n568);
or (n571,n572,n575);
and (n572,n573,n574);
xor (n573,n523,n524);
and (n574,n79,n546);
and (n575,n576,n577);
xor (n576,n573,n574);
or (n577,n578,n581);
and (n578,n579,n580);
xor (n579,n529,n530);
and (n580,n86,n546);
and (n581,n582,n583);
xor (n582,n579,n580);
or (n583,n584,n587);
and (n584,n585,n586);
xor (n585,n535,n536);
and (n586,n93,n546);
and (n587,n588,n589);
xor (n588,n585,n586);
and (n589,n590,n591);
xor (n590,n541,n542);
and (n591,n99,n546);
and (n592,n51,n593);
or (n594,n595,n598);
and (n595,n596,n597);
xor (n596,n552,n553);
and (n597,n58,n593);
and (n598,n599,n600);
xor (n599,n596,n597);
or (n600,n601,n604);
and (n601,n602,n603);
xor (n602,n558,n559);
and (n603,n65,n593);
and (n604,n605,n606);
xor (n605,n602,n603);
or (n606,n607,n610);
and (n607,n608,n609);
xor (n608,n564,n565);
and (n609,n72,n593);
and (n610,n611,n612);
xor (n611,n608,n609);
or (n612,n613,n616);
and (n613,n614,n615);
xor (n614,n570,n571);
and (n615,n79,n593);
and (n616,n617,n618);
xor (n617,n614,n615);
or (n618,n619,n622);
and (n619,n620,n621);
xor (n620,n576,n577);
and (n621,n86,n593);
and (n622,n623,n624);
xor (n623,n620,n621);
or (n624,n625,n628);
and (n625,n626,n627);
xor (n626,n582,n583);
and (n627,n93,n593);
and (n628,n629,n630);
xor (n629,n626,n627);
and (n630,n631,n632);
xor (n631,n588,n589);
and (n632,n99,n593);
and (n633,n58,n634);
or (n635,n636,n639);
and (n636,n637,n638);
xor (n637,n599,n600);
and (n638,n65,n634);
and (n639,n640,n641);
xor (n640,n637,n638);
or (n641,n642,n645);
and (n642,n643,n644);
xor (n643,n605,n606);
and (n644,n72,n634);
and (n645,n646,n647);
xor (n646,n643,n644);
or (n647,n648,n651);
and (n648,n649,n650);
xor (n649,n611,n612);
and (n650,n79,n634);
and (n651,n652,n653);
xor (n652,n649,n650);
or (n653,n654,n657);
and (n654,n655,n656);
xor (n655,n617,n618);
and (n656,n86,n634);
and (n657,n658,n659);
xor (n658,n655,n656);
or (n659,n660,n663);
and (n660,n661,n662);
xor (n661,n623,n624);
and (n662,n93,n634);
and (n663,n664,n665);
xor (n664,n661,n662);
and (n665,n666,n667);
xor (n666,n629,n630);
and (n667,n99,n634);
xor (n668,n669,n1302);
xor (n669,n670,n1300);
xor (n670,n671,n1261);
xor (n671,n672,n1259);
xor (n672,n673,n1214);
xor (n673,n674,n1212);
xor (n674,n675,n1161);
xor (n675,n676,n1159);
xor (n676,n677,n1102);
xor (n677,n678,n1100);
xor (n678,n679,n1037);
xor (n679,n680,n1035);
or (n680,n681,n970);
and (n681,n682,n968);
or (n682,n683,n903);
and (n683,n684,n901);
or (n684,n685,n836);
and (n685,n686,n834);
or (n686,n687,n769);
and (n687,n688,n767);
and (n688,n689,n692);
and (n689,n690,n691);
or (n692,n693,n698);
and (n693,n694,n696);
and (n694,n690,n695);
and (n696,n697,n691);
and (n698,n699,n700);
xor (n699,n694,n696);
or (n700,n701,n705);
and (n701,n702,n703);
and (n702,n697,n695);
and (n703,n704,n691);
and (n705,n706,n707);
xor (n706,n702,n703);
or (n707,n708,n712);
and (n708,n709,n710);
and (n709,n704,n695);
and (n710,n711,n691);
and (n712,n713,n714);
xor (n713,n709,n710);
or (n714,n715,n719);
and (n715,n716,n717);
and (n716,n711,n695);
and (n717,n718,n691);
and (n719,n720,n721);
xor (n720,n716,n717);
or (n721,n722,n726);
and (n722,n723,n724);
and (n723,n718,n695);
and (n724,n725,n691);
and (n726,n727,n728);
xor (n727,n723,n724);
or (n728,n729,n733);
and (n729,n730,n731);
and (n730,n725,n695);
and (n731,n732,n691);
and (n733,n734,n735);
xor (n734,n730,n731);
or (n735,n736,n740);
and (n736,n737,n738);
and (n737,n732,n695);
and (n738,n739,n691);
and (n740,n741,n742);
xor (n741,n737,n738);
or (n742,n743,n747);
and (n743,n744,n745);
and (n744,n739,n695);
and (n745,n746,n691);
and (n747,n748,n749);
xor (n748,n744,n745);
or (n749,n750,n754);
and (n750,n751,n752);
and (n751,n746,n695);
and (n752,n753,n691);
and (n754,n755,n756);
xor (n755,n751,n752);
or (n756,n757,n761);
and (n757,n758,n759);
and (n758,n753,n695);
and (n759,n760,n691);
and (n761,n762,n763);
xor (n762,n758,n759);
and (n763,n764,n765);
and (n764,n760,n695);
and (n765,n766,n691);
and (n767,n690,n768);
and (n769,n770,n771);
xor (n770,n688,n767);
or (n771,n772,n775);
and (n772,n773,n774);
xor (n773,n689,n692);
and (n774,n697,n768);
and (n775,n776,n777);
xor (n776,n773,n774);
or (n777,n778,n781);
and (n778,n779,n780);
xor (n779,n699,n700);
and (n780,n704,n768);
and (n781,n782,n783);
xor (n782,n779,n780);
or (n783,n784,n787);
and (n784,n785,n786);
xor (n785,n706,n707);
and (n786,n711,n768);
and (n787,n788,n789);
xor (n788,n785,n786);
or (n789,n790,n793);
and (n790,n791,n792);
xor (n791,n713,n714);
and (n792,n718,n768);
and (n793,n794,n795);
xor (n794,n791,n792);
or (n795,n796,n799);
and (n796,n797,n798);
xor (n797,n720,n721);
and (n798,n725,n768);
and (n799,n800,n801);
xor (n800,n797,n798);
or (n801,n802,n805);
and (n802,n803,n804);
xor (n803,n727,n728);
and (n804,n732,n768);
and (n805,n806,n807);
xor (n806,n803,n804);
or (n807,n808,n811);
and (n808,n809,n810);
xor (n809,n734,n735);
and (n810,n739,n768);
and (n811,n812,n813);
xor (n812,n809,n810);
or (n813,n814,n817);
and (n814,n815,n816);
xor (n815,n741,n742);
and (n816,n746,n768);
and (n817,n818,n819);
xor (n818,n815,n816);
or (n819,n820,n823);
and (n820,n821,n822);
xor (n821,n748,n749);
and (n822,n753,n768);
and (n823,n824,n825);
xor (n824,n821,n822);
or (n825,n826,n829);
and (n826,n827,n828);
xor (n827,n755,n756);
and (n828,n760,n768);
and (n829,n830,n831);
xor (n830,n827,n828);
and (n831,n832,n833);
xor (n832,n762,n763);
and (n833,n766,n768);
and (n834,n690,n835);
and (n836,n837,n838);
xor (n837,n686,n834);
or (n838,n839,n842);
and (n839,n840,n841);
xor (n840,n770,n771);
and (n841,n697,n835);
and (n842,n843,n844);
xor (n843,n840,n841);
or (n844,n845,n848);
and (n845,n846,n847);
xor (n846,n776,n777);
and (n847,n704,n835);
and (n848,n849,n850);
xor (n849,n846,n847);
or (n850,n851,n854);
and (n851,n852,n853);
xor (n852,n782,n783);
and (n853,n711,n835);
and (n854,n855,n856);
xor (n855,n852,n853);
or (n856,n857,n860);
and (n857,n858,n859);
xor (n858,n788,n789);
and (n859,n718,n835);
and (n860,n861,n862);
xor (n861,n858,n859);
or (n862,n863,n866);
and (n863,n864,n865);
xor (n864,n794,n795);
and (n865,n725,n835);
and (n866,n867,n868);
xor (n867,n864,n865);
or (n868,n869,n872);
and (n869,n870,n871);
xor (n870,n800,n801);
and (n871,n732,n835);
and (n872,n873,n874);
xor (n873,n870,n871);
or (n874,n875,n878);
and (n875,n876,n877);
xor (n876,n806,n807);
and (n877,n739,n835);
and (n878,n879,n880);
xor (n879,n876,n877);
or (n880,n881,n884);
and (n881,n882,n883);
xor (n882,n812,n813);
and (n883,n746,n835);
and (n884,n885,n886);
xor (n885,n882,n883);
or (n886,n887,n890);
and (n887,n888,n889);
xor (n888,n818,n819);
and (n889,n753,n835);
and (n890,n891,n892);
xor (n891,n888,n889);
or (n892,n893,n896);
and (n893,n894,n895);
xor (n894,n824,n825);
and (n895,n760,n835);
and (n896,n897,n898);
xor (n897,n894,n895);
and (n898,n899,n900);
xor (n899,n830,n831);
and (n900,n766,n835);
and (n901,n690,n902);
and (n903,n904,n905);
xor (n904,n684,n901);
or (n905,n906,n909);
and (n906,n907,n908);
xor (n907,n837,n838);
and (n908,n697,n902);
and (n909,n910,n911);
xor (n910,n907,n908);
or (n911,n912,n915);
and (n912,n913,n914);
xor (n913,n843,n844);
and (n914,n704,n902);
and (n915,n916,n917);
xor (n916,n913,n914);
or (n917,n918,n921);
and (n918,n919,n920);
xor (n919,n849,n850);
and (n920,n711,n902);
and (n921,n922,n923);
xor (n922,n919,n920);
or (n923,n924,n927);
and (n924,n925,n926);
xor (n925,n855,n856);
and (n926,n718,n902);
and (n927,n928,n929);
xor (n928,n925,n926);
or (n929,n930,n933);
and (n930,n931,n932);
xor (n931,n861,n862);
and (n932,n725,n902);
and (n933,n934,n935);
xor (n934,n931,n932);
or (n935,n936,n939);
and (n936,n937,n938);
xor (n937,n867,n868);
and (n938,n732,n902);
and (n939,n940,n941);
xor (n940,n937,n938);
or (n941,n942,n945);
and (n942,n943,n944);
xor (n943,n873,n874);
and (n944,n739,n902);
and (n945,n946,n947);
xor (n946,n943,n944);
or (n947,n948,n951);
and (n948,n949,n950);
xor (n949,n879,n880);
and (n950,n746,n902);
and (n951,n952,n953);
xor (n952,n949,n950);
or (n953,n954,n957);
and (n954,n955,n956);
xor (n955,n885,n886);
and (n956,n753,n902);
and (n957,n958,n959);
xor (n958,n955,n956);
or (n959,n960,n963);
and (n960,n961,n962);
xor (n961,n891,n892);
and (n962,n760,n902);
and (n963,n964,n965);
xor (n964,n961,n962);
and (n965,n966,n967);
xor (n966,n897,n898);
and (n967,n766,n902);
and (n968,n690,n969);
and (n970,n971,n972);
xor (n971,n682,n968);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n904,n905);
and (n975,n697,n969);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n910,n911);
and (n981,n704,n969);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n916,n917);
and (n987,n711,n969);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n922,n923);
and (n993,n718,n969);
and (n994,n995,n996);
xor (n995,n992,n993);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n928,n929);
and (n999,n725,n969);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n934,n935);
and (n1005,n732,n969);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n940,n941);
and (n1011,n739,n969);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
xor (n1016,n946,n947);
and (n1017,n746,n969);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1024);
and (n1021,n1022,n1023);
xor (n1022,n952,n953);
and (n1023,n753,n969);
and (n1024,n1025,n1026);
xor (n1025,n1022,n1023);
or (n1026,n1027,n1030);
and (n1027,n1028,n1029);
xor (n1028,n958,n959);
and (n1029,n760,n969);
and (n1030,n1031,n1032);
xor (n1031,n1028,n1029);
and (n1032,n1033,n1034);
xor (n1033,n964,n965);
and (n1034,n766,n969);
and (n1035,n690,n1036);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
xor (n1039,n971,n972);
and (n1040,n697,n1036);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1047);
and (n1044,n1045,n1046);
xor (n1045,n977,n978);
and (n1046,n704,n1036);
and (n1047,n1048,n1049);
xor (n1048,n1045,n1046);
or (n1049,n1050,n1053);
and (n1050,n1051,n1052);
xor (n1051,n983,n984);
and (n1052,n711,n1036);
and (n1053,n1054,n1055);
xor (n1054,n1051,n1052);
or (n1055,n1056,n1059);
and (n1056,n1057,n1058);
xor (n1057,n989,n990);
and (n1058,n718,n1036);
and (n1059,n1060,n1061);
xor (n1060,n1057,n1058);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n995,n996);
and (n1064,n725,n1036);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n1001,n1002);
and (n1070,n732,n1036);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n1007,n1008);
and (n1076,n739,n1036);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
or (n1079,n1080,n1083);
and (n1080,n1081,n1082);
xor (n1081,n1013,n1014);
and (n1082,n746,n1036);
and (n1083,n1084,n1085);
xor (n1084,n1081,n1082);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
xor (n1087,n1019,n1020);
and (n1088,n753,n1036);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
xor (n1093,n1025,n1026);
and (n1094,n760,n1036);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
and (n1097,n1098,n1099);
xor (n1098,n1031,n1032);
and (n1099,n766,n1036);
and (n1100,n697,n1101);
or (n1102,n1103,n1106);
and (n1103,n1104,n1105);
xor (n1104,n1042,n1043);
and (n1105,n704,n1101);
and (n1106,n1107,n1108);
xor (n1107,n1104,n1105);
or (n1108,n1109,n1112);
and (n1109,n1110,n1111);
xor (n1110,n1048,n1049);
and (n1111,n711,n1101);
and (n1112,n1113,n1114);
xor (n1113,n1110,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
xor (n1116,n1054,n1055);
and (n1117,n718,n1101);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1060,n1061);
and (n1123,n725,n1101);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1066,n1067);
and (n1129,n732,n1101);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
xor (n1134,n1072,n1073);
and (n1135,n739,n1101);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
xor (n1140,n1078,n1079);
and (n1141,n746,n1101);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1084,n1085);
and (n1147,n753,n1101);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1090,n1091);
and (n1153,n760,n1101);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
and (n1156,n1157,n1158);
xor (n1157,n1096,n1097);
and (n1158,n766,n1101);
and (n1159,n704,n1160);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n1107,n1108);
and (n1164,n711,n1160);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1113,n1114);
and (n1170,n718,n1160);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1119,n1120);
and (n1176,n725,n1160);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1125,n1126);
and (n1182,n732,n1160);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1131,n1132);
and (n1188,n739,n1160);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1137,n1138);
and (n1194,n746,n1160);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1143,n1144);
and (n1200,n753,n1160);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1149,n1150);
and (n1206,n760,n1160);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
and (n1209,n1210,n1211);
xor (n1210,n1155,n1156);
and (n1211,n766,n1160);
and (n1212,n711,n1213);
or (n1214,n1215,n1218);
and (n1215,n1216,n1217);
xor (n1216,n1166,n1167);
and (n1217,n718,n1213);
and (n1218,n1219,n1220);
xor (n1219,n1216,n1217);
or (n1220,n1221,n1224);
and (n1221,n1222,n1223);
xor (n1222,n1172,n1173);
and (n1223,n725,n1213);
and (n1224,n1225,n1226);
xor (n1225,n1222,n1223);
or (n1226,n1227,n1230);
and (n1227,n1228,n1229);
xor (n1228,n1178,n1179);
and (n1229,n732,n1213);
and (n1230,n1231,n1232);
xor (n1231,n1228,n1229);
or (n1232,n1233,n1236);
and (n1233,n1234,n1235);
xor (n1234,n1184,n1185);
and (n1235,n739,n1213);
and (n1236,n1237,n1238);
xor (n1237,n1234,n1235);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1190,n1191);
and (n1241,n746,n1213);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1196,n1197);
and (n1247,n753,n1213);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1254);
and (n1251,n1252,n1253);
xor (n1252,n1202,n1203);
and (n1253,n760,n1213);
and (n1254,n1255,n1256);
xor (n1255,n1252,n1253);
and (n1256,n1257,n1258);
xor (n1257,n1208,n1209);
and (n1258,n766,n1213);
and (n1259,n718,n1260);
or (n1261,n1262,n1265);
and (n1262,n1263,n1264);
xor (n1263,n1219,n1220);
and (n1264,n725,n1260);
and (n1265,n1266,n1267);
xor (n1266,n1263,n1264);
or (n1267,n1268,n1271);
and (n1268,n1269,n1270);
xor (n1269,n1225,n1226);
and (n1270,n732,n1260);
and (n1271,n1272,n1273);
xor (n1272,n1269,n1270);
or (n1273,n1274,n1277);
and (n1274,n1275,n1276);
xor (n1275,n1231,n1232);
and (n1276,n739,n1260);
and (n1277,n1278,n1279);
xor (n1278,n1275,n1276);
or (n1279,n1280,n1283);
and (n1280,n1281,n1282);
xor (n1281,n1237,n1238);
and (n1282,n746,n1260);
and (n1283,n1284,n1285);
xor (n1284,n1281,n1282);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1243,n1244);
and (n1288,n753,n1260);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1249,n1250);
and (n1294,n760,n1260);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
and (n1297,n1298,n1299);
xor (n1298,n1255,n1256);
and (n1299,n766,n1260);
and (n1300,n725,n1301);
or (n1302,n1303,n1306);
and (n1303,n1304,n1305);
xor (n1304,n1266,n1267);
and (n1305,n732,n1301);
and (n1306,n1307,n1308);
xor (n1307,n1304,n1305);
or (n1308,n1309,n1312);
and (n1309,n1310,n1311);
xor (n1310,n1272,n1273);
and (n1311,n739,n1301);
and (n1312,n1313,n1314);
xor (n1313,n1310,n1311);
or (n1314,n1315,n1318);
and (n1315,n1316,n1317);
xor (n1316,n1278,n1279);
and (n1317,n746,n1301);
and (n1318,n1319,n1320);
xor (n1319,n1316,n1317);
or (n1320,n1321,n1324);
and (n1321,n1322,n1323);
xor (n1322,n1284,n1285);
and (n1323,n753,n1301);
and (n1324,n1325,n1326);
xor (n1325,n1322,n1323);
or (n1326,n1327,n1330);
and (n1327,n1328,n1329);
xor (n1328,n1290,n1291);
and (n1329,n760,n1301);
and (n1330,n1331,n1332);
xor (n1331,n1328,n1329);
and (n1332,n1333,n1334);
xor (n1333,n1296,n1297);
and (n1334,n766,n1301);
xor (n1336,n1337,n1970);
xor (n1337,n1338,n1968);
xor (n1338,n1339,n1929);
xor (n1339,n1340,n1927);
xor (n1340,n1341,n1882);
xor (n1341,n1342,n1880);
xor (n1342,n1343,n1829);
xor (n1343,n1344,n1827);
xor (n1344,n1345,n1770);
xor (n1345,n1346,n1768);
xor (n1346,n1347,n1705);
xor (n1347,n1348,n1703);
or (n1348,n1349,n1638);
and (n1349,n1350,n1636);
or (n1350,n1351,n1571);
and (n1351,n1352,n1569);
or (n1352,n1353,n1504);
and (n1353,n1354,n1502);
or (n1354,n1355,n1437);
and (n1355,n1356,n1435);
and (n1356,n1357,n1360);
and (n1357,n1358,n1359);
wire s0n1358,s1n1358,notn1358;
or (n1358,s0n1358,s1n1358);
not(notn1358,n1335);
and (s0n1358,notn1358,n23);
and (s1n1358,n1335,n690);
wire s0n1359,s1n1359,notn1359;
or (n1359,s0n1359,s1n1359);
not(notn1359,n1335);
and (s0n1359,notn1359,n24);
and (s1n1359,n1335,n691);
or (n1360,n1361,n1366);
and (n1361,n1362,n1364);
and (n1362,n1358,n1363);
wire s0n1363,s1n1363,notn1363;
or (n1363,s0n1363,s1n1363);
not(notn1363,n1335);
and (s0n1363,notn1363,n28);
and (s1n1363,n1335,n695);
and (n1364,n1365,n1359);
wire s0n1365,s1n1365,notn1365;
or (n1365,s0n1365,s1n1365);
not(notn1365,n1335);
and (s0n1365,notn1365,n30);
and (s1n1365,n1335,n697);
and (n1366,n1367,n1368);
xor (n1367,n1362,n1364);
or (n1368,n1369,n1373);
and (n1369,n1370,n1371);
and (n1370,n1365,n1363);
and (n1371,n1372,n1359);
wire s0n1372,s1n1372,notn1372;
or (n1372,s0n1372,s1n1372);
not(notn1372,n1335);
and (s0n1372,notn1372,n37);
and (s1n1372,n1335,n704);
and (n1373,n1374,n1375);
xor (n1374,n1370,n1371);
or (n1375,n1376,n1380);
and (n1376,n1377,n1378);
and (n1377,n1372,n1363);
and (n1378,n1379,n1359);
wire s0n1379,s1n1379,notn1379;
or (n1379,s0n1379,s1n1379);
not(notn1379,n1335);
and (s0n1379,notn1379,n44);
and (s1n1379,n1335,n711);
and (n1380,n1381,n1382);
xor (n1381,n1377,n1378);
or (n1382,n1383,n1387);
and (n1383,n1384,n1385);
and (n1384,n1379,n1363);
and (n1385,n1386,n1359);
wire s0n1386,s1n1386,notn1386;
or (n1386,s0n1386,s1n1386);
not(notn1386,n1335);
and (s0n1386,notn1386,n51);
and (s1n1386,n1335,n718);
and (n1387,n1388,n1389);
xor (n1388,n1384,n1385);
or (n1389,n1390,n1394);
and (n1390,n1391,n1392);
and (n1391,n1386,n1363);
and (n1392,n1393,n1359);
wire s0n1393,s1n1393,notn1393;
or (n1393,s0n1393,s1n1393);
not(notn1393,n1335);
and (s0n1393,notn1393,n58);
and (s1n1393,n1335,n725);
and (n1394,n1395,n1396);
xor (n1395,n1391,n1392);
or (n1396,n1397,n1401);
and (n1397,n1398,n1399);
and (n1398,n1393,n1363);
and (n1399,n1400,n1359);
wire s0n1400,s1n1400,notn1400;
or (n1400,s0n1400,s1n1400);
not(notn1400,n1335);
and (s0n1400,notn1400,n65);
and (s1n1400,n1335,n732);
and (n1401,n1402,n1403);
xor (n1402,n1398,n1399);
or (n1403,n1404,n1408);
and (n1404,n1405,n1406);
and (n1405,n1400,n1363);
and (n1406,n1407,n1359);
wire s0n1407,s1n1407,notn1407;
or (n1407,s0n1407,s1n1407);
not(notn1407,n1335);
and (s0n1407,notn1407,n72);
and (s1n1407,n1335,n739);
and (n1408,n1409,n1410);
xor (n1409,n1405,n1406);
or (n1410,n1411,n1415);
and (n1411,n1412,n1413);
and (n1412,n1407,n1363);
and (n1413,n1414,n1359);
wire s0n1414,s1n1414,notn1414;
or (n1414,s0n1414,s1n1414);
not(notn1414,n1335);
and (s0n1414,notn1414,n79);
and (s1n1414,n1335,n746);
and (n1415,n1416,n1417);
xor (n1416,n1412,n1413);
or (n1417,n1418,n1422);
and (n1418,n1419,n1420);
and (n1419,n1414,n1363);
and (n1420,n1421,n1359);
wire s0n1421,s1n1421,notn1421;
or (n1421,s0n1421,s1n1421);
not(notn1421,n1335);
and (s0n1421,notn1421,n86);
and (s1n1421,n1335,n753);
and (n1422,n1423,n1424);
xor (n1423,n1419,n1420);
or (n1424,n1425,n1429);
and (n1425,n1426,n1427);
and (n1426,n1421,n1363);
and (n1427,n1428,n1359);
wire s0n1428,s1n1428,notn1428;
or (n1428,s0n1428,s1n1428);
not(notn1428,n1335);
and (s0n1428,notn1428,n93);
and (s1n1428,n1335,n760);
and (n1429,n1430,n1431);
xor (n1430,n1426,n1427);
and (n1431,n1432,n1433);
and (n1432,n1428,n1363);
and (n1433,n1434,n1359);
wire s0n1434,s1n1434,notn1434;
or (n1434,s0n1434,s1n1434);
not(notn1434,n1335);
and (s0n1434,notn1434,n99);
and (s1n1434,n1335,n766);
and (n1435,n1358,n1436);
wire s0n1436,s1n1436,notn1436;
or (n1436,s0n1436,s1n1436);
not(notn1436,n1335);
and (s0n1436,notn1436,n101);
and (s1n1436,n1335,n768);
and (n1437,n1438,n1439);
xor (n1438,n1356,n1435);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1357,n1360);
and (n1442,n1365,n1436);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1367,n1368);
and (n1448,n1372,n1436);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1374,n1375);
and (n1454,n1379,n1436);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
or (n1457,n1458,n1461);
and (n1458,n1459,n1460);
xor (n1459,n1381,n1382);
and (n1460,n1386,n1436);
and (n1461,n1462,n1463);
xor (n1462,n1459,n1460);
or (n1463,n1464,n1467);
and (n1464,n1465,n1466);
xor (n1465,n1388,n1389);
and (n1466,n1393,n1436);
and (n1467,n1468,n1469);
xor (n1468,n1465,n1466);
or (n1469,n1470,n1473);
and (n1470,n1471,n1472);
xor (n1471,n1395,n1396);
and (n1472,n1400,n1436);
and (n1473,n1474,n1475);
xor (n1474,n1471,n1472);
or (n1475,n1476,n1479);
and (n1476,n1477,n1478);
xor (n1477,n1402,n1403);
and (n1478,n1407,n1436);
and (n1479,n1480,n1481);
xor (n1480,n1477,n1478);
or (n1481,n1482,n1485);
and (n1482,n1483,n1484);
xor (n1483,n1409,n1410);
and (n1484,n1414,n1436);
and (n1485,n1486,n1487);
xor (n1486,n1483,n1484);
or (n1487,n1488,n1491);
and (n1488,n1489,n1490);
xor (n1489,n1416,n1417);
and (n1490,n1421,n1436);
and (n1491,n1492,n1493);
xor (n1492,n1489,n1490);
or (n1493,n1494,n1497);
and (n1494,n1495,n1496);
xor (n1495,n1423,n1424);
and (n1496,n1428,n1436);
and (n1497,n1498,n1499);
xor (n1498,n1495,n1496);
and (n1499,n1500,n1501);
xor (n1500,n1430,n1431);
and (n1501,n1434,n1436);
and (n1502,n1358,n1503);
wire s0n1503,s1n1503,notn1503;
or (n1503,s0n1503,s1n1503);
not(notn1503,n1335);
and (s0n1503,notn1503,n168);
and (s1n1503,n1335,n835);
and (n1504,n1505,n1506);
xor (n1505,n1354,n1502);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1438,n1439);
and (n1509,n1365,n1503);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1444,n1445);
and (n1515,n1372,n1503);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1450,n1451);
and (n1521,n1379,n1503);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1456,n1457);
and (n1527,n1386,n1503);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1462,n1463);
and (n1533,n1393,n1503);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1468,n1469);
and (n1539,n1400,n1503);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1474,n1475);
and (n1545,n1407,n1503);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1480,n1481);
and (n1551,n1414,n1503);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
xor (n1556,n1486,n1487);
and (n1557,n1421,n1503);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1492,n1493);
and (n1563,n1428,n1503);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
and (n1566,n1567,n1568);
xor (n1567,n1498,n1499);
and (n1568,n1434,n1503);
and (n1569,n1358,n1570);
wire s0n1570,s1n1570,notn1570;
or (n1570,s0n1570,s1n1570);
not(notn1570,n1335);
and (s0n1570,notn1570,n235);
and (s1n1570,n1335,n902);
and (n1571,n1572,n1573);
xor (n1572,n1352,n1569);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1505,n1506);
and (n1576,n1365,n1570);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1511,n1512);
and (n1582,n1372,n1570);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1517,n1518);
and (n1588,n1379,n1570);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1523,n1524);
and (n1594,n1386,n1570);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
or (n1597,n1598,n1601);
and (n1598,n1599,n1600);
xor (n1599,n1529,n1530);
and (n1600,n1393,n1570);
and (n1601,n1602,n1603);
xor (n1602,n1599,n1600);
or (n1603,n1604,n1607);
and (n1604,n1605,n1606);
xor (n1605,n1535,n1536);
and (n1606,n1400,n1570);
and (n1607,n1608,n1609);
xor (n1608,n1605,n1606);
or (n1609,n1610,n1613);
and (n1610,n1611,n1612);
xor (n1611,n1541,n1542);
and (n1612,n1407,n1570);
and (n1613,n1614,n1615);
xor (n1614,n1611,n1612);
or (n1615,n1616,n1619);
and (n1616,n1617,n1618);
xor (n1617,n1547,n1548);
and (n1618,n1414,n1570);
and (n1619,n1620,n1621);
xor (n1620,n1617,n1618);
or (n1621,n1622,n1625);
and (n1622,n1623,n1624);
xor (n1623,n1553,n1554);
and (n1624,n1421,n1570);
and (n1625,n1626,n1627);
xor (n1626,n1623,n1624);
or (n1627,n1628,n1631);
and (n1628,n1629,n1630);
xor (n1629,n1559,n1560);
and (n1630,n1428,n1570);
and (n1631,n1632,n1633);
xor (n1632,n1629,n1630);
and (n1633,n1634,n1635);
xor (n1634,n1565,n1566);
and (n1635,n1434,n1570);
and (n1636,n1358,n1637);
wire s0n1637,s1n1637,notn1637;
or (n1637,s0n1637,s1n1637);
not(notn1637,n1335);
and (s0n1637,notn1637,n302);
and (s1n1637,n1335,n969);
and (n1638,n1639,n1640);
xor (n1639,n1350,n1636);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1572,n1573);
and (n1643,n1365,n1637);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1578,n1579);
and (n1649,n1372,n1637);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1584,n1585);
and (n1655,n1379,n1637);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1590,n1591);
and (n1661,n1386,n1637);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1596,n1597);
and (n1667,n1393,n1637);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
or (n1670,n1671,n1674);
and (n1671,n1672,n1673);
xor (n1672,n1602,n1603);
and (n1673,n1400,n1637);
and (n1674,n1675,n1676);
xor (n1675,n1672,n1673);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1608,n1609);
and (n1679,n1407,n1637);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1614,n1615);
and (n1685,n1414,n1637);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1620,n1621);
and (n1691,n1421,n1637);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1626,n1627);
and (n1697,n1428,n1637);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
and (n1700,n1701,n1702);
xor (n1701,n1632,n1633);
and (n1702,n1434,n1637);
and (n1703,n1358,n1704);
wire s0n1704,s1n1704,notn1704;
or (n1704,s0n1704,s1n1704);
not(notn1704,n1335);
and (s0n1704,notn1704,n369);
and (s1n1704,n1335,n1036);
or (n1705,n1706,n1709);
and (n1706,n1707,n1708);
xor (n1707,n1639,n1640);
and (n1708,n1365,n1704);
and (n1709,n1710,n1711);
xor (n1710,n1707,n1708);
or (n1711,n1712,n1715);
and (n1712,n1713,n1714);
xor (n1713,n1645,n1646);
and (n1714,n1372,n1704);
and (n1715,n1716,n1717);
xor (n1716,n1713,n1714);
or (n1717,n1718,n1721);
and (n1718,n1719,n1720);
xor (n1719,n1651,n1652);
and (n1720,n1379,n1704);
and (n1721,n1722,n1723);
xor (n1722,n1719,n1720);
or (n1723,n1724,n1727);
and (n1724,n1725,n1726);
xor (n1725,n1657,n1658);
and (n1726,n1386,n1704);
and (n1727,n1728,n1729);
xor (n1728,n1725,n1726);
or (n1729,n1730,n1733);
and (n1730,n1731,n1732);
xor (n1731,n1663,n1664);
and (n1732,n1393,n1704);
and (n1733,n1734,n1735);
xor (n1734,n1731,n1732);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1669,n1670);
and (n1738,n1400,n1704);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
or (n1741,n1742,n1745);
and (n1742,n1743,n1744);
xor (n1743,n1675,n1676);
and (n1744,n1407,n1704);
and (n1745,n1746,n1747);
xor (n1746,n1743,n1744);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1681,n1682);
and (n1750,n1414,n1704);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1687,n1688);
and (n1756,n1421,n1704);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1693,n1694);
and (n1762,n1428,n1704);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
and (n1765,n1766,n1767);
xor (n1766,n1699,n1700);
and (n1767,n1434,n1704);
and (n1768,n1365,n1769);
wire s0n1769,s1n1769,notn1769;
or (n1769,s0n1769,s1n1769);
not(notn1769,n1335);
and (s0n1769,notn1769,n434);
and (s1n1769,n1335,n1101);
or (n1770,n1771,n1774);
and (n1771,n1772,n1773);
xor (n1772,n1710,n1711);
and (n1773,n1372,n1769);
and (n1774,n1775,n1776);
xor (n1775,n1772,n1773);
or (n1776,n1777,n1780);
and (n1777,n1778,n1779);
xor (n1778,n1716,n1717);
and (n1779,n1379,n1769);
and (n1780,n1781,n1782);
xor (n1781,n1778,n1779);
or (n1782,n1783,n1786);
and (n1783,n1784,n1785);
xor (n1784,n1722,n1723);
and (n1785,n1386,n1769);
and (n1786,n1787,n1788);
xor (n1787,n1784,n1785);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1728,n1729);
and (n1791,n1393,n1769);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1734,n1735);
and (n1797,n1400,n1769);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
xor (n1802,n1740,n1741);
and (n1803,n1407,n1769);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
xor (n1808,n1746,n1747);
and (n1809,n1414,n1769);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
xor (n1814,n1752,n1753);
and (n1815,n1421,n1769);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
xor (n1820,n1758,n1759);
and (n1821,n1428,n1769);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
and (n1824,n1825,n1826);
xor (n1825,n1764,n1765);
and (n1826,n1434,n1769);
and (n1827,n1372,n1828);
wire s0n1828,s1n1828,notn1828;
or (n1828,s0n1828,s1n1828);
not(notn1828,n1335);
and (s0n1828,notn1828,n493);
and (s1n1828,n1335,n1160);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1775,n1776);
and (n1832,n1379,n1828);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1781,n1782);
and (n1838,n1386,n1828);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
or (n1841,n1842,n1845);
and (n1842,n1843,n1844);
xor (n1843,n1787,n1788);
and (n1844,n1393,n1828);
and (n1845,n1846,n1847);
xor (n1846,n1843,n1844);
or (n1847,n1848,n1851);
and (n1848,n1849,n1850);
xor (n1849,n1793,n1794);
and (n1850,n1400,n1828);
and (n1851,n1852,n1853);
xor (n1852,n1849,n1850);
or (n1853,n1854,n1857);
and (n1854,n1855,n1856);
xor (n1855,n1799,n1800);
and (n1856,n1407,n1828);
and (n1857,n1858,n1859);
xor (n1858,n1855,n1856);
or (n1859,n1860,n1863);
and (n1860,n1861,n1862);
xor (n1861,n1805,n1806);
and (n1862,n1414,n1828);
and (n1863,n1864,n1865);
xor (n1864,n1861,n1862);
or (n1865,n1866,n1869);
and (n1866,n1867,n1868);
xor (n1867,n1811,n1812);
and (n1868,n1421,n1828);
and (n1869,n1870,n1871);
xor (n1870,n1867,n1868);
or (n1871,n1872,n1875);
and (n1872,n1873,n1874);
xor (n1873,n1817,n1818);
and (n1874,n1428,n1828);
and (n1875,n1876,n1877);
xor (n1876,n1873,n1874);
and (n1877,n1878,n1879);
xor (n1878,n1823,n1824);
and (n1879,n1434,n1828);
and (n1880,n1379,n1881);
wire s0n1881,s1n1881,notn1881;
or (n1881,s0n1881,s1n1881);
not(notn1881,n1335);
and (s0n1881,notn1881,n546);
and (s1n1881,n1335,n1213);
or (n1882,n1883,n1886);
and (n1883,n1884,n1885);
xor (n1884,n1834,n1835);
and (n1885,n1386,n1881);
and (n1886,n1887,n1888);
xor (n1887,n1884,n1885);
or (n1888,n1889,n1892);
and (n1889,n1890,n1891);
xor (n1890,n1840,n1841);
and (n1891,n1393,n1881);
and (n1892,n1893,n1894);
xor (n1893,n1890,n1891);
or (n1894,n1895,n1898);
and (n1895,n1896,n1897);
xor (n1896,n1846,n1847);
and (n1897,n1400,n1881);
and (n1898,n1899,n1900);
xor (n1899,n1896,n1897);
or (n1900,n1901,n1904);
and (n1901,n1902,n1903);
xor (n1902,n1852,n1853);
and (n1903,n1407,n1881);
and (n1904,n1905,n1906);
xor (n1905,n1902,n1903);
or (n1906,n1907,n1910);
and (n1907,n1908,n1909);
xor (n1908,n1858,n1859);
and (n1909,n1414,n1881);
and (n1910,n1911,n1912);
xor (n1911,n1908,n1909);
or (n1912,n1913,n1916);
and (n1913,n1914,n1915);
xor (n1914,n1864,n1865);
and (n1915,n1421,n1881);
and (n1916,n1917,n1918);
xor (n1917,n1914,n1915);
or (n1918,n1919,n1922);
and (n1919,n1920,n1921);
xor (n1920,n1870,n1871);
and (n1921,n1428,n1881);
and (n1922,n1923,n1924);
xor (n1923,n1920,n1921);
and (n1924,n1925,n1926);
xor (n1925,n1876,n1877);
and (n1926,n1434,n1881);
and (n1927,n1386,n1928);
wire s0n1928,s1n1928,notn1928;
or (n1928,s0n1928,s1n1928);
not(notn1928,n1335);
and (s0n1928,notn1928,n593);
and (s1n1928,n1335,n1260);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1887,n1888);
and (n1932,n1393,n1928);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1893,n1894);
and (n1938,n1400,n1928);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1899,n1900);
and (n1944,n1407,n1928);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1905,n1906);
and (n1950,n1414,n1928);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1911,n1912);
and (n1956,n1421,n1928);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1963);
and (n1960,n1961,n1962);
xor (n1961,n1917,n1918);
and (n1962,n1428,n1928);
and (n1963,n1964,n1965);
xor (n1964,n1961,n1962);
and (n1965,n1966,n1967);
xor (n1966,n1923,n1924);
and (n1967,n1434,n1928);
and (n1968,n1393,n1969);
wire s0n1969,s1n1969,notn1969;
or (n1969,s0n1969,s1n1969);
not(notn1969,n1335);
and (s0n1969,notn1969,n634);
and (s1n1969,n1335,n1301);
or (n1970,n1971,n1974);
and (n1971,n1972,n1973);
xor (n1972,n1934,n1935);
and (n1973,n1400,n1969);
and (n1974,n1975,n1976);
xor (n1975,n1972,n1973);
or (n1976,n1977,n1980);
and (n1977,n1978,n1979);
xor (n1978,n1940,n1941);
and (n1979,n1407,n1969);
and (n1980,n1981,n1982);
xor (n1981,n1978,n1979);
or (n1982,n1983,n1986);
and (n1983,n1984,n1985);
xor (n1984,n1946,n1947);
and (n1985,n1414,n1969);
and (n1986,n1987,n1988);
xor (n1987,n1984,n1985);
or (n1988,n1989,n1992);
and (n1989,n1990,n1991);
xor (n1990,n1952,n1953);
and (n1991,n1421,n1969);
and (n1992,n1993,n1994);
xor (n1993,n1990,n1991);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1958,n1959);
and (n1997,n1428,n1969);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
and (n2000,n2001,n2002);
xor (n2001,n1964,n1965);
and (n2002,n1434,n1969);
endmodule
