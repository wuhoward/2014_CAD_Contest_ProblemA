module top (out,n13,n16,n17,n21,n24,n25,n29,n37,n40
        ,n41,n45,n55,n58,n59,n63,n70,n73,n74,n78
        ,n86,n89,n90,n94,n104,n107,n108,n112,n117,n326
        ,n420,n491,n577);
output out;
input n13;
input n16;
input n17;
input n21;
input n24;
input n25;
input n29;
input n37;
input n40;
input n41;
input n45;
input n55;
input n58;
input n59;
input n63;
input n70;
input n73;
input n74;
input n78;
input n86;
input n89;
input n90;
input n94;
input n104;
input n107;
input n108;
input n112;
input n117;
input n326;
input n420;
input n491;
input n577;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n105;
wire n106;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
xor (out,n0,n1261);
buf (n0,n1);
xor (n1,n2,n369);
xor (n2,n3,n291);
xor (n3,n4,n242);
or (n4,n5,n193,n241);
and (n5,n6,n183);
or (n6,n7,n153,n182);
and (n7,n8,n119);
or (n8,n9,n99,n118);
and (n9,n10,n50);
or (n10,n11,n33,n49);
and (n11,n12,n18);
and (n12,n13,n14);
not (n14,n15);
and (n15,n16,n17);
xnor (n18,n19,n30);
nor (n19,n20,n28);
and (n20,n21,n22);
and (n22,n23,n26);
xor (n23,n24,n25);
not (n26,n27);
xor (n27,n25,n13);
and (n28,n29,n27);
and (n30,n24,n31);
not (n31,n32);
and (n32,n25,n13);
and (n33,n18,n34);
xnor (n34,n35,n46);
nor (n35,n36,n44);
and (n36,n37,n38);
and (n38,n39,n42);
xor (n39,n40,n41);
not (n42,n43);
xor (n43,n41,n24);
and (n44,n45,n43);
and (n46,n40,n47);
not (n47,n48);
and (n48,n41,n24);
and (n49,n12,n34);
or (n50,n51,n82,n98);
and (n51,n52,n67);
xnor (n52,n53,n64);
nor (n53,n54,n62);
and (n54,n55,n56);
and (n56,n57,n60);
xor (n57,n58,n59);
not (n60,n61);
xor (n61,n59,n40);
and (n62,n63,n61);
and (n64,n58,n65);
not (n65,n66);
and (n66,n59,n40);
xnor (n67,n68,n79);
nor (n68,n69,n77);
and (n69,n70,n71);
and (n71,n72,n75);
xor (n72,n73,n74);
not (n75,n76);
xor (n76,n74,n58);
and (n77,n78,n76);
and (n79,n73,n80);
not (n80,n81);
and (n81,n74,n58);
and (n82,n67,n83);
xnor (n83,n84,n95);
nor (n84,n85,n93);
and (n85,n86,n87);
and (n87,n88,n91);
xor (n88,n89,n90);
not (n91,n92);
xor (n92,n90,n73);
and (n93,n94,n92);
and (n95,n89,n96);
not (n96,n97);
and (n97,n90,n73);
and (n98,n52,n83);
and (n99,n50,n100);
or (n100,n101,n116);
xnor (n101,n102,n113);
nor (n102,n103,n111);
and (n103,n104,n105);
and (n105,n106,n109);
xor (n106,n107,n108);
not (n109,n110);
xor (n110,n108,n89);
and (n111,n112,n110);
and (n113,n107,n114);
not (n114,n115);
and (n115,n108,n89);
and (n116,n117,n107);
and (n118,n10,n100);
or (n119,n120,n145,n152);
and (n120,n121,n131);
xor (n121,n122,n127);
xor (n122,n123,n124);
not (n123,n12);
xnor (n124,n125,n30);
not (n125,n126);
and (n126,n29,n22);
xnor (n127,n128,n46);
nor (n128,n129,n130);
and (n129,n45,n38);
and (n130,n21,n43);
xor (n131,n132,n141);
xor (n132,n133,n137);
xnor (n133,n134,n64);
nor (n134,n135,n136);
and (n135,n63,n56);
and (n136,n37,n61);
xnor (n137,n138,n79);
nor (n138,n139,n140);
and (n139,n78,n71);
and (n140,n55,n76);
xnor (n141,n142,n95);
nor (n142,n143,n144);
and (n143,n94,n87);
and (n144,n70,n92);
and (n145,n131,n146);
xor (n146,n147,n151);
xnor (n147,n148,n113);
nor (n148,n149,n150);
and (n149,n112,n105);
and (n150,n86,n110);
and (n151,n104,n107);
and (n152,n121,n146);
and (n153,n119,n154);
xor (n154,n155,n168);
xor (n155,n156,n157);
and (n156,n112,n107);
xor (n157,n158,n164);
xor (n158,n159,n160);
not (n159,n30);
xnor (n160,n161,n46);
nor (n161,n162,n163);
and (n162,n21,n38);
and (n163,n29,n43);
xnor (n164,n165,n64);
nor (n165,n166,n167);
and (n166,n37,n56);
and (n167,n45,n61);
xor (n168,n169,n178);
xor (n169,n170,n174);
xnor (n170,n171,n79);
nor (n171,n172,n173);
and (n172,n55,n71);
and (n173,n63,n76);
xnor (n174,n175,n95);
nor (n175,n176,n177);
and (n176,n70,n87);
and (n177,n78,n92);
xnor (n178,n179,n113);
nor (n179,n180,n181);
and (n180,n86,n105);
and (n181,n94,n110);
and (n182,n8,n154);
xor (n183,n184,n156);
xor (n184,n185,n189);
or (n185,n186,n187,n188);
and (n186,n30,n160);
and (n187,n160,n164);
and (n188,n30,n164);
or (n189,n190,n191,n192);
and (n190,n170,n174);
and (n191,n174,n178);
and (n192,n170,n178);
and (n193,n183,n194);
xor (n194,n195,n215);
xor (n195,n196,n209);
or (n196,n197,n206,n208);
and (n197,n198,n202);
or (n198,n199,n200,n201);
and (n199,n123,n124);
and (n200,n124,n127);
and (n201,n123,n127);
or (n202,n203,n204,n205);
and (n203,n133,n137);
and (n204,n137,n141);
and (n205,n133,n141);
and (n206,n202,n207);
and (n207,n147,n151);
and (n208,n198,n207);
or (n209,n210,n212,n214);
and (n210,n211,n168);
not (n211,n157);
and (n212,n168,n213);
not (n213,n156);
and (n214,n211,n213);
xor (n215,n216,n232);
xor (n216,n217,n218);
and (n217,n86,n107);
xor (n218,n219,n228);
xor (n219,n220,n224);
xnor (n220,n221,n79);
nor (n221,n222,n223);
and (n222,n63,n71);
and (n223,n37,n76);
xnor (n224,n225,n95);
nor (n225,n226,n227);
and (n226,n78,n87);
and (n227,n55,n92);
xnor (n228,n229,n113);
nor (n229,n230,n231);
and (n230,n94,n105);
and (n231,n70,n110);
xor (n232,n233,n237);
xor (n233,n159,n234);
xnor (n234,n235,n46);
not (n235,n236);
and (n236,n29,n38);
xnor (n237,n238,n64);
nor (n238,n239,n240);
and (n239,n45,n56);
and (n240,n21,n61);
and (n241,n6,n194);
xor (n242,n243,n269);
xor (n243,n244,n248);
or (n244,n245,n246,n247);
and (n245,n196,n209);
and (n246,n209,n215);
and (n247,n196,n215);
xor (n248,n249,n258);
xor (n249,n250,n254);
or (n250,n251,n252,n253);
and (n251,n185,n189);
and (n252,n189,n156);
and (n253,n185,n156);
or (n254,n255,n256,n257);
and (n255,n217,n218);
and (n256,n218,n232);
and (n257,n217,n232);
xor (n258,n259,n268);
xor (n259,n260,n264);
xnor (n260,n261,n95);
nor (n261,n262,n263);
and (n262,n55,n87);
and (n263,n63,n92);
xnor (n264,n265,n113);
nor (n265,n266,n267);
and (n266,n70,n105);
and (n267,n78,n110);
and (n268,n94,n107);
xor (n269,n270,n282);
not (n270,n271);
xor (n271,n272,n278);
xor (n272,n273,n274);
not (n273,n46);
xnor (n274,n275,n64);
nor (n275,n276,n277);
and (n276,n21,n56);
and (n277,n29,n61);
xnor (n278,n279,n79);
nor (n279,n280,n281);
and (n280,n37,n71);
and (n281,n45,n76);
xnor (n282,n283,n287);
or (n283,n284,n285,n286);
and (n284,n220,n224);
and (n285,n224,n228);
and (n286,n220,n228);
or (n287,n288,n289,n290);
and (n288,n159,n234);
and (n289,n234,n237);
and (n290,n159,n237);
and (n291,n292,n367);
or (n292,n293,n363,n366);
and (n293,n294,n361);
or (n294,n295,n357,n360);
and (n295,n296,n346);
or (n296,n297,n328,n345);
and (n297,n298,n314);
or (n298,n299,n308,n313);
and (n299,n300,n301);
not (n300,n17);
xnor (n301,n302,n12);
not (n302,n303);
and (n303,n29,n304);
and (n304,n305,n306);
xor (n305,n13,n16);
not (n306,n307);
xor (n307,n16,n17);
and (n308,n301,n309);
xnor (n309,n310,n30);
nor (n310,n311,n312);
and (n311,n45,n22);
and (n312,n21,n27);
and (n313,n300,n309);
or (n314,n315,n324,n327);
and (n315,n316,n320);
xnor (n316,n317,n95);
nor (n317,n318,n319);
and (n318,n112,n87);
and (n319,n86,n92);
xnor (n320,n321,n113);
nor (n321,n322,n323);
and (n322,n117,n105);
and (n323,n104,n110);
and (n324,n320,n325);
and (n325,n326,n107);
and (n327,n316,n325);
and (n328,n314,n329);
or (n329,n330,n339,n344);
and (n330,n331,n335);
xnor (n331,n332,n46);
nor (n332,n333,n334);
and (n333,n63,n38);
and (n334,n37,n43);
xnor (n335,n336,n64);
nor (n336,n337,n338);
and (n337,n78,n56);
and (n338,n55,n61);
and (n339,n335,n340);
xnor (n340,n341,n79);
nor (n341,n342,n343);
and (n342,n94,n71);
and (n343,n70,n76);
and (n344,n331,n340);
and (n345,n298,n329);
or (n346,n347,n353,n356);
and (n347,n348,n351);
not (n348,n349);
xor (n349,n350,n34);
xor (n350,n123,n18);
xor (n351,n352,n83);
xor (n352,n52,n67);
and (n353,n351,n354);
not (n354,n355);
xor (n355,n101,n116);
and (n356,n348,n354);
and (n357,n346,n358);
xor (n358,n359,n146);
xor (n359,n121,n131);
and (n360,n296,n358);
xor (n361,n362,n207);
xor (n362,n198,n202);
and (n363,n361,n364);
xor (n364,n365,n154);
xor (n365,n8,n119);
and (n366,n294,n364);
xor (n367,n368,n194);
xor (n368,n6,n183);
or (n369,n370,n440);
and (n370,n371,n372);
xor (n371,n292,n367);
and (n372,n373,n438);
or (n373,n374,n434,n437);
and (n374,n375,n432);
or (n375,n376,n428,n431);
and (n376,n377,n423);
or (n377,n378,n407,n422);
and (n378,n379,n395);
or (n379,n380,n389,n394);
and (n380,n381,n385);
xnor (n381,n382,n46);
nor (n382,n383,n384);
and (n383,n55,n38);
and (n384,n63,n43);
xnor (n385,n386,n64);
nor (n386,n387,n388);
and (n387,n70,n56);
and (n388,n78,n61);
and (n389,n385,n390);
xnor (n390,n391,n79);
nor (n391,n392,n393);
and (n392,n86,n71);
and (n393,n94,n76);
and (n394,n381,n390);
or (n395,n396,n401,n406);
and (n396,n17,n397);
xnor (n397,n398,n12);
nor (n398,n399,n400);
and (n399,n21,n304);
and (n400,n29,n307);
and (n401,n397,n402);
xnor (n402,n403,n30);
nor (n403,n404,n405);
and (n404,n37,n22);
and (n405,n45,n27);
and (n406,n17,n402);
and (n407,n395,n408);
or (n408,n409,n418,n421);
and (n409,n410,n414);
xnor (n410,n411,n95);
nor (n411,n412,n413);
and (n412,n104,n87);
and (n413,n112,n92);
xnor (n414,n415,n113);
nor (n415,n416,n417);
and (n416,n326,n105);
and (n417,n117,n110);
and (n418,n414,n419);
and (n419,n420,n107);
and (n421,n410,n419);
and (n422,n379,n408);
or (n423,n424,n426);
xor (n424,n425,n325);
xor (n425,n316,n320);
xor (n426,n427,n340);
xor (n427,n331,n335);
and (n428,n423,n429);
xor (n429,n430,n355);
xor (n430,n349,n351);
and (n431,n377,n429);
xor (n432,n433,n100);
xor (n433,n10,n50);
and (n434,n432,n435);
xor (n435,n436,n358);
xor (n436,n296,n346);
and (n437,n375,n435);
xor (n438,n439,n364);
xor (n439,n294,n361);
and (n440,n441,n442);
xor (n441,n371,n372);
or (n442,n443,n523);
and (n443,n444,n445);
xor (n444,n373,n438);
and (n445,n446,n521);
or (n446,n447,n517,n520);
and (n447,n448,n513);
or (n448,n449,n509,n512);
and (n449,n450,n498);
or (n450,n451,n484,n497);
and (n451,n452,n468);
or (n452,n453,n462,n467);
and (n453,n454,n458);
xnor (n454,n455,n30);
nor (n455,n456,n457);
and (n456,n63,n22);
and (n457,n37,n27);
xnor (n458,n459,n46);
nor (n459,n460,n461);
and (n460,n78,n38);
and (n461,n55,n43);
and (n462,n458,n463);
xnor (n463,n464,n64);
nor (n464,n465,n466);
and (n465,n94,n56);
and (n466,n70,n61);
and (n467,n454,n463);
or (n468,n469,n478,n483);
and (n469,n470,n474);
xnor (n470,n471,n79);
nor (n471,n472,n473);
and (n472,n112,n71);
and (n473,n86,n76);
xnor (n474,n475,n95);
nor (n475,n476,n477);
and (n476,n117,n87);
and (n477,n104,n92);
and (n478,n474,n479);
xnor (n479,n480,n113);
nor (n480,n481,n482);
and (n481,n420,n105);
and (n482,n326,n110);
and (n483,n470,n479);
and (n484,n468,n485);
and (n485,n486,n493);
xnor (n486,n487,n17);
not (n487,n488);
and (n488,n29,n489);
and (n489,n490,n492);
xor (n490,n17,n491);
not (n492,n491);
xnor (n493,n494,n12);
nor (n494,n495,n496);
and (n495,n45,n304);
and (n496,n21,n307);
and (n497,n452,n485);
or (n498,n499,n505,n508);
and (n499,n500,n502);
xor (n500,n501,n390);
xor (n501,n381,n385);
not (n502,n503);
xor (n503,n504,n402);
xor (n504,n300,n397);
and (n505,n502,n506);
xor (n506,n507,n419);
xor (n507,n410,n414);
and (n508,n500,n506);
and (n509,n498,n510);
xor (n510,n511,n309);
xor (n511,n300,n301);
and (n512,n450,n510);
and (n513,n514,n516);
xor (n514,n515,n408);
xor (n515,n379,n395);
xnor (n516,n424,n426);
and (n517,n513,n518);
xor (n518,n519,n329);
xor (n519,n298,n314);
and (n520,n448,n518);
xor (n521,n522,n435);
xor (n522,n375,n432);
and (n523,n524,n525);
xor (n524,n444,n445);
or (n525,n526,n605);
and (n526,n527,n528);
xor (n527,n446,n521);
or (n528,n529,n601,n604);
and (n529,n530,n599);
or (n530,n531,n596,n598);
and (n531,n532,n594);
or (n532,n533,n590,n593);
and (n533,n534,n580);
or (n534,n535,n568,n579);
and (n535,n536,n552);
or (n536,n537,n546,n551);
and (n537,n538,n542);
xnor (n538,n539,n17);
nor (n539,n540,n541);
and (n540,n21,n489);
and (n541,n29,n491);
xnor (n542,n543,n12);
nor (n543,n544,n545);
and (n544,n37,n304);
and (n545,n45,n307);
and (n546,n542,n547);
xnor (n547,n548,n30);
nor (n548,n549,n550);
and (n549,n55,n22);
and (n550,n63,n27);
and (n551,n538,n547);
or (n552,n553,n562,n567);
and (n553,n554,n558);
xnor (n554,n555,n46);
nor (n555,n556,n557);
and (n556,n70,n38);
and (n557,n78,n43);
xnor (n558,n559,n64);
nor (n559,n560,n561);
and (n560,n86,n56);
and (n561,n94,n61);
and (n562,n558,n563);
xnor (n563,n564,n79);
nor (n564,n565,n566);
and (n565,n104,n71);
and (n566,n112,n76);
and (n567,n554,n563);
and (n568,n552,n569);
and (n569,n570,n574);
xnor (n570,n571,n95);
nor (n571,n572,n573);
and (n572,n326,n87);
and (n573,n117,n92);
xnor (n574,n575,n113);
nor (n575,n576,n578);
and (n576,n577,n105);
and (n578,n420,n110);
and (n579,n536,n569);
or (n580,n581,n586,n589);
and (n581,n582,n584);
not (n582,n583);
nand (n583,n577,n107);
xor (n584,n585,n463);
xor (n585,n454,n458);
and (n586,n584,n587);
xor (n587,n588,n479);
xor (n588,n470,n474);
and (n589,n582,n587);
and (n590,n580,n591);
xor (n591,n592,n506);
xor (n592,n500,n502);
and (n593,n534,n591);
xor (n594,n595,n510);
xor (n595,n450,n498);
and (n596,n594,n597);
xor (n597,n514,n516);
and (n598,n532,n597);
xor (n599,n600,n518);
xor (n600,n448,n513);
and (n601,n599,n602);
xor (n602,n603,n429);
xor (n603,n377,n423);
and (n604,n530,n602);
and (n605,n606,n607);
xor (n606,n527,n528);
or (n607,n608,n685);
and (n608,n609,n611);
xor (n609,n610,n602);
xor (n610,n530,n599);
and (n611,n612,n683);
or (n612,n613,n679,n682);
and (n613,n614,n674);
or (n614,n615,n671,n673);
and (n615,n616,n662);
or (n616,n617,n644,n661);
and (n617,n618,n632);
or (n618,n619,n628,n631);
and (n619,n620,n624);
xnor (n620,n621,n79);
nor (n621,n622,n623);
and (n622,n117,n71);
and (n623,n104,n76);
xnor (n624,n625,n95);
nor (n625,n626,n627);
and (n626,n420,n87);
and (n627,n326,n92);
and (n628,n624,n629);
xnor (n629,n630,n113);
nand (n630,n577,n110);
and (n631,n620,n629);
or (n632,n633,n642,n643);
and (n633,n634,n638);
xnor (n634,n635,n17);
nor (n635,n636,n637);
and (n636,n45,n489);
and (n637,n21,n491);
xnor (n638,n639,n12);
nor (n639,n640,n641);
and (n640,n63,n304);
and (n641,n37,n307);
and (n642,n638,n113);
and (n643,n634,n113);
and (n644,n632,n645);
or (n645,n646,n655,n660);
and (n646,n647,n651);
xnor (n647,n648,n30);
nor (n648,n649,n650);
and (n649,n78,n22);
and (n650,n55,n27);
xnor (n651,n652,n46);
nor (n652,n653,n654);
and (n653,n94,n38);
and (n654,n70,n43);
and (n655,n651,n656);
xnor (n656,n657,n64);
nor (n657,n658,n659);
and (n658,n112,n56);
and (n659,n86,n61);
and (n660,n647,n656);
and (n661,n618,n645);
or (n662,n663,n668,n670);
and (n663,n664,n666);
xor (n664,n665,n547);
xor (n665,n538,n542);
xor (n666,n667,n563);
xor (n667,n554,n558);
and (n668,n666,n669);
xor (n669,n570,n574);
and (n670,n664,n669);
and (n671,n662,n672);
xor (n672,n486,n493);
and (n673,n616,n672);
and (n674,n675,n677);
xor (n675,n676,n569);
xor (n676,n536,n552);
xor (n677,n678,n587);
xor (n678,n582,n584);
and (n679,n674,n680);
xor (n680,n681,n485);
xor (n681,n452,n468);
and (n682,n614,n680);
xor (n683,n684,n597);
xor (n684,n532,n594);
and (n685,n686,n687);
xor (n686,n609,n611);
or (n687,n688,n695);
and (n688,n689,n690);
xor (n689,n612,n683);
and (n690,n691,n693);
xor (n691,n692,n680);
xor (n692,n614,n674);
xor (n693,n694,n591);
xor (n694,n534,n580);
and (n695,n696,n728);
xor (n696,n697,n722);
xor (n697,n698,n702);
or (n698,n613,n699,n701);
and (n699,n674,n700);
xnor (n700,n500,n506);
and (n701,n614,n700);
xor (n702,n703,n712);
xor (n703,n704,n707);
or (n704,n533,n705,n706);
and (n705,n580,n503);
and (n706,n534,n503);
xor (n707,n708,n408);
xor (n708,n379,n709);
or (n709,n710,n401,n711);
and (n710,n300,n397);
and (n711,n300,n402);
xor (n712,n713,n715);
xor (n713,n450,n714);
or (n714,n500,n506);
xor (n715,n716,n721);
xor (n716,n717,n719);
xor (n717,n718,n331);
xor (n718,n301,n309);
xor (n719,n720,n316);
xor (n720,n335,n340);
xnor (n721,n320,n325);
or (n722,n723,n725,n727);
and (n723,n680,n724);
xor (n724,n694,n503);
and (n725,n724,n726);
xor (n726,n692,n700);
and (n727,n680,n726);
or (n728,n729,n788);
and (n729,n730,n732);
xor (n730,n731,n726);
xor (n731,n680,n724);
or (n732,n733,n785,n787);
and (n733,n734,n783);
or (n734,n735,n779,n782);
and (n735,n736,n774);
or (n736,n737,n770,n773);
and (n737,n738,n754);
or (n738,n739,n748,n753);
and (n739,n740,n744);
xnor (n740,n741,n17);
nor (n741,n742,n743);
and (n742,n37,n489);
and (n743,n45,n491);
xnor (n744,n745,n12);
nor (n745,n746,n747);
and (n746,n55,n304);
and (n747,n63,n307);
and (n748,n744,n749);
xnor (n749,n750,n30);
nor (n750,n751,n752);
and (n751,n70,n22);
and (n752,n78,n27);
and (n753,n740,n749);
or (n754,n755,n764,n769);
and (n755,n756,n760);
xnor (n756,n757,n46);
nor (n757,n758,n759);
and (n758,n86,n38);
and (n759,n94,n43);
xnor (n760,n761,n64);
nor (n761,n762,n763);
and (n762,n104,n56);
and (n763,n112,n61);
and (n764,n760,n765);
xnor (n765,n766,n79);
nor (n766,n767,n768);
and (n767,n326,n71);
and (n768,n117,n76);
and (n769,n756,n765);
and (n770,n754,n771);
xor (n771,n772,n629);
xor (n772,n620,n624);
and (n773,n738,n771);
and (n774,n775,n777);
xor (n775,n776,n113);
xor (n776,n634,n638);
xor (n777,n778,n656);
xor (n778,n647,n651);
and (n779,n774,n780);
xor (n780,n781,n669);
xor (n781,n664,n666);
and (n782,n736,n780);
xor (n783,n784,n672);
xor (n784,n616,n662);
and (n785,n783,n786);
xor (n786,n675,n677);
and (n787,n734,n786);
and (n788,n789,n790);
xor (n789,n730,n732);
or (n790,n791,n845);
and (n791,n792,n794);
xor (n792,n793,n786);
xor (n793,n734,n783);
or (n794,n795,n841,n844);
and (n795,n796,n839);
or (n796,n797,n836,n838);
and (n797,n798,n834);
or (n798,n799,n828,n833);
and (n799,n800,n812);
or (n800,n801,n810,n811);
and (n801,n802,n806);
xnor (n802,n803,n17);
nor (n803,n804,n805);
and (n804,n63,n489);
and (n805,n37,n491);
xnor (n806,n807,n12);
nor (n807,n808,n809);
and (n808,n78,n304);
and (n809,n55,n307);
and (n810,n806,n95);
and (n811,n802,n95);
or (n812,n813,n822,n827);
and (n813,n814,n818);
xnor (n814,n815,n30);
nor (n815,n816,n817);
and (n816,n94,n22);
and (n817,n70,n27);
xnor (n818,n819,n46);
nor (n819,n820,n821);
and (n820,n112,n38);
and (n821,n86,n43);
and (n822,n818,n823);
xnor (n823,n824,n64);
nor (n824,n825,n826);
and (n825,n117,n56);
and (n826,n104,n61);
and (n827,n814,n823);
and (n828,n812,n829);
xnor (n829,n830,n95);
nor (n830,n831,n832);
and (n831,n577,n87);
and (n832,n420,n92);
and (n833,n800,n829);
xor (n834,n835,n771);
xor (n835,n738,n754);
and (n836,n834,n837);
xor (n837,n775,n777);
and (n838,n798,n837);
xor (n839,n840,n645);
xor (n840,n618,n632);
and (n841,n839,n842);
xor (n842,n843,n780);
xor (n843,n736,n774);
and (n844,n796,n842);
and (n845,n846,n847);
xor (n846,n792,n794);
or (n847,n848,n918);
and (n848,n849,n851);
xor (n849,n850,n842);
xor (n850,n796,n839);
or (n851,n852,n914,n917);
and (n852,n853,n909);
or (n853,n854,n905,n908);
and (n854,n855,n895);
or (n855,n856,n889,n894);
and (n856,n857,n873);
or (n857,n858,n867,n872);
and (n858,n859,n863);
xnor (n859,n860,n46);
nor (n860,n861,n862);
and (n861,n104,n38);
and (n862,n112,n43);
xnor (n863,n864,n64);
nor (n864,n865,n866);
and (n865,n326,n56);
and (n866,n117,n61);
and (n867,n863,n868);
xnor (n868,n869,n79);
nor (n869,n870,n871);
and (n870,n577,n71);
and (n871,n420,n76);
and (n872,n859,n868);
or (n873,n874,n883,n888);
and (n874,n875,n879);
xnor (n875,n876,n17);
nor (n876,n877,n878);
and (n877,n55,n489);
and (n878,n63,n491);
xnor (n879,n880,n12);
nor (n880,n881,n882);
and (n881,n70,n304);
and (n882,n78,n307);
and (n883,n879,n884);
xnor (n884,n885,n30);
nor (n885,n886,n887);
and (n886,n86,n22);
and (n887,n94,n27);
and (n888,n875,n884);
and (n889,n873,n890);
xnor (n890,n891,n79);
nor (n891,n892,n893);
and (n892,n420,n71);
and (n893,n326,n76);
and (n894,n857,n890);
or (n895,n896,n901,n904);
and (n896,n897,n899);
xnor (n897,n898,n95);
nand (n898,n577,n92);
xor (n899,n900,n95);
xor (n900,n802,n806);
and (n901,n899,n902);
xor (n902,n903,n823);
xor (n903,n814,n818);
and (n904,n897,n902);
and (n905,n895,n906);
xor (n906,n907,n765);
xor (n907,n756,n760);
and (n908,n855,n906);
and (n909,n910,n912);
xor (n910,n911,n749);
xor (n911,n740,n744);
xor (n912,n913,n829);
xor (n913,n800,n812);
and (n914,n909,n915);
xor (n915,n916,n837);
xor (n916,n798,n834);
and (n917,n853,n915);
and (n918,n919,n920);
xor (n919,n849,n851);
or (n920,n921,n973);
and (n921,n922,n924);
xor (n922,n923,n915);
xor (n923,n853,n909);
or (n924,n925,n970,n972);
and (n925,n926,n968);
or (n926,n927,n964,n967);
and (n927,n928,n962);
or (n928,n929,n958,n961);
and (n929,n930,n946);
or (n930,n931,n940,n945);
and (n931,n932,n936);
xnor (n932,n933,n30);
nor (n933,n934,n935);
and (n934,n112,n22);
and (n935,n86,n27);
xnor (n936,n937,n46);
nor (n937,n938,n939);
and (n938,n117,n38);
and (n939,n104,n43);
and (n940,n936,n941);
xnor (n941,n942,n64);
nor (n942,n943,n944);
and (n943,n420,n56);
and (n944,n326,n61);
and (n945,n932,n941);
or (n946,n947,n956,n957);
and (n947,n948,n952);
xnor (n948,n949,n17);
nor (n949,n950,n951);
and (n950,n78,n489);
and (n951,n55,n491);
xnor (n952,n953,n12);
nor (n953,n954,n955);
and (n954,n94,n304);
and (n955,n70,n307);
and (n956,n952,n79);
and (n957,n948,n79);
and (n958,n946,n959);
xor (n959,n960,n868);
xor (n960,n859,n863);
and (n961,n930,n959);
xor (n962,n963,n890);
xor (n963,n857,n873);
and (n964,n962,n965);
xor (n965,n966,n902);
xor (n966,n897,n899);
and (n967,n928,n965);
xor (n968,n969,n906);
xor (n969,n855,n895);
and (n970,n968,n971);
xor (n971,n910,n912);
and (n972,n926,n971);
and (n973,n974,n975);
xor (n974,n922,n924);
or (n975,n976,n1014);
and (n976,n977,n979);
xor (n977,n978,n971);
xor (n978,n926,n968);
and (n979,n980,n1012);
or (n980,n981,n1008,n1011);
and (n981,n982,n1006);
or (n982,n983,n1002,n1005);
and (n983,n984,n1000);
or (n984,n985,n994,n999);
and (n985,n986,n990);
xnor (n986,n987,n17);
nor (n987,n988,n989);
and (n988,n70,n489);
and (n989,n78,n491);
xnor (n990,n991,n12);
nor (n991,n992,n993);
and (n992,n86,n304);
and (n993,n94,n307);
and (n994,n990,n995);
xnor (n995,n996,n30);
nor (n996,n997,n998);
and (n997,n104,n22);
and (n998,n112,n27);
and (n999,n986,n995);
xnor (n1000,n1001,n79);
nand (n1001,n577,n76);
and (n1002,n1000,n1003);
xor (n1003,n1004,n941);
xor (n1004,n932,n936);
and (n1005,n984,n1003);
xor (n1006,n1007,n884);
xor (n1007,n875,n879);
and (n1008,n1006,n1009);
xor (n1009,n1010,n959);
xor (n1010,n930,n946);
and (n1011,n982,n1009);
xor (n1012,n1013,n965);
xor (n1013,n928,n962);
and (n1014,n1015,n1016);
xor (n1015,n977,n979);
or (n1016,n1017,n1069);
and (n1017,n1018,n1019);
xor (n1018,n980,n1012);
and (n1019,n1020,n1067);
or (n1020,n1021,n1063,n1066);
and (n1021,n1022,n1056);
or (n1022,n1023,n1050,n1055);
and (n1023,n1024,n1038);
or (n1024,n1025,n1034,n1037);
and (n1025,n1026,n1030);
xnor (n1026,n1027,n30);
nor (n1027,n1028,n1029);
and (n1028,n117,n22);
and (n1029,n104,n27);
xnor (n1030,n1031,n46);
nor (n1031,n1032,n1033);
and (n1032,n420,n38);
and (n1033,n326,n43);
and (n1034,n1030,n1035);
xnor (n1035,n1036,n64);
nand (n1036,n577,n61);
and (n1037,n1026,n1035);
or (n1038,n1039,n1048,n1049);
and (n1039,n1040,n1044);
xnor (n1040,n1041,n17);
nor (n1041,n1042,n1043);
and (n1042,n94,n489);
and (n1043,n70,n491);
xnor (n1044,n1045,n12);
nor (n1045,n1046,n1047);
and (n1046,n112,n304);
and (n1047,n86,n307);
and (n1048,n1044,n64);
and (n1049,n1040,n64);
and (n1050,n1038,n1051);
xnor (n1051,n1052,n46);
nor (n1052,n1053,n1054);
and (n1053,n326,n38);
and (n1054,n117,n43);
and (n1055,n1024,n1051);
and (n1056,n1057,n1061);
xnor (n1057,n1058,n64);
nor (n1058,n1059,n1060);
and (n1059,n577,n56);
and (n1060,n420,n61);
xor (n1061,n1062,n995);
xor (n1062,n986,n990);
and (n1063,n1056,n1064);
xor (n1064,n1065,n79);
xor (n1065,n948,n952);
and (n1066,n1022,n1064);
xor (n1067,n1068,n1009);
xor (n1068,n982,n1006);
and (n1069,n1070,n1071);
xor (n1070,n1018,n1019);
or (n1071,n1072,n1079);
and (n1072,n1073,n1074);
xor (n1073,n1020,n1067);
and (n1074,n1075,n1077);
xor (n1075,n1076,n1003);
xor (n1076,n984,n1000);
xor (n1077,n1078,n1064);
xor (n1078,n1022,n1056);
and (n1079,n1080,n1081);
xor (n1080,n1073,n1074);
or (n1081,n1082,n1115);
and (n1082,n1083,n1084);
xor (n1083,n1075,n1077);
or (n1084,n1085,n1112,n1114);
and (n1085,n1086,n1110);
or (n1086,n1087,n1106,n1109);
and (n1087,n1088,n1104);
or (n1088,n1089,n1098,n1103);
and (n1089,n1090,n1094);
xnor (n1090,n1091,n17);
nor (n1091,n1092,n1093);
and (n1092,n86,n489);
and (n1093,n94,n491);
xnor (n1094,n1095,n12);
nor (n1095,n1096,n1097);
and (n1096,n104,n304);
and (n1097,n112,n307);
and (n1098,n1094,n1099);
xnor (n1099,n1100,n30);
nor (n1100,n1101,n1102);
and (n1101,n326,n22);
and (n1102,n117,n27);
and (n1103,n1090,n1099);
xor (n1104,n1105,n1035);
xor (n1105,n1026,n1030);
and (n1106,n1104,n1107);
xor (n1107,n1108,n64);
xor (n1108,n1040,n1044);
and (n1109,n1088,n1107);
xor (n1110,n1111,n1051);
xor (n1111,n1024,n1038);
and (n1112,n1110,n1113);
xor (n1113,n1057,n1061);
and (n1114,n1086,n1113);
and (n1115,n1116,n1117);
xor (n1116,n1083,n1084);
or (n1117,n1118,n1151);
and (n1118,n1119,n1121);
xor (n1119,n1120,n1113);
xor (n1120,n1086,n1110);
and (n1121,n1122,n1149);
or (n1122,n1123,n1143,n1148);
and (n1123,n1124,n1136);
or (n1124,n1125,n1134,n1135);
and (n1125,n1126,n1130);
xnor (n1126,n1127,n17);
nor (n1127,n1128,n1129);
and (n1128,n112,n489);
and (n1129,n86,n491);
xnor (n1130,n1131,n12);
nor (n1131,n1132,n1133);
and (n1132,n117,n304);
and (n1133,n104,n307);
and (n1134,n1130,n46);
and (n1135,n1126,n46);
and (n1136,n1137,n1141);
xnor (n1137,n1138,n30);
nor (n1138,n1139,n1140);
and (n1139,n420,n22);
and (n1140,n326,n27);
xnor (n1141,n1142,n46);
nand (n1142,n577,n43);
and (n1143,n1136,n1144);
xnor (n1144,n1145,n46);
nor (n1145,n1146,n1147);
and (n1146,n577,n38);
and (n1147,n420,n43);
and (n1148,n1124,n1144);
xor (n1149,n1150,n1107);
xor (n1150,n1088,n1104);
and (n1151,n1152,n1153);
xor (n1152,n1119,n1121);
or (n1153,n1154,n1161);
and (n1154,n1155,n1156);
xor (n1155,n1122,n1149);
and (n1156,n1157,n1159);
xor (n1157,n1158,n1099);
xor (n1158,n1090,n1094);
xor (n1159,n1160,n1144);
xor (n1160,n1124,n1136);
and (n1161,n1162,n1163);
xor (n1162,n1155,n1156);
or (n1163,n1164,n1189);
and (n1164,n1165,n1166);
xor (n1165,n1157,n1159);
or (n1166,n1167,n1186,n1188);
and (n1167,n1168,n1184);
or (n1168,n1169,n1178,n1183);
and (n1169,n1170,n1174);
xnor (n1170,n1171,n17);
nor (n1171,n1172,n1173);
and (n1172,n104,n489);
and (n1173,n112,n491);
xnor (n1174,n1175,n12);
nor (n1175,n1176,n1177);
and (n1176,n326,n304);
and (n1177,n117,n307);
and (n1178,n1174,n1179);
xnor (n1179,n1180,n30);
nor (n1180,n1181,n1182);
and (n1181,n577,n22);
and (n1182,n420,n27);
and (n1183,n1170,n1179);
xor (n1184,n1185,n46);
xor (n1185,n1126,n1130);
and (n1186,n1184,n1187);
xor (n1187,n1137,n1141);
and (n1188,n1168,n1187);
and (n1189,n1190,n1191);
xor (n1190,n1165,n1166);
or (n1191,n1192,n1210);
and (n1192,n1193,n1195);
xor (n1193,n1194,n1187);
xor (n1194,n1168,n1184);
and (n1195,n1196,n1208);
or (n1196,n1197,n1206,n1207);
and (n1197,n1198,n1202);
xnor (n1198,n1199,n17);
nor (n1199,n1200,n1201);
and (n1200,n117,n489);
and (n1201,n104,n491);
xnor (n1202,n1203,n12);
nor (n1203,n1204,n1205);
and (n1204,n420,n304);
and (n1205,n326,n307);
and (n1206,n1202,n30);
and (n1207,n1198,n30);
xor (n1208,n1209,n1179);
xor (n1209,n1170,n1174);
and (n1210,n1211,n1212);
xor (n1211,n1193,n1195);
or (n1212,n1213,n1220);
and (n1213,n1214,n1215);
xor (n1214,n1196,n1208);
and (n1215,n1216,n1218);
xnor (n1216,n1217,n30);
nand (n1217,n577,n27);
xor (n1218,n1219,n30);
xor (n1219,n1198,n1202);
and (n1220,n1221,n1222);
xor (n1221,n1214,n1215);
or (n1222,n1223,n1234);
and (n1223,n1224,n1225);
xor (n1224,n1216,n1218);
and (n1225,n1226,n1230);
xnor (n1226,n1227,n17);
nor (n1227,n1228,n1229);
and (n1228,n326,n489);
and (n1229,n117,n491);
xnor (n1230,n1231,n12);
nor (n1231,n1232,n1233);
and (n1232,n577,n304);
and (n1233,n420,n307);
and (n1234,n1235,n1236);
xor (n1235,n1224,n1225);
or (n1236,n1237,n1244);
and (n1237,n1238,n1239);
xor (n1238,n1226,n1230);
and (n1239,n1240,n12);
xnor (n1240,n1241,n17);
nor (n1241,n1242,n1243);
and (n1242,n420,n489);
and (n1243,n326,n491);
and (n1244,n1245,n1246);
xor (n1245,n1238,n1239);
or (n1246,n1247,n1251);
and (n1247,n1248,n1250);
xnor (n1248,n1249,n12);
nand (n1249,n577,n307);
xor (n1250,n1240,n12);
and (n1251,n1252,n1253);
xor (n1252,n1248,n1250);
and (n1253,n1254,n1258);
xnor (n1254,n1255,n17);
nor (n1255,n1256,n1257);
and (n1256,n577,n489);
and (n1257,n420,n491);
and (n1258,n1259,n17);
xnor (n1259,n1260,n17);
nand (n1260,n577,n491);
buf (n1261,n1262);
xor (n1262,n1263,n1366);
xor (n1263,n1264,n1334);
xor (n1264,n1265,n1316);
or (n1265,n1266,n1307,n1315);
and (n1266,n1267,n1288);
or (n1267,n1268,n1286,n1287);
and (n1268,n1269,n1277);
or (n1269,n1270,n1274,n1276);
and (n1270,n1271,n50);
or (n1271,n1272,n33,n1273);
and (n1272,n123,n18);
and (n1273,n123,n34);
and (n1274,n50,n1275);
and (n1275,n101,n116);
and (n1276,n1271,n1275);
or (n1277,n1278,n1283,n1285);
and (n1278,n1279,n1281);
xor (n1279,n1280,n133);
xor (n1280,n124,n127);
xor (n1281,n1282,n147);
xor (n1282,n137,n141);
and (n1283,n1281,n1284);
not (n1284,n151);
and (n1285,n1279,n1284);
and (n1286,n1277,n154);
and (n1287,n1269,n154);
xor (n1288,n1289,n1305);
xor (n1289,n1290,n1301);
or (n1290,n1291,n1298,n1300);
and (n1291,n1292,n1295);
or (n1292,n200,n1293,n1294);
and (n1293,n127,n133);
and (n1294,n124,n133);
or (n1295,n204,n1296,n1297);
and (n1296,n141,n147);
and (n1297,n137,n147);
and (n1298,n1295,n1299);
buf (n1299,n151);
and (n1300,n1292,n1299);
or (n1301,n1302,n1303,n1304);
and (n1302,n156,n157);
and (n1303,n157,n168);
and (n1304,n156,n168);
xor (n1305,n1306,n217);
xor (n1306,n224,n228);
and (n1307,n1288,n1308);
xor (n1308,n1309,n1311);
xor (n1309,n1310,n220);
xor (n1310,n234,n237);
xnor (n1311,n1312,n189);
or (n1312,n1313,n187,n1314);
and (n1313,n159,n160);
and (n1314,n159,n164);
and (n1315,n1267,n1308);
xor (n1316,n1317,n1323);
xor (n1317,n1318,n1322);
or (n1318,n1319,n1320,n1321);
and (n1319,n1290,n1301);
and (n1320,n1301,n1305);
and (n1321,n1290,n1305);
and (n1322,n1309,n1311);
xor (n1323,n1324,n1326);
xor (n1324,n1325,n271);
or (n1325,n1312,n189);
xor (n1326,n1327,n258);
xor (n1327,n1328,n1331);
or (n1328,n285,n1329,n1330);
and (n1329,n228,n217);
and (n1330,n224,n217);
or (n1331,n289,n1332,n1333);
and (n1332,n237,n220);
and (n1333,n234,n220);
and (n1334,n1335,n1364);
or (n1335,n1336,n1360,n1363);
and (n1336,n1337,n1358);
or (n1337,n1338,n1354,n1357);
and (n1338,n1339,n1350);
or (n1339,n1340,n1347,n1349);
and (n1340,n1341,n1344);
or (n1341,n308,n1342,n1343);
and (n1342,n309,n331);
and (n1343,n301,n331);
or (n1344,n339,n1345,n1346);
and (n1345,n340,n316);
and (n1346,n335,n316);
and (n1347,n1344,n1348);
or (n1348,n320,n325);
and (n1349,n1341,n1348);
or (n1350,n1351,n1352,n1353);
and (n1351,n349,n351);
and (n1352,n351,n355);
and (n1353,n349,n355);
and (n1354,n1350,n1355);
xor (n1355,n1356,n1284);
xor (n1356,n1279,n1281);
and (n1357,n1339,n1355);
xor (n1358,n1359,n1299);
xor (n1359,n1292,n1295);
and (n1360,n1358,n1361);
xor (n1361,n1362,n154);
xor (n1362,n1269,n1277);
and (n1363,n1337,n1361);
xor (n1364,n1365,n1308);
xor (n1365,n1267,n1288);
or (n1366,n1367,n1391);
and (n1367,n1368,n1369);
xor (n1368,n1335,n1364);
and (n1369,n1370,n1389);
or (n1370,n1371,n1385,n1388);
and (n1371,n1372,n1383);
or (n1372,n1373,n1381,n1382);
and (n1373,n1374,n1377);
or (n1374,n1375,n1376,n422);
and (n1375,n379,n709);
and (n1376,n709,n408);
or (n1377,n1378,n1379,n1380);
and (n1378,n717,n719);
and (n1379,n719,n721);
and (n1380,n717,n721);
and (n1381,n1377,n429);
and (n1382,n1374,n429);
xor (n1383,n1384,n1275);
xor (n1384,n1271,n50);
and (n1385,n1383,n1386);
xor (n1386,n1387,n1355);
xor (n1387,n1339,n1350);
and (n1388,n1372,n1386);
xor (n1389,n1390,n1361);
xor (n1390,n1337,n1358);
and (n1391,n1392,n1393);
xor (n1392,n1368,n1369);
or (n1393,n1394,n1411);
and (n1394,n1395,n1396);
xor (n1395,n1370,n1389);
and (n1396,n1397,n1409);
or (n1397,n1398,n1405,n1408);
and (n1398,n1399,n1403);
or (n1399,n1400,n1401,n1402);
and (n1400,n450,n714);
and (n1401,n714,n715);
and (n1402,n450,n715);
xor (n1403,n1404,n1348);
xor (n1404,n1341,n1344);
and (n1405,n1403,n1406);
xor (n1406,n1407,n429);
xor (n1407,n1374,n1377);
and (n1408,n1399,n1406);
xor (n1409,n1410,n1386);
xor (n1410,n1372,n1383);
and (n1411,n1412,n1413);
xor (n1412,n1395,n1396);
or (n1413,n1414,n1423);
and (n1414,n1415,n1416);
xor (n1415,n1397,n1409);
and (n1416,n1417,n1421);
or (n1417,n1418,n1419,n1420);
and (n1418,n704,n707);
and (n1419,n707,n712);
and (n1420,n704,n712);
xor (n1421,n1422,n1406);
xor (n1422,n1399,n1403);
and (n1423,n1424,n1425);
xor (n1424,n1415,n1416);
or (n1425,n1426,n1429);
and (n1426,n1427,n1428);
xor (n1427,n1417,n1421);
and (n1428,n698,n702);
and (n1429,n1430,n1431);
xor (n1430,n1427,n1428);
or (n1431,n1432,n695);
and (n1432,n697,n722);
endmodule
