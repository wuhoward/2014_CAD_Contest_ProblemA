module top (out,n13,n17,n20,n21,n31,n34,n35,n39,n49
        ,n52,n53,n56,n58,n65,n68,n69,n73,n79,n87
        ,n90,n91,n95,n102,n105,n106,n110,n118,n121,n125
        ,n363,n432,n518);
output out;
input n13;
input n17;
input n20;
input n21;
input n31;
input n34;
input n35;
input n39;
input n49;
input n52;
input n53;
input n56;
input n58;
input n65;
input n68;
input n69;
input n73;
input n79;
input n87;
input n90;
input n91;
input n95;
input n102;
input n105;
input n106;
input n110;
input n118;
input n121;
input n125;
input n363;
input n432;
input n518;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n16;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n51;
wire n54;
wire n55;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
xor (out,n0,n1202);
buf (n0,n1);
xor (n1,n2,n383);
xor (n2,n3,n315);
xor (n3,n4,n261);
or (n4,n5,n212,n260);
and (n5,n6,n201);
or (n6,n7,n168,n200);
and (n7,n8,n131);
or (n8,n9,n81,n130);
and (n9,n10,n44);
or (n10,n11,n27,n43);
and (n11,n12,n14);
not (n12,n13);
xnor (n14,n15,n24);
not (n15,n16);
and (n16,n17,n18);
and (n18,n19,n22);
xor (n19,n20,n21);
not (n22,n23);
xor (n23,n21,n13);
and (n24,n20,n25);
not (n25,n26);
and (n26,n21,n13);
and (n27,n14,n28);
xnor (n28,n29,n40);
nor (n29,n30,n38);
and (n30,n31,n32);
and (n32,n33,n36);
xor (n33,n34,n35);
not (n36,n37);
xor (n37,n35,n20);
and (n38,n39,n37);
and (n40,n34,n41);
not (n41,n42);
and (n42,n35,n20);
and (n43,n12,n28);
or (n44,n45,n77,n80);
and (n45,n46,n62);
xnor (n46,n47,n59);
nor (n47,n48,n57);
and (n48,n49,n50);
and (n50,n51,n54);
xor (n51,n52,n53);
not (n54,n55);
xor (n55,n53,n56);
and (n57,n58,n55);
and (n59,n52,n60);
not (n60,n61);
and (n61,n53,n56);
xnor (n62,n63,n74);
nor (n63,n64,n72);
and (n64,n65,n66);
and (n66,n67,n70);
xor (n67,n68,n69);
not (n70,n71);
xor (n71,n69,n52);
and (n72,n73,n71);
and (n74,n68,n75);
not (n75,n76);
and (n76,n69,n52);
and (n77,n62,n78);
and (n78,n79,n68);
and (n80,n46,n78);
and (n81,n44,n82);
or (n82,n83,n114,n129);
and (n83,n84,n99);
xnor (n84,n85,n96);
nor (n85,n86,n94);
and (n86,n87,n88);
and (n88,n89,n92);
xor (n89,n90,n91);
not (n92,n93);
xor (n93,n91,n34);
and (n94,n95,n93);
and (n96,n90,n97);
not (n97,n98);
and (n98,n91,n34);
xnor (n99,n100,n111);
nor (n100,n101,n109);
and (n101,n102,n103);
and (n103,n104,n107);
xor (n104,n105,n106);
not (n107,n108);
xor (n108,n106,n90);
and (n109,n110,n108);
and (n111,n105,n112);
not (n112,n113);
and (n113,n106,n90);
and (n114,n99,n115);
xnor (n115,n116,n126);
nor (n116,n117,n124);
and (n117,n118,n119);
and (n119,n120,n122);
xor (n120,n56,n121);
not (n122,n123);
xor (n123,n121,n105);
and (n124,n125,n123);
and (n126,n56,n127);
not (n127,n128);
and (n128,n121,n105);
and (n129,n84,n115);
and (n130,n10,n82);
or (n131,n132,n159,n167);
and (n132,n133,n145);
not (n133,n134);
xor (n134,n135,n141);
xor (n135,n136,n137);
not (n136,n24);
xnor (n137,n138,n40);
nor (n138,n139,n140);
and (n139,n39,n32);
and (n140,n17,n37);
xnor (n141,n142,n96);
nor (n142,n143,n144);
and (n143,n95,n88);
and (n144,n31,n93);
xor (n145,n146,n155);
xor (n146,n147,n151);
xnor (n147,n148,n111);
nor (n148,n149,n150);
and (n149,n110,n103);
and (n150,n87,n108);
xnor (n151,n152,n126);
nor (n152,n153,n154);
and (n153,n125,n119);
and (n154,n102,n123);
xnor (n155,n156,n59);
nor (n156,n157,n158);
and (n157,n58,n50);
and (n158,n118,n55);
and (n159,n145,n160);
not (n160,n161);
xor (n161,n162,n166);
xnor (n162,n163,n74);
nor (n163,n164,n165);
and (n164,n73,n66);
and (n165,n49,n71);
and (n166,n65,n68);
and (n167,n133,n160);
and (n168,n131,n169);
xor (n169,n170,n194);
xor (n170,n171,n180);
xor (n171,n172,n176);
xor (n172,n136,n173);
xnor (n173,n174,n40);
not (n174,n175);
and (n175,n17,n32);
xnor (n176,n177,n96);
nor (n177,n178,n179);
and (n178,n31,n88);
and (n179,n39,n93);
xor (n180,n181,n190);
xor (n181,n182,n186);
xnor (n182,n183,n111);
nor (n183,n184,n185);
and (n184,n87,n103);
and (n185,n95,n108);
xnor (n186,n187,n126);
nor (n187,n188,n189);
and (n188,n102,n119);
and (n189,n110,n123);
xnor (n190,n191,n59);
nor (n191,n192,n193);
and (n192,n118,n50);
and (n193,n125,n55);
xor (n194,n195,n199);
xnor (n195,n196,n74);
nor (n196,n197,n198);
and (n197,n49,n66);
and (n198,n58,n71);
and (n199,n73,n68);
and (n200,n8,n169);
xor (n201,n202,n211);
xor (n202,n203,n207);
or (n203,n204,n205,n206);
and (n204,n136,n173);
and (n205,n173,n176);
and (n206,n136,n176);
or (n207,n208,n209,n210);
and (n208,n182,n186);
and (n209,n186,n190);
and (n210,n182,n190);
and (n211,n195,n199);
and (n212,n201,n213);
xor (n213,n214,n232);
xor (n214,n215,n228);
or (n215,n216,n225,n227);
and (n216,n217,n221);
or (n217,n218,n219,n220);
and (n218,n24,n137);
and (n219,n137,n141);
and (n220,n24,n141);
or (n221,n222,n223,n224);
and (n222,n147,n151);
and (n223,n151,n155);
and (n224,n147,n155);
and (n225,n221,n226);
or (n226,n162,n166);
and (n227,n217,n226);
or (n228,n229,n230,n231);
and (n229,n171,n180);
and (n230,n180,n194);
and (n231,n171,n194);
xor (n232,n233,n246);
xor (n233,n234,n235);
and (n234,n49,n68);
xor (n235,n236,n242);
xor (n236,n237,n238);
not (n237,n40);
xnor (n238,n239,n96);
nor (n239,n240,n241);
and (n240,n39,n88);
and (n241,n17,n93);
xnor (n242,n243,n111);
nor (n243,n244,n245);
and (n244,n95,n103);
and (n245,n31,n108);
xor (n246,n247,n256);
xor (n247,n248,n252);
xnor (n248,n249,n126);
nor (n249,n250,n251);
and (n250,n110,n119);
and (n251,n87,n123);
xnor (n252,n253,n59);
nor (n253,n254,n255);
and (n254,n125,n50);
and (n255,n102,n55);
xnor (n256,n257,n74);
nor (n257,n258,n259);
and (n258,n58,n66);
and (n259,n118,n71);
and (n260,n6,n213);
xor (n261,n262,n277);
xor (n262,n263,n267);
or (n263,n264,n265,n266);
and (n264,n215,n228);
and (n265,n228,n232);
and (n266,n215,n232);
xor (n267,n268,n234);
xor (n268,n269,n273);
or (n269,n270,n271,n272);
and (n270,n40,n238);
and (n271,n238,n242);
and (n272,n40,n242);
or (n273,n274,n275,n276);
and (n274,n248,n252);
and (n275,n252,n256);
and (n276,n248,n256);
xor (n277,n278,n289);
xor (n278,n279,n283);
or (n279,n280,n281,n282);
and (n280,n203,n207);
and (n281,n207,n211);
and (n282,n203,n211);
or (n283,n284,n286,n288);
and (n284,n285,n246);
not (n285,n235);
and (n286,n246,n287);
not (n287,n234);
and (n288,n285,n287);
xor (n289,n290,n306);
xor (n290,n291,n292);
and (n291,n58,n68);
xor (n292,n293,n302);
xor (n293,n294,n298);
xnor (n294,n295,n126);
nor (n295,n296,n297);
and (n296,n87,n119);
and (n297,n95,n123);
xnor (n298,n299,n59);
nor (n299,n300,n301);
and (n300,n102,n50);
and (n301,n110,n55);
xnor (n302,n303,n74);
nor (n303,n304,n305);
and (n304,n118,n66);
and (n305,n125,n71);
xor (n306,n307,n311);
xor (n307,n237,n308);
xnor (n308,n309,n96);
not (n309,n310);
and (n310,n17,n88);
xnor (n311,n312,n111);
nor (n312,n313,n314);
and (n313,n31,n103);
and (n314,n39,n108);
and (n315,n316,n381);
or (n316,n317,n377,n380);
and (n317,n318,n375);
or (n318,n319,n371,n374);
and (n319,n320,n366);
or (n320,n321,n350,n365);
and (n321,n322,n338);
or (n322,n323,n332,n337);
and (n323,n324,n328);
xnor (n324,n325,n96);
nor (n325,n326,n327);
and (n326,n110,n88);
and (n327,n87,n93);
xnor (n328,n329,n111);
nor (n329,n330,n331);
and (n330,n125,n103);
and (n331,n102,n108);
and (n332,n328,n333);
xnor (n333,n334,n126);
nor (n334,n335,n336);
and (n335,n58,n119);
and (n336,n118,n123);
and (n337,n324,n333);
or (n338,n339,n344,n349);
and (n339,n13,n340);
xnor (n340,n341,n24);
nor (n341,n342,n343);
and (n342,n39,n18);
and (n343,n17,n23);
and (n344,n340,n345);
xnor (n345,n346,n40);
nor (n346,n347,n348);
and (n347,n95,n32);
and (n348,n31,n37);
and (n349,n13,n345);
and (n350,n338,n351);
or (n351,n352,n361,n364);
and (n352,n353,n357);
xnor (n353,n354,n59);
nor (n354,n355,n356);
and (n355,n73,n50);
and (n356,n49,n55);
xnor (n357,n358,n74);
nor (n358,n359,n360);
and (n359,n79,n66);
and (n360,n65,n71);
and (n361,n357,n362);
and (n362,n363,n68);
and (n364,n353,n362);
and (n365,n322,n351);
or (n366,n367,n369);
xor (n367,n368,n78);
xor (n368,n46,n62);
xor (n369,n370,n115);
xor (n370,n84,n99);
and (n371,n366,n372);
xor (n372,n373,n161);
xor (n373,n134,n145);
and (n374,n320,n372);
xor (n375,n376,n226);
xor (n376,n217,n221);
and (n377,n375,n378);
xor (n378,n379,n169);
xor (n379,n8,n131);
and (n380,n318,n378);
xor (n381,n382,n213);
xor (n382,n6,n201);
or (n383,n384,n464);
and (n384,n385,n386);
xor (n385,n316,n381);
and (n386,n387,n462);
or (n387,n388,n458,n461);
and (n388,n389,n454);
or (n389,n390,n450,n453);
and (n390,n391,n439);
or (n391,n392,n425,n438);
and (n392,n393,n409);
or (n393,n394,n403,n408);
and (n394,n395,n399);
xnor (n395,n396,n40);
nor (n396,n397,n398);
and (n397,n87,n32);
and (n398,n95,n37);
xnor (n399,n400,n96);
nor (n400,n401,n402);
and (n401,n102,n88);
and (n402,n110,n93);
and (n403,n399,n404);
xnor (n404,n405,n111);
nor (n405,n406,n407);
and (n406,n118,n103);
and (n407,n125,n108);
and (n408,n395,n404);
or (n409,n410,n419,n424);
and (n410,n411,n415);
xnor (n411,n412,n126);
nor (n412,n413,n414);
and (n413,n49,n119);
and (n414,n58,n123);
xnor (n415,n416,n59);
nor (n416,n417,n418);
and (n417,n65,n50);
and (n418,n73,n55);
and (n419,n415,n420);
xnor (n420,n421,n74);
nor (n421,n422,n423);
and (n422,n363,n66);
and (n423,n79,n71);
and (n424,n411,n420);
and (n425,n409,n426);
and (n426,n427,n434);
xnor (n427,n428,n13);
not (n428,n429);
and (n429,n17,n430);
and (n430,n431,n433);
xor (n431,n13,n432);
not (n433,n432);
xnor (n434,n435,n24);
nor (n435,n436,n437);
and (n436,n31,n18);
and (n437,n39,n23);
and (n438,n393,n426);
or (n439,n440,n446,n449);
and (n440,n441,n443);
xor (n441,n442,n333);
xor (n442,n324,n328);
not (n443,n444);
xor (n444,n445,n345);
xor (n445,n12,n340);
and (n446,n443,n447);
xor (n447,n448,n362);
xor (n448,n353,n357);
and (n449,n441,n447);
and (n450,n439,n451);
xor (n451,n452,n28);
xor (n452,n12,n14);
and (n453,n391,n451);
and (n454,n455,n457);
xor (n455,n456,n351);
xor (n456,n322,n338);
xnor (n457,n367,n369);
and (n458,n454,n459);
xor (n459,n460,n82);
xor (n460,n10,n44);
and (n461,n389,n459);
xor (n462,n463,n378);
xor (n463,n318,n375);
and (n464,n465,n466);
xor (n465,n385,n386);
or (n466,n467,n546);
and (n467,n468,n469);
xor (n468,n387,n462);
or (n469,n470,n542,n545);
and (n470,n471,n540);
or (n471,n472,n537,n539);
and (n472,n473,n535);
or (n473,n474,n531,n534);
and (n474,n475,n521);
or (n475,n476,n509,n520);
and (n476,n477,n493);
or (n477,n478,n487,n492);
and (n478,n479,n483);
xnor (n479,n480,n13);
nor (n480,n481,n482);
and (n481,n39,n430);
and (n482,n17,n432);
xnor (n483,n484,n24);
nor (n484,n485,n486);
and (n485,n95,n18);
and (n486,n31,n23);
and (n487,n483,n488);
xnor (n488,n489,n40);
nor (n489,n490,n491);
and (n490,n110,n32);
and (n491,n87,n37);
and (n492,n479,n488);
or (n493,n494,n503,n508);
and (n494,n495,n499);
xnor (n495,n496,n96);
nor (n496,n497,n498);
and (n497,n125,n88);
and (n498,n102,n93);
xnor (n499,n500,n111);
nor (n500,n501,n502);
and (n501,n58,n103);
and (n502,n118,n108);
and (n503,n499,n504);
xnor (n504,n505,n126);
nor (n505,n506,n507);
and (n506,n73,n119);
and (n507,n49,n123);
and (n508,n495,n504);
and (n509,n493,n510);
and (n510,n511,n515);
xnor (n511,n512,n59);
nor (n512,n513,n514);
and (n513,n79,n50);
and (n514,n65,n55);
xnor (n515,n516,n74);
nor (n516,n517,n519);
and (n517,n518,n66);
and (n519,n363,n71);
and (n520,n477,n510);
or (n521,n522,n527,n530);
and (n522,n523,n525);
not (n523,n524);
nand (n524,n518,n68);
xor (n525,n526,n404);
xor (n526,n395,n399);
and (n527,n525,n528);
xor (n528,n529,n420);
xor (n529,n411,n415);
and (n530,n523,n528);
and (n531,n521,n532);
xor (n532,n533,n447);
xor (n533,n441,n443);
and (n534,n475,n532);
xor (n535,n536,n451);
xor (n536,n391,n439);
and (n537,n535,n538);
xor (n538,n455,n457);
and (n539,n473,n538);
xor (n540,n541,n459);
xor (n541,n389,n454);
and (n542,n540,n543);
xor (n543,n544,n372);
xor (n544,n320,n366);
and (n545,n471,n543);
and (n546,n547,n548);
xor (n547,n468,n469);
or (n548,n549,n626);
and (n549,n550,n552);
xor (n550,n551,n543);
xor (n551,n471,n540);
and (n552,n553,n624);
or (n553,n554,n620,n623);
and (n554,n555,n615);
or (n555,n556,n612,n614);
and (n556,n557,n603);
or (n557,n558,n585,n602);
and (n558,n559,n573);
or (n559,n560,n569,n572);
and (n560,n561,n565);
xnor (n561,n562,n126);
nor (n562,n563,n564);
and (n563,n65,n119);
and (n564,n73,n123);
xnor (n565,n566,n59);
nor (n566,n567,n568);
and (n567,n363,n50);
and (n568,n79,n55);
and (n569,n565,n570);
xnor (n570,n571,n74);
nand (n571,n518,n71);
and (n572,n561,n570);
or (n573,n574,n583,n584);
and (n574,n575,n579);
xnor (n575,n576,n13);
nor (n576,n577,n578);
and (n577,n31,n430);
and (n578,n39,n432);
xnor (n579,n580,n24);
nor (n580,n581,n582);
and (n581,n87,n18);
and (n582,n95,n23);
and (n583,n579,n74);
and (n584,n575,n74);
and (n585,n573,n586);
or (n586,n587,n596,n601);
and (n587,n588,n592);
xnor (n588,n589,n40);
nor (n589,n590,n591);
and (n590,n102,n32);
and (n591,n110,n37);
xnor (n592,n593,n96);
nor (n593,n594,n595);
and (n594,n118,n88);
and (n595,n125,n93);
and (n596,n592,n597);
xnor (n597,n598,n111);
nor (n598,n599,n600);
and (n599,n49,n103);
and (n600,n58,n108);
and (n601,n588,n597);
and (n602,n559,n586);
or (n603,n604,n609,n611);
and (n604,n605,n607);
xor (n605,n606,n488);
xor (n606,n479,n483);
xor (n607,n608,n504);
xor (n608,n495,n499);
and (n609,n607,n610);
xor (n610,n511,n515);
and (n611,n605,n610);
and (n612,n603,n613);
xor (n613,n427,n434);
and (n614,n557,n613);
and (n615,n616,n618);
xor (n616,n617,n510);
xor (n617,n477,n493);
xor (n618,n619,n528);
xor (n619,n523,n525);
and (n620,n615,n621);
xor (n621,n622,n426);
xor (n622,n393,n409);
and (n623,n555,n621);
xor (n624,n625,n538);
xor (n625,n473,n535);
and (n626,n627,n628);
xor (n627,n550,n552);
or (n628,n629,n636);
and (n629,n630,n631);
xor (n630,n553,n624);
and (n631,n632,n634);
xor (n632,n633,n621);
xor (n633,n555,n615);
xor (n634,n635,n532);
xor (n635,n475,n521);
and (n636,n637,n669);
xor (n637,n638,n663);
xor (n638,n639,n643);
or (n639,n554,n640,n642);
and (n640,n615,n641);
xnor (n641,n441,n447);
and (n642,n555,n641);
xor (n643,n644,n653);
xor (n644,n645,n648);
or (n645,n474,n646,n647);
and (n646,n521,n444);
and (n647,n475,n444);
xor (n648,n649,n351);
xor (n649,n322,n650);
or (n650,n651,n344,n652);
and (n651,n12,n340);
and (n652,n12,n345);
xor (n653,n654,n656);
xor (n654,n391,n655);
or (n655,n441,n447);
xor (n656,n657,n662);
xor (n657,n658,n660);
xor (n658,n659,n84);
xor (n659,n14,n28);
xor (n660,n661,n46);
xor (n661,n99,n115);
xnor (n662,n62,n78);
or (n663,n664,n666,n668);
and (n664,n621,n665);
xor (n665,n635,n444);
and (n666,n665,n667);
xor (n667,n633,n641);
and (n668,n621,n667);
or (n669,n670,n729);
and (n670,n671,n673);
xor (n671,n672,n667);
xor (n672,n621,n665);
or (n673,n674,n726,n728);
and (n674,n675,n724);
or (n675,n676,n720,n723);
and (n676,n677,n715);
or (n677,n678,n711,n714);
and (n678,n679,n695);
or (n679,n680,n689,n694);
and (n680,n681,n685);
xnor (n681,n682,n13);
nor (n682,n683,n684);
and (n683,n95,n430);
and (n684,n31,n432);
xnor (n685,n686,n24);
nor (n686,n687,n688);
and (n687,n110,n18);
and (n688,n87,n23);
and (n689,n685,n690);
xnor (n690,n691,n40);
nor (n691,n692,n693);
and (n692,n125,n32);
and (n693,n102,n37);
and (n694,n681,n690);
or (n695,n696,n705,n710);
and (n696,n697,n701);
xnor (n697,n698,n96);
nor (n698,n699,n700);
and (n699,n58,n88);
and (n700,n118,n93);
xnor (n701,n702,n111);
nor (n702,n703,n704);
and (n703,n73,n103);
and (n704,n49,n108);
and (n705,n701,n706);
xnor (n706,n707,n126);
nor (n707,n708,n709);
and (n708,n79,n119);
and (n709,n65,n123);
and (n710,n697,n706);
and (n711,n695,n712);
xor (n712,n713,n570);
xor (n713,n561,n565);
and (n714,n679,n712);
and (n715,n716,n718);
xor (n716,n717,n74);
xor (n717,n575,n579);
xor (n718,n719,n597);
xor (n719,n588,n592);
and (n720,n715,n721);
xor (n721,n722,n610);
xor (n722,n605,n607);
and (n723,n677,n721);
xor (n724,n725,n613);
xor (n725,n557,n603);
and (n726,n724,n727);
xor (n727,n616,n618);
and (n728,n675,n727);
and (n729,n730,n731);
xor (n730,n671,n673);
or (n731,n732,n786);
and (n732,n733,n735);
xor (n733,n734,n727);
xor (n734,n675,n724);
or (n735,n736,n782,n785);
and (n736,n737,n780);
or (n737,n738,n777,n779);
and (n738,n739,n775);
or (n739,n740,n769,n774);
and (n740,n741,n753);
or (n741,n742,n751,n752);
and (n742,n743,n747);
xnor (n743,n744,n13);
nor (n744,n745,n746);
and (n745,n87,n430);
and (n746,n95,n432);
xnor (n747,n748,n24);
nor (n748,n749,n750);
and (n749,n102,n18);
and (n750,n110,n23);
and (n751,n747,n59);
and (n752,n743,n59);
or (n753,n754,n763,n768);
and (n754,n755,n759);
xnor (n755,n756,n40);
nor (n756,n757,n758);
and (n757,n118,n32);
and (n758,n125,n37);
xnor (n759,n760,n96);
nor (n760,n761,n762);
and (n761,n49,n88);
and (n762,n58,n93);
and (n763,n759,n764);
xnor (n764,n765,n111);
nor (n765,n766,n767);
and (n766,n65,n103);
and (n767,n73,n108);
and (n768,n755,n764);
and (n769,n753,n770);
xnor (n770,n771,n59);
nor (n771,n772,n773);
and (n772,n518,n50);
and (n773,n363,n55);
and (n774,n741,n770);
xor (n775,n776,n712);
xor (n776,n679,n695);
and (n777,n775,n778);
xor (n778,n716,n718);
and (n779,n739,n778);
xor (n780,n781,n586);
xor (n781,n559,n573);
and (n782,n780,n783);
xor (n783,n784,n721);
xor (n784,n677,n715);
and (n785,n737,n783);
and (n786,n787,n788);
xor (n787,n733,n735);
or (n788,n789,n859);
and (n789,n790,n792);
xor (n790,n791,n783);
xor (n791,n737,n780);
or (n792,n793,n855,n858);
and (n793,n794,n850);
or (n794,n795,n846,n849);
and (n795,n796,n836);
or (n796,n797,n830,n835);
and (n797,n798,n814);
or (n798,n799,n808,n813);
and (n799,n800,n804);
xnor (n800,n801,n96);
nor (n801,n802,n803);
and (n802,n73,n88);
and (n803,n49,n93);
xnor (n804,n805,n111);
nor (n805,n806,n807);
and (n806,n79,n103);
and (n807,n65,n108);
and (n808,n804,n809);
xnor (n809,n810,n126);
nor (n810,n811,n812);
and (n811,n518,n119);
and (n812,n363,n123);
and (n813,n800,n809);
or (n814,n815,n824,n829);
and (n815,n816,n820);
xnor (n816,n817,n13);
nor (n817,n818,n819);
and (n818,n110,n430);
and (n819,n87,n432);
xnor (n820,n821,n24);
nor (n821,n822,n823);
and (n822,n125,n18);
and (n823,n102,n23);
and (n824,n820,n825);
xnor (n825,n826,n40);
nor (n826,n827,n828);
and (n827,n58,n32);
and (n828,n118,n37);
and (n829,n816,n825);
and (n830,n814,n831);
xnor (n831,n832,n126);
nor (n832,n833,n834);
and (n833,n363,n119);
and (n834,n79,n123);
and (n835,n798,n831);
or (n836,n837,n842,n845);
and (n837,n838,n840);
xnor (n838,n839,n59);
nand (n839,n518,n55);
xor (n840,n841,n59);
xor (n841,n743,n747);
and (n842,n840,n843);
xor (n843,n844,n764);
xor (n844,n755,n759);
and (n845,n838,n843);
and (n846,n836,n847);
xor (n847,n848,n706);
xor (n848,n697,n701);
and (n849,n796,n847);
and (n850,n851,n853);
xor (n851,n852,n690);
xor (n852,n681,n685);
xor (n853,n854,n770);
xor (n854,n741,n753);
and (n855,n850,n856);
xor (n856,n857,n778);
xor (n857,n739,n775);
and (n858,n794,n856);
and (n859,n860,n861);
xor (n860,n790,n792);
or (n861,n862,n914);
and (n862,n863,n865);
xor (n863,n864,n856);
xor (n864,n794,n850);
or (n865,n866,n911,n913);
and (n866,n867,n909);
or (n867,n868,n905,n908);
and (n868,n869,n903);
or (n869,n870,n899,n902);
and (n870,n871,n887);
or (n871,n872,n881,n886);
and (n872,n873,n877);
xnor (n873,n874,n40);
nor (n874,n875,n876);
and (n875,n49,n32);
and (n876,n58,n37);
xnor (n877,n878,n96);
nor (n878,n879,n880);
and (n879,n65,n88);
and (n880,n73,n93);
and (n881,n877,n882);
xnor (n882,n883,n111);
nor (n883,n884,n885);
and (n884,n363,n103);
and (n885,n79,n108);
and (n886,n873,n882);
or (n887,n888,n897,n898);
and (n888,n889,n893);
xnor (n889,n890,n13);
nor (n890,n891,n892);
and (n891,n102,n430);
and (n892,n110,n432);
xnor (n893,n894,n24);
nor (n894,n895,n896);
and (n895,n118,n18);
and (n896,n125,n23);
and (n897,n893,n126);
and (n898,n889,n126);
and (n899,n887,n900);
xor (n900,n901,n809);
xor (n901,n800,n804);
and (n902,n871,n900);
xor (n903,n904,n831);
xor (n904,n798,n814);
and (n905,n903,n906);
xor (n906,n907,n843);
xor (n907,n838,n840);
and (n908,n869,n906);
xor (n909,n910,n847);
xor (n910,n796,n836);
and (n911,n909,n912);
xor (n912,n851,n853);
and (n913,n867,n912);
and (n914,n915,n916);
xor (n915,n863,n865);
or (n916,n917,n955);
and (n917,n918,n920);
xor (n918,n919,n912);
xor (n919,n867,n909);
and (n920,n921,n953);
or (n921,n922,n949,n952);
and (n922,n923,n947);
or (n923,n924,n943,n946);
and (n924,n925,n941);
or (n925,n926,n935,n940);
and (n926,n927,n931);
xnor (n927,n928,n13);
nor (n928,n929,n930);
and (n929,n125,n430);
and (n930,n102,n432);
xnor (n931,n932,n24);
nor (n932,n933,n934);
and (n933,n58,n18);
and (n934,n118,n23);
and (n935,n931,n936);
xnor (n936,n937,n40);
nor (n937,n938,n939);
and (n938,n73,n32);
and (n939,n49,n37);
and (n940,n927,n936);
xnor (n941,n942,n126);
nand (n942,n518,n123);
and (n943,n941,n944);
xor (n944,n945,n882);
xor (n945,n873,n877);
and (n946,n925,n944);
xor (n947,n948,n825);
xor (n948,n816,n820);
and (n949,n947,n950);
xor (n950,n951,n900);
xor (n951,n871,n887);
and (n952,n923,n950);
xor (n953,n954,n906);
xor (n954,n869,n903);
and (n955,n956,n957);
xor (n956,n918,n920);
or (n957,n958,n1010);
and (n958,n959,n960);
xor (n959,n921,n953);
and (n960,n961,n1008);
or (n961,n962,n1004,n1007);
and (n962,n963,n997);
or (n963,n964,n991,n996);
and (n964,n965,n979);
or (n965,n966,n975,n978);
and (n966,n967,n971);
xnor (n967,n968,n40);
nor (n968,n969,n970);
and (n969,n65,n32);
and (n970,n73,n37);
xnor (n971,n972,n96);
nor (n972,n973,n974);
and (n973,n363,n88);
and (n974,n79,n93);
and (n975,n971,n976);
xnor (n976,n977,n111);
nand (n977,n518,n108);
and (n978,n967,n976);
or (n979,n980,n989,n990);
and (n980,n981,n985);
xnor (n981,n982,n13);
nor (n982,n983,n984);
and (n983,n118,n430);
and (n984,n125,n432);
xnor (n985,n986,n24);
nor (n986,n987,n988);
and (n987,n49,n18);
and (n988,n58,n23);
and (n989,n985,n111);
and (n990,n981,n111);
and (n991,n979,n992);
xnor (n992,n993,n96);
nor (n993,n994,n995);
and (n994,n79,n88);
and (n995,n65,n93);
and (n996,n965,n992);
and (n997,n998,n1002);
xnor (n998,n999,n111);
nor (n999,n1000,n1001);
and (n1000,n518,n103);
and (n1001,n363,n108);
xor (n1002,n1003,n936);
xor (n1003,n927,n931);
and (n1004,n997,n1005);
xor (n1005,n1006,n126);
xor (n1006,n889,n893);
and (n1007,n963,n1005);
xor (n1008,n1009,n950);
xor (n1009,n923,n947);
and (n1010,n1011,n1012);
xor (n1011,n959,n960);
or (n1012,n1013,n1020);
and (n1013,n1014,n1015);
xor (n1014,n961,n1008);
and (n1015,n1016,n1018);
xor (n1016,n1017,n944);
xor (n1017,n925,n941);
xor (n1018,n1019,n1005);
xor (n1019,n963,n997);
and (n1020,n1021,n1022);
xor (n1021,n1014,n1015);
or (n1022,n1023,n1056);
and (n1023,n1024,n1025);
xor (n1024,n1016,n1018);
or (n1025,n1026,n1053,n1055);
and (n1026,n1027,n1051);
or (n1027,n1028,n1047,n1050);
and (n1028,n1029,n1045);
or (n1029,n1030,n1039,n1044);
and (n1030,n1031,n1035);
xnor (n1031,n1032,n13);
nor (n1032,n1033,n1034);
and (n1033,n58,n430);
and (n1034,n118,n432);
xnor (n1035,n1036,n24);
nor (n1036,n1037,n1038);
and (n1037,n73,n18);
and (n1038,n49,n23);
and (n1039,n1035,n1040);
xnor (n1040,n1041,n40);
nor (n1041,n1042,n1043);
and (n1042,n79,n32);
and (n1043,n65,n37);
and (n1044,n1031,n1040);
xor (n1045,n1046,n976);
xor (n1046,n967,n971);
and (n1047,n1045,n1048);
xor (n1048,n1049,n111);
xor (n1049,n981,n985);
and (n1050,n1029,n1048);
xor (n1051,n1052,n992);
xor (n1052,n965,n979);
and (n1053,n1051,n1054);
xor (n1054,n998,n1002);
and (n1055,n1027,n1054);
and (n1056,n1057,n1058);
xor (n1057,n1024,n1025);
or (n1058,n1059,n1092);
and (n1059,n1060,n1062);
xor (n1060,n1061,n1054);
xor (n1061,n1027,n1051);
and (n1062,n1063,n1090);
or (n1063,n1064,n1084,n1089);
and (n1064,n1065,n1077);
or (n1065,n1066,n1075,n1076);
and (n1066,n1067,n1071);
xnor (n1067,n1068,n13);
nor (n1068,n1069,n1070);
and (n1069,n49,n430);
and (n1070,n58,n432);
xnor (n1071,n1072,n24);
nor (n1072,n1073,n1074);
and (n1073,n65,n18);
and (n1074,n73,n23);
and (n1075,n1071,n96);
and (n1076,n1067,n96);
and (n1077,n1078,n1082);
xnor (n1078,n1079,n40);
nor (n1079,n1080,n1081);
and (n1080,n363,n32);
and (n1081,n79,n37);
xnor (n1082,n1083,n96);
nand (n1083,n518,n93);
and (n1084,n1077,n1085);
xnor (n1085,n1086,n96);
nor (n1086,n1087,n1088);
and (n1087,n518,n88);
and (n1088,n363,n93);
and (n1089,n1065,n1085);
xor (n1090,n1091,n1048);
xor (n1091,n1029,n1045);
and (n1092,n1093,n1094);
xor (n1093,n1060,n1062);
or (n1094,n1095,n1102);
and (n1095,n1096,n1097);
xor (n1096,n1063,n1090);
and (n1097,n1098,n1100);
xor (n1098,n1099,n1040);
xor (n1099,n1031,n1035);
xor (n1100,n1101,n1085);
xor (n1101,n1065,n1077);
and (n1102,n1103,n1104);
xor (n1103,n1096,n1097);
or (n1104,n1105,n1130);
and (n1105,n1106,n1107);
xor (n1106,n1098,n1100);
or (n1107,n1108,n1127,n1129);
and (n1108,n1109,n1125);
or (n1109,n1110,n1119,n1124);
and (n1110,n1111,n1115);
xnor (n1111,n1112,n13);
nor (n1112,n1113,n1114);
and (n1113,n73,n430);
and (n1114,n49,n432);
xnor (n1115,n1116,n24);
nor (n1116,n1117,n1118);
and (n1117,n79,n18);
and (n1118,n65,n23);
and (n1119,n1115,n1120);
xnor (n1120,n1121,n40);
nor (n1121,n1122,n1123);
and (n1122,n518,n32);
and (n1123,n363,n37);
and (n1124,n1111,n1120);
xor (n1125,n1126,n96);
xor (n1126,n1067,n1071);
and (n1127,n1125,n1128);
xor (n1128,n1078,n1082);
and (n1129,n1109,n1128);
and (n1130,n1131,n1132);
xor (n1131,n1106,n1107);
or (n1132,n1133,n1151);
and (n1133,n1134,n1136);
xor (n1134,n1135,n1128);
xor (n1135,n1109,n1125);
and (n1136,n1137,n1149);
or (n1137,n1138,n1147,n1148);
and (n1138,n1139,n1143);
xnor (n1139,n1140,n13);
nor (n1140,n1141,n1142);
and (n1141,n65,n430);
and (n1142,n73,n432);
xnor (n1143,n1144,n24);
nor (n1144,n1145,n1146);
and (n1145,n363,n18);
and (n1146,n79,n23);
and (n1147,n1143,n40);
and (n1148,n1139,n40);
xor (n1149,n1150,n1120);
xor (n1150,n1111,n1115);
and (n1151,n1152,n1153);
xor (n1152,n1134,n1136);
or (n1153,n1154,n1161);
and (n1154,n1155,n1156);
xor (n1155,n1137,n1149);
and (n1156,n1157,n1159);
xnor (n1157,n1158,n40);
nand (n1158,n518,n37);
xor (n1159,n1160,n40);
xor (n1160,n1139,n1143);
and (n1161,n1162,n1163);
xor (n1162,n1155,n1156);
or (n1163,n1164,n1175);
and (n1164,n1165,n1166);
xor (n1165,n1157,n1159);
and (n1166,n1167,n1171);
xnor (n1167,n1168,n13);
nor (n1168,n1169,n1170);
and (n1169,n79,n430);
and (n1170,n65,n432);
xnor (n1171,n1172,n24);
nor (n1172,n1173,n1174);
and (n1173,n518,n18);
and (n1174,n363,n23);
and (n1175,n1176,n1177);
xor (n1176,n1165,n1166);
or (n1177,n1178,n1185);
and (n1178,n1179,n1180);
xor (n1179,n1167,n1171);
and (n1180,n1181,n24);
xnor (n1181,n1182,n13);
nor (n1182,n1183,n1184);
and (n1183,n363,n430);
and (n1184,n79,n432);
and (n1185,n1186,n1187);
xor (n1186,n1179,n1180);
or (n1187,n1188,n1192);
and (n1188,n1189,n1191);
xnor (n1189,n1190,n24);
nand (n1190,n518,n23);
xor (n1191,n1181,n24);
and (n1192,n1193,n1194);
xor (n1193,n1189,n1191);
and (n1194,n1195,n1199);
xnor (n1195,n1196,n13);
nor (n1196,n1197,n1198);
and (n1197,n518,n430);
and (n1198,n363,n432);
and (n1199,n1200,n13);
xnor (n1200,n1201,n13);
nand (n1201,n518,n432);
buf (n1202,n1203);
xor (n1203,n1204,n1306);
xor (n1204,n1205,n1284);
xor (n1205,n1206,n1259);
or (n1206,n1207,n1243,n1258);
and (n1207,n1208,n1234);
or (n1208,n1209,n1225,n1233);
and (n1209,n1210,n1221);
or (n1210,n1211,n1218,n1220);
and (n1211,n1212,n1215);
or (n1212,n27,n1213,n1214);
and (n1213,n28,n84);
and (n1214,n14,n84);
or (n1215,n114,n1216,n1217);
and (n1216,n115,n46);
and (n1217,n99,n46);
and (n1218,n1215,n1219);
or (n1219,n62,n78);
and (n1220,n1212,n1219);
or (n1221,n1222,n1223,n1224);
and (n1222,n134,n145);
and (n1223,n145,n161);
and (n1224,n134,n161);
and (n1225,n1221,n1226);
xor (n1226,n1227,n1232);
xor (n1227,n1228,n1230);
xor (n1228,n1229,n182);
xor (n1229,n173,n176);
xor (n1230,n1231,n195);
xor (n1231,n186,n190);
not (n1232,n199);
and (n1233,n1210,n1226);
xor (n1234,n1235,n1242);
xor (n1235,n1236,n1239);
or (n1236,n205,n1237,n1238);
and (n1237,n176,n182);
and (n1238,n173,n182);
or (n1239,n209,n1240,n1241);
and (n1240,n190,n195);
and (n1241,n186,n195);
buf (n1242,n199);
and (n1243,n1234,n1244);
xor (n1244,n1245,n232);
xor (n1245,n1246,n1254);
or (n1246,n1247,n1251,n1253);
and (n1247,n1248,n221);
or (n1248,n1249,n219,n1250);
and (n1249,n136,n137);
and (n1250,n136,n141);
and (n1251,n221,n1252);
and (n1252,n162,n166);
and (n1253,n1248,n1252);
or (n1254,n1255,n1256,n1257);
and (n1255,n1228,n1230);
and (n1256,n1230,n1232);
and (n1257,n1228,n1232);
and (n1258,n1208,n1244);
xor (n1259,n1260,n1277);
xor (n1260,n1261,n1265);
or (n1261,n1262,n1263,n1264);
and (n1262,n1246,n1254);
and (n1263,n1254,n232);
and (n1264,n1246,n232);
xor (n1265,n1266,n1275);
xor (n1266,n1267,n1271);
or (n1267,n1268,n1269,n1270);
and (n1268,n1236,n1239);
and (n1269,n1239,n1242);
and (n1270,n1236,n1242);
or (n1271,n1272,n1273,n1274);
and (n1272,n234,n235);
and (n1273,n235,n246);
and (n1274,n234,n246);
xor (n1275,n1276,n291);
xor (n1276,n298,n302);
xor (n1277,n1278,n1280);
xor (n1278,n1279,n294);
xor (n1279,n308,n311);
xnor (n1280,n1281,n273);
or (n1281,n1282,n271,n1283);
and (n1282,n237,n238);
and (n1283,n237,n242);
and (n1284,n1285,n1304);
or (n1285,n1286,n1300,n1303);
and (n1286,n1287,n1298);
or (n1287,n1288,n1296,n1297);
and (n1288,n1289,n1292);
or (n1289,n1290,n1291,n365);
and (n1290,n322,n650);
and (n1291,n650,n351);
or (n1292,n1293,n1294,n1295);
and (n1293,n658,n660);
and (n1294,n660,n662);
and (n1295,n658,n662);
and (n1296,n1292,n372);
and (n1297,n1289,n372);
xor (n1298,n1299,n1252);
xor (n1299,n1248,n221);
and (n1300,n1298,n1301);
xor (n1301,n1302,n1226);
xor (n1302,n1210,n1221);
and (n1303,n1287,n1301);
xor (n1304,n1305,n1244);
xor (n1305,n1208,n1234);
or (n1306,n1307,n1324);
and (n1307,n1308,n1309);
xor (n1308,n1285,n1304);
and (n1309,n1310,n1322);
or (n1310,n1311,n1318,n1321);
and (n1311,n1312,n1316);
or (n1312,n1313,n1314,n1315);
and (n1313,n391,n655);
and (n1314,n655,n656);
and (n1315,n391,n656);
xor (n1316,n1317,n1219);
xor (n1317,n1212,n1215);
and (n1318,n1316,n1319);
xor (n1319,n1320,n372);
xor (n1320,n1289,n1292);
and (n1321,n1312,n1319);
xor (n1322,n1323,n1301);
xor (n1323,n1287,n1298);
and (n1324,n1325,n1326);
xor (n1325,n1308,n1309);
or (n1326,n1327,n1336);
and (n1327,n1328,n1329);
xor (n1328,n1310,n1322);
and (n1329,n1330,n1334);
or (n1330,n1331,n1332,n1333);
and (n1331,n645,n648);
and (n1332,n648,n653);
and (n1333,n645,n653);
xor (n1334,n1335,n1319);
xor (n1335,n1312,n1316);
and (n1336,n1337,n1338);
xor (n1337,n1328,n1329);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1330,n1334);
and (n1341,n639,n643);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n636);
and (n1345,n638,n663);
endmodule
