module top (out,n3,n4,n5,n23,n24,n29,n33,n40,n49
        ,n50,n56,n60,n66,n84,n91,n92,n102,n122,n124
        ,n130,n140,n158,n167,n177,n181,n188,n213);
output out;
input n3;
input n4;
input n5;
input n23;
input n24;
input n29;
input n33;
input n40;
input n49;
input n50;
input n56;
input n60;
input n66;
input n84;
input n91;
input n92;
input n102;
input n122;
input n124;
input n130;
input n140;
input n158;
input n167;
input n177;
input n181;
input n188;
input n213;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
xnor (out,n0,n552);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n549);
nand (n7,n8,n548);
or (n8,n9,n298);
not (n9,n10);
nand (n10,n11,n297);
nand (n11,n12,n262);
not (n12,n13);
xor (n13,n14,n216);
xor (n14,n15,n105);
xor (n15,n16,n69);
xor (n16,n17,n43);
nand (n17,n18,n37);
or (n18,n19,n31);
nand (n19,n20,n27);
nor (n20,n21,n25);
and (n21,n22,n24);
not (n22,n23);
and (n25,n23,n26);
not (n26,n24);
nand (n27,n28,n30);
or (n28,n26,n29);
nand (n30,n26,n29);
nor (n31,n32,n35);
and (n32,n33,n34);
not (n34,n29);
and (n35,n36,n29);
not (n36,n33);
or (n37,n20,n38);
nor (n38,n39,n41);
and (n39,n34,n40);
and (n41,n29,n42);
not (n42,n40);
nand (n43,n44,n63);
or (n44,n45,n58);
nand (n45,n46,n53);
nor (n46,n47,n51);
and (n47,n48,n50);
not (n48,n49);
and (n51,n49,n52);
not (n52,n50);
nand (n53,n54,n57);
or (n54,n50,n55);
not (n55,n56);
nand (n57,n55,n50);
nor (n58,n59,n61);
and (n59,n55,n60);
and (n61,n56,n62);
not (n62,n60);
or (n63,n46,n64);
nor (n64,n65,n67);
and (n65,n55,n66);
and (n67,n56,n68);
not (n68,n66);
nand (n69,n70,n104);
or (n70,n71,n77);
not (n71,n72);
nand (n72,n73,n29);
nand (n73,n74,n75);
or (n74,n23,n24);
nand (n75,n76,n36);
or (n76,n26,n22);
not (n77,n78);
nand (n78,n79,n98);
or (n79,n80,n86);
not (n80,n81);
nand (n81,n82,n85);
or (n82,n49,n83);
not (n83,n84);
or (n85,n48,n84);
not (n86,n87);
nor (n87,n88,n94);
nand (n88,n89,n93);
or (n89,n90,n92);
not (n90,n91);
nand (n93,n90,n92);
nor (n94,n95,n96);
and (n95,n48,n92);
and (n96,n49,n97);
not (n97,n92);
nand (n98,n88,n99);
nand (n99,n100,n103);
or (n100,n49,n101);
not (n101,n102);
or (n103,n48,n102);
or (n104,n78,n72);
xor (n105,n106,n193);
xor (n106,n107,n144);
or (n107,n108,n143);
and (n108,n109,n117);
xor (n109,n110,n111);
nor (n110,n20,n36);
nand (n111,n112,n116);
or (n112,n113,n86);
nor (n113,n114,n115);
and (n114,n68,n49);
and (n115,n66,n48);
nand (n116,n81,n88);
nand (n117,n118,n136);
or (n118,n119,n127);
not (n119,n120);
nand (n120,n121,n125);
or (n121,n122,n123);
not (n123,n124);
or (n125,n126,n124);
not (n126,n122);
nand (n127,n128,n132);
nand (n128,n129,n131);
or (n129,n130,n126);
nand (n131,n126,n130);
not (n132,n133);
nand (n133,n134,n135);
or (n134,n55,n130);
nand (n135,n55,n130);
nand (n136,n137,n133);
not (n137,n138);
nor (n138,n139,n141);
and (n139,n126,n140);
and (n141,n122,n142);
not (n142,n140);
and (n143,n110,n111);
or (n144,n145,n192);
and (n145,n146,n184);
xor (n146,n147,n170);
nand (n147,n148,n163);
or (n148,n149,n153);
not (n149,n150);
nand (n150,n151,n152);
or (n151,n23,n42);
or (n152,n22,n40);
not (n153,n154);
and (n154,n155,n160);
not (n155,n156);
nand (n156,n157,n159);
or (n157,n158,n126);
nand (n159,n158,n126);
nand (n160,n161,n162);
or (n161,n158,n22);
nand (n162,n22,n158);
nand (n163,n164,n156);
not (n164,n165);
nor (n165,n166,n168);
and (n166,n22,n167);
and (n168,n23,n169);
not (n169,n167);
nand (n170,n171,n178);
or (n171,n172,n175);
nor (n172,n173,n174);
and (n173,n90,n102);
and (n174,n91,n101);
nand (n175,n91,n176);
not (n176,n177);
or (n178,n179,n176);
nor (n179,n180,n182);
and (n180,n90,n181);
and (n182,n91,n183);
not (n183,n181);
nand (n184,n185,n191);
or (n185,n45,n186);
nor (n186,n187,n189);
and (n187,n55,n188);
and (n189,n56,n190);
not (n190,n188);
or (n191,n46,n58);
and (n192,n147,n170);
xor (n193,n194,n208);
xor (n194,n195,n201);
nand (n195,n196,n197);
or (n196,n127,n138);
or (n197,n132,n198);
nor (n198,n199,n200);
and (n199,n126,n188);
and (n200,n122,n190);
nand (n201,n202,n203);
or (n202,n153,n165);
or (n203,n155,n204);
not (n204,n205);
nor (n205,n206,n207);
and (n206,n123,n22);
and (n207,n23,n124);
nand (n208,n209,n210);
or (n209,n179,n175);
or (n210,n211,n176);
nor (n211,n212,n214);
and (n212,n90,n213);
and (n214,n91,n215);
not (n215,n213);
or (n216,n217,n261);
and (n217,n218,n260);
xor (n218,n219,n234);
and (n219,n220,n226);
and (n220,n221,n23);
nand (n221,n222,n223);
or (n222,n122,n158);
nand (n223,n224,n36);
or (n224,n225,n126);
not (n225,n158);
nand (n226,n227,n232);
or (n227,n228,n86);
not (n228,n229);
nand (n229,n230,n231);
or (n230,n49,n62);
or (n231,n48,n60);
or (n232,n233,n113);
not (n233,n88);
or (n234,n235,n259);
and (n235,n236,n252);
xor (n236,n237,n245);
nand (n237,n238,n239);
or (n238,n132,n119);
nand (n239,n240,n244);
not (n240,n241);
nor (n241,n242,n243);
and (n242,n169,n122);
and (n243,n167,n126);
not (n244,n127);
nand (n245,n246,n251);
or (n246,n247,n153);
not (n247,n248);
nand (n248,n249,n250);
or (n249,n23,n36);
or (n250,n22,n33);
nand (n251,n150,n156);
nand (n252,n253,n258);
or (n253,n254,n175);
not (n254,n255);
nor (n255,n256,n257);
and (n256,n83,n90);
and (n257,n91,n84);
or (n258,n172,n176);
and (n259,n237,n245);
xor (n260,n109,n117);
and (n261,n219,n234);
not (n262,n263);
or (n263,n264,n296);
and (n264,n265,n295);
xor (n265,n266,n267);
xor (n266,n146,n184);
or (n267,n268,n294);
and (n268,n269,n277);
xor (n269,n270,n276);
nand (n270,n271,n275);
or (n271,n45,n272);
nor (n272,n273,n274);
and (n273,n55,n140);
and (n274,n56,n142);
or (n275,n186,n46);
xor (n276,n220,n226);
or (n277,n278,n293);
and (n278,n279,n287);
xor (n279,n280,n281);
and (n280,n156,n33);
nand (n281,n282,n283);
or (n282,n176,n254);
or (n283,n284,n175);
nor (n284,n285,n286);
and (n285,n90,n66);
and (n286,n91,n68);
nand (n287,n288,n292);
or (n288,n127,n289);
nor (n289,n290,n291);
and (n290,n126,n40);
and (n291,n122,n42);
or (n292,n132,n241);
and (n293,n280,n281);
and (n294,n270,n276);
xor (n295,n218,n260);
and (n296,n266,n267);
nand (n297,n13,n263);
not (n298,n299);
nand (n299,n300,n547);
or (n300,n301,n542);
nor (n301,n302,n534);
and (n302,n303,n503);
or (n303,n304,n502);
and (n304,n305,n393);
xor (n305,n306,n357);
or (n306,n307,n356);
and (n307,n308,n335);
xor (n308,n309,n318);
nand (n309,n310,n314);
or (n310,n45,n311);
nor (n311,n312,n313);
and (n312,n55,n40);
and (n313,n56,n42);
or (n314,n46,n315);
nor (n315,n316,n317);
and (n316,n55,n167);
and (n317,n56,n169);
nor (n318,n319,n330);
not (n319,n320);
nand (n320,n321,n326);
or (n321,n175,n322);
not (n322,n323);
nor (n323,n324,n325);
and (n324,n91,n140);
and (n325,n142,n90);
nand (n326,n327,n177);
nand (n327,n328,n329);
or (n328,n188,n90);
nand (n329,n90,n188);
nand (n330,n331,n56);
nand (n331,n332,n333);
or (n332,n49,n50);
nand (n333,n334,n36);
or (n334,n52,n48);
xor (n335,n336,n346);
xor (n336,n337,n338);
and (n337,n133,n33);
nand (n338,n339,n344);
or (n339,n176,n340);
not (n340,n341);
nor (n341,n342,n343);
and (n342,n91,n60);
and (n343,n62,n90);
or (n344,n345,n175);
not (n345,n327);
nand (n346,n347,n352);
or (n347,n348,n86);
not (n348,n349);
nor (n349,n350,n351);
and (n350,n49,n124);
and (n351,n123,n48);
nand (n352,n88,n353);
nand (n353,n354,n355);
or (n354,n49,n142);
or (n355,n48,n140);
and (n356,n309,n318);
xor (n357,n358,n372);
xor (n358,n359,n369);
xor (n359,n360,n366);
nor (n360,n361,n126);
nor (n361,n362,n364);
and (n362,n363,n36);
nand (n363,n56,n130);
and (n364,n55,n365);
not (n365,n130);
nand (n366,n367,n368);
or (n367,n175,n340);
or (n368,n284,n176);
or (n369,n370,n371);
and (n370,n336,n346);
and (n371,n337,n338);
xor (n372,n373,n387);
xor (n373,n374,n380);
nand (n374,n375,n379);
or (n375,n127,n376);
nor (n376,n377,n378);
and (n377,n126,n33);
and (n378,n122,n36);
or (n379,n289,n132);
nand (n380,n381,n386);
or (n381,n382,n233);
not (n382,n383);
nand (n383,n384,n385);
or (n384,n49,n190);
or (n385,n48,n188);
nand (n386,n87,n353);
nand (n387,n388,n389);
or (n388,n45,n315);
or (n389,n46,n390);
nor (n390,n391,n392);
and (n391,n124,n55);
and (n392,n56,n123);
or (n393,n394,n501);
and (n394,n395,n419);
xor (n395,n396,n418);
or (n396,n397,n417);
and (n397,n398,n413);
xor (n398,n399,n406);
nand (n399,n400,n405);
or (n400,n401,n86);
not (n401,n402);
nand (n402,n403,n404);
or (n403,n49,n169);
or (n404,n48,n167);
nand (n405,n88,n349);
nand (n406,n407,n412);
or (n407,n408,n45);
not (n408,n409);
nand (n409,n410,n411);
or (n410,n36,n56);
or (n411,n55,n33);
or (n412,n46,n311);
nand (n413,n414,n416);
or (n414,n415,n319);
not (n415,n330);
or (n416,n320,n330);
and (n417,n399,n406);
xor (n418,n308,n335);
or (n419,n420,n500);
and (n420,n421,n442);
xor (n421,n422,n441);
or (n422,n423,n440);
and (n423,n424,n433);
xor (n424,n425,n426);
nor (n425,n46,n36);
nand (n426,n427,n432);
or (n427,n428,n86);
not (n428,n429);
nor (n429,n430,n431);
and (n430,n42,n48);
and (n431,n49,n40);
nand (n432,n88,n402);
nand (n433,n434,n439);
or (n434,n175,n435);
not (n435,n436);
nor (n436,n437,n438);
and (n437,n123,n90);
and (n438,n91,n124);
or (n439,n322,n176);
and (n440,n425,n426);
xor (n441,n398,n413);
or (n442,n443,n499);
and (n443,n444,n498);
xor (n444,n445,n459);
nor (n445,n446,n454);
not (n446,n447);
nand (n447,n448,n449);
or (n448,n176,n435);
nand (n449,n450,n453);
nor (n450,n451,n452);
and (n451,n169,n90);
and (n452,n91,n167);
not (n453,n175);
nand (n454,n455,n49);
nand (n455,n456,n457);
or (n456,n92,n91);
or (n457,n458,n33);
and (n458,n91,n92);
nand (n459,n460,n497);
or (n460,n461,n485);
not (n461,n462);
nand (n462,n463,n484);
or (n463,n464,n473);
nor (n464,n465,n466);
and (n465,n88,n33);
nand (n466,n467,n469);
or (n467,n176,n468);
not (n468,n450);
nand (n469,n470,n453);
nand (n470,n471,n472);
or (n471,n42,n91);
or (n472,n90,n40);
nand (n473,n474,n477);
not (n474,n475);
nand (n475,n476,n91);
nand (n476,n33,n177);
nand (n477,n478,n480);
or (n478,n176,n479);
not (n479,n470);
nand (n480,n481,n453);
nor (n481,n482,n483);
and (n482,n36,n90);
and (n483,n91,n33);
nand (n484,n465,n466);
not (n485,n486);
nand (n486,n487,n491);
nor (n487,n488,n489);
and (n488,n454,n447);
and (n489,n490,n446);
not (n490,n454);
nor (n491,n492,n496);
and (n492,n87,n493);
nand (n493,n494,n495);
or (n494,n49,n36);
or (n495,n48,n33);
and (n496,n88,n429);
or (n497,n487,n491);
xor (n498,n424,n433);
and (n499,n445,n459);
and (n500,n422,n441);
and (n501,n396,n418);
and (n502,n306,n357);
nor (n503,n504,n529);
nor (n504,n505,n520);
xor (n505,n506,n519);
xor (n506,n507,n508);
xor (n507,n236,n252);
or (n508,n509,n518);
and (n509,n510,n517);
xor (n510,n511,n514);
nand (n511,n512,n513);
or (n512,n382,n86);
nand (n513,n88,n229);
nand (n514,n515,n516);
or (n515,n45,n390);
or (n516,n46,n272);
and (n517,n360,n366);
and (n518,n511,n514);
xor (n519,n269,n277);
or (n520,n521,n528);
and (n521,n522,n527);
xor (n522,n523,n526);
or (n523,n524,n525);
and (n524,n373,n387);
and (n525,n374,n380);
xor (n526,n279,n287);
xor (n527,n510,n517);
and (n528,n523,n526);
nor (n529,n530,n531);
xor (n530,n522,n527);
or (n531,n532,n533);
and (n532,n358,n372);
and (n533,n359,n369);
not (n534,n535);
nand (n535,n536,n541);
or (n536,n537,n539);
not (n537,n538);
nand (n538,n530,n531);
not (n539,n540);
nand (n540,n505,n520);
not (n541,n504);
nor (n542,n543,n544);
xor (n543,n265,n295);
or (n544,n545,n546);
and (n545,n506,n519);
and (n546,n507,n508);
nand (n547,n543,n544);
or (n548,n299,n10);
not (n549,n550);
nand (n550,n551,n3);
not (n551,n4);
wire s0n552,s1n552,notn552;
or (n552,s0n552,s1n552);
not(notn552,n4);
and (s0n552,notn552,n553);
and (s1n552,n4,1'b0);
wire s0n553,s1n553,notn553;
or (n553,s0n553,s1n553);
not(notn553,n3);
and (s0n553,notn553,n5);
and (s1n553,n3,n554);
xor (n554,n555,n878);
xor (n555,n556,n875);
xor (n556,n557,n874);
xor (n557,n558,n865);
xor (n558,n559,n864);
xor (n559,n560,n850);
xor (n560,n561,n849);
xor (n561,n562,n828);
xor (n562,n563,n827);
xor (n563,n564,n801);
xor (n564,n565,n800);
xor (n565,n566,n767);
xor (n566,n567,n766);
xor (n567,n568,n728);
xor (n568,n569,n727);
xor (n569,n570,n684);
xor (n570,n571,n683);
xor (n571,n572,n633);
xor (n572,n573,n632);
xor (n573,n574,n577);
xor (n574,n575,n576);
and (n575,n29,n33);
and (n576,n24,n40);
or (n577,n578,n581);
and (n578,n579,n580);
and (n579,n24,n33);
and (n580,n23,n40);
and (n581,n582,n583);
xor (n582,n579,n580);
or (n583,n584,n587);
and (n584,n585,n586);
and (n585,n23,n33);
and (n586,n158,n40);
and (n587,n588,n589);
xor (n588,n585,n586);
or (n589,n590,n593);
and (n590,n591,n592);
and (n591,n158,n33);
and (n592,n122,n40);
and (n593,n594,n595);
xor (n594,n591,n592);
or (n595,n596,n599);
and (n596,n597,n598);
and (n597,n122,n33);
and (n598,n130,n40);
and (n599,n600,n601);
xor (n600,n597,n598);
or (n601,n602,n605);
and (n602,n603,n604);
and (n603,n130,n33);
and (n604,n56,n40);
and (n605,n606,n607);
xor (n606,n603,n604);
or (n607,n608,n611);
and (n608,n609,n610);
and (n609,n56,n33);
and (n610,n50,n40);
and (n611,n612,n613);
xor (n612,n609,n610);
or (n613,n614,n616);
and (n614,n615,n431);
and (n615,n50,n33);
and (n616,n617,n618);
xor (n617,n615,n431);
or (n618,n619,n622);
and (n619,n620,n621);
and (n620,n49,n33);
and (n621,n92,n40);
and (n622,n623,n624);
xor (n623,n620,n621);
or (n624,n625,n628);
and (n625,n626,n627);
and (n626,n92,n33);
and (n627,n91,n40);
and (n628,n629,n630);
xor (n629,n626,n627);
and (n630,n483,n631);
and (n631,n177,n40);
and (n632,n23,n167);
or (n633,n634,n637);
and (n634,n635,n636);
xor (n635,n582,n583);
and (n636,n158,n167);
and (n637,n638,n639);
xor (n638,n635,n636);
or (n639,n640,n643);
and (n640,n641,n642);
xor (n641,n588,n589);
and (n642,n122,n167);
and (n643,n644,n645);
xor (n644,n641,n642);
or (n645,n646,n649);
and (n646,n647,n648);
xor (n647,n594,n595);
and (n648,n130,n167);
and (n649,n650,n651);
xor (n650,n647,n648);
or (n651,n652,n655);
and (n652,n653,n654);
xor (n653,n600,n601);
and (n654,n56,n167);
and (n655,n656,n657);
xor (n656,n653,n654);
or (n657,n658,n661);
and (n658,n659,n660);
xor (n659,n606,n607);
and (n660,n50,n167);
and (n661,n662,n663);
xor (n662,n659,n660);
or (n663,n664,n667);
and (n664,n665,n666);
xor (n665,n612,n613);
and (n666,n49,n167);
and (n667,n668,n669);
xor (n668,n665,n666);
or (n669,n670,n673);
and (n670,n671,n672);
xor (n671,n617,n618);
and (n672,n92,n167);
and (n673,n674,n675);
xor (n674,n671,n672);
or (n675,n676,n678);
and (n676,n677,n452);
xor (n677,n623,n624);
and (n678,n679,n680);
xor (n679,n677,n452);
and (n680,n681,n682);
xor (n681,n629,n630);
and (n682,n177,n167);
and (n683,n158,n124);
or (n684,n685,n688);
and (n685,n686,n687);
xor (n686,n638,n639);
and (n687,n122,n124);
and (n688,n689,n690);
xor (n689,n686,n687);
or (n690,n691,n694);
and (n691,n692,n693);
xor (n692,n644,n645);
and (n693,n130,n124);
and (n694,n695,n696);
xor (n695,n692,n693);
or (n696,n697,n700);
and (n697,n698,n699);
xor (n698,n650,n651);
and (n699,n56,n124);
and (n700,n701,n702);
xor (n701,n698,n699);
or (n702,n703,n706);
and (n703,n704,n705);
xor (n704,n656,n657);
and (n705,n50,n124);
and (n706,n707,n708);
xor (n707,n704,n705);
or (n708,n709,n711);
and (n709,n710,n350);
xor (n710,n662,n663);
and (n711,n712,n713);
xor (n712,n710,n350);
or (n713,n714,n717);
and (n714,n715,n716);
xor (n715,n668,n669);
and (n716,n92,n124);
and (n717,n718,n719);
xor (n718,n715,n716);
or (n719,n720,n722);
and (n720,n721,n438);
xor (n721,n674,n675);
and (n722,n723,n724);
xor (n723,n721,n438);
and (n724,n725,n726);
xor (n725,n679,n680);
and (n726,n177,n124);
and (n727,n122,n140);
or (n728,n729,n732);
and (n729,n730,n731);
xor (n730,n689,n690);
and (n731,n130,n140);
and (n732,n733,n734);
xor (n733,n730,n731);
or (n734,n735,n738);
and (n735,n736,n737);
xor (n736,n695,n696);
and (n737,n56,n140);
and (n738,n739,n740);
xor (n739,n736,n737);
or (n740,n741,n744);
and (n741,n742,n743);
xor (n742,n701,n702);
and (n743,n50,n140);
and (n744,n745,n746);
xor (n745,n742,n743);
or (n746,n747,n750);
and (n747,n748,n749);
xor (n748,n707,n708);
and (n749,n49,n140);
and (n750,n751,n752);
xor (n751,n748,n749);
or (n752,n753,n756);
and (n753,n754,n755);
xor (n754,n712,n713);
and (n755,n92,n140);
and (n756,n757,n758);
xor (n757,n754,n755);
or (n758,n759,n761);
and (n759,n760,n324);
xor (n760,n718,n719);
and (n761,n762,n763);
xor (n762,n760,n324);
and (n763,n764,n765);
xor (n764,n723,n724);
and (n765,n177,n140);
and (n766,n130,n188);
or (n767,n768,n771);
and (n768,n769,n770);
xor (n769,n733,n734);
and (n770,n56,n188);
and (n771,n772,n773);
xor (n772,n769,n770);
or (n773,n774,n777);
and (n774,n775,n776);
xor (n775,n739,n740);
and (n776,n50,n188);
and (n777,n778,n779);
xor (n778,n775,n776);
or (n779,n780,n783);
and (n780,n781,n782);
xor (n781,n745,n746);
and (n782,n49,n188);
and (n783,n784,n785);
xor (n784,n781,n782);
or (n785,n786,n789);
and (n786,n787,n788);
xor (n787,n751,n752);
and (n788,n92,n188);
and (n789,n790,n791);
xor (n790,n787,n788);
or (n791,n792,n795);
and (n792,n793,n794);
xor (n793,n757,n758);
and (n794,n91,n188);
and (n795,n796,n797);
xor (n796,n793,n794);
and (n797,n798,n799);
xor (n798,n762,n763);
and (n799,n177,n188);
and (n800,n56,n60);
or (n801,n802,n805);
and (n802,n803,n804);
xor (n803,n772,n773);
and (n804,n50,n60);
and (n805,n806,n807);
xor (n806,n803,n804);
or (n807,n808,n811);
and (n808,n809,n810);
xor (n809,n778,n779);
and (n810,n49,n60);
and (n811,n812,n813);
xor (n812,n809,n810);
or (n813,n814,n817);
and (n814,n815,n816);
xor (n815,n784,n785);
and (n816,n92,n60);
and (n817,n818,n819);
xor (n818,n815,n816);
or (n819,n820,n822);
and (n820,n821,n342);
xor (n821,n790,n791);
and (n822,n823,n824);
xor (n823,n821,n342);
and (n824,n825,n826);
xor (n825,n796,n797);
and (n826,n177,n60);
and (n827,n50,n66);
or (n828,n829,n832);
and (n829,n830,n831);
xor (n830,n806,n807);
and (n831,n49,n66);
and (n832,n833,n834);
xor (n833,n830,n831);
or (n834,n835,n838);
and (n835,n836,n837);
xor (n836,n812,n813);
and (n837,n92,n66);
and (n838,n839,n840);
xor (n839,n836,n837);
or (n840,n841,n844);
and (n841,n842,n843);
xor (n842,n818,n819);
and (n843,n91,n66);
and (n844,n845,n846);
xor (n845,n842,n843);
and (n846,n847,n848);
xor (n847,n823,n824);
and (n848,n177,n66);
and (n849,n49,n84);
or (n850,n851,n854);
and (n851,n852,n853);
xor (n852,n833,n834);
and (n853,n92,n84);
and (n854,n855,n856);
xor (n855,n852,n853);
or (n856,n857,n859);
and (n857,n858,n257);
xor (n858,n839,n840);
and (n859,n860,n861);
xor (n860,n858,n257);
and (n861,n862,n863);
xor (n862,n845,n846);
and (n863,n177,n84);
and (n864,n92,n102);
or (n865,n866,n869);
and (n866,n867,n868);
xor (n867,n855,n856);
and (n868,n91,n102);
and (n869,n870,n871);
xor (n870,n867,n868);
and (n871,n872,n873);
xor (n872,n860,n861);
and (n873,n177,n102);
and (n874,n91,n181);
and (n875,n876,n877);
xor (n876,n870,n871);
and (n877,n177,n181);
and (n878,n177,n213);
endmodule
