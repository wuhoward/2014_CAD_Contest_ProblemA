module top (out,n5,n21,n23,n24,n33,n34,n36,n37,n47
        ,n56,n60,n70,n71,n73,n74,n81,n87,n99,n100
        ,n102,n103,n106,n112,n124,n125,n134,n139,n167,n206
        ,n285,n291,n300,n310,n316,n1025);
output out;
input n5;
input n21;
input n23;
input n24;
input n33;
input n34;
input n36;
input n37;
input n47;
input n56;
input n60;
input n70;
input n71;
input n73;
input n74;
input n81;
input n87;
input n99;
input n100;
input n102;
input n103;
input n106;
input n112;
input n124;
input n125;
input n134;
input n139;
input n167;
input n206;
input n285;
input n291;
input n300;
input n310;
input n316;
input n1025;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n35;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n101;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
xor (out,n0,n1027);
and (n0,n1,n1026);
or (n1,n2,n1025);
nand (n2,n3,n766);
or (n3,n4,n6);
not (n4,n5);
not (n6,n7);
xor (n7,n8,n264);
and (n8,n9,n262);
not (n9,n10);
nor (n10,n11,n217);
or (n11,n12,n216);
and (n12,n13,n176);
xor (n13,n14,n90);
xor (n14,n15,n62);
xor (n15,n16,n50);
nand (n16,n17,n43);
or (n17,n18,n28);
not (n18,n19);
nor (n19,n20,n25);
and (n20,n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n5);
and (s0n22,notn22,n23);
and (s1n22,n5,n24);
and (n25,n26,n27);
not (n26,n21);
not (n27,n22);
nand (n28,n29,n40);
nor (n29,n30,n38);
and (n30,n31,n35);
not (n31,n32);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n5);
and (s0n32,notn32,n33);
and (s1n32,n5,n34);
wire s0n35,s1n35,notn35;
or (n35,s0n35,s1n35);
not(notn35,n5);
and (s0n35,notn35,n36);
and (s1n35,n5,n37);
and (n38,n32,n39);
not (n39,n35);
nand (n40,n41,n42);
or (n41,n31,n22);
nand (n42,n22,n31);
nand (n43,n44,n45);
not (n44,n29);
nor (n45,n46,n48);
and (n46,n47,n22);
and (n48,n49,n27);
not (n49,n47);
nor (n50,n51,n57);
nand (n51,n22,n52);
not (n52,n53);
wire s0n53,s1n53,notn53;
or (n53,s0n53,s1n53);
not(notn53,n5);
and (s0n53,notn53,1'b0);
and (s1n53,n5,n55);
and (n55,n56,n24);
nor (n57,n58,n61);
and (n58,n53,n59);
not (n59,n60);
and (n61,n52,n60);
nand (n62,n63,n84);
or (n63,n64,n79);
nand (n64,n65,n76);
not (n65,n66);
nand (n66,n67,n75);
or (n67,n68,n72);
not (n68,n69);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n5);
and (s0n69,notn69,n70);
and (s1n69,n5,n71);
wire s0n72,s1n72,notn72;
or (n72,s0n72,s1n72);
not(notn72,n5);
and (s0n72,notn72,n73);
and (s1n72,n5,n74);
nand (n75,n72,n68);
nand (n76,n77,n78);
or (n77,n68,n35);
nand (n78,n35,n68);
nor (n79,n80,n82);
and (n80,n39,n81);
and (n82,n35,n83);
not (n83,n81);
or (n84,n65,n85);
nor (n85,n86,n88);
and (n86,n39,n87);
and (n88,n35,n89);
not (n89,n87);
xor (n90,n91,n154);
xor (n91,n92,n140);
xor (n92,n93,n116);
nand (n93,n94,n109);
or (n94,n95,n104);
not (n95,n96);
nor (n96,n97,n101);
not (n97,n98);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n5);
and (s0n98,notn98,n99);
and (s1n98,n5,n100);
wire s0n101,s1n101,notn101;
or (n101,s0n101,s1n101);
not(notn101,n5);
and (s0n101,notn101,n102);
and (s1n101,n5,n103);
nor (n104,n105,n107);
and (n105,n97,n106);
and (n107,n98,n108);
not (n108,n106);
or (n109,n110,n115);
nor (n110,n111,n113);
and (n111,n97,n112);
and (n113,n98,n114);
not (n114,n112);
not (n115,n101);
nand (n116,n117,n137);
or (n117,n118,n131);
not (n118,n119);
and (n119,n120,n127);
nand (n120,n121,n126);
or (n121,n122,n72);
not (n122,n123);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n5);
and (s0n123,notn123,n124);
and (s1n123,n5,n125);
nand (n126,n72,n122);
not (n127,n128);
nand (n128,n129,n130);
or (n129,n122,n98);
nand (n130,n98,n122);
nor (n131,n132,n135);
and (n132,n133,n134);
not (n133,n72);
and (n135,n72,n136);
not (n136,n134);
or (n137,n138,n127);
xor (n138,n139,n133);
and (n140,n141,n148);
nand (n141,n142,n147);
or (n142,n95,n143);
nor (n143,n144,n145);
and (n144,n97,n139);
and (n145,n98,n146);
not (n146,n139);
or (n147,n104,n115);
nand (n148,n149,n153);
or (n149,n118,n150);
nor (n150,n151,n152);
and (n151,n133,n87);
and (n152,n72,n89);
or (n153,n127,n131);
or (n154,n155,n175);
and (n155,n156,n169);
xor (n156,n157,n163);
nand (n157,n158,n162);
or (n158,n159,n28);
nor (n159,n160,n161);
and (n160,n60,n27);
and (n161,n59,n22);
nand (n162,n44,n19);
nor (n163,n51,n164);
nor (n164,n165,n168);
and (n165,n53,n166);
not (n166,n167);
and (n168,n52,n167);
nand (n169,n170,n174);
or (n170,n64,n171);
nor (n171,n172,n173);
and (n172,n39,n47);
and (n173,n35,n49);
or (n174,n65,n79);
and (n175,n157,n163);
or (n176,n177,n215);
and (n177,n178,n193);
xor (n178,n179,n180);
xor (n179,n141,n148);
and (n180,n181,n187);
nand (n181,n182,n186);
or (n182,n95,n183);
nor (n183,n184,n185);
and (n184,n97,n134);
and (n185,n98,n136);
or (n186,n143,n115);
nand (n187,n188,n192);
or (n188,n118,n189);
nor (n189,n190,n191);
and (n190,n133,n81);
and (n191,n72,n83);
or (n192,n150,n127);
or (n193,n194,n214);
and (n194,n195,n208);
xor (n195,n196,n202);
nand (n196,n197,n201);
or (n197,n28,n198);
nor (n198,n199,n200);
and (n199,n27,n167);
and (n200,n22,n166);
or (n201,n29,n159);
nor (n202,n51,n203);
nor (n203,n204,n207);
and (n204,n53,n205);
not (n205,n206);
and (n207,n52,n206);
nand (n208,n209,n210);
or (n209,n171,n65);
or (n210,n64,n211);
nor (n211,n212,n213);
and (n212,n39,n21);
and (n213,n35,n26);
and (n214,n196,n202);
and (n215,n179,n180);
and (n216,n14,n90);
xor (n217,n218,n259);
xor (n218,n219,n238);
xor (n219,n220,n232);
xor (n220,n221,n228);
nand (n221,n222,n224);
or (n222,n223,n28);
not (n223,n45);
or (n224,n29,n225);
nor (n225,n226,n227);
and (n226,n27,n81);
and (n227,n22,n83);
nor (n228,n51,n229);
nor (n229,n230,n231);
and (n230,n53,n26);
and (n231,n52,n21);
nand (n232,n233,n234);
or (n233,n64,n85);
or (n234,n65,n235);
nor (n235,n236,n237);
and (n236,n39,n134);
and (n237,n35,n136);
xor (n238,n239,n256);
xor (n239,n240,n255);
xor (n240,n241,n249);
nand (n241,n242,n243);
or (n242,n95,n110);
or (n243,n244,n115);
nor (n244,n245,n247);
and (n245,n97,n246);
and (n246,n56,n112);
and (n247,n98,n248);
not (n248,n246);
nand (n249,n250,n251);
or (n250,n138,n118);
nand (n251,n128,n252);
nand (n252,n253,n254);
or (n253,n72,n108);
or (n254,n133,n106);
and (n255,n93,n116);
or (n256,n257,n258);
and (n257,n15,n62);
and (n258,n16,n50);
or (n259,n260,n261);
and (n260,n91,n154);
and (n261,n92,n140);
not (n262,n263);
and (n263,n11,n217);
nand (n264,n265,n755,n765);
nand (n265,n266,n676);
nand (n266,n267,n531,n675);
nand (n267,n268,n484);
nand (n268,n269,n483);
or (n269,n270,n438);
nor (n270,n271,n437);
and (n271,n272,n409);
not (n272,n273);
nor (n273,n274,n369);
or (n274,n275,n368);
and (n275,n276,n339);
xor (n276,n277,n320);
or (n277,n278,n319);
and (n278,n279,n306);
xor (n279,n280,n294);
nand (n280,n281,n288);
or (n281,n282,n28);
not (n282,n283);
nand (n283,n284,n286);
or (n284,n27,n285);
or (n286,n22,n287);
not (n287,n285);
or (n288,n29,n289);
nor (n289,n290,n292);
and (n290,n291,n27);
and (n292,n293,n22);
not (n293,n291);
nand (n294,n295,n302);
or (n295,n296,n118);
not (n296,n297);
nand (n297,n298,n301);
or (n298,n72,n299);
not (n299,n300);
or (n301,n133,n300);
nand (n302,n128,n303);
nor (n303,n304,n305);
and (n304,n206,n72);
and (n305,n205,n133);
nand (n306,n307,n313);
or (n307,n64,n308);
nor (n308,n309,n311);
and (n309,n39,n310);
and (n311,n35,n312);
not (n312,n310);
or (n313,n65,n314);
nor (n314,n315,n317);
and (n315,n39,n316);
and (n317,n35,n318);
not (n318,n316);
and (n319,n280,n294);
xor (n320,n321,n333);
xor (n321,n322,n324);
and (n322,n323,n285);
not (n323,n51);
nand (n324,n325,n329);
or (n325,n95,n326);
nor (n326,n327,n328);
and (n327,n59,n98);
and (n328,n60,n97);
or (n329,n330,n115);
nor (n330,n331,n332);
and (n331,n97,n21);
and (n332,n98,n26);
nand (n333,n334,n335);
or (n334,n28,n289);
or (n335,n29,n336);
nor (n336,n337,n338);
and (n337,n310,n27);
and (n338,n312,n22);
xor (n339,n340,n354);
xor (n340,n341,n348);
nand (n341,n342,n344);
or (n342,n118,n343);
not (n343,n303);
or (n344,n127,n345);
nor (n345,n346,n347);
and (n346,n133,n167);
and (n347,n72,n166);
nand (n348,n349,n350);
or (n349,n64,n314);
or (n350,n65,n351);
nor (n351,n352,n353);
and (n352,n39,n300);
and (n353,n35,n299);
and (n354,n355,n360);
nor (n355,n356,n27);
nor (n356,n357,n359);
and (n357,n39,n358);
nand (n358,n32,n285);
and (n359,n31,n287);
nand (n360,n361,n366);
or (n361,n362,n95);
not (n362,n363);
nor (n363,n364,n365);
and (n364,n167,n98);
and (n365,n166,n97);
nand (n366,n367,n101);
not (n367,n326);
and (n368,n277,n320);
xor (n369,n370,n392);
xor (n370,n371,n389);
xor (n371,n372,n383);
xor (n372,n373,n379);
nand (n373,n374,n375);
or (n374,n336,n28);
nand (n375,n376,n44);
nor (n376,n377,n378);
and (n377,n316,n22);
and (n378,n318,n27);
nor (n379,n51,n380);
nor (n380,n381,n382);
and (n381,n53,n293);
and (n382,n52,n291);
nand (n383,n384,n385);
or (n384,n95,n330);
or (n385,n386,n115);
nor (n386,n387,n388);
and (n387,n97,n47);
and (n388,n98,n49);
or (n389,n390,n391);
and (n390,n340,n354);
and (n391,n341,n348);
xor (n392,n393,n406);
xor (n393,n394,n400);
nand (n394,n395,n396);
or (n395,n64,n351);
or (n396,n65,n397);
nor (n397,n398,n399);
and (n398,n39,n206);
and (n399,n35,n205);
nand (n400,n401,n402);
or (n401,n118,n345);
or (n402,n403,n127);
nor (n403,n404,n405);
and (n404,n133,n60);
and (n405,n72,n59);
or (n406,n407,n408);
and (n407,n321,n333);
and (n408,n322,n324);
not (n409,n410);
nand (n410,n411,n412);
xor (n411,n276,n339);
or (n412,n413,n436);
and (n413,n414,n435);
xor (n414,n415,n416);
xor (n415,n355,n360);
or (n416,n417,n434);
and (n417,n418,n427);
xor (n418,n419,n420);
and (n419,n44,n285);
nand (n420,n421,n422);
or (n421,n115,n362);
nand (n422,n423,n96);
not (n423,n424);
nor (n424,n425,n426);
and (n425,n206,n97);
and (n426,n205,n98);
nand (n427,n428,n433);
or (n428,n429,n118);
not (n429,n430);
nor (n430,n431,n432);
and (n431,n316,n72);
and (n432,n133,n318);
nand (n433,n128,n297);
and (n434,n419,n420);
xor (n435,n279,n306);
and (n436,n415,n416);
and (n437,n274,n369);
nor (n438,n439,n480);
xor (n439,n440,n477);
xor (n440,n441,n460);
xor (n441,n442,n454);
xor (n442,n443,n450);
nand (n443,n444,n446);
or (n444,n445,n28);
not (n445,n376);
nand (n446,n44,n447);
nor (n447,n448,n449);
and (n448,n300,n22);
and (n449,n299,n27);
nor (n450,n51,n451);
nor (n451,n452,n453);
and (n452,n53,n312);
and (n453,n52,n310);
nand (n454,n455,n456);
or (n455,n64,n397);
or (n456,n65,n457);
nor (n457,n458,n459);
and (n458,n39,n167);
and (n459,n35,n166);
xor (n460,n461,n474);
xor (n461,n462,n468);
nand (n462,n463,n464);
or (n463,n95,n386);
or (n464,n465,n115);
nor (n465,n466,n467);
and (n466,n97,n81);
and (n467,n98,n83);
nand (n468,n469,n470);
or (n469,n118,n403);
or (n470,n471,n127);
nor (n471,n472,n473);
and (n472,n133,n21);
and (n473,n72,n26);
or (n474,n475,n476);
and (n475,n372,n383);
and (n476,n373,n379);
or (n477,n478,n479);
and (n478,n393,n406);
and (n479,n394,n400);
or (n480,n481,n482);
and (n481,n370,n392);
and (n482,n371,n389);
nand (n483,n439,n480);
nand (n484,n485,n527);
not (n485,n486);
xor (n486,n487,n526);
xor (n487,n488,n507);
xor (n488,n489,n501);
xor (n489,n490,n497);
nand (n490,n491,n493);
or (n491,n492,n28);
not (n492,n447);
nand (n493,n44,n494);
nor (n494,n495,n496);
and (n495,n206,n22);
and (n496,n205,n27);
nor (n497,n51,n498);
nor (n498,n499,n500);
and (n499,n53,n318);
and (n500,n52,n316);
nand (n501,n502,n503);
or (n502,n64,n457);
or (n503,n65,n504);
nor (n504,n505,n506);
and (n505,n39,n60);
and (n506,n35,n59);
xor (n507,n508,n523);
xor (n508,n509,n522);
xor (n509,n510,n516);
nand (n510,n511,n512);
or (n511,n95,n465);
or (n512,n513,n115);
nor (n513,n514,n515);
and (n514,n97,n87);
and (n515,n98,n89);
nand (n516,n517,n518);
or (n517,n118,n471);
or (n518,n127,n519);
nor (n519,n520,n521);
and (n520,n133,n47);
and (n521,n72,n49);
and (n522,n462,n468);
or (n523,n524,n525);
and (n524,n442,n454);
and (n525,n443,n450);
and (n526,n461,n474);
not (n527,n528);
or (n528,n529,n530);
and (n529,n440,n477);
and (n530,n441,n460);
nand (n531,n484,n532,n674);
nor (n532,n533,n671);
nor (n533,n534,n669);
and (n534,n535,n664);
or (n535,n536,n663);
and (n536,n537,n579);
xor (n537,n538,n572);
or (n538,n539,n571);
and (n539,n540,n559);
xor (n540,n541,n548);
nand (n541,n542,n547);
or (n542,n543,n118);
not (n543,n544);
nor (n544,n545,n546);
and (n545,n312,n133);
and (n546,n310,n72);
nand (n547,n128,n430);
nand (n548,n549,n554);
or (n549,n550,n65);
not (n550,n551);
nor (n551,n552,n553);
and (n552,n291,n35);
and (n553,n293,n39);
nand (n554,n555,n556);
not (n555,n64);
nand (n556,n557,n558);
or (n557,n39,n285);
or (n558,n35,n287);
xor (n559,n560,n565);
and (n560,n561,n35);
nand (n561,n562,n564);
or (n562,n72,n563);
and (n563,n285,n69);
or (n564,n69,n285);
nand (n565,n566,n570);
or (n566,n95,n567);
nor (n567,n568,n569);
and (n568,n97,n300);
and (n569,n98,n299);
or (n570,n424,n115);
and (n571,n541,n548);
xor (n572,n573,n578);
xor (n573,n574,n577);
nand (n574,n575,n576);
or (n575,n550,n64);
or (n576,n65,n308);
and (n577,n560,n565);
xor (n578,n418,n427);
or (n579,n580,n662);
and (n580,n581,n602);
xor (n581,n582,n601);
or (n582,n583,n600);
and (n583,n584,n593);
xor (n584,n585,n586);
and (n585,n66,n285);
nand (n586,n587,n592);
or (n587,n588,n118);
not (n588,n589);
nor (n589,n590,n591);
and (n590,n291,n72);
and (n591,n293,n133);
nand (n592,n544,n128);
nand (n593,n594,n599);
or (n594,n95,n595);
not (n595,n596);
nor (n596,n597,n598);
and (n597,n318,n97);
and (n598,n316,n98);
or (n599,n567,n115);
and (n600,n585,n586);
xor (n601,n540,n559);
or (n602,n603,n661);
and (n603,n604,n660);
xor (n604,n605,n619);
nor (n605,n606,n614);
not (n606,n607);
nand (n607,n608,n613);
or (n608,n609,n95);
not (n609,n610);
nand (n610,n611,n612);
or (n611,n312,n98);
nand (n612,n98,n312);
nand (n613,n596,n101);
nand (n614,n615,n72);
nand (n615,n616,n618);
or (n616,n98,n617);
and (n617,n285,n123);
or (n618,n123,n285);
nand (n619,n620,n658);
or (n620,n621,n644);
not (n621,n622);
nand (n622,n623,n643);
or (n623,n624,n633);
nor (n624,n625,n632);
nand (n625,n626,n631);
or (n626,n627,n95);
not (n627,n628);
nand (n628,n629,n630);
or (n629,n293,n98);
nand (n630,n98,n293);
nand (n631,n610,n101);
nor (n632,n127,n287);
nand (n633,n634,n641);
nand (n634,n635,n640);
or (n635,n636,n95);
not (n636,n637);
nand (n637,n638,n639);
or (n638,n97,n285);
or (n639,n98,n287);
nand (n640,n628,n101);
nor (n641,n642,n97);
and (n642,n285,n101);
nand (n643,n625,n632);
not (n644,n645);
nand (n645,n646,n654);
not (n646,n647);
nand (n647,n648,n653);
or (n648,n649,n118);
not (n649,n650);
nand (n650,n651,n652);
or (n651,n133,n285);
or (n652,n72,n287);
nand (n653,n128,n589);
nor (n654,n655,n657);
and (n655,n606,n656);
not (n656,n614);
and (n657,n607,n614);
nand (n658,n659,n647);
not (n659,n654);
xor (n660,n584,n593);
and (n661,n605,n619);
and (n662,n582,n601);
and (n663,n538,n572);
or (n664,n665,n666);
xor (n665,n414,n435);
or (n666,n667,n668);
and (n667,n573,n578);
and (n668,n574,n577);
not (n669,n670);
nand (n670,n665,n666);
nand (n671,n672,n272);
not (n672,n673);
nor (n673,n411,n412);
not (n674,n438);
nand (n675,n486,n528);
nor (n676,n677,n734);
nand (n677,n678,n727);
not (n678,n679);
nor (n679,n680,n718);
xor (n680,n681,n709);
xor (n681,n682,n683);
xor (n682,n195,n208);
xor (n683,n684,n693);
xor (n684,n685,n686);
xor (n685,n181,n187);
and (n686,n687,n690);
nand (n687,n688,n689);
or (n688,n95,n513);
or (n689,n183,n115);
nand (n690,n691,n692);
or (n691,n118,n519);
or (n692,n189,n127);
or (n693,n694,n708);
and (n694,n695,n705);
xor (n695,n696,n701);
nand (n696,n697,n699);
or (n697,n698,n28);
not (n698,n494);
nand (n699,n700,n44);
not (n700,n198);
nor (n701,n51,n702);
nor (n702,n703,n704);
and (n703,n53,n299);
and (n704,n52,n300);
nand (n705,n706,n707);
or (n706,n64,n504);
or (n707,n65,n211);
and (n708,n696,n701);
or (n709,n710,n717);
and (n710,n711,n714);
xor (n711,n712,n713);
xor (n712,n687,n690);
and (n713,n510,n516);
or (n714,n715,n716);
and (n715,n489,n501);
and (n716,n490,n497);
and (n717,n712,n713);
or (n718,n719,n726);
and (n719,n720,n723);
xor (n720,n721,n722);
xor (n721,n695,n705);
xor (n722,n711,n714);
or (n723,n724,n725);
and (n724,n508,n523);
and (n725,n509,n522);
and (n726,n721,n722);
nand (n727,n728,n730);
not (n728,n729);
xor (n729,n720,n723);
not (n730,n731);
or (n731,n732,n733);
and (n732,n487,n526);
and (n733,n488,n507);
nand (n734,n735,n748);
nand (n735,n736,n744);
not (n736,n737);
xor (n737,n738,n741);
xor (n738,n739,n740);
xor (n739,n156,n169);
xor (n740,n178,n193);
or (n741,n742,n743);
and (n742,n684,n693);
and (n743,n685,n686);
not (n744,n745);
or (n745,n746,n747);
and (n746,n681,n709);
and (n747,n682,n683);
nand (n748,n749,n751);
not (n749,n750);
xor (n750,n13,n176);
not (n751,n752);
or (n752,n753,n754);
and (n753,n738,n741);
and (n754,n739,n740);
nand (n755,n756,n748);
nand (n756,n757,n764);
or (n757,n758,n759);
not (n758,n735);
not (n759,n760);
nand (n760,n761,n763);
or (n761,n679,n762);
nand (n762,n729,n731);
nand (n763,n680,n718);
nand (n764,n737,n745);
nand (n765,n752,n750);
not (n766,n767);
and (n767,n768,n4,n56);
nand (n768,n769,n1024);
or (n769,n770,n823);
not (n770,n771);
nor (n771,n772,n822);
and (n772,n773,n811);
not (n773,n774);
or (n774,n775,n810);
and (n775,n776,n791);
xor (n776,n777,n787);
nand (n777,n778,n783);
or (n778,n779,n29);
not (n779,n780);
nand (n780,n781,n782);
or (n781,n22,n248);
or (n782,n27,n246);
or (n783,n28,n784);
nor (n784,n785,n786);
and (n785,n27,n112);
and (n786,n22,n114);
nand (n787,n788,n789,n323);
or (n788,n53,n106);
not (n789,n790);
and (n790,n106,n53);
or (n791,n792,n809);
and (n792,n793,n805);
xor (n793,n794,n799);
nand (n794,n795,n796);
or (n795,n555,n66);
nand (n796,n797,n798);
or (n797,n35,n248);
or (n798,n39,n246);
nand (n799,n800,n804);
or (n800,n28,n801);
nor (n801,n802,n803);
and (n802,n27,n106);
and (n803,n22,n108);
or (n804,n29,n784);
nor (n805,n51,n806);
nor (n806,n807,n808);
and (n807,n53,n146);
and (n808,n52,n139);
and (n809,n794,n799);
and (n810,n777,n787);
not (n811,n812);
xor (n812,n813,n821);
xor (n813,n814,n817);
nand (n814,n815,n780);
or (n815,n816,n44);
not (n816,n28);
nor (n817,n51,n818);
nor (n818,n819,n820);
and (n819,n53,n114);
and (n820,n52,n112);
not (n821,n787);
and (n822,n774,n812);
nand (n823,n824,n1001,n1023);
nand (n824,n264,n825);
and (n825,n826,n957,n996);
and (n826,n827,n879,n951);
nor (n827,n10,n828);
not (n828,n829);
nand (n829,n830,n875);
not (n830,n831);
xor (n831,n832,n851);
xor (n832,n833,n848);
xor (n833,n834,n842);
xor (n834,n835,n839);
nor (n835,n51,n836);
nor (n836,n837,n838);
and (n837,n53,n49);
and (n838,n52,n47);
nand (n839,n840,n841);
or (n840,n101,n96);
not (n841,n244);
nand (n842,n843,n847);
or (n843,n844,n65);
nor (n844,n845,n846);
and (n845,n139,n39);
and (n846,n146,n35);
or (n847,n64,n235);
or (n848,n849,n850);
and (n849,n239,n256);
and (n850,n240,n255);
xor (n851,n852,n857);
xor (n852,n853,n854);
and (n853,n241,n249);
or (n854,n855,n856);
and (n855,n220,n232);
and (n856,n221,n228);
nand (n857,n858,n874);
or (n858,n859,n867);
not (n859,n860);
nand (n860,n861,n863);
or (n861,n118,n862);
not (n862,n252);
or (n863,n127,n864);
nor (n864,n865,n866);
and (n865,n133,n112);
and (n866,n72,n114);
not (n867,n868);
nand (n868,n869,n870);
or (n869,n28,n225);
or (n870,n29,n871);
nor (n871,n872,n873);
and (n872,n27,n87);
and (n873,n22,n89);
or (n874,n868,n860);
not (n875,n876);
or (n876,n877,n878);
and (n877,n218,n259);
and (n878,n219,n238);
nand (n879,n880,n941);
not (n880,n881);
xor (n881,n882,n933);
xor (n882,n883,n903);
xor (n883,n884,n899);
xor (n884,n885,n890);
nand (n885,n886,n887);
or (n886,n119,n128);
nand (n887,n888,n889);
or (n888,n72,n248);
or (n889,n133,n246);
nand (n890,n891,n895);
or (n891,n64,n892);
nor (n892,n893,n894);
and (n893,n39,n106);
and (n894,n35,n108);
or (n895,n65,n896);
nor (n896,n897,n898);
and (n897,n39,n112);
and (n898,n35,n114);
nor (n899,n51,n900);
nor (n900,n901,n902);
and (n901,n53,n89);
and (n902,n52,n87);
xor (n903,n904,n919);
xor (n904,n905,n914);
nand (n905,n906,n910);
or (n906,n28,n907);
nor (n907,n908,n909);
and (n908,n27,n134);
and (n909,n22,n136);
or (n910,n29,n911);
nor (n911,n912,n913);
and (n912,n27,n139);
and (n913,n22,n146);
nand (n914,n915,n917);
or (n915,n916,n127);
not (n916,n887);
nand (n917,n918,n119);
not (n918,n864);
or (n919,n920,n932);
and (n920,n921,n929);
xor (n921,n922,n926);
nor (n922,n51,n923);
nor (n923,n924,n925);
and (n924,n53,n83);
and (n925,n52,n81);
nand (n926,n927,n928);
or (n927,n64,n844);
or (n928,n65,n892);
nand (n929,n930,n931);
or (n930,n28,n871);
or (n931,n29,n907);
and (n932,n922,n926);
or (n933,n934,n940);
and (n934,n935,n937);
xor (n935,n936,n874);
not (n936,n914);
or (n937,n938,n939);
and (n938,n834,n842);
and (n939,n835,n839);
and (n940,n936,n874);
not (n941,n942);
or (n942,n943,n950);
and (n943,n944,n947);
xor (n944,n945,n946);
xor (n945,n921,n929);
xor (n946,n935,n937);
or (n947,n948,n949);
and (n948,n852,n857);
and (n949,n853,n854);
and (n950,n945,n946);
not (n951,n952);
nor (n952,n953,n954);
xor (n953,n944,n947);
or (n954,n955,n956);
and (n955,n832,n851);
and (n956,n833,n848);
nor (n957,n958,n983);
nor (n958,n959,n962);
or (n959,n960,n961);
and (n960,n882,n933);
and (n961,n883,n903);
xor (n962,n963,n980);
xor (n963,n964,n967);
or (n964,n965,n966);
and (n965,n884,n899);
and (n966,n885,n890);
xor (n967,n968,n976);
xor (n968,n969,n972);
nand (n969,n970,n971);
or (n970,n28,n911);
or (n971,n29,n801);
nor (n972,n51,n973);
nor (n973,n974,n975);
and (n974,n53,n136);
and (n975,n52,n134);
nor (n976,n977,n979);
and (n977,n555,n978);
not (n978,n896);
and (n979,n66,n796);
or (n980,n981,n982);
and (n981,n904,n919);
and (n982,n905,n914);
and (n983,n984,n988);
not (n984,n985);
or (n985,n986,n987);
and (n986,n963,n980);
and (n987,n964,n967);
not (n988,n989);
xor (n989,n990,n993);
xor (n990,n991,n992);
not (n991,n976);
xor (n992,n793,n805);
or (n993,n994,n995);
and (n994,n968,n976);
and (n995,n969,n972);
or (n996,n997,n1000);
or (n997,n998,n999);
and (n998,n990,n993);
and (n999,n991,n992);
xor (n1000,n776,n791);
nand (n1001,n1002,n996);
nand (n1002,n1003,n1017);
or (n1003,n1004,n1005);
not (n1004,n957);
not (n1005,n1006);
nand (n1006,n1007,n1016);
or (n1007,n1008,n1009);
not (n1008,n879);
not (n1009,n1010);
nand (n1010,n1011,n1015);
or (n1011,n1012,n952);
nor (n1012,n1013,n1014);
and (n1013,n263,n829);
nor (n1014,n830,n875);
nand (n1015,n953,n954);
or (n1016,n880,n941);
nor (n1017,n1018,n1022);
and (n1018,n1019,n1021);
not (n1019,n1020);
nand (n1020,n959,n962);
not (n1021,n983);
nor (n1022,n984,n988);
nand (n1023,n997,n1000);
nand (n1024,n770,n823);
nand (n1026,n2,n1025);
xor (n1027,n1025,n1028);
wire s0n1028,s1n1028,notn1028;
or (n1028,s0n1028,s1n1028);
not(notn1028,n5);
and (s0n1028,notn1028,n1029);
and (s1n1028,n5,n2329);
and (n1029,n56,n1030);
xor (n1030,n1031,n1845);
xor (n1031,n1032,n2327);
xor (n1032,n1033,n1840);
xor (n1033,n1034,n2320);
xor (n1034,n1035,n1834);
xor (n1035,n1036,n2308);
xor (n1036,n1037,n1828);
xor (n1037,n1038,n2291);
xor (n1038,n1039,n1822);
xor (n1039,n1040,n2269);
xor (n1040,n1041,n1816);
xor (n1041,n1042,n2242);
xor (n1042,n1043,n1810);
xor (n1043,n1044,n2210);
xor (n1044,n1045,n1804);
xor (n1045,n1046,n2173);
xor (n1046,n1047,n1798);
xor (n1047,n1048,n2131);
xor (n1048,n1049,n1792);
xor (n1049,n1050,n2084);
xor (n1050,n1051,n1786);
xor (n1051,n1052,n2032);
xor (n1052,n1053,n1780);
xor (n1053,n1054,n1975);
xor (n1054,n1055,n1774);
xor (n1055,n1056,n1913);
xor (n1056,n1057,n1768);
xor (n1057,n1058,n1846);
xor (n1058,n1059,n790);
xor (n1059,n1060,n1760);
xor (n1060,n1061,n1759);
xor (n1061,n1062,n1671);
xor (n1062,n1063,n1670);
xor (n1063,n1064,n1572);
xor (n1064,n1065,n1571);
xor (n1065,n1066,n1469);
xor (n1066,n1067,n1468);
xor (n1067,n1068,n1361);
xor (n1068,n1069,n1360);
xor (n1069,n1070,n1081);
xor (n1070,n1071,n1080);
xor (n1071,n1072,n1079);
xor (n1072,n1073,n1078);
xor (n1073,n1074,n1077);
xor (n1074,n1075,n1076);
and (n1075,n246,n101);
and (n1076,n246,n98);
and (n1077,n1075,n1076);
and (n1078,n246,n123);
and (n1079,n1073,n1078);
and (n1080,n246,n72);
or (n1081,n1082,n1083);
and (n1082,n1071,n1080);
and (n1083,n1070,n1084);
or (n1084,n1082,n1085);
and (n1085,n1070,n1086);
or (n1086,n1082,n1087);
and (n1087,n1070,n1088);
or (n1088,n1082,n1089);
and (n1089,n1070,n1090);
or (n1090,n1091,n1275);
and (n1091,n1092,n1274);
xor (n1092,n1072,n1093);
or (n1093,n1094,n1186);
and (n1094,n1095,n1185);
xor (n1095,n1074,n1096);
or (n1096,n1077,n1097);
and (n1097,n1098,n1100);
xor (n1098,n1075,n1099);
and (n1099,n112,n98);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
and (n1102,n112,n101);
and (n1103,n106,n98);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
and (n1108,n106,n101);
and (n1109,n139,n98);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
and (n1114,n139,n101);
and (n1115,n134,n98);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
and (n1120,n134,n101);
and (n1121,n87,n98);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
and (n1126,n87,n101);
and (n1127,n81,n98);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
and (n1132,n81,n101);
and (n1133,n47,n98);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
and (n1138,n47,n101);
and (n1139,n21,n98);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
and (n1144,n21,n101);
and (n1145,n60,n98);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1151);
and (n1149,n1150,n364);
and (n1150,n60,n101);
and (n1151,n1152,n1153);
xor (n1152,n1150,n364);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
and (n1155,n167,n101);
and (n1156,n206,n98);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1163);
and (n1160,n1161,n1162);
and (n1161,n206,n101);
and (n1162,n300,n98);
and (n1163,n1164,n1165);
xor (n1164,n1161,n1162);
or (n1165,n1166,n1168);
and (n1166,n1167,n598);
and (n1167,n300,n101);
and (n1168,n1169,n1170);
xor (n1169,n1167,n598);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
and (n1172,n316,n101);
and (n1173,n310,n98);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
and (n1178,n310,n101);
and (n1179,n291,n98);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
and (n1182,n1183,n1184);
and (n1183,n291,n101);
and (n1184,n285,n98);
and (n1185,n112,n123);
and (n1186,n1187,n1188);
xor (n1187,n1095,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1098,n1100);
and (n1191,n106,n123);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1105,n1106);
and (n1197,n139,n123);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1111,n1112);
and (n1203,n134,n123);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1117,n1118);
and (n1209,n87,n123);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1123,n1124);
and (n1215,n81,n123);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1129,n1130);
and (n1221,n47,n123);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1135,n1136);
and (n1227,n21,n123);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1141,n1142);
and (n1233,n60,n123);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1147,n1148);
and (n1239,n167,n123);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1246);
and (n1243,n1244,n1245);
xor (n1244,n1152,n1153);
and (n1245,n206,n123);
and (n1246,n1247,n1248);
xor (n1247,n1244,n1245);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1158,n1159);
and (n1251,n300,n123);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1164,n1165);
and (n1257,n316,n123);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1169,n1170);
and (n1263,n310,n123);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
or (n1266,n1267,n1270);
and (n1267,n1268,n1269);
xor (n1268,n1175,n1176);
and (n1269,n291,n123);
and (n1270,n1271,n1272);
xor (n1271,n1268,n1269);
and (n1272,n1273,n617);
xor (n1273,n1181,n1182);
and (n1274,n112,n72);
and (n1275,n1276,n1277);
xor (n1276,n1092,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1187,n1188);
and (n1280,n106,n72);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1193,n1194);
and (n1286,n139,n72);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1199,n1200);
and (n1292,n134,n72);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1205,n1206);
and (n1298,n87,n72);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1211,n1212);
and (n1304,n81,n72);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1217,n1218);
and (n1310,n47,n72);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1223,n1224);
and (n1316,n21,n72);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1229,n1230);
and (n1322,n60,n72);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
or (n1325,n1326,n1329);
and (n1326,n1327,n1328);
xor (n1327,n1235,n1236);
and (n1328,n167,n72);
and (n1329,n1330,n1331);
xor (n1330,n1327,n1328);
or (n1331,n1332,n1334);
and (n1332,n1333,n304);
xor (n1333,n1241,n1242);
and (n1334,n1335,n1336);
xor (n1335,n1333,n304);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1247,n1248);
and (n1339,n300,n72);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1345);
and (n1343,n1344,n431);
xor (n1344,n1253,n1254);
and (n1345,n1346,n1347);
xor (n1346,n1344,n431);
or (n1347,n1348,n1350);
and (n1348,n1349,n546);
xor (n1349,n1259,n1260);
and (n1350,n1351,n1352);
xor (n1351,n1349,n546);
or (n1352,n1353,n1355);
and (n1353,n1354,n590);
xor (n1354,n1265,n1266);
and (n1355,n1356,n1357);
xor (n1356,n1354,n590);
and (n1357,n1358,n1359);
xor (n1358,n1271,n1272);
and (n1359,n285,n72);
and (n1360,n246,n69);
or (n1361,n1362,n1364);
and (n1362,n1363,n1360);
xor (n1363,n1070,n1084);
and (n1364,n1365,n1366);
xor (n1365,n1363,n1360);
or (n1366,n1367,n1369);
and (n1367,n1368,n1360);
xor (n1368,n1070,n1086);
and (n1369,n1370,n1371);
xor (n1370,n1368,n1360);
or (n1371,n1372,n1374);
and (n1372,n1373,n1360);
xor (n1373,n1070,n1088);
and (n1374,n1375,n1376);
xor (n1375,n1373,n1360);
or (n1376,n1377,n1380);
and (n1377,n1378,n1379);
xor (n1378,n1070,n1090);
and (n1379,n112,n69);
and (n1380,n1381,n1382);
xor (n1381,n1378,n1379);
or (n1382,n1383,n1386);
and (n1383,n1384,n1385);
xor (n1384,n1276,n1277);
and (n1385,n106,n69);
and (n1386,n1387,n1388);
xor (n1387,n1384,n1385);
or (n1388,n1389,n1392);
and (n1389,n1390,n1391);
xor (n1390,n1282,n1283);
and (n1391,n139,n69);
and (n1392,n1393,n1394);
xor (n1393,n1390,n1391);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1288,n1289);
and (n1397,n134,n69);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
or (n1400,n1401,n1404);
and (n1401,n1402,n1403);
xor (n1402,n1294,n1295);
and (n1403,n87,n69);
and (n1404,n1405,n1406);
xor (n1405,n1402,n1403);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1300,n1301);
and (n1409,n81,n69);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1306,n1307);
and (n1415,n47,n69);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1312,n1313);
and (n1421,n21,n69);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1318,n1319);
and (n1427,n60,n69);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1324,n1325);
and (n1433,n167,n69);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1330,n1331);
and (n1439,n206,n69);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1335,n1336);
and (n1445,n300,n69);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1341,n1342);
and (n1451,n316,n69);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1346,n1347);
and (n1457,n310,n69);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1351,n1352);
and (n1463,n291,n69);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
and (n1466,n1467,n563);
xor (n1467,n1356,n1357);
and (n1468,n246,n35);
or (n1469,n1470,n1472);
and (n1470,n1471,n1468);
xor (n1471,n1365,n1366);
and (n1472,n1473,n1474);
xor (n1473,n1471,n1468);
or (n1474,n1475,n1477);
and (n1475,n1476,n1468);
xor (n1476,n1370,n1371);
and (n1477,n1478,n1479);
xor (n1478,n1476,n1468);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1375,n1376);
and (n1482,n112,n35);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1381,n1382);
and (n1488,n106,n35);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1387,n1388);
and (n1494,n139,n35);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1393,n1394);
and (n1500,n134,n35);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1399,n1400);
and (n1506,n87,n35);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1405,n1406);
and (n1512,n81,n35);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1411,n1412);
and (n1518,n47,n35);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1417,n1418);
and (n1524,n21,n35);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1423,n1424);
and (n1530,n60,n35);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1429,n1430);
and (n1536,n167,n35);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1435,n1436);
and (n1542,n206,n35);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1441,n1442);
and (n1548,n300,n35);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1447,n1448);
and (n1554,n316,n35);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1453,n1454);
and (n1560,n310,n35);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1566);
and (n1564,n1565,n552);
xor (n1565,n1459,n1460);
and (n1566,n1567,n1568);
xor (n1567,n1565,n552);
and (n1568,n1569,n1570);
xor (n1569,n1465,n1466);
and (n1570,n285,n35);
and (n1571,n246,n32);
or (n1572,n1573,n1575);
and (n1573,n1574,n1571);
xor (n1574,n1473,n1474);
and (n1575,n1576,n1577);
xor (n1576,n1574,n1571);
or (n1577,n1578,n1581);
and (n1578,n1579,n1580);
xor (n1579,n1478,n1479);
and (n1580,n112,n32);
and (n1581,n1582,n1583);
xor (n1582,n1579,n1580);
or (n1583,n1584,n1587);
and (n1584,n1585,n1586);
xor (n1585,n1484,n1485);
and (n1586,n106,n32);
and (n1587,n1588,n1589);
xor (n1588,n1585,n1586);
or (n1589,n1590,n1593);
and (n1590,n1591,n1592);
xor (n1591,n1490,n1491);
and (n1592,n139,n32);
and (n1593,n1594,n1595);
xor (n1594,n1591,n1592);
or (n1595,n1596,n1599);
and (n1596,n1597,n1598);
xor (n1597,n1496,n1497);
and (n1598,n134,n32);
and (n1599,n1600,n1601);
xor (n1600,n1597,n1598);
or (n1601,n1602,n1605);
and (n1602,n1603,n1604);
xor (n1603,n1502,n1503);
and (n1604,n87,n32);
and (n1605,n1606,n1607);
xor (n1606,n1603,n1604);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1508,n1509);
and (n1610,n81,n32);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1514,n1515);
and (n1616,n47,n32);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1520,n1521);
and (n1622,n21,n32);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1526,n1527);
and (n1628,n60,n32);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1532,n1533);
and (n1634,n167,n32);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1538,n1539);
and (n1640,n206,n32);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1544,n1545);
and (n1646,n300,n32);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1550,n1551);
and (n1652,n316,n32);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1556,n1557);
and (n1658,n310,n32);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1562,n1563);
and (n1664,n291,n32);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
and (n1667,n1668,n1669);
xor (n1668,n1567,n1568);
not (n1669,n358);
and (n1670,n246,n22);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1576,n1577);
and (n1674,n112,n22);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1582,n1583);
and (n1680,n106,n22);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
xor (n1685,n1588,n1589);
and (n1686,n139,n22);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
or (n1689,n1690,n1693);
and (n1690,n1691,n1692);
xor (n1691,n1594,n1595);
and (n1692,n134,n22);
and (n1693,n1694,n1695);
xor (n1694,n1691,n1692);
or (n1695,n1696,n1699);
and (n1696,n1697,n1698);
xor (n1697,n1600,n1601);
and (n1698,n87,n22);
and (n1699,n1700,n1701);
xor (n1700,n1697,n1698);
or (n1701,n1702,n1705);
and (n1702,n1703,n1704);
xor (n1703,n1606,n1607);
and (n1704,n81,n22);
and (n1705,n1706,n1707);
xor (n1706,n1703,n1704);
or (n1707,n1708,n1710);
and (n1708,n1709,n46);
xor (n1709,n1612,n1613);
and (n1710,n1711,n1712);
xor (n1711,n1709,n46);
or (n1712,n1713,n1715);
and (n1713,n1714,n20);
xor (n1714,n1618,n1619);
and (n1715,n1716,n1717);
xor (n1716,n1714,n20);
or (n1717,n1718,n1721);
and (n1718,n1719,n1720);
xor (n1719,n1624,n1625);
and (n1720,n60,n22);
and (n1721,n1722,n1723);
xor (n1722,n1719,n1720);
or (n1723,n1724,n1727);
and (n1724,n1725,n1726);
xor (n1725,n1630,n1631);
and (n1726,n167,n22);
and (n1727,n1728,n1729);
xor (n1728,n1725,n1726);
or (n1729,n1730,n1732);
and (n1730,n1731,n495);
xor (n1731,n1636,n1637);
and (n1732,n1733,n1734);
xor (n1733,n1731,n495);
or (n1734,n1735,n1737);
and (n1735,n1736,n448);
xor (n1736,n1642,n1643);
and (n1737,n1738,n1739);
xor (n1738,n1736,n448);
or (n1739,n1740,n1742);
and (n1740,n1741,n377);
xor (n1741,n1648,n1649);
and (n1742,n1743,n1744);
xor (n1743,n1741,n377);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1654,n1655);
and (n1747,n310,n22);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
or (n1750,n1751,n1754);
and (n1751,n1752,n1753);
xor (n1752,n1660,n1661);
and (n1753,n291,n22);
and (n1754,n1755,n1756);
xor (n1755,n1752,n1753);
and (n1756,n1757,n1758);
xor (n1757,n1666,n1667);
and (n1758,n285,n22);
and (n1759,n112,n53);
or (n1760,n1761,n1763);
and (n1761,n1762,n790);
xor (n1762,n1676,n1677);
and (n1763,n1764,n1765);
xor (n1764,n1762,n790);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1682,n1683);
and (n1768,n139,n53);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1688,n1689);
and (n1774,n134,n53);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1694,n1695);
and (n1780,n87,n53);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1700,n1701);
and (n1786,n81,n53);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1706,n1707);
and (n1792,n47,n53);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1711,n1712);
and (n1798,n21,n53);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1716,n1717);
and (n1804,n60,n53);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1722,n1723);
and (n1810,n167,n53);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1728,n1729);
and (n1816,n206,n53);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1733,n1734);
and (n1822,n300,n53);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
xor (n1827,n1738,n1739);
and (n1828,n316,n53);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
or (n1831,n1832,n1835);
and (n1832,n1833,n1834);
xor (n1833,n1743,n1744);
and (n1834,n310,n53);
and (n1835,n1836,n1837);
xor (n1836,n1833,n1834);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
xor (n1839,n1749,n1750);
and (n1840,n291,n53);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
and (n1843,n1844,n1845);
xor (n1844,n1755,n1756);
and (n1845,n285,n53);
or (n1846,n1847,n1849);
and (n1847,n1848,n1768);
xor (n1848,n1764,n1765);
and (n1849,n1850,n1851);
xor (n1850,n1848,n1768);
or (n1851,n1852,n1854);
and (n1852,n1853,n1774);
xor (n1853,n1770,n1771);
and (n1854,n1855,n1856);
xor (n1855,n1853,n1774);
or (n1856,n1857,n1859);
and (n1857,n1858,n1780);
xor (n1858,n1776,n1777);
and (n1859,n1860,n1861);
xor (n1860,n1858,n1780);
or (n1861,n1862,n1864);
and (n1862,n1863,n1786);
xor (n1863,n1782,n1783);
and (n1864,n1865,n1866);
xor (n1865,n1863,n1786);
or (n1866,n1867,n1869);
and (n1867,n1868,n1792);
xor (n1868,n1788,n1789);
and (n1869,n1870,n1871);
xor (n1870,n1868,n1792);
or (n1871,n1872,n1874);
and (n1872,n1873,n1798);
xor (n1873,n1794,n1795);
and (n1874,n1875,n1876);
xor (n1875,n1873,n1798);
or (n1876,n1877,n1879);
and (n1877,n1878,n1804);
xor (n1878,n1800,n1801);
and (n1879,n1880,n1881);
xor (n1880,n1878,n1804);
or (n1881,n1882,n1884);
and (n1882,n1883,n1810);
xor (n1883,n1806,n1807);
and (n1884,n1885,n1886);
xor (n1885,n1883,n1810);
or (n1886,n1887,n1889);
and (n1887,n1888,n1816);
xor (n1888,n1812,n1813);
and (n1889,n1890,n1891);
xor (n1890,n1888,n1816);
or (n1891,n1892,n1894);
and (n1892,n1893,n1822);
xor (n1893,n1818,n1819);
and (n1894,n1895,n1896);
xor (n1895,n1893,n1822);
or (n1896,n1897,n1899);
and (n1897,n1898,n1828);
xor (n1898,n1824,n1825);
and (n1899,n1900,n1901);
xor (n1900,n1898,n1828);
or (n1901,n1902,n1904);
and (n1902,n1903,n1834);
xor (n1903,n1830,n1831);
and (n1904,n1905,n1906);
xor (n1905,n1903,n1834);
or (n1906,n1907,n1909);
and (n1907,n1908,n1840);
xor (n1908,n1836,n1837);
and (n1909,n1910,n1911);
xor (n1910,n1908,n1840);
and (n1911,n1912,n1845);
xor (n1912,n1842,n1843);
or (n1913,n1914,n1916);
and (n1914,n1915,n1774);
xor (n1915,n1850,n1851);
and (n1916,n1917,n1918);
xor (n1917,n1915,n1774);
or (n1918,n1919,n1921);
and (n1919,n1920,n1780);
xor (n1920,n1855,n1856);
and (n1921,n1922,n1923);
xor (n1922,n1920,n1780);
or (n1923,n1924,n1926);
and (n1924,n1925,n1786);
xor (n1925,n1860,n1861);
and (n1926,n1927,n1928);
xor (n1927,n1925,n1786);
or (n1928,n1929,n1931);
and (n1929,n1930,n1792);
xor (n1930,n1865,n1866);
and (n1931,n1932,n1933);
xor (n1932,n1930,n1792);
or (n1933,n1934,n1936);
and (n1934,n1935,n1798);
xor (n1935,n1870,n1871);
and (n1936,n1937,n1938);
xor (n1937,n1935,n1798);
or (n1938,n1939,n1941);
and (n1939,n1940,n1804);
xor (n1940,n1875,n1876);
and (n1941,n1942,n1943);
xor (n1942,n1940,n1804);
or (n1943,n1944,n1946);
and (n1944,n1945,n1810);
xor (n1945,n1880,n1881);
and (n1946,n1947,n1948);
xor (n1947,n1945,n1810);
or (n1948,n1949,n1951);
and (n1949,n1950,n1816);
xor (n1950,n1885,n1886);
and (n1951,n1952,n1953);
xor (n1952,n1950,n1816);
or (n1953,n1954,n1956);
and (n1954,n1955,n1822);
xor (n1955,n1890,n1891);
and (n1956,n1957,n1958);
xor (n1957,n1955,n1822);
or (n1958,n1959,n1961);
and (n1959,n1960,n1828);
xor (n1960,n1895,n1896);
and (n1961,n1962,n1963);
xor (n1962,n1960,n1828);
or (n1963,n1964,n1966);
and (n1964,n1965,n1834);
xor (n1965,n1900,n1901);
and (n1966,n1967,n1968);
xor (n1967,n1965,n1834);
or (n1968,n1969,n1971);
and (n1969,n1970,n1840);
xor (n1970,n1905,n1906);
and (n1971,n1972,n1973);
xor (n1972,n1970,n1840);
and (n1973,n1974,n1845);
xor (n1974,n1910,n1911);
or (n1975,n1976,n1978);
and (n1976,n1977,n1780);
xor (n1977,n1917,n1918);
and (n1978,n1979,n1980);
xor (n1979,n1977,n1780);
or (n1980,n1981,n1983);
and (n1981,n1982,n1786);
xor (n1982,n1922,n1923);
and (n1983,n1984,n1985);
xor (n1984,n1982,n1786);
or (n1985,n1986,n1988);
and (n1986,n1987,n1792);
xor (n1987,n1927,n1928);
and (n1988,n1989,n1990);
xor (n1989,n1987,n1792);
or (n1990,n1991,n1993);
and (n1991,n1992,n1798);
xor (n1992,n1932,n1933);
and (n1993,n1994,n1995);
xor (n1994,n1992,n1798);
or (n1995,n1996,n1998);
and (n1996,n1997,n1804);
xor (n1997,n1937,n1938);
and (n1998,n1999,n2000);
xor (n1999,n1997,n1804);
or (n2000,n2001,n2003);
and (n2001,n2002,n1810);
xor (n2002,n1942,n1943);
and (n2003,n2004,n2005);
xor (n2004,n2002,n1810);
or (n2005,n2006,n2008);
and (n2006,n2007,n1816);
xor (n2007,n1947,n1948);
and (n2008,n2009,n2010);
xor (n2009,n2007,n1816);
or (n2010,n2011,n2013);
and (n2011,n2012,n1822);
xor (n2012,n1952,n1953);
and (n2013,n2014,n2015);
xor (n2014,n2012,n1822);
or (n2015,n2016,n2018);
and (n2016,n2017,n1828);
xor (n2017,n1957,n1958);
and (n2018,n2019,n2020);
xor (n2019,n2017,n1828);
or (n2020,n2021,n2023);
and (n2021,n2022,n1834);
xor (n2022,n1962,n1963);
and (n2023,n2024,n2025);
xor (n2024,n2022,n1834);
or (n2025,n2026,n2028);
and (n2026,n2027,n1840);
xor (n2027,n1967,n1968);
and (n2028,n2029,n2030);
xor (n2029,n2027,n1840);
and (n2030,n2031,n1845);
xor (n2031,n1972,n1973);
or (n2032,n2033,n2035);
and (n2033,n2034,n1786);
xor (n2034,n1979,n1980);
and (n2035,n2036,n2037);
xor (n2036,n2034,n1786);
or (n2037,n2038,n2040);
and (n2038,n2039,n1792);
xor (n2039,n1984,n1985);
and (n2040,n2041,n2042);
xor (n2041,n2039,n1792);
or (n2042,n2043,n2045);
and (n2043,n2044,n1798);
xor (n2044,n1989,n1990);
and (n2045,n2046,n2047);
xor (n2046,n2044,n1798);
or (n2047,n2048,n2050);
and (n2048,n2049,n1804);
xor (n2049,n1994,n1995);
and (n2050,n2051,n2052);
xor (n2051,n2049,n1804);
or (n2052,n2053,n2055);
and (n2053,n2054,n1810);
xor (n2054,n1999,n2000);
and (n2055,n2056,n2057);
xor (n2056,n2054,n1810);
or (n2057,n2058,n2060);
and (n2058,n2059,n1816);
xor (n2059,n2004,n2005);
and (n2060,n2061,n2062);
xor (n2061,n2059,n1816);
or (n2062,n2063,n2065);
and (n2063,n2064,n1822);
xor (n2064,n2009,n2010);
and (n2065,n2066,n2067);
xor (n2066,n2064,n1822);
or (n2067,n2068,n2070);
and (n2068,n2069,n1828);
xor (n2069,n2014,n2015);
and (n2070,n2071,n2072);
xor (n2071,n2069,n1828);
or (n2072,n2073,n2075);
and (n2073,n2074,n1834);
xor (n2074,n2019,n2020);
and (n2075,n2076,n2077);
xor (n2076,n2074,n1834);
or (n2077,n2078,n2080);
and (n2078,n2079,n1840);
xor (n2079,n2024,n2025);
and (n2080,n2081,n2082);
xor (n2081,n2079,n1840);
and (n2082,n2083,n1845);
xor (n2083,n2029,n2030);
or (n2084,n2085,n2087);
and (n2085,n2086,n1792);
xor (n2086,n2036,n2037);
and (n2087,n2088,n2089);
xor (n2088,n2086,n1792);
or (n2089,n2090,n2092);
and (n2090,n2091,n1798);
xor (n2091,n2041,n2042);
and (n2092,n2093,n2094);
xor (n2093,n2091,n1798);
or (n2094,n2095,n2097);
and (n2095,n2096,n1804);
xor (n2096,n2046,n2047);
and (n2097,n2098,n2099);
xor (n2098,n2096,n1804);
or (n2099,n2100,n2102);
and (n2100,n2101,n1810);
xor (n2101,n2051,n2052);
and (n2102,n2103,n2104);
xor (n2103,n2101,n1810);
or (n2104,n2105,n2107);
and (n2105,n2106,n1816);
xor (n2106,n2056,n2057);
and (n2107,n2108,n2109);
xor (n2108,n2106,n1816);
or (n2109,n2110,n2112);
and (n2110,n2111,n1822);
xor (n2111,n2061,n2062);
and (n2112,n2113,n2114);
xor (n2113,n2111,n1822);
or (n2114,n2115,n2117);
and (n2115,n2116,n1828);
xor (n2116,n2066,n2067);
and (n2117,n2118,n2119);
xor (n2118,n2116,n1828);
or (n2119,n2120,n2122);
and (n2120,n2121,n1834);
xor (n2121,n2071,n2072);
and (n2122,n2123,n2124);
xor (n2123,n2121,n1834);
or (n2124,n2125,n2127);
and (n2125,n2126,n1840);
xor (n2126,n2076,n2077);
and (n2127,n2128,n2129);
xor (n2128,n2126,n1840);
and (n2129,n2130,n1845);
xor (n2130,n2081,n2082);
or (n2131,n2132,n2134);
and (n2132,n2133,n1798);
xor (n2133,n2088,n2089);
and (n2134,n2135,n2136);
xor (n2135,n2133,n1798);
or (n2136,n2137,n2139);
and (n2137,n2138,n1804);
xor (n2138,n2093,n2094);
and (n2139,n2140,n2141);
xor (n2140,n2138,n1804);
or (n2141,n2142,n2144);
and (n2142,n2143,n1810);
xor (n2143,n2098,n2099);
and (n2144,n2145,n2146);
xor (n2145,n2143,n1810);
or (n2146,n2147,n2149);
and (n2147,n2148,n1816);
xor (n2148,n2103,n2104);
and (n2149,n2150,n2151);
xor (n2150,n2148,n1816);
or (n2151,n2152,n2154);
and (n2152,n2153,n1822);
xor (n2153,n2108,n2109);
and (n2154,n2155,n2156);
xor (n2155,n2153,n1822);
or (n2156,n2157,n2159);
and (n2157,n2158,n1828);
xor (n2158,n2113,n2114);
and (n2159,n2160,n2161);
xor (n2160,n2158,n1828);
or (n2161,n2162,n2164);
and (n2162,n2163,n1834);
xor (n2163,n2118,n2119);
and (n2164,n2165,n2166);
xor (n2165,n2163,n1834);
or (n2166,n2167,n2169);
and (n2167,n2168,n1840);
xor (n2168,n2123,n2124);
and (n2169,n2170,n2171);
xor (n2170,n2168,n1840);
and (n2171,n2172,n1845);
xor (n2172,n2128,n2129);
or (n2173,n2174,n2176);
and (n2174,n2175,n1804);
xor (n2175,n2135,n2136);
and (n2176,n2177,n2178);
xor (n2177,n2175,n1804);
or (n2178,n2179,n2181);
and (n2179,n2180,n1810);
xor (n2180,n2140,n2141);
and (n2181,n2182,n2183);
xor (n2182,n2180,n1810);
or (n2183,n2184,n2186);
and (n2184,n2185,n1816);
xor (n2185,n2145,n2146);
and (n2186,n2187,n2188);
xor (n2187,n2185,n1816);
or (n2188,n2189,n2191);
and (n2189,n2190,n1822);
xor (n2190,n2150,n2151);
and (n2191,n2192,n2193);
xor (n2192,n2190,n1822);
or (n2193,n2194,n2196);
and (n2194,n2195,n1828);
xor (n2195,n2155,n2156);
and (n2196,n2197,n2198);
xor (n2197,n2195,n1828);
or (n2198,n2199,n2201);
and (n2199,n2200,n1834);
xor (n2200,n2160,n2161);
and (n2201,n2202,n2203);
xor (n2202,n2200,n1834);
or (n2203,n2204,n2206);
and (n2204,n2205,n1840);
xor (n2205,n2165,n2166);
and (n2206,n2207,n2208);
xor (n2207,n2205,n1840);
and (n2208,n2209,n1845);
xor (n2209,n2170,n2171);
or (n2210,n2211,n2213);
and (n2211,n2212,n1810);
xor (n2212,n2177,n2178);
and (n2213,n2214,n2215);
xor (n2214,n2212,n1810);
or (n2215,n2216,n2218);
and (n2216,n2217,n1816);
xor (n2217,n2182,n2183);
and (n2218,n2219,n2220);
xor (n2219,n2217,n1816);
or (n2220,n2221,n2223);
and (n2221,n2222,n1822);
xor (n2222,n2187,n2188);
and (n2223,n2224,n2225);
xor (n2224,n2222,n1822);
or (n2225,n2226,n2228);
and (n2226,n2227,n1828);
xor (n2227,n2192,n2193);
and (n2228,n2229,n2230);
xor (n2229,n2227,n1828);
or (n2230,n2231,n2233);
and (n2231,n2232,n1834);
xor (n2232,n2197,n2198);
and (n2233,n2234,n2235);
xor (n2234,n2232,n1834);
or (n2235,n2236,n2238);
and (n2236,n2237,n1840);
xor (n2237,n2202,n2203);
and (n2238,n2239,n2240);
xor (n2239,n2237,n1840);
and (n2240,n2241,n1845);
xor (n2241,n2207,n2208);
or (n2242,n2243,n2245);
and (n2243,n2244,n1816);
xor (n2244,n2214,n2215);
and (n2245,n2246,n2247);
xor (n2246,n2244,n1816);
or (n2247,n2248,n2250);
and (n2248,n2249,n1822);
xor (n2249,n2219,n2220);
and (n2250,n2251,n2252);
xor (n2251,n2249,n1822);
or (n2252,n2253,n2255);
and (n2253,n2254,n1828);
xor (n2254,n2224,n2225);
and (n2255,n2256,n2257);
xor (n2256,n2254,n1828);
or (n2257,n2258,n2260);
and (n2258,n2259,n1834);
xor (n2259,n2229,n2230);
and (n2260,n2261,n2262);
xor (n2261,n2259,n1834);
or (n2262,n2263,n2265);
and (n2263,n2264,n1840);
xor (n2264,n2234,n2235);
and (n2265,n2266,n2267);
xor (n2266,n2264,n1840);
and (n2267,n2268,n1845);
xor (n2268,n2239,n2240);
or (n2269,n2270,n2272);
and (n2270,n2271,n1822);
xor (n2271,n2246,n2247);
and (n2272,n2273,n2274);
xor (n2273,n2271,n1822);
or (n2274,n2275,n2277);
and (n2275,n2276,n1828);
xor (n2276,n2251,n2252);
and (n2277,n2278,n2279);
xor (n2278,n2276,n1828);
or (n2279,n2280,n2282);
and (n2280,n2281,n1834);
xor (n2281,n2256,n2257);
and (n2282,n2283,n2284);
xor (n2283,n2281,n1834);
or (n2284,n2285,n2287);
and (n2285,n2286,n1840);
xor (n2286,n2261,n2262);
and (n2287,n2288,n2289);
xor (n2288,n2286,n1840);
and (n2289,n2290,n1845);
xor (n2290,n2266,n2267);
or (n2291,n2292,n2294);
and (n2292,n2293,n1828);
xor (n2293,n2273,n2274);
and (n2294,n2295,n2296);
xor (n2295,n2293,n1828);
or (n2296,n2297,n2299);
and (n2297,n2298,n1834);
xor (n2298,n2278,n2279);
and (n2299,n2300,n2301);
xor (n2300,n2298,n1834);
or (n2301,n2302,n2304);
and (n2302,n2303,n1840);
xor (n2303,n2283,n2284);
and (n2304,n2305,n2306);
xor (n2305,n2303,n1840);
and (n2306,n2307,n1845);
xor (n2307,n2288,n2289);
or (n2308,n2309,n2311);
and (n2309,n2310,n1834);
xor (n2310,n2295,n2296);
and (n2311,n2312,n2313);
xor (n2312,n2310,n1834);
or (n2313,n2314,n2316);
and (n2314,n2315,n1840);
xor (n2315,n2300,n2301);
and (n2316,n2317,n2318);
xor (n2317,n2315,n1840);
and (n2318,n2319,n1845);
xor (n2319,n2305,n2306);
or (n2320,n2321,n2323);
and (n2321,n2322,n1840);
xor (n2322,n2312,n2313);
and (n2323,n2324,n2325);
xor (n2324,n2322,n1840);
and (n2325,n2326,n1845);
xor (n2326,n2317,n2318);
and (n2327,n2328,n1845);
xor (n2328,n2324,n2325);
xor (n2329,n2241,n1845);
endmodule
