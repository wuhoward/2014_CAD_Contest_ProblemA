module top (out,n16,n18,n19,n21,n24,n28,n30,n32,n35
        ,n39,n41,n43,n46,n52,n54,n56,n59,n63,n65
        ,n67,n70,n75,n77,n78,n92,n106,n107,n179,n188
        ,n189,n225,n297,n327,n328,n631,n635,n637,n663,n664
        ,n771,n788,n789,n975,n979,n981,n992,n1004,n1018);
output out;
input n16;
input n18;
input n19;
input n21;
input n24;
input n28;
input n30;
input n32;
input n35;
input n39;
input n41;
input n43;
input n46;
input n52;
input n54;
input n56;
input n59;
input n63;
input n65;
input n67;
input n70;
input n75;
input n77;
input n78;
input n92;
input n106;
input n107;
input n179;
input n188;
input n189;
input n225;
input n297;
input n327;
input n328;
input n631;
input n635;
input n637;
input n663;
input n664;
input n771;
input n788;
input n789;
input n975;
input n979;
input n981;
input n992;
input n1004;
input n1018;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n17;
wire n20;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n40;
wire n42;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n64;
wire n66;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n632;
wire n633;
wire n634;
wire n636;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n976;
wire n977;
wire n978;
wire n980;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
xor (out,n0,n2962);
xnor (n0,n1,n2914);
nand (n1,n2,n952);
nor (n2,n3,n937);
nor (n3,n4,n530);
nand (n4,n5,n425);
nor (n5,n6,n370);
nor (n6,n7,n247);
xor (n7,n8,n204);
xor (n8,n9,n95);
xor (n9,n10,n82);
xor (n10,n11,n47);
xor (n11,n12,n36);
xor (n12,n13,n25);
xor (n13,n14,n24);
or (n14,n15,n20);
and (n15,n16,n17);
xor (n17,n18,n19);
and (n20,n21,n22);
nor (n22,n17,n23);
xnor (n23,n24,n18);
xor (n25,n26,n35);
or (n26,n27,n31);
and (n27,n28,n29);
xor (n29,n30,n24);
and (n31,n32,n33);
nor (n33,n29,n34);
xnor (n34,n35,n30);
xor (n36,n37,n46);
or (n37,n38,n42);
and (n38,n39,n40);
xor (n40,n41,n35);
and (n42,n43,n44);
nor (n44,n40,n45);
xnor (n45,n46,n41);
xor (n47,n48,n71);
xor (n48,n49,n60);
xor (n49,n50,n59);
or (n50,n51,n55);
and (n51,n52,n53);
xor (n53,n54,n46);
and (n55,n56,n57);
nor (n57,n53,n58);
xnor (n58,n59,n54);
xor (n60,n61,n70);
or (n61,n62,n66);
and (n62,n63,n64);
xor (n64,n65,n59);
and (n66,n67,n68);
nor (n68,n64,n69);
xnor (n69,n70,n65);
not (n71,n72);
xor (n72,n73,n19);
or (n73,n74,n79);
and (n74,n75,n76);
xor (n76,n77,n78);
and (n79,n75,n80);
nor (n80,n76,n81);
xnor (n81,n19,n77);
nand (n82,n83,n93,n94);
nand (n83,n84,n88);
xor (n84,n85,n59);
or (n85,n86,n87);
and (n86,n56,n53);
and (n87,n63,n57);
xor (n88,n89,n70);
or (n89,n90,n91);
and (n90,n67,n64);
and (n91,n92,n68);
nand (n93,n70,n88);
nand (n94,n84,n70);
xor (n95,n96,n166);
xor (n96,n97,n132);
xor (n97,n98,n120);
xor (n98,n70,n99);
nand (n99,n100,n114,n119);
nand (n100,n101,n111);
not (n101,n102);
xor (n102,n103,n78);
or (n103,n104,n108);
and (n104,n75,n105);
xor (n105,n106,n107);
and (n108,n75,n109);
nor (n109,n105,n110);
xnor (n110,n78,n106);
xor (n111,n112,n19);
or (n112,n74,n113);
and (n113,n16,n80);
nand (n114,n115,n111);
xor (n115,n116,n35);
or (n116,n117,n118);
and (n117,n32,n29);
and (n118,n39,n33);
nand (n119,n101,n115);
nand (n120,n121,n126,n131);
nand (n121,n122,n102);
xor (n122,n123,n24);
or (n123,n124,n125);
and (n124,n21,n17);
and (n125,n28,n22);
nand (n126,n127,n102);
xor (n127,n128,n46);
or (n128,n129,n130);
and (n129,n43,n40);
and (n130,n52,n44);
nand (n131,n122,n127);
nand (n132,n133,n152,n165);
nand (n133,n134,n136);
xor (n134,n135,n115);
xor (n135,n101,n111);
nand (n136,n137,n146,n151);
nand (n137,n138,n142);
xor (n138,n139,n19);
or (n139,n140,n141);
and (n140,n16,n76);
and (n141,n21,n80);
xor (n142,n143,n35);
or (n143,n144,n145);
and (n144,n39,n29);
and (n145,n43,n33);
nand (n146,n147,n142);
xor (n147,n148,n24);
or (n148,n149,n150);
and (n149,n28,n17);
and (n150,n32,n22);
nand (n151,n138,n147);
nand (n152,n153,n136);
nand (n153,n154,n159,n164);
nand (n154,n101,n155);
xor (n155,n156,n46);
or (n156,n157,n158);
and (n157,n52,n40);
and (n158,n56,n44);
nand (n159,n160,n155);
xor (n160,n161,n59);
or (n161,n162,n163);
and (n162,n63,n53);
and (n163,n67,n57);
nand (n164,n101,n160);
nand (n165,n134,n153);
nand (n166,n167,n172,n203);
nand (n167,n168,n170);
xor (n168,n169,n70);
xor (n169,n84,n88);
xor (n170,n171,n127);
xor (n171,n122,n102);
nand (n172,n173,n170);
nand (n173,n174,n180,n202);
nand (n174,n175,n70);
xor (n175,n176,n70);
or (n176,n177,n178);
and (n177,n92,n64);
and (n178,n179,n68);
nand (n180,n181,n70);
nand (n181,n182,n196,n201);
nand (n182,n183,n193);
not (n183,n184);
xor (n184,n185,n107);
or (n185,n186,n190);
and (n186,n75,n187);
xor (n187,n188,n189);
and (n190,n75,n191);
nor (n191,n187,n192);
xnor (n192,n107,n188);
xor (n193,n194,n78);
or (n194,n104,n195);
and (n195,n16,n109);
nand (n196,n197,n193);
xor (n197,n198,n19);
or (n198,n199,n200);
and (n199,n21,n76);
and (n200,n28,n80);
nand (n201,n183,n197);
nand (n202,n175,n181);
nand (n203,n168,n173);
nand (n204,n205,n243,n246);
nand (n205,n206,n241);
nand (n206,n207,n227,n240);
nand (n207,n208,n210);
xor (n208,n209,n147);
xor (n209,n138,n142);
nand (n210,n211,n220,n226);
nand (n211,n212,n216);
xor (n212,n213,n24);
or (n213,n214,n215);
and (n214,n32,n17);
and (n215,n39,n22);
xor (n216,n217,n35);
or (n217,n218,n219);
and (n218,n43,n29);
and (n219,n52,n33);
nand (n220,n221,n216);
xor (n221,n222,n70);
or (n222,n223,n224);
and (n223,n179,n64);
and (n224,n225,n68);
nand (n226,n212,n221);
nand (n227,n228,n210);
nand (n228,n229,n234,n239);
nand (n229,n184,n230);
xor (n230,n231,n46);
or (n231,n232,n233);
and (n232,n56,n40);
and (n233,n63,n44);
nand (n234,n235,n230);
xor (n235,n236,n59);
or (n236,n237,n238);
and (n237,n67,n53);
and (n238,n92,n57);
nand (n239,n184,n235);
nand (n240,n208,n228);
xor (n241,n242,n153);
xor (n242,n134,n136);
nand (n243,n244,n241);
xor (n244,n245,n173);
xor (n245,n168,n170);
nand (n246,n206,n244);
nand (n247,n248,n280,n369);
nand (n248,n249,n278);
nand (n249,n250,n254,n277);
nand (n250,n251,n253);
xor (n251,n252,n160);
xor (n252,n101,n155);
xor (n253,n176,n181);
nand (n254,n255,n253);
nand (n255,n256,n259,n276);
nand (n256,n70,n257);
xor (n257,n258,n197);
xor (n258,n183,n193);
nand (n259,n260,n257);
nand (n260,n261,n270,n275);
nand (n261,n262,n266);
xor (n262,n263,n78);
or (n263,n264,n265);
and (n264,n16,n105);
and (n265,n21,n109);
xor (n266,n267,n19);
or (n267,n268,n269);
and (n268,n28,n76);
and (n269,n32,n80);
nand (n270,n271,n266);
xor (n271,n272,n24);
or (n272,n273,n274);
and (n273,n39,n17);
and (n274,n43,n22);
nand (n275,n262,n271);
nand (n276,n70,n260);
nand (n277,n251,n255);
xor (n278,n279,n244);
xor (n279,n206,n241);
nand (n280,n281,n278);
nand (n281,n282,n306,n368);
nand (n282,n283,n285);
xor (n283,n284,n228);
xor (n284,n208,n210);
nand (n285,n286,n302,n305);
nand (n286,n287,n300);
nand (n287,n288,n298,n299);
nand (n288,n289,n293);
xor (n289,n290,n35);
or (n290,n291,n292);
and (n291,n52,n29);
and (n292,n56,n33);
xor (n293,n294,n70);
or (n294,n295,n296);
and (n295,n225,n64);
and (n296,n297,n68);
nand (n298,n183,n293);
nand (n299,n289,n183);
xor (n300,n301,n221);
xor (n301,n212,n216);
nand (n302,n303,n300);
xor (n303,n304,n235);
xor (n304,n184,n230);
nand (n305,n287,n303);
nand (n306,n307,n285);
nand (n307,n308,n364,n367);
nand (n308,n309,n342);
nand (n309,n310,n319,n341);
nand (n310,n311,n315);
xor (n311,n312,n46);
or (n312,n313,n314);
and (n313,n63,n40);
and (n314,n67,n44);
xor (n315,n316,n59);
or (n316,n317,n318);
and (n317,n92,n53);
and (n318,n179,n57);
nand (n319,n320,n315);
nand (n320,n321,n335,n340);
nand (n321,n322,n332);
not (n322,n323);
xor (n323,n324,n189);
or (n324,n325,n329);
and (n325,n75,n326);
xor (n326,n327,n328);
and (n329,n75,n330);
nor (n330,n326,n331);
xnor (n331,n189,n327);
xor (n332,n333,n107);
or (n333,n186,n334);
and (n334,n16,n191);
nand (n335,n336,n332);
xor (n336,n337,n19);
or (n337,n338,n339);
and (n338,n32,n76);
and (n339,n39,n80);
nand (n340,n322,n336);
nand (n341,n311,n320);
nand (n342,n343,n346,n363);
nand (n343,n70,n344);
xor (n344,n345,n271);
xor (n345,n262,n266);
nand (n346,n347,n344);
nand (n347,n348,n357,n362);
nand (n348,n349,n353);
xor (n349,n350,n78);
or (n350,n351,n352);
and (n351,n21,n105);
and (n352,n28,n109);
xor (n353,n354,n24);
or (n354,n355,n356);
and (n355,n43,n17);
and (n356,n52,n22);
nand (n357,n358,n353);
xor (n358,n359,n35);
or (n359,n360,n361);
and (n360,n56,n29);
and (n361,n63,n33);
nand (n362,n349,n358);
nand (n363,n70,n347);
nand (n364,n365,n342);
xor (n365,n366,n260);
xor (n366,n70,n257);
nand (n367,n309,n365);
nand (n368,n283,n307);
nand (n369,n249,n281);
nor (n370,n371,n375);
nand (n371,n372,n373,n374);
nand (n372,n9,n95);
nand (n373,n204,n95);
nand (n374,n9,n204);
xor (n375,n376,n421);
xor (n376,n377,n381);
nand (n377,n378,n379,n380);
nand (n378,n11,n47);
nand (n379,n82,n47);
nand (n380,n11,n82);
xor (n381,n382,n395);
xor (n382,n383,n387);
nand (n383,n384,n385,n386);
nand (n384,n70,n99);
nand (n385,n120,n99);
nand (n386,n70,n120);
xor (n387,n388,n391);
or (n388,n389,n390);
and (n389,n56,n64);
and (n390,n63,n68);
nand (n391,n392,n393,n394);
nand (n392,n13,n25);
nand (n393,n36,n25);
nand (n394,n13,n36);
xor (n395,n396,n411);
xor (n396,n397,n401);
nand (n397,n398,n399,n400);
nand (n398,n49,n60);
nand (n399,n71,n60);
nand (n400,n49,n71);
xor (n401,n402,n407);
xor (n402,n71,n403);
xor (n403,n404,n24);
or (n404,n405,n406);
and (n405,n75,n17);
and (n406,n16,n22);
xor (n407,n408,n35);
or (n408,n409,n410);
and (n409,n21,n29);
and (n410,n28,n33);
xor (n411,n412,n417);
xor (n412,n413,n72);
xor (n413,n414,n46);
or (n414,n415,n416);
and (n415,n32,n40);
and (n416,n39,n44);
xor (n417,n418,n59);
or (n418,n419,n420);
and (n419,n43,n53);
and (n420,n52,n57);
nand (n421,n422,n423,n424);
nand (n422,n97,n132);
nand (n423,n166,n132);
nand (n424,n97,n166);
nor (n425,n426,n482);
nor (n426,n427,n431);
nand (n427,n428,n429,n430);
nand (n428,n377,n381);
nand (n429,n421,n381);
nand (n430,n377,n421);
xor (n431,n432,n478);
xor (n432,n433,n456);
xor (n433,n434,n443);
xor (n434,n435,n439);
nand (n435,n436,n437,n438);
nand (n436,n71,n403);
nand (n437,n407,n403);
nand (n438,n71,n407);
nand (n439,n440,n441,n442);
nand (n440,n413,n72);
nand (n441,n417,n72);
nand (n442,n413,n417);
xor (n443,n444,n452);
xor (n444,n445,n448);
xor (n445,n446,n24);
or (n446,n405,n447);
and (n447,n75,n22);
xor (n448,n449,n59);
or (n449,n450,n451);
and (n450,n39,n53);
and (n451,n43,n57);
xor (n452,n453,n70);
or (n453,n454,n455);
and (n454,n52,n64);
and (n455,n56,n68);
xor (n456,n457,n474);
xor (n457,n458,n469);
xor (n458,n459,n70);
xor (n459,n460,n464);
xor (n460,n461,n46);
or (n461,n462,n463);
and (n462,n28,n40);
and (n463,n32,n44);
not (n464,n465);
xor (n465,n466,n35);
or (n466,n467,n468);
and (n467,n16,n29);
and (n468,n21,n33);
nand (n469,n470,n472,n473);
nand (n470,n471,n70);
xor (n471,n388,n70);
nand (n472,n391,n70);
nand (n473,n471,n391);
nand (n474,n475,n476,n477);
nand (n475,n397,n401);
nand (n476,n411,n401);
nand (n477,n397,n411);
nand (n478,n479,n480,n481);
nand (n479,n383,n387);
nand (n480,n395,n387);
nand (n481,n383,n395);
nor (n482,n483,n487);
nand (n483,n484,n485,n486);
nand (n484,n433,n456);
nand (n485,n478,n456);
nand (n486,n433,n478);
xor (n487,n488,n526);
xor (n488,n489,n493);
nand (n489,n490,n491,n492);
nand (n490,n435,n439);
nand (n491,n443,n439);
nand (n492,n435,n443);
xor (n493,n494,n509);
xor (n494,n495,n499);
nand (n495,n496,n497,n498);
nand (n496,n460,n464);
nand (n497,n70,n464);
nand (n498,n460,n70);
xor (n499,n500,n70);
xor (n500,n501,n505);
xor (n501,n502,n70);
or (n502,n503,n504);
and (n503,n43,n64);
and (n504,n52,n68);
xor (n505,n506,n46);
or (n506,n507,n508);
and (n507,n21,n40);
and (n508,n28,n44);
xor (n509,n510,n515);
xor (n510,n465,n511);
nand (n511,n512,n513,n514);
nand (n512,n445,n448);
nand (n513,n452,n448);
nand (n514,n445,n452);
xor (n515,n516,n522);
xor (n516,n517,n518);
not (n517,n445);
xor (n518,n519,n35);
or (n519,n520,n521);
and (n520,n75,n29);
and (n521,n16,n33);
xor (n522,n523,n59);
or (n523,n524,n525);
and (n524,n32,n53);
and (n525,n39,n57);
nand (n526,n527,n528,n529);
nand (n527,n458,n469);
nand (n528,n474,n469);
nand (n529,n458,n474);
nor (n530,n531,n931);
nor (n531,n532,n907);
nor (n532,n533,n905);
nor (n533,n534,n880);
nand (n534,n535,n842);
nand (n535,n536,n758,n841);
nand (n536,n537,n621);
xor (n537,n538,n611);
xor (n538,n539,n561);
xor (n539,n540,n545);
xor (n540,n541,n70);
xor (n541,n542,n46);
or (n542,n543,n544);
and (n543,n67,n40);
and (n544,n92,n44);
nand (n545,n546,n555,n560);
nand (n546,n547,n551);
xor (n547,n548,n19);
or (n548,n549,n550);
and (n549,n39,n76);
and (n550,n43,n80);
xor (n551,n552,n107);
or (n552,n553,n554);
and (n553,n16,n187);
and (n554,n21,n191);
nand (n555,n556,n551);
xor (n556,n557,n78);
or (n557,n558,n559);
and (n558,n28,n105);
and (n559,n32,n109);
nand (n560,n547,n556);
nand (n561,n562,n593,n610);
nand (n562,n563,n579);
nand (n563,n564,n573,n578);
nand (n564,n565,n569);
xor (n565,n566,n19);
or (n566,n567,n568);
and (n567,n43,n76);
and (n568,n52,n80);
xor (n569,n570,n107);
or (n570,n571,n572);
and (n571,n21,n187);
and (n572,n28,n191);
nand (n573,n574,n569);
xor (n574,n575,n24);
or (n575,n576,n577);
and (n576,n56,n17);
and (n577,n63,n22);
nand (n578,n565,n574);
xor (n579,n580,n589);
xor (n580,n581,n585);
xor (n581,n582,n24);
or (n582,n583,n584);
and (n583,n52,n17);
and (n584,n56,n22);
xor (n585,n586,n35);
or (n586,n587,n588);
and (n587,n63,n29);
and (n588,n67,n33);
xor (n589,n590,n59);
or (n590,n591,n592);
and (n591,n225,n53);
and (n592,n297,n57);
nand (n593,n594,n579);
nand (n594,n595,n604,n609);
nand (n595,n596,n600);
xor (n596,n597,n189);
or (n597,n598,n599);
and (n598,n16,n326);
and (n599,n21,n330);
xor (n600,n601,n35);
or (n601,n602,n603);
and (n602,n67,n29);
and (n603,n92,n33);
nand (n604,n605,n600);
xor (n605,n606,n46);
or (n606,n607,n608);
and (n607,n179,n40);
and (n608,n225,n44);
nand (n609,n596,n605);
nand (n610,n563,n594);
xor (n611,n612,n617);
xor (n612,n613,n615);
xor (n613,n614,n336);
xor (n614,n322,n332);
xor (n615,n616,n358);
xor (n616,n349,n353);
nand (n617,n618,n619,n620);
nand (n618,n581,n585);
nand (n619,n589,n585);
nand (n620,n581,n589);
xor (n621,n622,n697);
xor (n622,n623,n677);
nand (n623,n624,n650,n676);
nand (n624,n625,n640);
nand (n625,n626,n638,n639);
nand (n626,n627,n632);
xor (n627,n628,n59);
or (n628,n629,n630);
and (n629,n297,n53);
and (n630,n631,n57);
xor (n632,n633,n70);
or (n633,n634,n636);
and (n634,n635,n64);
and (n636,n637,n68);
nand (n638,n70,n632);
nand (n639,n627,n70);
xor (n640,n641,n646);
xor (n641,n642,n322);
xor (n642,n643,n70);
or (n643,n644,n645);
and (n644,n631,n64);
and (n645,n635,n68);
xor (n646,n647,n46);
or (n647,n648,n649);
and (n648,n92,n40);
and (n649,n179,n44);
nand (n650,n651,n640);
xor (n651,n652,n674);
xor (n652,n70,n653);
nand (n653,n654,n668,n673);
nand (n654,n655,n658);
xor (n655,n656,n189);
or (n656,n325,n657);
and (n657,n16,n330);
not (n658,n659);
xor (n659,n660,n328);
or (n660,n661,n665);
and (n661,n75,n662);
xor (n662,n663,n664);
and (n665,n75,n666);
nor (n666,n662,n667);
xnor (n667,n328,n663);
nand (n668,n669,n658);
xor (n669,n670,n78);
or (n670,n671,n672);
and (n671,n32,n105);
and (n672,n39,n109);
nand (n673,n655,n669);
xor (n674,n675,n556);
xor (n675,n547,n551);
nand (n676,n625,n651);
xor (n677,n678,n693);
xor (n678,n679,n683);
nand (n679,n680,n681,n682);
nand (n680,n642,n322);
nand (n681,n646,n322);
nand (n682,n642,n646);
xor (n683,n684,n323);
xor (n684,n685,n689);
xor (n685,n686,n59);
or (n686,n687,n688);
and (n687,n179,n53);
and (n688,n225,n57);
xor (n689,n690,n70);
or (n690,n691,n692);
and (n691,n297,n64);
and (n692,n631,n68);
nand (n693,n694,n695,n696);
nand (n694,n70,n653);
nand (n695,n674,n653);
nand (n696,n70,n674);
nand (n697,n698,n754,n757);
nand (n698,n699,n719);
nand (n699,n700,n715,n718);
nand (n700,n701,n713);
nand (n701,n702,n707,n712);
nand (n702,n659,n703);
xor (n703,n704,n78);
or (n704,n705,n706);
and (n705,n39,n105);
and (n706,n43,n109);
nand (n707,n708,n703);
xor (n708,n709,n19);
or (n709,n710,n711);
and (n710,n52,n76);
and (n711,n56,n80);
nand (n712,n659,n708);
xor (n713,n714,n574);
xor (n714,n565,n569);
nand (n715,n716,n713);
xor (n716,n717,n669);
xor (n717,n655,n658);
nand (n718,n701,n716);
nand (n719,n720,n750,n753);
nand (n720,n721,n734);
nand (n721,n722,n728,n733);
nand (n722,n723,n727);
xor (n723,n724,n107);
or (n724,n725,n726);
and (n725,n28,n187);
and (n726,n32,n191);
not (n727,n596);
nand (n728,n729,n727);
xor (n729,n730,n24);
or (n730,n731,n732);
and (n731,n63,n17);
and (n732,n67,n22);
nand (n733,n723,n729);
nand (n734,n735,n744,n749);
nand (n735,n736,n740);
xor (n736,n737,n35);
or (n737,n738,n739);
and (n738,n92,n29);
and (n739,n179,n33);
xor (n740,n741,n46);
or (n741,n742,n743);
and (n742,n225,n40);
and (n743,n297,n44);
nand (n744,n745,n740);
xor (n745,n746,n59);
or (n746,n747,n748);
and (n747,n631,n53);
and (n748,n635,n57);
nand (n749,n736,n745);
nand (n750,n751,n734);
xor (n751,n752,n605);
xor (n752,n596,n600);
nand (n753,n721,n751);
nand (n754,n755,n719);
xor (n755,n756,n594);
xor (n756,n563,n579);
nand (n757,n699,n755);
nand (n758,n759,n621);
nand (n759,n760,n837,n840);
nand (n760,n761,n763);
xor (n761,n762,n651);
xor (n762,n625,n640);
nand (n763,n764,n797,n836);
nand (n764,n765,n795);
nand (n765,n766,n772,n794);
nand (n766,n767,n70);
xor (n767,n768,n70);
or (n768,n769,n770);
and (n769,n637,n64);
and (n770,n771,n68);
nand (n772,n773,n70);
nand (n773,n774,n782,n793);
nand (n774,n775,n778);
xor (n775,n776,n328);
or (n776,n661,n777);
and (n777,n16,n666);
xor (n778,n779,n189);
or (n779,n780,n781);
and (n780,n21,n326);
and (n781,n28,n330);
nand (n782,n783,n778);
not (n783,n784);
xor (n784,n785,n664);
or (n785,n786,n790);
and (n786,n75,n787);
xor (n787,n788,n789);
and (n790,n75,n791);
nor (n791,n787,n792);
xnor (n792,n664,n788);
nand (n793,n775,n783);
nand (n794,n767,n773);
xor (n795,n796,n70);
xor (n796,n627,n632);
nand (n797,n798,n795);
nand (n798,n799,n818,n835);
nand (n799,n800,n816);
nand (n800,n801,n810,n815);
nand (n801,n802,n806);
xor (n802,n803,n107);
or (n803,n804,n805);
and (n804,n32,n187);
and (n805,n39,n191);
xor (n806,n807,n78);
or (n807,n808,n809);
and (n808,n43,n105);
and (n809,n52,n109);
nand (n810,n811,n806);
xor (n811,n812,n19);
or (n812,n813,n814);
and (n813,n56,n76);
and (n814,n63,n80);
nand (n815,n802,n811);
xor (n816,n817,n708);
xor (n817,n659,n703);
nand (n818,n819,n816);
nand (n819,n820,n829,n834);
nand (n820,n821,n825);
xor (n821,n822,n35);
or (n822,n823,n824);
and (n823,n179,n29);
and (n824,n225,n33);
xor (n825,n826,n328);
or (n826,n827,n828);
and (n827,n16,n662);
and (n828,n21,n666);
nand (n829,n830,n825);
xor (n830,n831,n24);
or (n831,n832,n833);
and (n832,n67,n17);
and (n833,n92,n22);
nand (n834,n821,n830);
nand (n835,n800,n819);
nand (n836,n765,n798);
nand (n837,n838,n763);
xor (n838,n839,n755);
xor (n839,n699,n719);
nand (n840,n761,n838);
nand (n841,n537,n759);
xor (n842,n843,n876);
xor (n843,n844,n848);
nand (n844,n845,n846,n847);
nand (n845,n539,n561);
nand (n846,n611,n561);
nand (n847,n539,n611);
xor (n848,n849,n864);
xor (n849,n850,n854);
nand (n850,n851,n852,n853);
nand (n851,n679,n683);
nand (n852,n693,n683);
nand (n853,n679,n693);
xor (n854,n855,n862);
xor (n855,n856,n860);
nand (n856,n857,n858,n859);
nand (n857,n685,n689);
nand (n858,n323,n689);
nand (n859,n685,n323);
xor (n860,n861,n320);
xor (n861,n311,n315);
xor (n862,n863,n183);
xor (n863,n289,n293);
xor (n864,n865,n872);
xor (n865,n866,n870);
nand (n866,n867,n868,n869);
nand (n867,n541,n70);
nand (n868,n545,n70);
nand (n869,n541,n545);
xor (n870,n871,n347);
xor (n871,n70,n344);
nand (n872,n873,n874,n875);
nand (n873,n613,n615);
nand (n874,n617,n615);
nand (n875,n613,n617);
nand (n876,n877,n878,n879);
nand (n877,n623,n677);
nand (n878,n697,n677);
nand (n879,n623,n697);
nor (n880,n881,n885);
nand (n881,n882,n883,n884);
nand (n882,n844,n848);
nand (n883,n876,n848);
nand (n884,n844,n876);
xor (n885,n886,n901);
xor (n886,n887,n889);
xor (n887,n888,n365);
xor (n888,n309,n342);
xor (n889,n890,n897);
xor (n890,n891,n893);
xor (n891,n892,n303);
xor (n892,n287,n300);
nand (n893,n894,n895,n896);
nand (n894,n856,n860);
nand (n895,n862,n860);
nand (n896,n856,n862);
nand (n897,n898,n899,n900);
nand (n898,n866,n870);
nand (n899,n872,n870);
nand (n900,n866,n872);
nand (n901,n902,n903,n904);
nand (n902,n850,n854);
nand (n903,n864,n854);
nand (n904,n850,n864);
not (n905,n906);
nand (n906,n881,n885);
not (n907,n908);
nor (n908,n909,n924);
nor (n909,n910,n914);
nand (n910,n911,n912,n913);
nand (n911,n887,n889);
nand (n912,n901,n889);
nand (n913,n887,n901);
xor (n914,n915,n920);
xor (n915,n916,n918);
xor (n916,n917,n255);
xor (n917,n251,n253);
xor (n918,n919,n307);
xor (n919,n283,n285);
nand (n920,n921,n922,n923);
nand (n921,n891,n893);
nand (n922,n897,n893);
nand (n923,n891,n897);
nor (n924,n925,n929);
nand (n925,n926,n927,n928);
nand (n926,n916,n918);
nand (n927,n920,n918);
nand (n928,n916,n920);
xor (n929,n930,n281);
xor (n930,n249,n278);
not (n931,n932);
nor (n932,n933,n935);
nor (n933,n934,n924);
nand (n934,n910,n914);
not (n935,n936);
nand (n936,n925,n929);
not (n937,n938);
nor (n938,n939,n946);
nor (n939,n940,n945);
nor (n940,n941,n943);
nor (n941,n942,n370);
nand (n942,n7,n247);
not (n943,n944);
nand (n944,n371,n375);
not (n945,n425);
not (n946,n947);
nor (n947,n948,n950);
nor (n948,n949,n482);
nand (n949,n427,n431);
not (n950,n951);
nand (n951,n483,n487);
nand (n952,n953,n957);
nor (n953,n954,n4);
nand (n954,n955,n908);
nor (n955,n956,n880);
nor (n956,n535,n842);
nand (n957,n958,n2488);
nor (n958,n959,n2456);
nor (n959,n960,n1929);
nor (n960,n961,n1914);
nor (n961,n962,n1635);
nand (n962,n963,n1418);
nor (n963,n964,n1317);
nor (n964,n965,n1227);
nand (n965,n966,n1142,n1226);
nand (n966,n967,n1044);
xor (n967,n968,n1020);
xor (n968,n969,n994);
xor (n969,n970,n982);
xor (n970,n971,n976);
xor (n971,n972,n24);
or (n972,n973,n974);
and (n973,n771,n17);
and (n974,n975,n22);
xor (n976,n977,n35);
or (n977,n978,n980);
and (n978,n979,n29);
and (n980,n981,n33);
xor (n982,n983,n987);
xor (n983,n984,n664);
or (n984,n985,n986);
and (n985,n43,n787);
and (n986,n52,n791);
xnor (n987,n988,n789);
nor (n988,n989,n993);
and (n989,n39,n990);
and (n990,n991,n789);
not (n991,n992);
and (n993,n32,n992);
nand (n994,n995,n1005,n1019);
nand (n995,n996,n1000);
xor (n996,n997,n24);
or (n997,n998,n999);
and (n998,n975,n17);
and (n999,n979,n22);
xor (n1000,n1001,n35);
or (n1001,n1002,n1003);
and (n1002,n981,n29);
and (n1003,n1004,n33);
nand (n1005,n1006,n1000);
xor (n1006,n1007,n1016);
xor (n1007,n1008,n1012);
xor (n1008,n1009,n664);
or (n1009,n1010,n1011);
and (n1010,n52,n787);
and (n1011,n56,n791);
xor (n1012,n1013,n189);
or (n1013,n1014,n1015);
and (n1014,n92,n326);
and (n1015,n179,n330);
xnor (n1016,n1017,n46);
nand (n1017,n1018,n40);
nand (n1019,n996,n1006);
xor (n1020,n1021,n1030);
xor (n1021,n1022,n1026);
xor (n1022,n1023,n46);
or (n1023,n1024,n1025);
and (n1024,n1004,n40);
and (n1025,n1018,n44);
nand (n1026,n1027,n1028,n1029);
nand (n1027,n1008,n1012);
nand (n1028,n1016,n1012);
nand (n1029,n1008,n1016);
xor (n1030,n1031,n1040);
xor (n1031,n1032,n1036);
xor (n1032,n1033,n189);
or (n1033,n1034,n1035);
and (n1034,n67,n326);
and (n1035,n92,n330);
xor (n1036,n1037,n328);
or (n1037,n1038,n1039);
and (n1038,n56,n662);
and (n1039,n63,n666);
xor (n1040,n1041,n107);
or (n1041,n1042,n1043);
and (n1042,n179,n187);
and (n1043,n225,n191);
nand (n1044,n1045,n1099,n1141);
nand (n1045,n1046,n1048);
xor (n1046,n1047,n1006);
xor (n1047,n996,n1000);
xor (n1048,n1049,n1088);
xor (n1049,n1050,n1066);
nand (n1050,n1051,n1060,n1065);
nand (n1051,n1052,n1056);
xor (n1052,n1053,n189);
or (n1053,n1054,n1055);
and (n1054,n179,n326);
and (n1055,n225,n330);
xor (n1056,n1057,n328);
or (n1057,n1058,n1059);
and (n1058,n67,n662);
and (n1059,n92,n666);
nand (n1060,n1061,n1056);
xor (n1061,n1062,n107);
or (n1062,n1063,n1064);
and (n1063,n297,n187);
and (n1064,n631,n191);
nand (n1065,n1052,n1061);
nand (n1066,n1067,n1082,n1087);
nand (n1067,n1068,n1077);
xor (n1068,n1069,n1073);
xnor (n1069,n1070,n789);
nor (n1070,n1071,n1072);
and (n1071,n52,n990);
and (n1072,n43,n992);
xor (n1073,n1074,n664);
or (n1074,n1075,n1076);
and (n1075,n56,n787);
and (n1076,n63,n791);
and (n1077,n1078,n35);
xnor (n1078,n1079,n789);
nor (n1079,n1080,n1081);
and (n1080,n56,n990);
and (n1081,n52,n992);
nand (n1082,n1083,n1077);
xor (n1083,n1084,n78);
or (n1084,n1085,n1086);
and (n1085,n635,n105);
and (n1086,n637,n109);
nand (n1087,n1068,n1083);
xor (n1088,n1089,n1095);
xor (n1089,n1090,n1094);
xor (n1090,n1091,n78);
or (n1091,n1092,n1093);
and (n1092,n631,n105);
and (n1093,n635,n109);
and (n1094,n1069,n1073);
xor (n1095,n1096,n19);
or (n1096,n1097,n1098);
and (n1097,n637,n76);
and (n1098,n771,n80);
nand (n1099,n1100,n1048);
nand (n1100,n1101,n1125,n1140);
nand (n1101,n1102,n1123);
nand (n1102,n1103,n1117,n1122);
nand (n1103,n1104,n1113);
and (n1104,n1105,n1109);
xnor (n1105,n1106,n789);
nor (n1106,n1107,n1108);
and (n1107,n63,n990);
and (n1108,n56,n992);
xor (n1109,n1110,n664);
or (n1110,n1111,n1112);
and (n1111,n67,n787);
and (n1112,n92,n791);
xor (n1113,n1114,n78);
or (n1114,n1115,n1116);
and (n1115,n637,n105);
and (n1116,n771,n109);
nand (n1117,n1118,n1113);
xor (n1118,n1119,n19);
or (n1119,n1120,n1121);
and (n1120,n975,n76);
and (n1121,n979,n80);
nand (n1122,n1104,n1118);
xor (n1123,n1124,n1083);
xor (n1124,n1068,n1077);
nand (n1125,n1126,n1123);
xor (n1126,n1127,n1136);
xor (n1127,n1128,n1132);
xor (n1128,n1129,n19);
or (n1129,n1130,n1131);
and (n1130,n771,n76);
and (n1131,n975,n80);
xor (n1132,n1133,n24);
or (n1133,n1134,n1135);
and (n1134,n979,n17);
and (n1135,n981,n22);
xor (n1136,n1137,n35);
or (n1137,n1138,n1139);
and (n1138,n1004,n29);
and (n1139,n1018,n33);
nand (n1140,n1102,n1126);
nand (n1141,n1046,n1100);
nand (n1142,n1143,n1044);
xor (n1143,n1144,n1183);
xor (n1144,n1145,n1149);
nand (n1145,n1146,n1147,n1148);
nand (n1146,n1050,n1066);
nand (n1147,n1088,n1066);
nand (n1148,n1050,n1088);
xor (n1149,n1150,n1172);
xor (n1150,n1151,n1168);
nand (n1151,n1152,n1162,n1167);
nand (n1152,n1153,n1157);
xor (n1153,n1154,n328);
or (n1154,n1155,n1156);
and (n1155,n63,n662);
and (n1156,n67,n666);
xor (n1157,n1158,n46);
xnor (n1158,n1159,n789);
nor (n1159,n1160,n1161);
and (n1160,n43,n990);
and (n1161,n39,n992);
nand (n1162,n1163,n1157);
xor (n1163,n1164,n107);
or (n1164,n1165,n1166);
and (n1165,n225,n187);
and (n1166,n297,n191);
nand (n1167,n1153,n1163);
nand (n1168,n1169,n1170,n1171);
nand (n1169,n1090,n1094);
nand (n1170,n1095,n1094);
nand (n1171,n1090,n1095);
xor (n1172,n1173,n1179);
xor (n1173,n1174,n1175);
and (n1174,n1158,n46);
xor (n1175,n1176,n78);
or (n1176,n1177,n1178);
and (n1177,n297,n105);
and (n1178,n631,n109);
xor (n1179,n1180,n19);
or (n1180,n1181,n1182);
and (n1181,n635,n76);
and (n1182,n637,n80);
nand (n1183,n1184,n1191,n1225);
nand (n1184,n1185,n1189);
nand (n1185,n1186,n1187,n1188);
nand (n1186,n1128,n1132);
nand (n1187,n1136,n1132);
nand (n1188,n1128,n1136);
xor (n1189,n1190,n1163);
xor (n1190,n1153,n1157);
nand (n1191,n1192,n1189);
nand (n1192,n1193,n1210,n1224);
nand (n1193,n1194,n1208);
nand (n1194,n1195,n1204,n1207);
nand (n1195,n1196,n1200);
xor (n1196,n1197,n664);
or (n1197,n1198,n1199);
and (n1198,n63,n787);
and (n1199,n67,n791);
xor (n1200,n1201,n189);
or (n1201,n1202,n1203);
and (n1202,n225,n326);
and (n1203,n297,n330);
nand (n1204,n1205,n1200);
xnor (n1205,n1206,n35);
nand (n1206,n1018,n29);
nand (n1207,n1196,n1205);
xor (n1208,n1209,n1061);
xor (n1209,n1052,n1056);
nand (n1210,n1211,n1208);
nand (n1211,n1212,n1218,n1223);
nand (n1212,n1213,n1217);
xor (n1213,n1214,n328);
or (n1214,n1215,n1216);
and (n1215,n92,n662);
and (n1216,n179,n666);
xor (n1217,n1078,n35);
nand (n1218,n1219,n1217);
xor (n1219,n1220,n107);
or (n1220,n1221,n1222);
and (n1221,n631,n187);
and (n1222,n635,n191);
nand (n1223,n1213,n1219);
nand (n1224,n1194,n1211);
nand (n1225,n1185,n1192);
nand (n1226,n967,n1143);
xor (n1227,n1228,n1313);
xor (n1228,n1229,n1250);
xor (n1229,n1230,n1246);
xor (n1230,n1231,n1242);
xor (n1231,n1232,n1238);
xor (n1232,n1233,n1237);
xor (n1233,n1234,n35);
or (n1234,n1235,n1236);
and (n1235,n975,n29);
and (n1236,n979,n33);
and (n1237,n983,n987);
xor (n1238,n1239,n46);
or (n1239,n1240,n1241);
and (n1240,n981,n40);
and (n1241,n1004,n44);
nand (n1242,n1243,n1244,n1245);
nand (n1243,n1022,n1026);
nand (n1244,n1030,n1026);
nand (n1245,n1022,n1030);
nand (n1246,n1247,n1248,n1249);
nand (n1247,n1151,n1168);
nand (n1248,n1172,n1168);
nand (n1249,n1151,n1172);
xor (n1250,n1251,n1309);
xor (n1251,n1252,n1276);
xor (n1252,n1253,n1272);
xor (n1253,n1254,n1258);
nand (n1254,n1255,n1256,n1257);
nand (n1255,n1174,n1175);
nand (n1256,n1179,n1175);
nand (n1257,n1174,n1179);
xor (n1258,n1259,n1268);
xor (n1259,n1260,n1264);
xnor (n1260,n1261,n789);
nor (n1261,n1262,n1263);
and (n1262,n32,n990);
and (n1263,n28,n992);
xor (n1264,n1265,n189);
or (n1265,n1266,n1267);
and (n1266,n63,n326);
and (n1267,n67,n330);
xor (n1268,n1269,n328);
or (n1269,n1270,n1271);
and (n1270,n52,n662);
and (n1271,n56,n666);
nand (n1272,n1273,n1274,n1275);
nand (n1273,n1032,n1036);
nand (n1274,n1040,n1036);
nand (n1275,n1032,n1040);
xor (n1276,n1277,n1295);
xor (n1277,n1278,n1282);
nand (n1278,n1279,n1280,n1281);
nand (n1279,n971,n976);
nand (n1280,n982,n976);
nand (n1281,n971,n982);
xor (n1282,n1283,n1293);
xor (n1283,n1284,n1288);
xor (n1284,n1285,n107);
or (n1285,n1286,n1287);
and (n1286,n92,n187);
and (n1287,n179,n191);
xor (n1288,n59,n1289);
xor (n1289,n1290,n664);
or (n1290,n1291,n1292);
and (n1291,n39,n787);
and (n1292,n43,n791);
xnor (n1293,n1294,n59);
nand (n1294,n1018,n53);
xor (n1295,n1296,n1305);
xor (n1296,n1297,n1301);
xor (n1297,n1298,n78);
or (n1298,n1299,n1300);
and (n1299,n225,n105);
and (n1300,n297,n109);
xor (n1301,n1302,n19);
or (n1302,n1303,n1304);
and (n1303,n631,n76);
and (n1304,n635,n80);
xor (n1305,n1306,n24);
or (n1306,n1307,n1308);
and (n1307,n637,n17);
and (n1308,n771,n22);
nand (n1309,n1310,n1311,n1312);
nand (n1310,n969,n994);
nand (n1311,n1020,n994);
nand (n1312,n969,n1020);
nand (n1313,n1314,n1315,n1316);
nand (n1314,n1145,n1149);
nand (n1315,n1183,n1149);
nand (n1316,n1145,n1183);
nor (n1317,n1318,n1322);
nand (n1318,n1319,n1320,n1321);
nand (n1319,n1229,n1250);
nand (n1320,n1313,n1250);
nand (n1321,n1229,n1313);
xor (n1322,n1323,n1332);
xor (n1323,n1324,n1328);
nand (n1324,n1325,n1326,n1327);
nand (n1325,n1231,n1242);
nand (n1326,n1246,n1242);
nand (n1327,n1231,n1246);
nand (n1328,n1329,n1330,n1331);
nand (n1329,n1252,n1276);
nand (n1330,n1309,n1276);
nand (n1331,n1252,n1309);
xor (n1332,n1333,n1394);
xor (n1333,n1334,n1365);
xor (n1334,n1335,n1354);
xor (n1335,n1336,n1350);
xor (n1336,n1337,n1346);
xor (n1337,n1338,n1342);
xor (n1338,n1339,n189);
or (n1339,n1340,n1341);
and (n1340,n56,n326);
and (n1341,n63,n330);
xor (n1342,n1343,n328);
or (n1343,n1344,n1345);
and (n1344,n43,n662);
and (n1345,n52,n666);
xor (n1346,n1347,n107);
or (n1347,n1348,n1349);
and (n1348,n67,n187);
and (n1349,n92,n191);
nand (n1350,n1351,n1352,n1353);
nand (n1351,n1284,n1288);
nand (n1352,n1293,n1288);
nand (n1353,n1284,n1293);
xor (n1354,n1355,n1361);
xor (n1355,n1356,n1360);
xor (n1356,n1357,n78);
or (n1357,n1358,n1359);
and (n1358,n179,n105);
and (n1359,n225,n109);
and (n1360,n59,n1289);
xor (n1361,n1362,n19);
or (n1362,n1363,n1364);
and (n1363,n297,n76);
and (n1364,n631,n80);
xor (n1365,n1366,n1390);
xor (n1366,n1367,n1371);
nand (n1367,n1368,n1369,n1370);
nand (n1368,n1297,n1301);
nand (n1369,n1305,n1301);
nand (n1370,n1297,n1305);
xor (n1371,n1372,n1381);
xor (n1372,n1373,n1377);
xor (n1373,n1374,n24);
or (n1374,n1375,n1376);
and (n1375,n635,n17);
and (n1376,n637,n22);
xor (n1377,n1378,n35);
or (n1378,n1379,n1380);
and (n1379,n771,n29);
and (n1380,n975,n33);
xor (n1381,n1382,n1386);
xnor (n1382,n1383,n789);
nor (n1383,n1384,n1385);
and (n1384,n28,n990);
and (n1385,n21,n992);
xor (n1386,n1387,n664);
or (n1387,n1388,n1389);
and (n1388,n32,n787);
and (n1389,n39,n791);
nand (n1390,n1391,n1392,n1393);
nand (n1391,n1233,n1237);
nand (n1392,n1238,n1237);
nand (n1393,n1233,n1238);
xor (n1394,n1395,n1414);
xor (n1395,n1396,n1410);
xor (n1396,n1397,n1406);
xor (n1397,n1398,n1402);
xor (n1398,n1399,n46);
or (n1399,n1400,n1401);
and (n1400,n979,n40);
and (n1401,n981,n44);
xor (n1402,n1403,n59);
or (n1403,n1404,n1405);
and (n1404,n1004,n53);
and (n1405,n1018,n57);
nand (n1406,n1407,n1408,n1409);
nand (n1407,n1260,n1264);
nand (n1408,n1268,n1264);
nand (n1409,n1260,n1268);
nand (n1410,n1411,n1412,n1413);
nand (n1411,n1254,n1258);
nand (n1412,n1272,n1258);
nand (n1413,n1254,n1272);
nand (n1414,n1415,n1416,n1417);
nand (n1415,n1278,n1282);
nand (n1416,n1295,n1282);
nand (n1417,n1278,n1295);
nor (n1418,n1419,n1524);
nor (n1419,n1420,n1424);
nand (n1420,n1421,n1422,n1423);
nand (n1421,n1324,n1328);
nand (n1422,n1332,n1328);
nand (n1423,n1324,n1332);
xor (n1424,n1425,n1520);
xor (n1425,n1426,n1460);
xor (n1426,n1427,n1456);
xor (n1427,n1428,n1432);
nand (n1428,n1429,n1430,n1431);
nand (n1429,n1336,n1350);
nand (n1430,n1354,n1350);
nand (n1431,n1336,n1354);
xor (n1432,n1433,n1442);
xor (n1433,n1434,n1438);
xor (n1434,n1435,n59);
or (n1435,n1436,n1437);
and (n1436,n981,n53);
and (n1437,n1004,n57);
nand (n1438,n1439,n1440,n1441);
nand (n1439,n1356,n1360);
nand (n1440,n1361,n1360);
nand (n1441,n1356,n1361);
xor (n1442,n1443,n1452);
xor (n1443,n1444,n1448);
xor (n1444,n1445,n189);
or (n1445,n1446,n1447);
and (n1446,n52,n326);
and (n1447,n56,n330);
xnor (n1448,n1449,n789);
nor (n1449,n1450,n1451);
and (n1450,n21,n990);
and (n1451,n16,n992);
xor (n1452,n1453,n328);
or (n1453,n1454,n1455);
and (n1454,n39,n662);
and (n1455,n43,n666);
nand (n1456,n1457,n1458,n1459);
nand (n1457,n1367,n1371);
nand (n1458,n1390,n1371);
nand (n1459,n1367,n1390);
xor (n1460,n1461,n1516);
xor (n1461,n1462,n1484);
xor (n1462,n1463,n1472);
xor (n1463,n1464,n1468);
nand (n1464,n1465,n1466,n1467);
nand (n1465,n1338,n1342);
nand (n1466,n1346,n1342);
nand (n1467,n1338,n1346);
nand (n1468,n1469,n1470,n1471);
nand (n1469,n1373,n1377);
nand (n1470,n1381,n1377);
nand (n1471,n1373,n1381);
xor (n1472,n1473,n1480);
xor (n1473,n1474,n1478);
xor (n1474,n1475,n107);
or (n1475,n1476,n1477);
and (n1476,n63,n187);
and (n1477,n67,n191);
xnor (n1478,n1479,n70);
nand (n1479,n1018,n64);
xor (n1480,n1481,n78);
or (n1481,n1482,n1483);
and (n1482,n92,n105);
and (n1483,n179,n109);
xor (n1484,n1485,n1504);
xor (n1485,n1486,n1490);
nand (n1486,n1487,n1488,n1489);
nand (n1487,n1398,n1402);
nand (n1488,n1406,n1402);
nand (n1489,n1398,n1406);
xor (n1490,n1491,n1500);
xor (n1491,n1492,n1496);
xor (n1492,n1493,n19);
or (n1493,n1494,n1495);
and (n1494,n225,n76);
and (n1495,n297,n80);
xor (n1496,n1497,n24);
or (n1497,n1498,n1499);
and (n1498,n631,n17);
and (n1499,n635,n22);
xor (n1500,n1501,n35);
or (n1501,n1502,n1503);
and (n1502,n637,n29);
and (n1503,n771,n33);
xor (n1504,n1505,n1512);
xor (n1505,n1506,n1511);
xor (n1506,n70,n1507);
xor (n1507,n1508,n664);
or (n1508,n1509,n1510);
and (n1509,n28,n787);
and (n1510,n32,n791);
and (n1511,n1382,n1386);
xor (n1512,n1513,n46);
or (n1513,n1514,n1515);
and (n1514,n975,n40);
and (n1515,n979,n44);
nand (n1516,n1517,n1518,n1519);
nand (n1517,n1396,n1410);
nand (n1518,n1414,n1410);
nand (n1519,n1396,n1414);
nand (n1520,n1521,n1522,n1523);
nand (n1521,n1334,n1365);
nand (n1522,n1394,n1365);
nand (n1523,n1334,n1394);
nor (n1524,n1525,n1529);
nand (n1525,n1526,n1527,n1528);
nand (n1526,n1426,n1460);
nand (n1527,n1520,n1460);
nand (n1528,n1426,n1520);
xor (n1529,n1530,n1539);
xor (n1530,n1531,n1535);
nand (n1531,n1532,n1533,n1534);
nand (n1532,n1428,n1432);
nand (n1533,n1456,n1432);
nand (n1534,n1428,n1456);
nand (n1535,n1536,n1537,n1538);
nand (n1536,n1462,n1484);
nand (n1537,n1516,n1484);
nand (n1538,n1462,n1516);
xor (n1539,n1540,n1601);
xor (n1540,n1541,n1565);
xor (n1541,n1542,n1561);
xor (n1542,n1543,n1547);
nand (n1543,n1544,n1545,n1546);
nand (n1544,n1492,n1496);
nand (n1545,n1500,n1496);
nand (n1546,n1492,n1500);
xor (n1547,n1548,n1557);
xor (n1548,n1549,n1553);
xor (n1549,n1550,n78);
or (n1550,n1551,n1552);
and (n1551,n67,n105);
and (n1552,n92,n109);
xor (n1553,n1554,n19);
or (n1554,n1555,n1556);
and (n1555,n179,n76);
and (n1556,n225,n80);
xor (n1557,n1558,n24);
or (n1558,n1559,n1560);
and (n1559,n297,n17);
and (n1560,n631,n22);
nand (n1561,n1562,n1563,n1564);
nand (n1562,n1506,n1511);
nand (n1563,n1512,n1511);
nand (n1564,n1506,n1512);
xor (n1565,n1566,n1587);
xor (n1566,n1567,n1583);
xor (n1567,n1568,n1582);
xor (n1568,n1569,n1573);
xor (n1569,n1570,n35);
or (n1570,n1571,n1572);
and (n1571,n635,n29);
and (n1572,n637,n33);
xor (n1573,n1574,n1578);
xnor (n1574,n1575,n789);
nor (n1575,n1576,n1577);
and (n1576,n16,n990);
and (n1577,n75,n992);
xor (n1578,n1579,n664);
or (n1579,n1580,n1581);
and (n1580,n21,n787);
and (n1581,n28,n791);
and (n1582,n70,n1507);
nand (n1583,n1584,n1585,n1586);
nand (n1584,n1434,n1438);
nand (n1585,n1442,n1438);
nand (n1586,n1434,n1442);
xor (n1587,n1588,n1597);
xor (n1588,n1589,n1593);
xor (n1589,n1590,n46);
or (n1590,n1591,n1592);
and (n1591,n771,n40);
and (n1592,n975,n44);
xor (n1593,n1594,n70);
or (n1594,n1595,n1596);
and (n1595,n1004,n64);
and (n1596,n1018,n68);
xor (n1597,n1598,n59);
or (n1598,n1599,n1600);
and (n1599,n979,n53);
and (n1600,n981,n57);
xor (n1601,n1602,n1631);
xor (n1602,n1603,n1627);
xor (n1603,n1604,n1623);
xor (n1604,n1605,n1609);
nand (n1605,n1606,n1607,n1608);
nand (n1606,n1444,n1448);
nand (n1607,n1452,n1448);
nand (n1608,n1444,n1452);
xor (n1609,n1610,n1619);
xor (n1610,n1611,n1615);
xor (n1611,n1612,n189);
or (n1612,n1613,n1614);
and (n1613,n43,n326);
and (n1614,n52,n330);
xor (n1615,n1616,n328);
or (n1616,n1617,n1618);
and (n1617,n32,n662);
and (n1618,n39,n666);
xor (n1619,n1620,n107);
or (n1620,n1621,n1622);
and (n1621,n56,n187);
and (n1622,n63,n191);
nand (n1623,n1624,n1625,n1626);
nand (n1624,n1474,n1478);
nand (n1625,n1480,n1478);
nand (n1626,n1474,n1480);
nand (n1627,n1628,n1629,n1630);
nand (n1628,n1464,n1468);
nand (n1629,n1472,n1468);
nand (n1630,n1464,n1472);
nand (n1631,n1632,n1633,n1634);
nand (n1632,n1486,n1490);
nand (n1633,n1504,n1490);
nand (n1634,n1486,n1504);
nor (n1635,n1636,n1908);
nor (n1636,n1637,n1884);
nor (n1637,n1638,n1882);
nor (n1638,n1639,n1857);
nand (n1639,n1640,n1819);
nand (n1640,n1641,n1766,n1818);
nand (n1641,n1642,n1693);
xor (n1642,n1643,n1680);
xor (n1643,n1644,n1665);
nand (n1644,n1645,n1659,n1664);
nand (n1645,n1646,n1655);
and (n1646,n1647,n1651);
xnor (n1647,n1648,n789);
nor (n1648,n1649,n1650);
and (n1649,n92,n990);
and (n1650,n67,n992);
xor (n1651,n1652,n664);
or (n1652,n1653,n1654);
and (n1653,n179,n787);
and (n1654,n225,n791);
xor (n1655,n1656,n78);
or (n1656,n1657,n1658);
and (n1657,n975,n105);
and (n1658,n979,n109);
nand (n1659,n1660,n1655);
xor (n1660,n1661,n19);
or (n1661,n1662,n1663);
and (n1662,n981,n76);
and (n1663,n1004,n80);
nand (n1664,n1646,n1660);
xor (n1665,n1666,n1675);
xor (n1666,n1667,n1671);
xor (n1667,n1668,n189);
or (n1668,n1669,n1670);
and (n1669,n297,n326);
and (n1670,n631,n330);
xor (n1671,n1672,n328);
or (n1672,n1673,n1674);
and (n1673,n179,n662);
and (n1674,n225,n666);
and (n1675,n1676,n24);
xnor (n1676,n1677,n789);
nor (n1677,n1678,n1679);
and (n1678,n67,n990);
and (n1679,n63,n992);
nand (n1680,n1681,n1687,n1692);
nand (n1681,n1682,n1686);
xor (n1682,n1683,n328);
or (n1683,n1684,n1685);
and (n1684,n225,n662);
and (n1685,n297,n666);
xor (n1686,n1676,n24);
nand (n1687,n1688,n1686);
xor (n1688,n1689,n107);
or (n1689,n1690,n1691);
and (n1690,n637,n187);
and (n1691,n771,n191);
nand (n1692,n1682,n1688);
xor (n1693,n1694,n1730);
xor (n1694,n1695,n1706);
xor (n1695,n1696,n1702);
xor (n1696,n1697,n1701);
xor (n1697,n1698,n107);
or (n1698,n1699,n1700);
and (n1699,n635,n187);
and (n1700,n637,n191);
xor (n1701,n1105,n1109);
xor (n1702,n1703,n78);
or (n1703,n1704,n1705);
and (n1704,n771,n105);
and (n1705,n975,n109);
xor (n1706,n1707,n1716);
xor (n1707,n1708,n1712);
xor (n1708,n1709,n19);
or (n1709,n1710,n1711);
and (n1710,n979,n76);
and (n1711,n981,n80);
xor (n1712,n1713,n24);
or (n1713,n1714,n1715);
and (n1714,n1004,n17);
and (n1715,n1018,n22);
nand (n1716,n1717,n1724,n1729);
nand (n1717,n1718,n1722);
xor (n1718,n1719,n664);
or (n1719,n1720,n1721);
and (n1720,n92,n787);
and (n1721,n179,n791);
xnor (n1722,n1723,n24);
nand (n1723,n1018,n17);
nand (n1724,n1725,n1722);
xor (n1725,n1726,n189);
or (n1726,n1727,n1728);
and (n1727,n631,n326);
and (n1728,n635,n330);
nand (n1729,n1718,n1725);
nand (n1730,n1731,n1751,n1765);
nand (n1731,n1732,n1734);
xor (n1732,n1733,n1725);
xor (n1733,n1718,n1722);
nand (n1734,n1735,n1744,n1750);
nand (n1735,n1736,n1740);
xor (n1736,n1737,n189);
or (n1737,n1738,n1739);
and (n1738,n635,n326);
and (n1739,n637,n330);
xor (n1740,n1741,n328);
or (n1741,n1742,n1743);
and (n1742,n297,n662);
and (n1743,n631,n666);
nand (n1744,n1745,n1740);
and (n1745,n1746,n19);
xnor (n1746,n1747,n789);
nor (n1747,n1748,n1749);
and (n1748,n179,n990);
and (n1749,n92,n992);
nand (n1750,n1736,n1745);
nand (n1751,n1752,n1734);
nand (n1752,n1753,n1759,n1764);
nand (n1753,n1754,n1758);
xor (n1754,n1755,n107);
or (n1755,n1756,n1757);
and (n1756,n771,n187);
and (n1757,n975,n191);
xor (n1758,n1647,n1651);
nand (n1759,n1760,n1758);
xor (n1760,n1761,n78);
or (n1761,n1762,n1763);
and (n1762,n979,n105);
and (n1763,n981,n109);
nand (n1764,n1754,n1760);
nand (n1765,n1732,n1752);
nand (n1766,n1767,n1693);
nand (n1767,n1768,n1773,n1817);
nand (n1768,n1769,n1771);
xor (n1769,n1770,n1660);
xor (n1770,n1646,n1655);
xor (n1771,n1772,n1688);
xor (n1772,n1682,n1686);
nand (n1773,n1774,n1771);
nand (n1774,n1775,n1794,n1816);
nand (n1775,n1776,n1780);
xor (n1776,n1777,n19);
or (n1777,n1778,n1779);
and (n1778,n1004,n76);
and (n1779,n1018,n80);
nand (n1780,n1781,n1788,n1793);
nand (n1781,n1782,n1786);
xor (n1782,n1783,n664);
or (n1783,n1784,n1785);
and (n1784,n225,n787);
and (n1785,n297,n791);
xnor (n1786,n1787,n19);
nand (n1787,n1018,n76);
nand (n1788,n1789,n1786);
xor (n1789,n1790,n189);
or (n1790,n1791,n1792);
and (n1791,n637,n326);
and (n1792,n771,n330);
nand (n1793,n1782,n1789);
nand (n1794,n1795,n1780);
nand (n1795,n1796,n1810,n1815);
nand (n1796,n1797,n1801);
xor (n1797,n1798,n328);
or (n1798,n1799,n1800);
and (n1799,n631,n662);
and (n1800,n635,n666);
and (n1801,n1802,n1806);
xnor (n1802,n1803,n789);
nor (n1803,n1804,n1805);
and (n1804,n225,n990);
and (n1805,n179,n992);
xor (n1806,n1807,n664);
or (n1807,n1808,n1809);
and (n1808,n297,n787);
and (n1809,n631,n791);
nand (n1810,n1811,n1801);
xor (n1811,n1812,n107);
or (n1812,n1813,n1814);
and (n1813,n975,n187);
and (n1814,n979,n191);
nand (n1815,n1797,n1811);
nand (n1816,n1776,n1795);
nand (n1817,n1769,n1774);
nand (n1818,n1642,n1767);
xor (n1819,n1820,n1835);
xor (n1820,n1821,n1831);
xor (n1821,n1822,n1829);
xor (n1822,n1823,n1827);
nand (n1823,n1824,n1825,n1826);
nand (n1824,n1667,n1671);
nand (n1825,n1675,n1671);
nand (n1826,n1667,n1675);
xor (n1827,n1828,n1118);
xor (n1828,n1104,n1113);
xor (n1829,n1830,n1219);
xor (n1830,n1213,n1217);
nand (n1831,n1832,n1833,n1834);
nand (n1832,n1695,n1706);
nand (n1833,n1730,n1706);
nand (n1834,n1695,n1730);
xor (n1835,n1836,n1845);
xor (n1836,n1837,n1841);
nand (n1837,n1838,n1839,n1840);
nand (n1838,n1708,n1712);
nand (n1839,n1716,n1712);
nand (n1840,n1708,n1716);
nand (n1841,n1842,n1843,n1844);
nand (n1842,n1644,n1665);
nand (n1843,n1680,n1665);
nand (n1844,n1644,n1680);
xor (n1845,n1846,n1855);
xor (n1846,n1847,n1851);
xor (n1847,n1848,n24);
or (n1848,n1849,n1850);
and (n1849,n981,n17);
and (n1850,n1004,n22);
nand (n1851,n1852,n1853,n1854);
nand (n1852,n1697,n1701);
nand (n1853,n1702,n1701);
nand (n1854,n1697,n1702);
xor (n1855,n1856,n1205);
xor (n1856,n1196,n1200);
nor (n1857,n1858,n1862);
nand (n1858,n1859,n1860,n1861);
nand (n1859,n1821,n1831);
nand (n1860,n1835,n1831);
nand (n1861,n1821,n1835);
xor (n1862,n1863,n1870);
xor (n1863,n1864,n1866);
xor (n1864,n1865,n1126);
xor (n1865,n1102,n1123);
nand (n1866,n1867,n1868,n1869);
nand (n1867,n1837,n1841);
nand (n1868,n1845,n1841);
nand (n1869,n1837,n1845);
xor (n1870,n1871,n1880);
xor (n1871,n1872,n1876);
nand (n1872,n1873,n1874,n1875);
nand (n1873,n1847,n1851);
nand (n1874,n1855,n1851);
nand (n1875,n1847,n1855);
nand (n1876,n1877,n1878,n1879);
nand (n1877,n1823,n1827);
nand (n1878,n1829,n1827);
nand (n1879,n1823,n1829);
xor (n1880,n1881,n1211);
xor (n1881,n1194,n1208);
not (n1882,n1883);
nand (n1883,n1858,n1862);
not (n1884,n1885);
nor (n1885,n1886,n1901);
nor (n1886,n1887,n1891);
nand (n1887,n1888,n1889,n1890);
nand (n1888,n1864,n1866);
nand (n1889,n1870,n1866);
nand (n1890,n1864,n1870);
xor (n1891,n1892,n1899);
xor (n1892,n1893,n1895);
xor (n1893,n1894,n1192);
xor (n1894,n1185,n1189);
nand (n1895,n1896,n1897,n1898);
nand (n1896,n1872,n1876);
nand (n1897,n1880,n1876);
nand (n1898,n1872,n1880);
xor (n1899,n1900,n1100);
xor (n1900,n1046,n1048);
nor (n1901,n1902,n1906);
nand (n1902,n1903,n1904,n1905);
nand (n1903,n1893,n1895);
nand (n1904,n1899,n1895);
nand (n1905,n1893,n1899);
xor (n1906,n1907,n1143);
xor (n1907,n967,n1044);
not (n1908,n1909);
nor (n1909,n1910,n1912);
nor (n1910,n1911,n1901);
nand (n1911,n1887,n1891);
not (n1912,n1913);
nand (n1913,n1902,n1906);
not (n1914,n1915);
nor (n1915,n1916,n1923);
nor (n1916,n1917,n1922);
nor (n1917,n1918,n1920);
nor (n1918,n1919,n1317);
nand (n1919,n965,n1227);
not (n1920,n1921);
nand (n1921,n1318,n1322);
not (n1922,n1418);
not (n1923,n1924);
nor (n1924,n1925,n1927);
nor (n1925,n1926,n1524);
nand (n1926,n1420,n1424);
not (n1927,n1928);
nand (n1928,n1525,n1529);
not (n1929,n1930);
nor (n1930,n1931,n2346);
nand (n1931,n1932,n2159);
nor (n1932,n1933,n2045);
nor (n1933,n1934,n1938);
nand (n1934,n1935,n1936,n1937);
nand (n1935,n1531,n1535);
nand (n1936,n1539,n1535);
nand (n1937,n1531,n1539);
xor (n1938,n1939,n2041);
xor (n1939,n1940,n1973);
xor (n1940,n1941,n1969);
xor (n1941,n1942,n1965);
xor (n1942,n1943,n1961);
xor (n1943,n1944,n1957);
xor (n1944,n1945,n1954);
xor (n1945,n1946,n1950);
xor (n1946,n1947,n664);
or (n1947,n1948,n1949);
and (n1948,n16,n787);
and (n1949,n21,n791);
xor (n1950,n1951,n328);
or (n1951,n1952,n1953);
and (n1952,n28,n662);
and (n1953,n32,n666);
xnor (n1954,n1955,n789);
nor (n1955,n1956,n1577);
and (n1956,n75,n990);
nand (n1957,n1958,n1959,n1960);
nand (n1958,n1549,n1553);
nand (n1959,n1557,n1553);
nand (n1960,n1549,n1557);
nand (n1961,n1962,n1963,n1964);
nand (n1962,n1569,n1573);
nand (n1963,n1582,n1573);
nand (n1964,n1569,n1582);
nand (n1965,n1966,n1967,n1968);
nand (n1966,n1543,n1547);
nand (n1967,n1561,n1547);
nand (n1968,n1543,n1561);
nand (n1969,n1970,n1971,n1972);
nand (n1970,n1567,n1583);
nand (n1971,n1587,n1583);
nand (n1972,n1567,n1587);
xor (n1973,n1974,n2037);
xor (n1974,n1975,n2013);
xor (n1975,n1976,n1998);
xor (n1976,n1977,n1991);
xor (n1977,n1978,n1987);
xor (n1978,n1979,n1983);
xor (n1979,n1980,n107);
or (n1980,n1981,n1982);
and (n1981,n52,n187);
and (n1982,n56,n191);
xor (n1983,n1984,n78);
or (n1984,n1985,n1986);
and (n1985,n63,n105);
and (n1986,n67,n109);
xor (n1987,n1988,n19);
or (n1988,n1989,n1990);
and (n1989,n92,n76);
and (n1990,n179,n80);
xor (n1991,n1992,n1994);
xor (n1992,n70,n1993);
and (n1993,n1574,n1578);
xor (n1994,n1995,n46);
or (n1995,n1996,n1997);
and (n1996,n637,n40);
and (n1997,n771,n44);
xor (n1998,n1999,n2008);
xor (n1999,n2000,n2004);
xor (n2000,n2001,n24);
or (n2001,n2002,n2003);
and (n2002,n225,n17);
and (n2003,n297,n22);
xor (n2004,n2005,n35);
or (n2005,n2006,n2007);
and (n2006,n631,n29);
and (n2007,n635,n33);
xor (n2008,n70,n2009);
xor (n2009,n2010,n189);
or (n2010,n2011,n2012);
and (n2011,n39,n326);
and (n2012,n43,n330);
xor (n2013,n2014,n2023);
xor (n2014,n2015,n2019);
nand (n2015,n2016,n2017,n2018);
nand (n2016,n1589,n1593);
nand (n2017,n1597,n1593);
nand (n2018,n1589,n1597);
nand (n2019,n2020,n2021,n2022);
nand (n2020,n1605,n1609);
nand (n2021,n1623,n1609);
nand (n2022,n1605,n1623);
xor (n2023,n2024,n2033);
xor (n2024,n2025,n2029);
xor (n2025,n2026,n59);
or (n2026,n2027,n2028);
and (n2027,n975,n53);
and (n2028,n979,n57);
xor (n2029,n2030,n70);
or (n2030,n2031,n2032);
and (n2031,n981,n64);
and (n2032,n1004,n68);
nand (n2033,n2034,n2035,n2036);
nand (n2034,n1611,n1615);
nand (n2035,n1619,n1615);
nand (n2036,n1611,n1619);
nand (n2037,n2038,n2039,n2040);
nand (n2038,n1603,n1627);
nand (n2039,n1631,n1627);
nand (n2040,n1603,n1631);
nand (n2041,n2042,n2043,n2044);
nand (n2042,n1541,n1565);
nand (n2043,n1601,n1565);
nand (n2044,n1541,n1601);
nor (n2045,n2046,n2050);
nand (n2046,n2047,n2048,n2049);
nand (n2047,n1940,n1973);
nand (n2048,n2041,n1973);
nand (n2049,n1940,n2041);
xor (n2050,n2051,n2060);
xor (n2051,n2052,n2056);
nand (n2052,n2053,n2054,n2055);
nand (n2053,n1942,n1965);
nand (n2054,n1969,n1965);
nand (n2055,n1942,n1969);
nand (n2056,n2057,n2058,n2059);
nand (n2057,n1975,n2013);
nand (n2058,n2037,n2013);
nand (n2059,n1975,n2037);
xor (n2060,n2061,n2118);
xor (n2061,n2062,n2093);
xor (n2062,n2063,n2079);
xor (n2063,n2064,n2068);
nand (n2064,n2065,n2066,n2067);
nand (n2065,n70,n1993);
nand (n2066,n1994,n1993);
nand (n2067,n70,n1994);
xor (n2068,n2069,n2075);
xor (n2069,n2070,n2074);
xor (n2070,n2071,n35);
or (n2071,n2072,n2073);
and (n2072,n297,n29);
and (n2073,n631,n33);
and (n2074,n70,n2009);
xor (n2075,n2076,n46);
or (n2076,n2077,n2078);
and (n2077,n635,n40);
and (n2078,n637,n44);
xor (n2079,n2080,n2089);
xor (n2080,n2081,n2085);
xor (n2081,n2082,n59);
or (n2082,n2083,n2084);
and (n2083,n771,n53);
and (n2084,n975,n57);
xor (n2085,n2086,n70);
or (n2086,n2087,n2088);
and (n2087,n979,n64);
and (n2088,n981,n68);
nand (n2089,n2090,n2091,n2092);
nand (n2090,n1946,n1950);
nand (n2091,n1954,n1950);
nand (n2092,n1946,n1954);
xor (n2093,n2094,n2103);
xor (n2094,n2095,n2099);
nand (n2095,n2096,n2097,n2098);
nand (n2096,n2025,n2029);
nand (n2097,n2033,n2029);
nand (n2098,n2025,n2033);
nand (n2099,n2100,n2101,n2102);
nand (n2100,n1944,n1957);
nand (n2101,n1961,n1957);
nand (n2102,n1944,n1961);
xor (n2103,n2104,n70);
xor (n2104,n2105,n2109);
nand (n2105,n2106,n2107,n2108);
nand (n2106,n1979,n1983);
nand (n2107,n1987,n1983);
nand (n2108,n1979,n1987);
xor (n2109,n2110,n2115);
not (n2110,n2111);
xor (n2111,n2112,n189);
or (n2112,n2113,n2114);
and (n2113,n32,n326);
and (n2114,n39,n330);
xor (n2115,n2116,n664);
or (n2116,n786,n2117);
and (n2117,n16,n791);
xor (n2118,n2119,n2155);
xor (n2119,n2120,n2124);
nand (n2120,n2121,n2122,n2123);
nand (n2121,n1977,n1991);
nand (n2122,n1998,n1991);
nand (n2123,n1977,n1998);
xor (n2124,n2125,n2144);
xor (n2125,n2126,n2130);
nand (n2126,n2127,n2128,n2129);
nand (n2127,n2000,n2004);
nand (n2128,n2008,n2004);
nand (n2129,n2000,n2008);
xor (n2130,n2131,n2140);
xor (n2131,n2132,n2136);
xor (n2132,n2133,n78);
or (n2133,n2134,n2135);
and (n2134,n56,n105);
and (n2135,n63,n109);
xor (n2136,n2137,n19);
or (n2137,n2138,n2139);
and (n2138,n67,n76);
and (n2139,n92,n80);
xor (n2140,n2141,n24);
or (n2141,n2142,n2143);
and (n2142,n179,n17);
and (n2143,n225,n22);
xor (n2144,n2145,n2151);
xor (n2145,n2146,n2150);
xor (n2146,n2147,n328);
or (n2147,n2148,n2149);
and (n2148,n21,n662);
and (n2149,n28,n666);
not (n2150,n1954);
xor (n2151,n2152,n107);
or (n2152,n2153,n2154);
and (n2153,n43,n187);
and (n2154,n52,n191);
nand (n2155,n2156,n2157,n2158);
nand (n2156,n2015,n2019);
nand (n2157,n2023,n2019);
nand (n2158,n2015,n2023);
nor (n2159,n2160,n2267);
nor (n2160,n2161,n2165);
nand (n2161,n2162,n2163,n2164);
nand (n2162,n2052,n2056);
nand (n2163,n2060,n2056);
nand (n2164,n2052,n2060);
xor (n2165,n2166,n2263);
xor (n2166,n2167,n2207);
xor (n2167,n2168,n2203);
xor (n2168,n2169,n2199);
xor (n2169,n2170,n2195);
xor (n2170,n2171,n2185);
xor (n2171,n2172,n2181);
xor (n2172,n2173,n2177);
xor (n2173,n2174,n78);
or (n2174,n2175,n2176);
and (n2175,n52,n105);
and (n2176,n56,n109);
xor (n2177,n2178,n19);
or (n2178,n2179,n2180);
and (n2179,n63,n76);
and (n2180,n67,n80);
xor (n2181,n2182,n35);
or (n2182,n2183,n2184);
and (n2183,n225,n29);
and (n2184,n297,n33);
xor (n2185,n2186,n2191);
xor (n2186,n2187,n784);
xor (n2187,n2188,n189);
or (n2188,n2189,n2190);
and (n2189,n28,n326);
and (n2190,n32,n330);
xor (n2191,n2192,n107);
or (n2192,n2193,n2194);
and (n2193,n39,n187);
and (n2194,n43,n191);
nand (n2195,n2196,n2197,n2198);
nand (n2196,n2070,n2074);
nand (n2197,n2075,n2074);
nand (n2198,n2070,n2075);
nand (n2199,n2200,n2201,n2202);
nand (n2200,n2064,n2068);
nand (n2201,n2079,n2068);
nand (n2202,n2064,n2079);
nand (n2203,n2204,n2205,n2206);
nand (n2204,n2095,n2099);
nand (n2205,n2103,n2099);
nand (n2206,n2095,n2103);
xor (n2207,n2208,n2259);
xor (n2208,n2209,n2230);
xor (n2209,n2210,n2226);
xor (n2210,n2211,n2222);
xor (n2211,n2212,n2218);
xor (n2212,n2213,n2214);
not (n2213,n825);
xor (n2214,n2215,n24);
or (n2215,n2216,n2217);
and (n2216,n92,n17);
and (n2217,n179,n22);
xor (n2218,n2219,n46);
or (n2219,n2220,n2221);
and (n2220,n631,n40);
and (n2221,n635,n44);
nand (n2222,n2223,n2224,n2225);
nand (n2223,n2081,n2085);
nand (n2224,n2089,n2085);
nand (n2225,n2081,n2089);
nand (n2226,n2227,n2228,n2229);
nand (n2227,n2105,n2109);
nand (n2228,n70,n2109);
nand (n2229,n2105,n70);
xor (n2230,n2231,n2255);
xor (n2231,n2232,n2245);
xor (n2232,n2233,n2242);
xor (n2233,n2234,n2238);
xor (n2234,n2235,n59);
or (n2235,n2236,n2237);
and (n2236,n637,n53);
and (n2237,n771,n57);
xor (n2238,n2239,n70);
or (n2239,n2240,n2241);
and (n2240,n975,n64);
and (n2241,n979,n68);
nand (n2242,n2110,n2243,n2244);
nand (n2243,n2115,n2111);
not (n2244,n2115);
xor (n2245,n2246,n2251);
xor (n2246,n70,n2247);
nand (n2247,n2248,n2249,n2250);
nand (n2248,n2146,n2150);
nand (n2249,n2151,n2150);
nand (n2250,n2146,n2151);
nand (n2251,n2252,n2253,n2254);
nand (n2252,n2132,n2136);
nand (n2253,n2140,n2136);
nand (n2254,n2132,n2140);
nand (n2255,n2256,n2257,n2258);
nand (n2256,n2126,n2130);
nand (n2257,n2144,n2130);
nand (n2258,n2126,n2144);
nand (n2259,n2260,n2261,n2262);
nand (n2260,n2120,n2124);
nand (n2261,n2155,n2124);
nand (n2262,n2120,n2155);
nand (n2263,n2264,n2265,n2266);
nand (n2264,n2062,n2093);
nand (n2265,n2118,n2093);
nand (n2266,n2062,n2118);
nor (n2267,n2268,n2272);
nand (n2268,n2269,n2270,n2271);
nand (n2269,n2167,n2207);
nand (n2270,n2263,n2207);
nand (n2271,n2167,n2263);
xor (n2272,n2273,n2282);
xor (n2273,n2274,n2278);
nand (n2274,n2275,n2276,n2277);
nand (n2275,n2169,n2199);
nand (n2276,n2203,n2199);
nand (n2277,n2169,n2203);
nand (n2278,n2279,n2280,n2281);
nand (n2279,n2209,n2230);
nand (n2280,n2259,n2230);
nand (n2281,n2209,n2259);
xor (n2282,n2283,n2314);
xor (n2283,n2284,n2288);
nand (n2284,n2285,n2286,n2287);
nand (n2285,n2232,n2245);
nand (n2286,n2255,n2245);
nand (n2287,n2232,n2255);
xor (n2288,n2289,n2302);
xor (n2289,n2290,n2294);
nand (n2290,n2291,n2292,n2293);
nand (n2291,n70,n2247);
nand (n2292,n2251,n2247);
nand (n2293,n70,n2251);
xor (n2294,n2295,n2298);
xor (n2295,n2296,n70);
xor (n2296,n2297,n783);
xor (n2297,n775,n778);
nand (n2298,n2299,n2300,n2301);
nand (n2299,n2187,n784);
nand (n2300,n2191,n784);
nand (n2301,n2187,n2191);
xor (n2302,n2303,n2310);
xor (n2303,n2304,n2306);
xor (n2304,n2305,n811);
xor (n2305,n802,n806);
nand (n2306,n2307,n2308,n2309);
nand (n2307,n2173,n2177);
nand (n2308,n2181,n2177);
nand (n2309,n2173,n2181);
nand (n2310,n2311,n2312,n2313);
nand (n2311,n2234,n2238);
nand (n2312,n2242,n2238);
nand (n2313,n2234,n2242);
xor (n2314,n2315,n2324);
xor (n2315,n2316,n2320);
nand (n2316,n2317,n2318,n2319);
nand (n2317,n2171,n2185);
nand (n2318,n2195,n2185);
nand (n2319,n2171,n2195);
nand (n2320,n2321,n2322,n2323);
nand (n2321,n2211,n2222);
nand (n2322,n2226,n2222);
nand (n2323,n2211,n2226);
xor (n2324,n2325,n2332);
xor (n2325,n2326,n2330);
nand (n2326,n2327,n2328,n2329);
nand (n2327,n2213,n2214);
nand (n2328,n2218,n2214);
nand (n2329,n2213,n2218);
xor (n2330,n2331,n830);
xor (n2331,n821,n825);
xor (n2332,n2333,n2342);
xor (n2333,n2334,n2338);
xor (n2334,n2335,n46);
or (n2335,n2336,n2337);
and (n2336,n297,n40);
and (n2337,n631,n44);
xor (n2338,n2339,n59);
or (n2339,n2340,n2341);
and (n2340,n635,n53);
and (n2341,n637,n57);
xor (n2342,n2343,n70);
or (n2343,n2344,n2345);
and (n2344,n771,n64);
and (n2345,n975,n68);
nand (n2346,n2347,n2431);
nor (n2347,n2348,n2398);
nor (n2348,n2349,n2353);
nand (n2349,n2350,n2351,n2352);
nand (n2350,n2274,n2278);
nand (n2351,n2282,n2278);
nand (n2352,n2274,n2282);
xor (n2353,n2354,n2394);
xor (n2354,n2355,n2375);
xor (n2355,n2356,n2363);
xor (n2356,n2357,n2359);
xor (n2357,n2358,n819);
xor (n2358,n800,n816);
nand (n2359,n2360,n2361,n2362);
nand (n2360,n2326,n2330);
nand (n2361,n2332,n2330);
nand (n2362,n2326,n2332);
xor (n2363,n2364,n2371);
xor (n2364,n2365,n2369);
nand (n2365,n2366,n2367,n2368);
nand (n2366,n2334,n2338);
nand (n2367,n2342,n2338);
nand (n2368,n2334,n2342);
xor (n2369,n2370,n729);
xor (n2370,n723,n727);
nand (n2371,n2372,n2373,n2374);
nand (n2372,n2296,n70);
nand (n2373,n2298,n70);
nand (n2374,n2296,n2298);
xor (n2375,n2376,n2390);
xor (n2376,n2377,n2381);
nand (n2377,n2378,n2379,n2380);
nand (n2378,n2290,n2294);
nand (n2379,n2302,n2294);
nand (n2380,n2290,n2302);
xor (n2381,n2382,n2386);
xor (n2382,n2383,n2385);
xor (n2383,n2384,n745);
xor (n2384,n736,n740);
xor (n2385,n768,n773);
nand (n2386,n2387,n2388,n2389);
nand (n2387,n2304,n2306);
nand (n2388,n2310,n2306);
nand (n2389,n2304,n2310);
nand (n2390,n2391,n2392,n2393);
nand (n2391,n2316,n2320);
nand (n2392,n2324,n2320);
nand (n2393,n2316,n2324);
nand (n2394,n2395,n2396,n2397);
nand (n2395,n2284,n2288);
nand (n2396,n2314,n2288);
nand (n2397,n2284,n2314);
nor (n2398,n2399,n2403);
nand (n2399,n2400,n2401,n2402);
nand (n2400,n2355,n2375);
nand (n2401,n2394,n2375);
nand (n2402,n2355,n2394);
xor (n2403,n2404,n2427);
xor (n2404,n2405,n2415);
xor (n2405,n2406,n2413);
xor (n2406,n2407,n2409);
xor (n2407,n2408,n716);
xor (n2408,n701,n713);
nand (n2409,n2410,n2411,n2412);
nand (n2410,n2365,n2369);
nand (n2411,n2371,n2369);
nand (n2412,n2365,n2371);
xor (n2413,n2414,n751);
xor (n2414,n721,n734);
xor (n2415,n2416,n2423);
xor (n2416,n2417,n2419);
xor (n2417,n2418,n798);
xor (n2418,n765,n795);
nand (n2419,n2420,n2421,n2422);
nand (n2420,n2383,n2385);
nand (n2421,n2386,n2385);
nand (n2422,n2383,n2386);
nand (n2423,n2424,n2425,n2426);
nand (n2424,n2357,n2359);
nand (n2425,n2363,n2359);
nand (n2426,n2357,n2363);
nand (n2427,n2428,n2429,n2430);
nand (n2428,n2377,n2381);
nand (n2429,n2390,n2381);
nand (n2430,n2377,n2390);
nor (n2431,n2432,n2449);
nor (n2432,n2433,n2437);
nand (n2433,n2434,n2435,n2436);
nand (n2434,n2405,n2415);
nand (n2435,n2427,n2415);
nand (n2436,n2405,n2427);
xor (n2437,n2438,n2445);
xor (n2438,n2439,n2443);
nand (n2439,n2440,n2441,n2442);
nand (n2440,n2407,n2409);
nand (n2441,n2413,n2409);
nand (n2442,n2407,n2413);
xor (n2443,n2444,n838);
xor (n2444,n761,n763);
nand (n2445,n2446,n2447,n2448);
nand (n2446,n2417,n2419);
nand (n2447,n2423,n2419);
nand (n2448,n2417,n2423);
nor (n2449,n2450,n2454);
nand (n2450,n2451,n2452,n2453);
nand (n2451,n2439,n2443);
nand (n2452,n2445,n2443);
nand (n2453,n2439,n2445);
xor (n2454,n2455,n759);
xor (n2455,n537,n621);
not (n2456,n2457);
nor (n2457,n2458,n2473);
nor (n2458,n2346,n2459);
nor (n2459,n2460,n2467);
nor (n2460,n2461,n2466);
nor (n2461,n2462,n2464);
nor (n2462,n2463,n2045);
nand (n2463,n1934,n1938);
not (n2464,n2465);
nand (n2465,n2046,n2050);
not (n2466,n2159);
not (n2467,n2468);
nor (n2468,n2469,n2471);
nor (n2469,n2470,n2267);
nand (n2470,n2161,n2165);
not (n2471,n2472);
nand (n2472,n2268,n2272);
not (n2473,n2474);
nor (n2474,n2475,n2482);
nor (n2475,n2476,n2481);
nor (n2476,n2477,n2479);
nor (n2477,n2478,n2398);
nand (n2478,n2349,n2353);
not (n2479,n2480);
nand (n2480,n2399,n2403);
not (n2481,n2431);
not (n2482,n2483);
nor (n2483,n2484,n2486);
nor (n2484,n2485,n2449);
nand (n2485,n2433,n2437);
not (n2486,n2487);
nand (n2487,n2450,n2454);
nand (n2488,n2489,n2908);
nand (n2489,n2490,n2801);
nor (n2490,n2491,n2786);
nor (n2491,n2492,n2657);
nand (n2492,n2493,n2634);
nor (n2493,n2494,n2611);
nor (n2494,n2495,n2584);
nand (n2495,n2496,n2541,n2583);
nand (n2496,n2497,n2509);
xor (n2497,n2498,n2504);
xor (n2498,n2499,n2500);
xor (n2499,n1802,n1806);
xor (n2500,n2501,n78);
or (n2501,n2502,n2503);
and (n2502,n1004,n105);
and (n2503,n1018,n109);
and (n2504,n78,n2505);
xor (n2505,n2506,n664);
or (n2506,n2507,n2508);
and (n2507,n631,n787);
and (n2508,n635,n791);
nand (n2509,n2510,n2527,n2540);
nand (n2510,n2511,n2512);
xor (n2511,n78,n2505);
nand (n2512,n2513,n2522,n2526);
nand (n2513,n2514,n2518);
xor (n2514,n2515,n189);
or (n2515,n2516,n2517);
and (n2516,n979,n326);
and (n2517,n981,n330);
xor (n2518,n2519,n328);
or (n2519,n2520,n2521);
and (n2520,n771,n662);
and (n2521,n975,n666);
nand (n2522,n2523,n2518);
and (n2523,n107,n2524);
xnor (n2524,n2525,n107);
nand (n2525,n1018,n187);
nand (n2526,n2514,n2523);
nand (n2527,n2528,n2512);
xor (n2528,n2529,n2536);
xor (n2529,n2530,n2534);
xnor (n2530,n2531,n789);
nor (n2531,n2532,n2533);
and (n2532,n297,n990);
and (n2533,n225,n992);
xnor (n2534,n2535,n78);
nand (n2535,n1018,n105);
xor (n2536,n2537,n189);
or (n2537,n2538,n2539);
and (n2538,n975,n326);
and (n2539,n979,n330);
nand (n2540,n2511,n2528);
nand (n2541,n2542,n2509);
xor (n2542,n2543,n2562);
xor (n2543,n2544,n2548);
nand (n2544,n2545,n2546,n2547);
nand (n2545,n2530,n2534);
nand (n2546,n2536,n2534);
nand (n2547,n2530,n2536);
xor (n2548,n2549,n2558);
xor (n2549,n2550,n2554);
xor (n2550,n2551,n189);
or (n2551,n2552,n2553);
and (n2552,n771,n326);
and (n2553,n975,n330);
xor (n2554,n2555,n328);
or (n2555,n2556,n2557);
and (n2556,n635,n662);
and (n2557,n637,n666);
xor (n2558,n2559,n107);
or (n2559,n2560,n2561);
and (n2560,n979,n187);
and (n2561,n981,n191);
nand (n2562,n2563,n2577,n2582);
nand (n2563,n2564,n2568);
xor (n2564,n2565,n328);
or (n2565,n2566,n2567);
and (n2566,n637,n662);
and (n2567,n771,n666);
and (n2568,n2569,n2573);
xnor (n2569,n2570,n789);
nor (n2570,n2571,n2572);
and (n2571,n631,n990);
and (n2572,n297,n992);
xor (n2573,n2574,n664);
or (n2574,n2575,n2576);
and (n2575,n635,n787);
and (n2576,n637,n791);
nand (n2577,n2578,n2568);
xor (n2578,n2579,n107);
or (n2579,n2580,n2581);
and (n2580,n981,n187);
and (n2581,n1004,n191);
nand (n2582,n2564,n2578);
nand (n2583,n2497,n2542);
xor (n2584,n2585,n2599);
xor (n2585,n2586,n2595);
xor (n2586,n2587,n2593);
xor (n2587,n2588,n2592);
xor (n2588,n2589,n78);
or (n2589,n2590,n2591);
and (n2590,n981,n105);
and (n2591,n1004,n109);
xor (n2592,n1746,n19);
xor (n2593,n2594,n1789);
xor (n2594,n1782,n1786);
nand (n2595,n2596,n2597,n2598);
nand (n2596,n2544,n2548);
nand (n2597,n2562,n2548);
nand (n2598,n2544,n2562);
xor (n2599,n2600,n2609);
xor (n2600,n2601,n2605);
nand (n2601,n2602,n2603,n2604);
nand (n2602,n2499,n2500);
nand (n2603,n2504,n2500);
nand (n2604,n2499,n2504);
nand (n2605,n2606,n2607,n2608);
nand (n2606,n2550,n2554);
nand (n2607,n2558,n2554);
nand (n2608,n2550,n2558);
xor (n2609,n2610,n1811);
xor (n2610,n1797,n1801);
nor (n2611,n2612,n2616);
nand (n2612,n2613,n2614,n2615);
nand (n2613,n2586,n2595);
nand (n2614,n2599,n2595);
nand (n2615,n2586,n2599);
xor (n2616,n2617,n2624);
xor (n2617,n2618,n2620);
xor (n2618,n2619,n1795);
xor (n2619,n1776,n1780);
nand (n2620,n2621,n2622,n2623);
nand (n2621,n2601,n2605);
nand (n2622,n2609,n2605);
nand (n2623,n2601,n2609);
xor (n2624,n2625,n2630);
xor (n2625,n2626,n2628);
xor (n2626,n2627,n1745);
xor (n2627,n1736,n1740);
xor (n2628,n2629,n1760);
xor (n2629,n1754,n1758);
nand (n2630,n2631,n2632,n2633);
nand (n2631,n2588,n2592);
nand (n2632,n2593,n2592);
nand (n2633,n2588,n2593);
nor (n2634,n2635,n2650);
nor (n2635,n2636,n2640);
nand (n2636,n2637,n2638,n2639);
nand (n2637,n2618,n2620);
nand (n2638,n2624,n2620);
nand (n2639,n2618,n2624);
xor (n2640,n2641,n2648);
xor (n2641,n2642,n2644);
xor (n2642,n2643,n1752);
xor (n2643,n1732,n1734);
nand (n2644,n2645,n2646,n2647);
nand (n2645,n2626,n2628);
nand (n2646,n2630,n2628);
nand (n2647,n2626,n2630);
xor (n2648,n2649,n1774);
xor (n2649,n1769,n1771);
nor (n2650,n2651,n2655);
nand (n2651,n2652,n2653,n2654);
nand (n2652,n2642,n2644);
nand (n2653,n2648,n2644);
nand (n2654,n2642,n2648);
xor (n2655,n2656,n1767);
xor (n2656,n1642,n1693);
nor (n2657,n2658,n2780);
nor (n2658,n2659,n2756);
nor (n2659,n2660,n2753);
nor (n2660,n2661,n2729);
nand (n2661,n2662,n2701);
or (n2662,n2663,n2687,n2700);
and (n2663,n2664,n2673);
xor (n2664,n2665,n2669);
xnor (n2665,n2666,n789);
nor (n2666,n2667,n2668);
and (n2667,n637,n990);
and (n2668,n635,n992);
xnor (n2669,n2670,n664);
nor (n2670,n2671,n2672);
and (n2671,n975,n791);
and (n2672,n771,n787);
or (n2673,n2674,n2681,n2686);
and (n2674,n2675,n2677);
not (n2675,n2676);
nand (n2676,n1018,n326);
xnor (n2677,n2678,n789);
nor (n2678,n2679,n2680);
and (n2679,n771,n990);
and (n2680,n637,n992);
and (n2681,n2677,n2682);
xnor (n2682,n2683,n664);
nor (n2683,n2684,n2685);
and (n2684,n979,n791);
and (n2685,n975,n787);
and (n2686,n2675,n2682);
and (n2687,n2673,n2688);
xor (n2688,n2689,n2696);
xor (n2689,n2690,n2692);
and (n2690,n189,n2691);
xnor (n2691,n2676,n189);
xnor (n2692,n2693,n328);
nor (n2693,n2694,n2695);
and (n2694,n981,n666);
and (n2695,n979,n662);
xnor (n2696,n2697,n189);
nor (n2697,n2698,n2699);
and (n2698,n1018,n330);
and (n2699,n1004,n326);
and (n2700,n2664,n2688);
xor (n2701,n2702,n2718);
xor (n2702,n2703,n2707);
or (n2703,n2704,n2705,n2706);
and (n2704,n2690,n2692);
and (n2705,n2692,n2696);
and (n2706,n2690,n2696);
xor (n2707,n2708,n2714);
xor (n2708,n2709,n2710);
and (n2709,n2665,n2669);
xnor (n2710,n2711,n328);
nor (n2711,n2712,n2713);
and (n2712,n979,n666);
and (n2713,n975,n662);
xnor (n2714,n2715,n189);
nor (n2715,n2716,n2717);
and (n2716,n1004,n330);
and (n2717,n981,n326);
xor (n2718,n2719,n2725);
xor (n2719,n2720,n2721);
not (n2720,n2525);
xnor (n2721,n2722,n789);
nor (n2722,n2723,n2724);
and (n2723,n635,n990);
and (n2724,n631,n992);
xnor (n2725,n2726,n664);
nor (n2726,n2727,n2728);
and (n2727,n771,n791);
and (n2728,n637,n787);
nor (n2729,n2730,n2734);
or (n2730,n2731,n2732,n2733);
and (n2731,n2703,n2707);
and (n2732,n2707,n2718);
and (n2733,n2703,n2718);
xor (n2734,n2735,n2742);
xor (n2735,n2736,n2740);
or (n2736,n2737,n2738,n2739);
and (n2737,n2709,n2710);
and (n2738,n2710,n2714);
and (n2739,n2709,n2714);
xor (n2740,n2741,n2523);
xor (n2741,n2514,n2518);
xor (n2742,n2743,n2749);
xor (n2743,n2744,n2748);
xor (n2744,n2745,n107);
or (n2745,n2746,n2747);
and (n2746,n1004,n187);
and (n2747,n1018,n191);
xor (n2748,n2569,n2573);
or (n2749,n2750,n2751,n2752);
and (n2750,n2720,n2721);
and (n2751,n2721,n2725);
and (n2752,n2720,n2725);
not (n2753,n2754);
not (n2754,n2755);
and (n2755,n2730,n2734);
not (n2756,n2757);
nor (n2757,n2758,n2773);
nor (n2758,n2759,n2763);
nand (n2759,n2760,n2761,n2762);
nand (n2760,n2736,n2740);
nand (n2761,n2742,n2740);
nand (n2762,n2736,n2742);
xor (n2763,n2764,n2771);
xor (n2764,n2765,n2767);
xor (n2765,n2766,n2578);
xor (n2766,n2564,n2568);
nand (n2767,n2768,n2769,n2770);
nand (n2768,n2744,n2748);
nand (n2769,n2749,n2748);
nand (n2770,n2744,n2749);
xor (n2771,n2772,n2528);
xor (n2772,n2511,n2512);
nor (n2773,n2774,n2778);
nand (n2774,n2775,n2776,n2777);
nand (n2775,n2765,n2767);
nand (n2776,n2771,n2767);
nand (n2777,n2765,n2771);
xor (n2778,n2779,n2542);
xor (n2779,n2497,n2509);
not (n2780,n2781);
nor (n2781,n2782,n2784);
nor (n2782,n2783,n2773);
nand (n2783,n2759,n2763);
not (n2784,n2785);
nand (n2785,n2774,n2778);
not (n2786,n2787);
nor (n2787,n2788,n2795);
nor (n2788,n2789,n2794);
nor (n2789,n2790,n2792);
nor (n2790,n2791,n2611);
nand (n2791,n2495,n2584);
not (n2792,n2793);
nand (n2793,n2612,n2616);
not (n2794,n2634);
not (n2795,n2796);
nor (n2796,n2797,n2799);
nor (n2797,n2798,n2650);
nand (n2798,n2636,n2640);
not (n2799,n2800);
nand (n2800,n2651,n2655);
nand (n2801,n2802,n2806);
nor (n2802,n2803,n2492);
nand (n2803,n2804,n2757);
nor (n2804,n2805,n2729);
nor (n2805,n2662,n2701);
or (n2806,n2807,n2829);
and (n2807,n2808,n2810);
xor (n2808,n2809,n2688);
xor (n2809,n2664,n2673);
or (n2810,n2811,n2825,n2828);
and (n2811,n2812,n2821);
and (n2812,n2813,n2817);
xnor (n2813,n2814,n789);
nor (n2814,n2815,n2816);
and (n2815,n975,n990);
and (n2816,n771,n992);
xnor (n2817,n2818,n664);
nor (n2818,n2819,n2820);
and (n2819,n981,n791);
and (n2820,n979,n787);
xnor (n2821,n2822,n328);
nor (n2822,n2823,n2824);
and (n2823,n1004,n666);
and (n2824,n981,n662);
and (n2825,n2821,n2826);
xor (n2826,n2827,n2682);
xor (n2827,n2675,n2677);
and (n2828,n2812,n2826);
and (n2829,n2830,n2831);
xor (n2830,n2808,n2810);
or (n2831,n2832,n2847);
and (n2832,n2833,n2845);
or (n2833,n2834,n2839,n2844);
and (n2834,n2835,n2836);
xor (n2835,n2813,n2817);
and (n2836,n328,n2837);
xnor (n2837,n2838,n328);
nand (n2838,n1018,n662);
and (n2839,n2836,n2840);
xnor (n2840,n2841,n328);
nor (n2841,n2842,n2843);
and (n2842,n1018,n666);
and (n2843,n1004,n662);
and (n2844,n2835,n2840);
xor (n2845,n2846,n2826);
xor (n2846,n2812,n2821);
and (n2847,n2848,n2849);
xor (n2848,n2833,n2845);
or (n2849,n2850,n2866);
and (n2850,n2851,n2853);
xor (n2851,n2852,n2840);
xor (n2852,n2835,n2836);
or (n2853,n2854,n2860,n2865);
and (n2854,n2855,n2856);
not (n2855,n2838);
xnor (n2856,n2857,n789);
nor (n2857,n2858,n2859);
and (n2858,n979,n990);
and (n2859,n975,n992);
and (n2860,n2856,n2861);
xnor (n2861,n2862,n664);
nor (n2862,n2863,n2864);
and (n2863,n1004,n791);
and (n2864,n981,n787);
and (n2865,n2855,n2861);
and (n2866,n2867,n2868);
xor (n2867,n2851,n2853);
or (n2868,n2869,n2880);
and (n2869,n2870,n2872);
xor (n2870,n2871,n2861);
xor (n2871,n2855,n2856);
and (n2872,n2873,n2876);
and (n2873,n664,n2874);
xnor (n2874,n2875,n664);
nand (n2875,n1018,n787);
xnor (n2876,n2877,n789);
nor (n2877,n2878,n2879);
and (n2878,n981,n990);
and (n2879,n979,n992);
and (n2880,n2881,n2882);
xor (n2881,n2870,n2872);
or (n2882,n2883,n2889);
and (n2883,n2884,n2888);
xnor (n2884,n2885,n664);
nor (n2885,n2886,n2887);
and (n2886,n1018,n791);
and (n2887,n1004,n787);
xor (n2888,n2873,n2876);
and (n2889,n2890,n2891);
xor (n2890,n2884,n2888);
or (n2891,n2892,n2898);
and (n2892,n2893,n2897);
xnor (n2893,n2894,n789);
nor (n2894,n2895,n2896);
and (n2895,n1004,n990);
and (n2896,n981,n992);
not (n2897,n2875);
and (n2898,n2899,n2900);
xor (n2899,n2893,n2897);
and (n2900,n2901,n2905);
xnor (n2901,n2902,n789);
nor (n2902,n2903,n2904);
and (n2903,n1018,n990);
and (n2904,n1004,n992);
and (n2905,n2906,n789);
xnor (n2906,n2907,n789);
nand (n2907,n1018,n992);
not (n2908,n2909);
nand (n2909,n2910,n1930);
nor (n2910,n2911,n962);
nand (n2911,n2912,n1885);
nor (n2912,n2913,n1857);
nor (n2913,n1640,n1819);
nand (n2914,n2915,n2961);
not (n2915,n2916);
nor (n2916,n2917,n2921);
nand (n2917,n2918,n2919,n2920);
nand (n2918,n489,n493);
nand (n2919,n526,n493);
nand (n2920,n489,n526);
xor (n2921,n2922,n2957);
xor (n2922,n2923,n2927);
nand (n2923,n2924,n2925,n2926);
nand (n2924,n465,n511);
nand (n2925,n515,n511);
nand (n2926,n465,n515);
xor (n2927,n2928,n2947);
xor (n2928,n2929,n2943);
xor (n2929,n2930,n2939);
xor (n2930,n2931,n2935);
xor (n2931,n2932,n46);
or (n2932,n2933,n2934);
and (n2933,n16,n40);
and (n2934,n21,n44);
xor (n2935,n2936,n70);
or (n2936,n2937,n2938);
and (n2937,n39,n64);
and (n2938,n43,n68);
xor (n2939,n2940,n59);
or (n2940,n2941,n2942);
and (n2941,n28,n53);
and (n2942,n32,n57);
nand (n2943,n2944,n2945,n2946);
nand (n2944,n501,n505);
nand (n2945,n70,n505);
nand (n2946,n501,n70);
xor (n2947,n2948,n2953);
xor (n2948,n2949,n70);
not (n2949,n2950);
xor (n2950,n2951,n35);
or (n2951,n520,n2952);
and (n2952,n75,n33);
nand (n2953,n2954,n2955,n2956);
nand (n2954,n517,n518);
nand (n2955,n522,n518);
nand (n2956,n517,n522);
nand (n2957,n2958,n2959,n2960);
nand (n2958,n495,n499);
nand (n2959,n509,n499);
nand (n2960,n495,n509);
nand (n2961,n2917,n2921);
xor (n2962,n2963,n3200);
xor (n2963,n2964,n3088);
xor (n2964,n2965,n3003);
xor (n2965,n2966,n2990);
xor (n2966,n2967,n2976);
or (n2967,n2968,n2973,n2975);
and (n2968,n2969,n465);
or (n2969,n2970,n2971,n2972);
and (n2970,n517,n448);
not (n2971,n513);
and (n2972,n517,n452);
and (n2973,n465,n2974);
not (n2974,n515);
and (n2975,n2969,n2974);
xor (n2976,n2977,n2987);
xor (n2977,n2978,n2982);
or (n2978,n2979,n2980,n2981);
and (n2979,n445,n518);
not (n2980,n2955);
and (n2981,n445,n522);
or (n2982,n2983,n2984,n2986);
and (n2983,n517,n500);
and (n2984,n500,n2985);
not (n2985,n496);
and (n2986,n517,n2985);
xor (n2987,n2988,n2989);
xor (n2988,n2950,n2929);
not (n2989,n2944);
or (n2990,n2991,n2999,n3002);
and (n2991,n2992,n2997);
or (n2992,n2993,n2995,n2996);
and (n2993,n2994,n459);
not (n2994,n443);
and (n2995,n459,n435);
and (n2996,n2994,n435);
xor (n2997,n2998,n2985);
xor (n2998,n517,n500);
and (n2999,n2997,n3000);
xor (n3000,n3001,n2974);
xor (n3001,n2969,n465);
and (n3002,n2992,n3000);
or (n3003,n3004,n3025,n3087);
and (n3004,n3005,n3023);
or (n3005,n3006,n3019,n3022);
and (n3006,n3007,n3011);
or (n3007,n3008,n3009,n3010);
not (n3008,n442);
and (n3009,n417,n471);
and (n3010,n413,n471);
or (n3011,n3012,n3017,n3018);
and (n3012,n391,n3013);
or (n3013,n3014,n3015,n3016);
and (n3014,n72,n49);
not (n3015,n398);
and (n3016,n72,n60);
and (n3017,n3013,n401);
and (n3018,n391,n401);
and (n3019,n3011,n3020);
xor (n3020,n3021,n435);
xor (n3021,n2994,n459);
and (n3022,n3007,n3020);
xor (n3023,n3024,n3000);
xor (n3024,n2992,n2997);
and (n3025,n3023,n3026);
or (n3026,n3027,n3040,n3086);
and (n3027,n3028,n3038);
or (n3028,n3029,n3034,n3037);
and (n3029,n3030,n3032);
xor (n3030,n3031,n471);
xor (n3031,n413,n417);
and (n3032,n11,n3033);
not (n3033,n47);
and (n3034,n3032,n3035);
xor (n3035,n3036,n401);
xor (n3036,n391,n3013);
and (n3037,n3030,n3035);
xor (n3038,n3039,n3020);
xor (n3039,n3007,n3011);
and (n3040,n3038,n3041);
or (n3041,n3042,n3055,n3085);
and (n3042,n3043,n3053);
or (n3043,n3044,n3050,n3052);
and (n3044,n3045,n3046);
not (n3045,n83);
or (n3046,n3047,n3048,n3049);
not (n3047,n100);
and (n3048,n111,n122);
and (n3049,n101,n122);
and (n3050,n3046,n3051);
not (n3051,n10);
and (n3052,n3045,n3051);
xor (n3053,n3054,n3035);
xor (n3054,n3030,n3032);
and (n3055,n3053,n3056);
or (n3056,n3057,n3071,n3084);
and (n3057,n3058,n3062);
or (n3058,n3059,n3060,n3061);
and (n3059,n115,n127);
and (n3060,n127,n169);
and (n3061,n115,n169);
or (n3062,n3063,n3068,n3070);
and (n3063,n136,n3064);
or (n3064,n3065,n3066,n3067);
and (n3065,n102,n155);
not (n3066,n159);
and (n3067,n102,n160);
and (n3068,n3064,n3069);
xor (n3069,n135,n122);
and (n3070,n136,n3069);
and (n3071,n3062,n3072);
or (n3072,n3073,n3080,n3083);
and (n3073,n3074,n3075);
not (n3074,n207);
or (n3075,n3076,n3078,n3079);
and (n3076,n175,n3077);
not (n3077,n251);
and (n3078,n3077,n181);
not (n3079,n202);
and (n3080,n3075,n3081);
xor (n3081,n3082,n169);
xor (n3082,n115,n127);
and (n3083,n3074,n3081);
and (n3084,n3058,n3072);
and (n3085,n3043,n3056);
and (n3086,n3028,n3041);
and (n3087,n3005,n3026);
or (n3088,n3089,n3091);
xor (n3089,n3090,n3026);
xor (n3090,n3005,n3023);
or (n3091,n3092,n3094);
xor (n3092,n3093,n3041);
xor (n3093,n3028,n3038);
or (n3094,n3095,n3127,n3199);
and (n3095,n3096,n3125);
or (n3096,n3097,n3121,n3124);
and (n3097,n3098,n3100);
xor (n3098,n3099,n3051);
xor (n3099,n3045,n3046);
or (n3100,n3101,n3117,n3120);
and (n3101,n3102,n3104);
xor (n3102,n3103,n3069);
xor (n3103,n136,n3064);
or (n3104,n3105,n3111,n3116);
and (n3105,n284,n3106);
and (n3106,n3107,n300);
or (n3107,n3108,n3109,n3110);
and (n3108,n184,n289);
not (n3109,n288);
and (n3110,n184,n293);
and (n3111,n3106,n3112);
or (n3112,n3113,n3114,n3115);
not (n3113,n234);
and (n3114,n235,n260);
and (n3115,n230,n260);
and (n3116,n284,n3112);
and (n3117,n3104,n3118);
xor (n3118,n3119,n3081);
xor (n3119,n3074,n3075);
and (n3120,n3102,n3118);
and (n3121,n3100,n3122);
xor (n3122,n3123,n3072);
xor (n3123,n3058,n3062);
and (n3124,n3098,n3122);
xor (n3125,n3126,n3056);
xor (n3126,n3043,n3053);
and (n3127,n3125,n3128);
or (n3128,n3129,n3131);
xor (n3129,n3130,n3122);
xor (n3130,n3098,n3100);
or (n3131,n3132,n3163,n3198);
and (n3132,n3133,n3161);
or (n3133,n3134,n3143,n3160);
and (n3134,n3135,n3137);
xor (n3135,n3136,n181);
xor (n3136,n175,n3077);
or (n3137,n3138,n3140,n3142);
and (n3138,n3139,n257);
not (n3139,n310);
and (n3140,n257,n3141);
xor (n3141,n3107,n300);
and (n3142,n3139,n3141);
and (n3143,n3137,n3144);
or (n3144,n3145,n3156,n3159);
and (n3145,n3146,n3151);
or (n3146,n3147,n3149,n3150);
and (n3147,n344,n3148);
not (n3148,n862);
and (n3149,n3148,n861);
and (n3150,n344,n861);
or (n3151,n3152,n3154,n3155);
and (n3152,n347,n3153);
not (n3153,n857);
and (n3154,n3153,n320);
and (n3155,n347,n320);
and (n3156,n3151,n3157);
xor (n3157,n3158,n260);
xor (n3158,n230,n235);
and (n3159,n3146,n3157);
and (n3160,n3135,n3144);
xor (n3161,n3162,n3118);
xor (n3162,n3102,n3104);
and (n3163,n3161,n3164);
or (n3164,n3165,n3194,n3197);
and (n3165,n3166,n3168);
xor (n3166,n3167,n3112);
xor (n3167,n284,n3106);
or (n3168,n3169,n3190,n3193);
and (n3169,n3170,n3188);
or (n3170,n3171,n3184,n3187);
and (n3171,n3172,n3176);
or (n3172,n3173,n3174,n3175);
and (n3173,n541,n615);
and (n3174,n615,n684);
and (n3175,n541,n684);
or (n3176,n3177,n3178,n3183);
and (n3177,n545,n617);
and (n3178,n617,n3179);
or (n3179,n3180,n3181,n3182);
and (n3180,n323,n646);
not (n3181,n682);
and (n3182,n323,n642);
and (n3183,n545,n3179);
and (n3184,n3176,n3185);
xor (n3185,n3186,n861);
xor (n3186,n344,n3148);
and (n3187,n3172,n3185);
xor (n3188,n3189,n3141);
xor (n3189,n3139,n257);
and (n3190,n3188,n3191);
xor (n3191,n3192,n3157);
xor (n3192,n3146,n3151);
and (n3193,n3170,n3191);
and (n3194,n3168,n3195);
xor (n3195,n3196,n3144);
xor (n3196,n3135,n3137);
and (n3197,n3166,n3195);
and (n3198,n3133,n3164);
and (n3199,n3096,n3128);
and (n3200,n3201,n3202);
xnor (n3201,n3089,n3091);
and (n3202,n3203,n3204);
xnor (n3203,n3092,n3094);
and (n3204,n3205,n3207);
xor (n3205,n3206,n3128);
xor (n3206,n3096,n3125);
and (n3207,n3208,n3209);
xnor (n3208,n3129,n3131);
or (n3209,n3210,n3290);
and (n3210,n3211,n3213);
xor (n3211,n3212,n3164);
xor (n3212,n3133,n3161);
or (n3213,n3214,n3216);
xor (n3214,n3215,n3195);
xor (n3215,n3166,n3168);
or (n3216,n3217,n3240,n3289);
and (n3217,n3218,n3238);
or (n3218,n3219,n3234,n3237);
and (n3219,n3220,n3222);
xor (n3220,n3221,n320);
xor (n3221,n347,n3153);
or (n3222,n3223,n3230,n3233);
and (n3223,n613,n3224);
or (n3224,n3225,n3227,n3229);
and (n3225,n674,n3226);
not (n3226,n640);
and (n3227,n3226,n3228);
not (n3228,n626);
and (n3229,n674,n3228);
and (n3230,n3224,n3231);
xor (n3231,n3232,n684);
xor (n3232,n541,n615);
and (n3233,n613,n3231);
and (n3234,n3222,n3235);
xor (n3235,n3236,n3185);
xor (n3236,n3172,n3176);
and (n3237,n3220,n3235);
xor (n3238,n3239,n3191);
xor (n3239,n3170,n3188);
and (n3240,n3238,n3241);
or (n3241,n3242,n3253,n3288);
and (n3242,n3243,n3251);
or (n3243,n3244,n3247,n3250);
and (n3244,n3245,n561);
xor (n3245,n3246,n3179);
xor (n3246,n545,n617);
and (n3247,n561,n3248);
xor (n3248,n3249,n3231);
xor (n3249,n613,n3224);
and (n3250,n3245,n3248);
xor (n3251,n3252,n3235);
xor (n3252,n3220,n3222);
and (n3253,n3251,n3254);
or (n3254,n3255,n3284,n3287);
and (n3255,n3256,n3269);
or (n3256,n3257,n3267,n3268);
and (n3257,n3258,n719);
or (n3258,n3259,n3264,n3266);
and (n3259,n3260,n713);
or (n3260,n3261,n3262,n3263);
and (n3261,n658,n703);
not (n3262,n707);
and (n3263,n658,n708);
and (n3264,n713,n3265);
not (n3265,n716);
and (n3266,n3260,n3265);
not (n3267,n754);
and (n3268,n3258,n755);
or (n3269,n3270,n3277,n3283);
and (n3270,n3271,n3275);
or (n3271,n3272,n3273,n3274);
and (n3272,n659,n655);
not (n3273,n673);
and (n3274,n659,n669);
xor (n3275,n3276,n3228);
xor (n3276,n674,n3226);
and (n3277,n3275,n3278);
or (n3278,n3279,n3280,n3282);
and (n3279,n658,n796);
and (n3280,n796,n3281);
not (n3281,n2410);
and (n3282,n658,n3281);
and (n3283,n3271,n3278);
and (n3284,n3269,n3285);
xor (n3285,n3286,n3248);
xor (n3286,n3245,n561);
and (n3287,n3256,n3285);
and (n3288,n3243,n3254);
and (n3289,n3218,n3241);
and (n3290,n3291,n3292);
xor (n3291,n3211,n3213);
and (n3292,n3293,n3294);
xnor (n3293,n3214,n3216);
or (n3294,n3295,n3380);
and (n3295,n3296,n3298);
xor (n3296,n3297,n3241);
xor (n3297,n3218,n3238);
or (n3298,n3299,n3301);
xor (n3299,n3300,n3254);
xor (n3300,n3243,n3251);
or (n3301,n3302,n3324,n3379);
and (n3302,n3303,n3322);
or (n3303,n3304,n3318,n3321);
and (n3304,n3305,n3307);
xor (n3305,n3306,n755);
xor (n3306,n3258,n719);
or (n3307,n3308,n3311,n3317);
and (n3308,n3309,n2413);
xor (n3309,n3310,n3265);
xor (n3310,n3260,n713);
and (n3311,n2413,n3312);
or (n3312,n3313,n3314,n3316);
not (n3313,n835);
and (n3314,n819,n3315);
not (n3315,n816);
and (n3316,n800,n3315);
and (n3317,n3309,n3312);
and (n3318,n3307,n3319);
xor (n3319,n3320,n3278);
xor (n3320,n3271,n3275);
and (n3321,n3305,n3319);
xor (n3322,n3323,n3285);
xor (n3323,n3256,n3269);
and (n3324,n3322,n3325);
or (n3325,n3326,n3341,n3378);
and (n3326,n3327,n3339);
or (n3327,n3328,n3335,n3338);
and (n3328,n3329,n3333);
or (n3329,n3330,n3331,n3332);
and (n3330,n767,n2383);
and (n3331,n2383,n2364);
and (n3332,n767,n2364);
xor (n3333,n3334,n3281);
xor (n3334,n658,n796);
and (n3335,n3333,n3336);
and (n3336,n2359,n3337);
not (n3337,n2357);
and (n3338,n3329,n3336);
xor (n3339,n3340,n3319);
xor (n3340,n3305,n3307);
and (n3341,n3339,n3342);
or (n3342,n3343,n3363,n3377);
and (n3343,n3344,n3361);
or (n3344,n3345,n3350,n3360);
and (n3345,n3346,n2386);
or (n3346,n3347,n3348,n3349);
and (n3347,n784,n775);
not (n3348,n774);
and (n3349,n784,n778);
and (n3350,n2386,n3351);
or (n3351,n3352,n3357,n3359);
and (n3352,n783,n3353);
or (n3353,n3354,n3355,n3356);
and (n3354,n783,n2187);
not (n3355,n2301);
and (n3356,n783,n2191);
and (n3357,n3353,n3358);
not (n3358,n2296);
and (n3359,n783,n3358);
and (n3360,n3346,n3351);
xor (n3361,n3362,n3312);
xor (n3362,n3309,n2413);
and (n3363,n3361,n3364);
or (n3364,n3365,n3369,n3376);
and (n3365,n3366,n3368);
xor (n3366,n3367,n2364);
xor (n3367,n767,n2383);
not (n3368,n2356);
and (n3369,n3368,n3370);
or (n3370,n3371,n3374,n3375);
and (n3371,n3372,n2302);
and (n3372,n2171,n3373);
not (n3373,n2185);
and (n3374,n2302,n2324);
and (n3375,n3372,n2324);
and (n3376,n3366,n3370);
and (n3377,n3344,n3364);
and (n3378,n3327,n3342);
and (n3379,n3303,n3325);
and (n3380,n3381,n3382);
xor (n3381,n3296,n3298);
and (n3382,n3383,n3384);
xnor (n3383,n3299,n3301);
or (n3384,n3385,n3589);
and (n3385,n3386,n3388);
xor (n3386,n3387,n3325);
xor (n3387,n3303,n3322);
or (n3388,n3389,n3464,n3588);
and (n3389,n3390,n3462);
or (n3390,n3391,n3458,n3461);
and (n3391,n3392,n3394);
xor (n3392,n3393,n3336);
xor (n3393,n3329,n3333);
or (n3394,n3395,n3429,n3457);
and (n3395,n3396,n3427);
or (n3396,n3397,n3415,n3426);
and (n3397,n3398,n3407);
and (n3398,n3399,n2211);
or (n3399,n3400,n3405,n3406);
and (n3400,n3401,n2081);
or (n3401,n3402,n3403,n3404);
and (n3402,n2150,n1946);
not (n3403,n2090);
and (n3404,n2150,n1950);
not (n3405,n2223);
and (n3406,n3401,n2085);
or (n3407,n3408,n3413,n3414);
and (n3408,n2251,n3409);
or (n3409,n3410,n3411,n3412);
and (n3410,n2150,n2070);
not (n3411,n2198);
and (n3412,n2150,n2075);
and (n3413,n3409,n2232);
and (n3414,n2251,n2232);
and (n3415,n3407,n3416);
or (n3416,n3417,n3423,n3425);
and (n3417,n3418,n3419);
not (n3418,n2170);
or (n3419,n3420,n3421,n3422);
and (n3420,n1954,n2146);
not (n3421,n2250);
and (n3422,n1954,n2151);
and (n3423,n3419,n3424);
not (n3424,n2227);
and (n3425,n3418,n3424);
and (n3426,n3398,n3416);
xor (n3427,n3428,n3351);
xor (n3428,n3346,n2386);
and (n3429,n3427,n3430);
or (n3430,n3431,n3453,n3456);
and (n3431,n3432,n3434);
xor (n3432,n3433,n3358);
xor (n3433,n783,n3353);
or (n3434,n3435,n3444,n3452);
and (n3435,n3436,n3443);
or (n3436,n3437,n3439,n3442);
and (n3437,n2130,n3438);
not (n3438,n2127);
and (n3439,n3438,n3440);
xor (n3440,n3441,n2075);
xor (n3441,n2150,n2070);
and (n3442,n2130,n3440);
xor (n3443,n3399,n2211);
and (n3444,n3443,n3445);
or (n3445,n3446,n3450,n3451);
and (n3446,n3447,n3448);
not (n3447,n2144);
xor (n3448,n3449,n2085);
xor (n3449,n3401,n2081);
and (n3450,n3448,n2104);
and (n3451,n3447,n2104);
and (n3452,n3436,n3445);
and (n3453,n3434,n3454);
xor (n3454,n3455,n2324);
xor (n3455,n3372,n2302);
and (n3456,n3432,n3454);
and (n3457,n3396,n3430);
and (n3458,n3394,n3459);
xor (n3459,n3460,n3364);
xor (n3460,n3344,n3361);
and (n3461,n3392,n3459);
xor (n3462,n3463,n3342);
xor (n3463,n3327,n3339);
and (n3464,n3462,n3465);
or (n3465,n3466,n3499,n3587);
and (n3466,n3467,n3497);
or (n3467,n3468,n3493,n3496);
and (n3468,n3469,n3471);
xor (n3469,n3470,n3370);
xor (n3470,n3366,n3368);
or (n3471,n3472,n3489,n3492);
and (n3472,n3473,n3475);
xor (n3473,n3474,n3416);
xor (n3474,n3398,n3407);
or (n3475,n3476,n3481,n3488);
and (n3476,n3477,n3479);
xor (n3477,n3478,n2232);
xor (n3478,n2251,n3409);
xor (n3479,n3480,n3424);
xor (n3480,n3418,n3419);
and (n3481,n3479,n3482);
and (n3482,n2095,n3483);
or (n3483,n3484,n3485,n3487);
not (n3484,n2101);
and (n3485,n1961,n3486);
not (n3486,n1944);
and (n3487,n1957,n3486);
and (n3488,n3477,n3482);
and (n3489,n3475,n3490);
xor (n3490,n3491,n3454);
xor (n3491,n3432,n3434);
and (n3492,n3473,n3490);
and (n3493,n3471,n3494);
xor (n3494,n3495,n3430);
xor (n3495,n3396,n3427);
and (n3496,n3469,n3494);
xor (n3497,n3498,n3459);
xor (n3498,n3392,n3394);
and (n3499,n3497,n3500);
or (n3500,n3501,n3558,n3586);
and (n3501,n3502,n3504);
xor (n3502,n3503,n3494);
xor (n3503,n3469,n3471);
or (n3504,n3505,n3537,n3557);
and (n3505,n3506,n3535);
or (n3506,n3507,n3520,n3534);
and (n3507,n3508,n3518);
or (n3508,n3509,n3516,n3517);
and (n3509,n3510,n3514);
or (n3510,n3511,n3512,n3513);
and (n3511,n2009,n1994);
and (n3512,n1994,n1977);
and (n3513,n2009,n1977);
xor (n3514,n3515,n3440);
xor (n3515,n2130,n3438);
and (n3516,n3514,n2155);
and (n3517,n3510,n2155);
xor (n3518,n3519,n3445);
xor (n3519,n3436,n3443);
and (n3520,n3518,n3521);
or (n3521,n3522,n3531,n3533);
and (n3522,n3523,n3529);
or (n3523,n3524,n3525,n3528);
and (n3524,n1999,n1993);
and (n3525,n1993,n3526);
xor (n3526,n3527,n1977);
xor (n3527,n2009,n1994);
and (n3528,n1999,n3526);
xor (n3529,n3530,n2104);
xor (n3530,n3447,n3448);
and (n3531,n3529,n3532);
xor (n3532,n2095,n3483);
and (n3533,n3523,n3532);
and (n3534,n3508,n3521);
xor (n3535,n3536,n3490);
xor (n3536,n3473,n3475);
and (n3537,n3535,n3538);
or (n3538,n3539,n3553,n3556);
and (n3539,n3540,n3542);
xor (n3540,n3541,n3482);
xor (n3541,n3477,n3479);
or (n3542,n3543,n3551,n3552);
and (n3543,n3544,n3546);
xor (n3544,n3545,n2155);
xor (n3545,n3510,n3514);
or (n3546,n3547,n3548,n3550);
not (n3547,n2054);
and (n3548,n1969,n3549);
not (n3549,n1942);
and (n3550,n1965,n3549);
and (n3551,n3546,n2056);
and (n3552,n3544,n2056);
and (n3553,n3542,n3554);
xor (n3554,n3555,n3521);
xor (n3555,n3508,n3518);
and (n3556,n3540,n3554);
and (n3557,n3506,n3538);
and (n3558,n3504,n3559);
or (n3559,n3560,n3562);
xor (n3560,n3561,n3538);
xor (n3561,n3506,n3535);
or (n3562,n3563,n3579,n3585);
and (n3563,n3564,n3577);
or (n3564,n3565,n3573,n3576);
and (n3565,n3566,n3568);
xor (n3566,n3567,n3532);
xor (n3567,n3523,n3529);
or (n3568,n3569,n3571,n3572);
and (n3569,n3570,n2041);
not (n3570,n1940);
not (n3571,n2048);
and (n3572,n3570,n1973);
and (n3573,n3568,n3574);
xor (n3574,n3575,n2056);
xor (n3575,n3544,n3546);
and (n3576,n3566,n3574);
xor (n3577,n3578,n3554);
xor (n3578,n3540,n3542);
and (n3579,n3577,n3580);
or (n3580,n3581,n3583);
or (n3581,n1934,n3582);
not (n3582,n1938);
xor (n3583,n3584,n3574);
xor (n3584,n3566,n3568);
and (n3585,n3564,n3580);
and (n3586,n3502,n3559);
and (n3587,n3467,n3500);
and (n3588,n3390,n3465);
and (n3589,n3590,n3591);
xor (n3590,n3386,n3388);
and (n3591,n3592,n3594);
xor (n3592,n3593,n3465);
xor (n3593,n3390,n3462);
or (n3594,n3595,n3597);
xor (n3595,n3596,n3500);
xor (n3596,n3467,n3497);
and (n3597,n3598,n3599);
not (n3598,n3595);
and (n3599,n3600,n3602);
xor (n3600,n3601,n3559);
xor (n3601,n3502,n3504);
and (n3602,n3603,n3604);
xnor (n3603,n3560,n3562);
and (n3604,n3605,n3607);
xor (n3605,n3606,n3580);
xor (n3606,n3564,n3577);
and (n3607,n3608,n3609);
xnor (n3608,n3581,n3583);
and (n3609,n3610,n3613);
not (n3610,n3611);
nand (n3611,n3612,n2463);
not (n3612,n1933);
nand (n3613,n960,n3614);
nand (n3614,n2910,n2489);
endmodule
