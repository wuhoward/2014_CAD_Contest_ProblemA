module top (out,n7,n19,n21,n22,n24,n26,n27,n32,n39
        ,n46,n52,n55,n56,n74,n75,n87,n88,n94,n95
        ,n114,n115,n121,n122,n127,n133,n142,n151,n166,n179
        ,n185,n204,n210,n670,n682,n697,n704,n708,n713,n718
        ,n724,n730,n735,n757,n768,n783,n794);
output out;
input n7;
input n19;
input n21;
input n22;
input n24;
input n26;
input n27;
input n32;
input n39;
input n46;
input n52;
input n55;
input n56;
input n74;
input n75;
input n87;
input n88;
input n94;
input n95;
input n114;
input n115;
input n121;
input n122;
input n127;
input n133;
input n142;
input n151;
input n166;
input n179;
input n185;
input n204;
input n210;
input n670;
input n682;
input n697;
input n704;
input n708;
input n713;
input n718;
input n724;
input n730;
input n735;
input n757;
input n768;
input n783;
input n794;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n20;
wire n23;
wire n25;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n123;
wire n124;
wire n125;
wire n126;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n705;
wire n706;
wire n707;
wire n709;
wire n710;
wire n711;
wire n712;
wire n714;
wire n715;
wire n716;
wire n717;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n731;
wire n732;
wire n733;
wire n734;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
xnor (out,n0,n811);
nor (n0,n1,n795,n807);
and (n1,n2,n683);
nor (n2,n3,n671);
nor (n3,n4,n670);
nand (n4,n5,n96);
or (n5,n6,n8);
not (n6,n7);
not (n8,n9);
xor (n9,n10,n92);
xor (n10,n11,n89);
xor (n11,n12,n85);
xor (n12,n13,n76);
xor (n13,n14,n72);
xor (n14,n15,n57);
xor (n15,n16,n53);
xor (n16,n17,n28);
xor (n17,n18,n23);
and (n18,n19,n20);
wire s0n20,s1n20,notn20;
or (n20,s0n20,s1n20);
not(notn20,n7);
and (s0n20,notn20,n21);
and (s1n20,n7,n22);
and (n23,n24,n25);
wire s0n25,s1n25,notn25;
or (n25,s0n25,s1n25);
not(notn25,n7);
and (s0n25,notn25,n26);
and (s1n25,n7,n27);
or (n28,n29,n33);
and (n29,n30,n31);
and (n30,n24,n20);
and (n31,n32,n25);
and (n33,n34,n35);
xor (n34,n30,n31);
or (n35,n36,n40);
and (n36,n37,n38);
and (n37,n32,n20);
and (n38,n39,n25);
and (n40,n41,n42);
xor (n41,n37,n38);
or (n42,n43,n47);
and (n43,n44,n45);
and (n44,n39,n20);
and (n45,n46,n25);
and (n47,n48,n49);
xor (n48,n44,n45);
and (n49,n50,n51);
and (n50,n46,n20);
and (n51,n52,n25);
and (n53,n32,n54);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n7);
and (s0n54,notn54,n55);
and (s1n54,n7,n56);
or (n57,n58,n61);
and (n58,n59,n60);
xor (n59,n34,n35);
and (n60,n39,n54);
and (n61,n62,n63);
xor (n62,n59,n60);
or (n63,n64,n67);
and (n64,n65,n66);
xor (n65,n41,n42);
and (n66,n46,n54);
and (n67,n68,n69);
xor (n68,n65,n66);
and (n69,n70,n71);
xor (n70,n48,n49);
and (n71,n52,n54);
and (n72,n39,n73);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n7);
and (s0n73,notn73,n74);
and (s1n73,n7,n75);
or (n76,n77,n80);
and (n77,n78,n79);
xor (n78,n62,n63);
and (n79,n46,n73);
and (n80,n81,n82);
xor (n81,n78,n79);
and (n82,n83,n84);
xor (n83,n68,n69);
and (n84,n52,n73);
and (n85,n46,n86);
wire s0n86,s1n86,notn86;
or (n86,s0n86,s1n86);
not(notn86,n7);
and (s0n86,notn86,n87);
and (s1n86,n7,n88);
and (n89,n90,n91);
xor (n90,n81,n82);
and (n91,n52,n86);
and (n92,n52,n93);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n7);
and (s0n93,notn93,n94);
and (s1n93,n7,n95);
nand (n96,n97,n6);
nand (n97,n98,n669);
or (n98,n99,n337);
not (n99,n100);
nand (n100,n101,n336);
not (n101,n102);
nor (n102,n103,n290);
xor (n103,n104,n250);
xor (n104,n105,n169);
xor (n105,n106,n147);
xor (n106,n107,n136);
nand (n107,n108,n130);
or (n108,n109,n124);
nand (n109,n110,n118);
nor (n110,n111,n116);
and (n111,n112,n93);
not (n112,n113);
wire s0n113,s1n113,notn113;
or (n113,s0n113,s1n113);
not(notn113,n7);
and (s0n113,notn113,n114);
and (s1n113,n7,n115);
and (n116,n113,n117);
not (n117,n93);
nand (n118,n119,n123);
or (n119,n112,n120);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n7);
and (s0n120,notn120,n121);
and (s1n120,n7,n122);
nand (n123,n120,n112);
nor (n124,n125,n128);
and (n125,n126,n127);
not (n126,n120);
and (n128,n120,n129);
not (n129,n127);
or (n130,n110,n131);
nor (n131,n132,n134);
and (n132,n133,n126);
and (n134,n135,n120);
not (n135,n133);
nor (n136,n137,n143);
nand (n137,n120,n138);
not (n138,n139);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n7);
and (s0n139,notn139,1'b0);
and (s1n139,n7,n141);
and (n141,n142,n122);
nor (n143,n144,n146);
and (n144,n139,n145);
not (n145,n19);
and (n146,n138,n19);
nand (n147,n148,n159);
or (n148,n149,n154);
nor (n149,n150,n152);
and (n150,n117,n151);
and (n152,n93,n153);
not (n153,n151);
not (n154,n155);
nand (n155,n156,n158);
or (n156,n157,n73);
not (n157,n86);
nand (n158,n73,n157);
or (n159,n160,n164);
nand (n160,n154,n161);
nand (n161,n162,n163);
or (n162,n157,n93);
nand (n163,n93,n157);
nor (n164,n165,n167);
and (n165,n117,n166);
and (n167,n93,n168);
not (n168,n166);
xor (n169,n170,n226);
xor (n170,n171,n213);
xor (n171,n172,n189);
nand (n172,n173,n182);
or (n173,n174,n177);
not (n174,n175);
nor (n175,n176,n20);
not (n176,n25);
nor (n177,n178,n180);
and (n178,n176,n179);
and (n180,n25,n181);
not (n181,n179);
or (n182,n183,n188);
nor (n183,n184,n186);
and (n184,n176,n185);
and (n186,n25,n187);
not (n187,n185);
not (n188,n20);
nand (n189,n190,n207);
or (n190,n191,n201);
not (n191,n192);
and (n192,n193,n197);
nand (n193,n194,n196);
or (n194,n195,n73);
not (n195,n54);
nand (n196,n73,n195);
not (n197,n198);
nand (n198,n199,n200);
or (n199,n195,n25);
nand (n200,n25,n195);
nor (n201,n202,n205);
and (n202,n203,n204);
not (n203,n73);
and (n205,n73,n206);
not (n206,n204);
or (n207,n208,n197);
nor (n208,n209,n211);
and (n209,n203,n210);
and (n211,n73,n212);
not (n212,n210);
and (n213,n214,n220);
nand (n214,n215,n219);
or (n215,n174,n216);
nor (n216,n217,n218);
and (n217,n176,n210);
and (n218,n25,n212);
or (n219,n177,n188);
nand (n220,n221,n225);
or (n221,n191,n222);
nor (n222,n223,n224);
and (n223,n203,n151);
and (n224,n73,n153);
or (n225,n201,n197);
or (n226,n227,n249);
and (n227,n228,n243);
xor (n228,n229,n238);
nand (n229,n230,n235);
or (n230,n231,n109);
not (n231,n232);
nor (n232,n233,n234);
and (n233,n19,n120);
and (n234,n145,n126);
nand (n235,n236,n237);
not (n236,n124);
not (n237,n110);
nor (n238,n137,n239);
nor (n239,n240,n242);
and (n240,n139,n241);
not (n241,n24);
and (n242,n138,n24);
nand (n243,n244,n248);
or (n244,n160,n245);
nor (n245,n246,n247);
and (n246,n117,n133);
and (n247,n93,n135);
or (n248,n154,n164);
and (n249,n229,n238);
or (n250,n251,n289);
and (n251,n252,n267);
xor (n252,n253,n254);
xor (n253,n214,n220);
and (n254,n255,n261);
nand (n255,n256,n260);
or (n256,n174,n257);
nor (n257,n258,n259);
and (n258,n176,n204);
and (n259,n25,n206);
or (n260,n216,n188);
nand (n261,n262,n266);
or (n262,n191,n263);
nor (n263,n264,n265);
and (n264,n203,n166);
and (n265,n73,n168);
or (n266,n197,n222);
or (n267,n268,n288);
and (n268,n269,n282);
xor (n269,n270,n277);
nand (n270,n271,n276);
or (n271,n272,n109);
not (n272,n273);
nor (n273,n274,n275);
and (n274,n24,n120);
and (n275,n241,n126);
nand (n276,n237,n232);
nor (n277,n137,n278);
nor (n278,n279,n281);
and (n279,n139,n280);
not (n280,n32);
and (n281,n138,n32);
nand (n282,n283,n287);
or (n283,n160,n284);
nor (n284,n285,n286);
and (n285,n117,n127);
and (n286,n93,n129);
or (n287,n154,n245);
and (n288,n270,n277);
and (n289,n253,n254);
or (n290,n291,n335);
and (n291,n292,n295);
xor (n292,n293,n294);
xor (n293,n228,n243);
xor (n294,n252,n267);
or (n295,n296,n334);
and (n296,n297,n312);
xor (n297,n298,n299);
xor (n298,n255,n261);
and (n299,n300,n306);
nand (n300,n301,n305);
or (n301,n174,n302);
nor (n302,n303,n304);
and (n303,n176,n151);
and (n304,n25,n153);
or (n305,n257,n188);
nand (n306,n307,n311);
or (n307,n191,n308);
nor (n308,n309,n310);
and (n309,n203,n133);
and (n310,n73,n135);
or (n311,n263,n197);
or (n312,n313,n333);
and (n313,n314,n327);
xor (n314,n315,n322);
nand (n315,n316,n321);
or (n316,n317,n109);
not (n317,n318);
nor (n318,n319,n320);
and (n319,n32,n120);
and (n320,n280,n126);
nand (n321,n237,n273);
nor (n322,n137,n323);
nor (n323,n324,n326);
and (n324,n139,n325);
not (n325,n39);
and (n326,n138,n39);
nand (n327,n328,n332);
or (n328,n160,n329);
nor (n329,n330,n331);
and (n330,n117,n19);
and (n331,n93,n145);
or (n332,n154,n284);
and (n333,n315,n322);
and (n334,n298,n299);
and (n335,n293,n294);
nand (n336,n103,n290);
not (n337,n338);
nand (n338,n339,n668);
or (n339,n340,n374);
not (n340,n341);
nand (n341,n342,n344);
not (n342,n343);
xor (n343,n292,n295);
not (n344,n345);
or (n345,n346,n373);
and (n346,n347,n350);
xor (n347,n348,n349);
xor (n348,n269,n282);
xor (n349,n297,n312);
and (n350,n351,n352);
xor (n351,n300,n306);
or (n352,n353,n372);
and (n353,n354,n366);
xor (n354,n355,n361);
nand (n355,n356,n360);
or (n356,n357,n109);
nor (n357,n358,n359);
and (n358,n39,n126);
and (n359,n325,n120);
nand (n360,n318,n237);
nor (n361,n137,n362);
nor (n362,n363,n365);
and (n363,n139,n364);
not (n364,n46);
and (n365,n138,n46);
nand (n366,n367,n371);
or (n367,n174,n368);
nor (n368,n369,n370);
and (n369,n176,n166);
and (n370,n25,n168);
or (n371,n302,n188);
and (n372,n355,n361);
and (n373,n348,n349);
not (n374,n375);
nand (n375,n376,n528,n667);
nand (n376,n377,n521);
nand (n377,n378,n520);
or (n378,n379,n509);
nor (n379,n380,n508);
and (n380,n381,n480);
not (n381,n382);
nor (n382,n383,n463);
or (n383,n384,n462);
and (n384,n385,n433);
xor (n385,n386,n420);
or (n386,n387,n419);
and (n387,n388,n410);
xor (n388,n389,n400);
nand (n389,n390,n396);
or (n390,n391,n109);
not (n391,n392);
nand (n392,n393,n394);
or (n393,n126,n52);
or (n394,n120,n395);
not (n395,n52);
or (n396,n110,n397);
nor (n397,n398,n399);
and (n398,n46,n126);
and (n399,n364,n120);
nand (n400,n401,n406);
or (n401,n402,n191);
not (n402,n403);
nand (n403,n404,n405);
or (n404,n73,n241);
or (n405,n203,n24);
nand (n406,n198,n407);
nor (n407,n408,n409);
and (n408,n19,n73);
and (n409,n145,n203);
nand (n410,n411,n415);
or (n411,n160,n412);
nor (n412,n413,n414);
and (n413,n117,n39);
and (n414,n93,n325);
or (n415,n154,n416);
nor (n416,n417,n418);
and (n417,n117,n32);
and (n418,n93,n280);
and (n419,n389,n400);
xor (n420,n421,n430);
xor (n421,n422,n424);
and (n422,n423,n52);
not (n423,n137);
nand (n424,n425,n429);
or (n425,n174,n426);
nor (n426,n427,n428);
and (n427,n135,n25);
and (n428,n133,n176);
or (n429,n368,n188);
nand (n430,n431,n432);
or (n431,n109,n397);
or (n432,n110,n357);
xor (n433,n434,n448);
xor (n434,n435,n442);
nand (n435,n436,n438);
or (n436,n191,n437);
not (n437,n407);
or (n438,n197,n439);
nor (n439,n440,n441);
and (n440,n203,n127);
and (n441,n73,n129);
nand (n442,n443,n444);
or (n443,n160,n416);
or (n444,n154,n445);
nor (n445,n446,n447);
and (n446,n117,n24);
and (n447,n93,n241);
and (n448,n449,n454);
nor (n449,n450,n126);
nor (n450,n451,n453);
and (n451,n117,n452);
nand (n452,n113,n52);
and (n453,n112,n395);
nand (n454,n455,n460);
or (n455,n456,n174);
not (n456,n457);
nor (n457,n458,n459);
and (n458,n127,n25);
and (n459,n129,n176);
nand (n460,n461,n20);
not (n461,n426);
and (n462,n386,n420);
xor (n463,n464,n469);
xor (n464,n465,n466);
xor (n465,n354,n366);
or (n466,n467,n468);
and (n467,n434,n448);
and (n468,n435,n442);
xor (n469,n470,n477);
xor (n470,n471,n474);
nand (n471,n472,n473);
or (n472,n160,n445);
or (n473,n154,n329);
nand (n474,n475,n476);
or (n475,n191,n439);
or (n476,n308,n197);
or (n477,n478,n479);
and (n478,n421,n430);
and (n479,n422,n424);
not (n480,n481);
nand (n481,n482,n483);
xor (n482,n385,n433);
or (n483,n484,n507);
and (n484,n485,n506);
xor (n485,n486,n487);
xor (n486,n449,n454);
or (n487,n488,n505);
and (n488,n489,n498);
xor (n489,n490,n491);
and (n490,n237,n52);
nand (n491,n492,n493);
or (n492,n188,n456);
nand (n493,n494,n175);
not (n494,n495);
nor (n495,n496,n497);
and (n496,n19,n176);
and (n497,n145,n25);
nand (n498,n499,n504);
or (n499,n500,n191);
not (n500,n501);
nor (n501,n502,n503);
and (n502,n32,n73);
and (n503,n203,n280);
nand (n504,n198,n403);
and (n505,n490,n491);
xor (n506,n388,n410);
and (n507,n486,n487);
and (n508,n383,n463);
nor (n509,n510,n517);
xor (n510,n511,n514);
xor (n511,n512,n513);
xor (n512,n314,n327);
xor (n513,n351,n352);
or (n514,n515,n516);
and (n515,n470,n477);
and (n516,n471,n474);
or (n517,n518,n519);
and (n518,n464,n469);
and (n519,n465,n466);
nand (n520,n510,n517);
nand (n521,n522,n524);
not (n522,n523);
xor (n523,n347,n350);
not (n524,n525);
or (n525,n526,n527);
and (n526,n511,n514);
and (n527,n512,n513);
nand (n528,n521,n529,n666);
nor (n529,n530,n663);
nor (n530,n531,n661);
and (n531,n532,n656);
or (n532,n533,n655);
and (n533,n534,n574);
xor (n534,n535,n567);
or (n535,n536,n566);
and (n536,n537,n555);
xor (n537,n538,n544);
nand (n538,n539,n543);
or (n539,n540,n191);
not (n540,n541);
nor (n541,n542,n72);
and (n542,n325,n203);
nand (n543,n198,n501);
nand (n544,n545,n550);
or (n545,n546,n154);
not (n546,n547);
nor (n547,n548,n549);
and (n548,n46,n93);
and (n549,n364,n117);
nand (n550,n551,n552);
not (n551,n160);
nand (n552,n553,n554);
or (n553,n117,n52);
or (n554,n93,n395);
xor (n555,n556,n560);
and (n556,n557,n93);
nand (n557,n558,n559);
or (n558,n73,n91);
or (n559,n86,n52);
nand (n560,n561,n565);
or (n561,n174,n562);
nor (n562,n563,n564);
and (n563,n176,n24);
and (n564,n25,n241);
or (n565,n495,n188);
and (n566,n538,n544);
xor (n567,n568,n573);
xor (n568,n569,n572);
nand (n569,n570,n571);
or (n570,n546,n160);
or (n571,n154,n412);
and (n572,n556,n560);
xor (n573,n489,n498);
or (n574,n575,n654);
and (n575,n576,n595);
xor (n576,n577,n594);
or (n577,n578,n593);
and (n578,n579,n587);
xor (n579,n580,n581);
and (n580,n155,n52);
nand (n581,n582,n586);
or (n582,n583,n191);
not (n583,n584);
nor (n584,n79,n585);
and (n585,n364,n203);
nand (n586,n541,n198);
nand (n587,n588,n592);
or (n588,n174,n589);
not (n589,n590);
nor (n590,n591,n31);
and (n591,n280,n176);
or (n592,n562,n188);
and (n593,n580,n581);
xor (n594,n537,n555);
or (n595,n596,n653);
and (n596,n597,n652);
xor (n597,n598,n611);
nor (n598,n599,n607);
not (n599,n600);
nand (n600,n601,n606);
or (n601,n602,n174);
not (n602,n603);
nand (n603,n604,n605);
or (n604,n325,n25);
nand (n605,n25,n325);
nand (n606,n590,n20);
nand (n607,n608,n73);
nand (n608,n609,n610);
or (n609,n25,n71);
or (n610,n54,n52);
nand (n611,n612,n650);
or (n612,n613,n636);
not (n613,n614);
nand (n614,n615,n635);
or (n615,n616,n625);
nor (n616,n617,n624);
nand (n617,n618,n623);
or (n618,n619,n174);
not (n619,n620);
nand (n620,n621,n622);
or (n621,n364,n25);
nand (n622,n25,n364);
nand (n623,n603,n20);
nor (n624,n197,n395);
nand (n625,n626,n633);
nand (n626,n627,n632);
or (n627,n628,n174);
not (n628,n629);
nand (n629,n630,n631);
or (n630,n176,n52);
or (n631,n25,n395);
nand (n632,n620,n20);
nor (n633,n634,n176);
and (n634,n52,n20);
nand (n635,n617,n624);
not (n636,n637);
nand (n637,n638,n646);
not (n638,n639);
nand (n639,n640,n645);
or (n640,n641,n191);
not (n641,n642);
nand (n642,n643,n644);
or (n643,n203,n52);
or (n644,n73,n395);
nand (n645,n198,n584);
nor (n646,n647,n649);
and (n647,n599,n648);
not (n648,n607);
and (n649,n600,n607);
nand (n650,n651,n639);
not (n651,n646);
xor (n652,n579,n587);
and (n653,n598,n611);
and (n654,n577,n594);
and (n655,n535,n567);
or (n656,n657,n658);
xor (n657,n485,n506);
or (n658,n659,n660);
and (n659,n568,n573);
and (n660,n569,n572);
not (n661,n662);
nand (n662,n657,n658);
nand (n663,n664,n381);
not (n664,n665);
nor (n665,n482,n483);
not (n666,n509);
nand (n667,n523,n525);
nand (n668,n343,n345);
or (n669,n338,n100);
nor (n671,n672,n682);
nand (n672,n673,n676);
or (n673,n6,n674);
not (n674,n675);
xor (n675,n90,n91);
nand (n676,n677,n6);
nand (n677,n678,n681);
or (n678,n679,n374);
not (n679,n680);
nand (n680,n341,n668);
or (n681,n375,n680);
not (n683,n684);
nand (n684,n685,n744,n769);
not (n685,n686);
not (n686,n687);
or (n687,n688,n698,n743);
not (n688,n689);
nand (n689,n690,n697);
and (n690,n691,n6);
nand (n691,n692,n696);
or (n692,n693,n694);
not (n693,n532);
not (n694,n695);
nand (n695,n656,n662);
or (n696,n695,n532);
and (n698,n690,n699);
or (n699,n700,n705,n742);
not (n700,n701);
nand (n701,n702,n704);
and (n702,n703,n6);
xor (n703,n534,n574);
and (n705,n702,n706);
or (n706,n707,n710,n741);
and (n707,n708,n709);
wire s0n709,s1n709,notn709;
or (n709,s0n709,s1n709);
not(notn709,n7);
and (s0n709,notn709,n9);
and (s1n709,n7,1'b0);
and (n710,n709,n711);
or (n711,n712,n715,n740);
and (n712,n713,n714);
wire s0n714,s1n714,notn714;
or (n714,s0n714,s1n714);
not(notn714,n7);
and (s0n714,notn714,n675);
and (s1n714,n7,1'b0);
and (n715,n714,n716);
or (n716,n717,n721,n739);
and (n717,n718,n719);
wire s0n719,s1n719,notn719;
or (n719,s0n719,s1n719);
not(notn719,n7);
and (s0n719,notn719,n720);
and (s1n719,n7,1'b0);
xor (n720,n83,n84);
and (n721,n719,n722);
or (n722,n723,n727,n738);
and (n723,n724,n725);
wire s0n725,s1n725,notn725;
or (n725,s0n725,s1n725);
not(notn725,n7);
and (s0n725,notn725,n726);
and (s1n725,n7,1'b0);
xor (n726,n70,n71);
and (n727,n725,n728);
or (n728,n729,n733,n737);
and (n729,n730,n731);
wire s0n731,s1n731,notn731;
or (n731,s0n731,s1n731);
not(notn731,n7);
and (s0n731,notn731,n732);
and (s1n731,n7,1'b0);
xor (n732,n50,n51);
and (n733,n731,n734);
and (n734,n735,n736);
wire s0n736,s1n736,notn736;
or (n736,s0n736,s1n736);
not(notn736,n7);
and (s0n736,notn736,n634);
and (s1n736,n7,1'b0);
and (n737,n730,n734);
and (n738,n724,n728);
and (n739,n718,n722);
and (n740,n713,n716);
and (n741,n708,n711);
and (n742,n704,n706);
and (n743,n697,n699);
nor (n744,n745,n758);
nor (n745,n746,n757);
nand (n746,n747,n749);
or (n747,n6,n748);
not (n748,n720);
nand (n749,n750,n6);
xnor (n750,n751,n752);
nand (n751,n521,n667);
nand (n752,n753,n520);
or (n753,n509,n754);
not (n754,n755);
nand (n755,n756,n379);
not (n756,n529);
nor (n758,n759,n768);
nand (n759,n760,n762);
or (n760,n6,n761);
not (n761,n726);
nand (n762,n763,n6);
nand (n763,n764,n767);
or (n764,n765,n754);
not (n765,n766);
nand (n766,n666,n520);
or (n767,n755,n766);
nor (n769,n770,n784);
nor (n770,n771,n783);
nand (n771,n772,n774);
or (n772,n6,n773);
not (n773,n732);
nand (n774,n775,n6);
nand (n775,n776,n782);
or (n776,n777,n779);
not (n777,n778);
or (n778,n508,n382);
not (n779,n780);
nand (n780,n781,n481);
or (n781,n530,n665);
or (n782,n780,n778);
nor (n784,n785,n794);
or (n785,n786,n787);
and (n786,n7,n634);
and (n787,n6,n788);
nand (n788,n789,n793);
or (n789,n790,n791);
not (n790,n530);
not (n791,n792);
nor (n792,n480,n665);
or (n793,n792,n530);
and (n795,n2,n796);
not (n796,n797);
nor (n797,n798,n803);
and (n798,n744,n799);
nand (n799,n800,n802);
or (n800,n770,n801);
nand (n801,n785,n794);
nand (n802,n771,n783);
nand (n803,n804,n806);
or (n804,n745,n805);
nand (n805,n759,n768);
nand (n806,n746,n757);
nand (n807,n808,n810);
or (n808,n3,n809);
nand (n809,n672,n682);
nand (n810,n4,n670);
or (n811,n812,n1201,n1232);
and (n812,n670,n813);
wire s0n813,s1n813,notn813;
or (n813,s0n813,s1n813);
not(notn813,n7);
and (s0n813,notn813,n814);
and (s1n813,n7,n9);
xor (n814,n815,n1162);
xor (n815,n816,n1199);
xor (n816,n817,n1157);
xor (n817,n818,n1192);
xor (n818,n819,n1151);
xor (n819,n820,n1180);
xor (n820,n821,n1145);
xor (n821,n822,n1163);
xor (n822,n823,n1139);
xor (n823,n824,n1136);
xor (n824,n825,n1135);
xor (n825,n826,n1105);
xor (n826,n827,n1104);
xor (n827,n828,n1065);
xor (n828,n829,n1064);
xor (n829,n830,n1022);
xor (n830,n831,n1021);
xor (n831,n832,n976);
xor (n832,n833,n975);
xor (n833,n834,n932);
xor (n834,n835,n931);
xor (n835,n836,n886);
xor (n836,n837,n885);
xor (n837,n838,n841);
xor (n838,n839,n840);
and (n839,n185,n20);
and (n840,n179,n25);
or (n841,n842,n845);
and (n842,n843,n844);
and (n843,n179,n20);
and (n844,n210,n25);
and (n845,n846,n847);
xor (n846,n843,n844);
or (n847,n848,n851);
and (n848,n849,n850);
and (n849,n210,n20);
and (n850,n204,n25);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n857);
and (n854,n855,n856);
and (n855,n204,n20);
and (n856,n151,n25);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n863);
and (n860,n861,n862);
and (n861,n151,n20);
and (n862,n166,n25);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n869);
and (n866,n867,n868);
and (n867,n166,n20);
and (n868,n133,n25);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n874);
and (n872,n873,n458);
and (n873,n133,n20);
and (n874,n875,n876);
xor (n875,n873,n458);
or (n876,n877,n880);
and (n877,n878,n879);
and (n878,n127,n20);
and (n879,n19,n25);
and (n880,n881,n882);
xor (n881,n878,n879);
or (n882,n883,n884);
and (n883,n18,n23);
and (n884,n17,n28);
and (n885,n210,n54);
or (n886,n887,n890);
and (n887,n888,n889);
xor (n888,n846,n847);
and (n889,n204,n54);
and (n890,n891,n892);
xor (n891,n888,n889);
or (n892,n893,n896);
and (n893,n894,n895);
xor (n894,n852,n853);
and (n895,n151,n54);
and (n896,n897,n898);
xor (n897,n894,n895);
or (n898,n899,n902);
and (n899,n900,n901);
xor (n900,n858,n859);
and (n901,n166,n54);
and (n902,n903,n904);
xor (n903,n900,n901);
or (n904,n905,n908);
and (n905,n906,n907);
xor (n906,n864,n865);
and (n907,n133,n54);
and (n908,n909,n910);
xor (n909,n906,n907);
or (n910,n911,n914);
and (n911,n912,n913);
xor (n912,n870,n871);
and (n913,n127,n54);
and (n914,n915,n916);
xor (n915,n912,n913);
or (n916,n917,n920);
and (n917,n918,n919);
xor (n918,n875,n876);
and (n919,n19,n54);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
xor (n924,n881,n882);
and (n925,n24,n54);
and (n926,n927,n928);
xor (n927,n924,n925);
or (n928,n929,n930);
and (n929,n16,n53);
and (n930,n15,n57);
and (n931,n204,n73);
or (n932,n933,n936);
and (n933,n934,n935);
xor (n934,n891,n892);
and (n935,n151,n73);
and (n936,n937,n938);
xor (n937,n934,n935);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n897,n898);
and (n941,n166,n73);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n903,n904);
and (n947,n133,n73);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n909,n910);
and (n953,n127,n73);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n959);
and (n957,n958,n408);
xor (n958,n915,n916);
and (n959,n960,n961);
xor (n960,n958,n408);
or (n961,n962,n965);
and (n962,n963,n964);
xor (n963,n921,n922);
and (n964,n24,n73);
and (n965,n966,n967);
xor (n966,n963,n964);
or (n967,n968,n970);
and (n968,n969,n502);
xor (n969,n927,n928);
and (n970,n971,n972);
xor (n971,n969,n502);
or (n972,n973,n974);
and (n973,n14,n72);
and (n974,n13,n76);
and (n975,n151,n86);
or (n976,n977,n980);
and (n977,n978,n979);
xor (n978,n937,n938);
and (n979,n166,n86);
and (n980,n981,n982);
xor (n981,n978,n979);
or (n982,n983,n986);
and (n983,n984,n985);
xor (n984,n943,n944);
and (n985,n133,n86);
and (n986,n987,n988);
xor (n987,n984,n985);
or (n988,n989,n992);
and (n989,n990,n991);
xor (n990,n949,n950);
and (n991,n127,n86);
and (n992,n993,n994);
xor (n993,n990,n991);
or (n994,n995,n998);
and (n995,n996,n997);
xor (n996,n955,n956);
and (n997,n19,n86);
and (n998,n999,n1000);
xor (n999,n996,n997);
or (n1000,n1001,n1004);
and (n1001,n1002,n1003);
xor (n1002,n960,n961);
and (n1003,n24,n86);
and (n1004,n1005,n1006);
xor (n1005,n1002,n1003);
or (n1006,n1007,n1010);
and (n1007,n1008,n1009);
xor (n1008,n966,n967);
and (n1009,n32,n86);
and (n1010,n1011,n1012);
xor (n1011,n1008,n1009);
or (n1012,n1013,n1016);
and (n1013,n1014,n1015);
xor (n1014,n971,n972);
and (n1015,n39,n86);
and (n1016,n1017,n1018);
xor (n1017,n1014,n1015);
or (n1018,n1019,n1020);
and (n1019,n12,n85);
and (n1020,n11,n89);
and (n1021,n166,n93);
or (n1022,n1023,n1026);
and (n1023,n1024,n1025);
xor (n1024,n981,n982);
and (n1025,n133,n93);
and (n1026,n1027,n1028);
xor (n1027,n1024,n1025);
or (n1028,n1029,n1032);
and (n1029,n1030,n1031);
xor (n1030,n987,n988);
and (n1031,n127,n93);
and (n1032,n1033,n1034);
xor (n1033,n1030,n1031);
or (n1034,n1035,n1038);
and (n1035,n1036,n1037);
xor (n1036,n993,n994);
and (n1037,n19,n93);
and (n1038,n1039,n1040);
xor (n1039,n1036,n1037);
or (n1040,n1041,n1044);
and (n1041,n1042,n1043);
xor (n1042,n999,n1000);
and (n1043,n24,n93);
and (n1044,n1045,n1046);
xor (n1045,n1042,n1043);
or (n1046,n1047,n1050);
and (n1047,n1048,n1049);
xor (n1048,n1005,n1006);
and (n1049,n32,n93);
and (n1050,n1051,n1052);
xor (n1051,n1048,n1049);
or (n1052,n1053,n1056);
and (n1053,n1054,n1055);
xor (n1054,n1011,n1012);
and (n1055,n39,n93);
and (n1056,n1057,n1058);
xor (n1057,n1054,n1055);
or (n1058,n1059,n1061);
and (n1059,n1060,n548);
xor (n1060,n1017,n1018);
and (n1061,n1062,n1063);
xor (n1062,n1060,n548);
and (n1063,n10,n92);
and (n1064,n133,n113);
or (n1065,n1066,n1069);
and (n1066,n1067,n1068);
xor (n1067,n1027,n1028);
and (n1068,n127,n113);
and (n1069,n1070,n1071);
xor (n1070,n1067,n1068);
or (n1071,n1072,n1075);
and (n1072,n1073,n1074);
xor (n1073,n1033,n1034);
and (n1074,n19,n113);
and (n1075,n1076,n1077);
xor (n1076,n1073,n1074);
or (n1077,n1078,n1081);
and (n1078,n1079,n1080);
xor (n1079,n1039,n1040);
and (n1080,n24,n113);
and (n1081,n1082,n1083);
xor (n1082,n1079,n1080);
or (n1083,n1084,n1087);
and (n1084,n1085,n1086);
xor (n1085,n1045,n1046);
and (n1086,n32,n113);
and (n1087,n1088,n1089);
xor (n1088,n1085,n1086);
or (n1089,n1090,n1093);
and (n1090,n1091,n1092);
xor (n1091,n1051,n1052);
and (n1092,n39,n113);
and (n1093,n1094,n1095);
xor (n1094,n1091,n1092);
or (n1095,n1096,n1099);
and (n1096,n1097,n1098);
xor (n1097,n1057,n1058);
and (n1098,n46,n113);
and (n1099,n1100,n1101);
xor (n1100,n1097,n1098);
and (n1101,n1102,n1103);
xor (n1102,n1062,n1063);
not (n1103,n452);
and (n1104,n127,n120);
or (n1105,n1106,n1108);
and (n1106,n1107,n233);
xor (n1107,n1070,n1071);
and (n1108,n1109,n1110);
xor (n1109,n1107,n233);
or (n1110,n1111,n1113);
and (n1111,n1112,n274);
xor (n1112,n1076,n1077);
and (n1113,n1114,n1115);
xor (n1114,n1112,n274);
or (n1115,n1116,n1118);
and (n1116,n1117,n319);
xor (n1117,n1082,n1083);
and (n1118,n1119,n1120);
xor (n1119,n1117,n319);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1088,n1089);
and (n1123,n39,n120);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1094,n1095);
and (n1129,n46,n120);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
and (n1132,n1133,n1134);
xor (n1133,n1100,n1101);
and (n1134,n52,n120);
and (n1135,n19,n139);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1109,n1110);
and (n1139,n24,n139);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1114,n1115);
and (n1145,n32,n139);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1119,n1120);
and (n1151,n39,n139);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1125,n1126);
and (n1157,n46,n139);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
and (n1160,n1161,n1162);
xor (n1161,n1131,n1132);
and (n1162,n52,n139);
or (n1163,n1164,n1166);
and (n1164,n1165,n1145);
xor (n1165,n1141,n1142);
and (n1166,n1167,n1168);
xor (n1167,n1165,n1145);
or (n1168,n1169,n1171);
and (n1169,n1170,n1151);
xor (n1170,n1147,n1148);
and (n1171,n1172,n1173);
xor (n1172,n1170,n1151);
or (n1173,n1174,n1176);
and (n1174,n1175,n1157);
xor (n1175,n1153,n1154);
and (n1176,n1177,n1178);
xor (n1177,n1175,n1157);
and (n1178,n1179,n1162);
xor (n1179,n1159,n1160);
or (n1180,n1181,n1183);
and (n1181,n1182,n1151);
xor (n1182,n1167,n1168);
and (n1183,n1184,n1185);
xor (n1184,n1182,n1151);
or (n1185,n1186,n1188);
and (n1186,n1187,n1157);
xor (n1187,n1172,n1173);
and (n1188,n1189,n1190);
xor (n1189,n1187,n1157);
and (n1190,n1191,n1162);
xor (n1191,n1177,n1178);
or (n1192,n1193,n1195);
and (n1193,n1194,n1157);
xor (n1194,n1184,n1185);
and (n1195,n1196,n1197);
xor (n1196,n1194,n1157);
and (n1197,n1198,n1162);
xor (n1198,n1189,n1190);
and (n1199,n1200,n1162);
xor (n1200,n1196,n1197);
and (n1201,n813,n1202);
or (n1202,n1203,n1206,n1231);
and (n1203,n682,n1204);
wire s0n1204,s1n1204,notn1204;
or (n1204,s0n1204,s1n1204);
not(notn1204,n7);
and (s0n1204,notn1204,n1205);
and (s1n1204,n7,n675);
xor (n1205,n1200,n1162);
and (n1206,n1204,n1207);
or (n1207,n1208,n1211,n1230);
and (n1208,n757,n1209);
wire s0n1209,s1n1209,notn1209;
or (n1209,s0n1209,s1n1209);
not(notn1209,n7);
and (s0n1209,notn1209,n1210);
and (s1n1209,n7,n720);
xor (n1210,n1198,n1162);
and (n1211,n1209,n1212);
or (n1212,n1213,n1216,n1229);
and (n1213,n768,n1214);
wire s0n1214,s1n1214,notn1214;
or (n1214,s0n1214,s1n1214);
not(notn1214,n7);
and (s0n1214,notn1214,n1215);
and (s1n1214,n7,n726);
xor (n1215,n1191,n1162);
and (n1216,n1214,n1217);
or (n1217,n1218,n1221,n1228);
and (n1218,n783,n1219);
wire s0n1219,s1n1219,notn1219;
or (n1219,s0n1219,s1n1219);
not(notn1219,n7);
and (s0n1219,notn1219,n1220);
and (s1n1219,n7,n732);
xor (n1220,n1179,n1162);
and (n1221,n1219,n1222);
or (n1222,n1223,n1226,n1227);
and (n1223,n794,n1224);
wire s0n1224,s1n1224,notn1224;
or (n1224,s0n1224,s1n1224);
not(notn1224,n7);
and (s0n1224,notn1224,n1225);
and (s1n1224,n7,n634);
xor (n1225,n1161,n1162);
and (n1226,n1224,n687);
and (n1227,n794,n687);
and (n1228,n783,n1222);
and (n1229,n768,n1217);
and (n1230,n757,n1212);
and (n1231,n682,n1207);
and (n1232,n670,n1202);
endmodule
