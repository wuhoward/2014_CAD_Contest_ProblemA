module top (out,n15,n17,n25,n27,n36,n44,n45,n50,n54
        ,n63,n64,n70,n74,n80,n90,n102,n113,n124,n136
        ,n147,n174,n195);
output out;
input n15;
input n17;
input n25;
input n27;
input n36;
input n44;
input n45;
input n50;
input n54;
input n63;
input n64;
input n70;
input n74;
input n80;
input n90;
input n102;
input n113;
input n124;
input n136;
input n147;
input n174;
input n195;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n16;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
xor (out,n0,n458);
nand (n0,n1,n457);
or (n1,n2,n249);
not (n2,n3);
nor (n3,n4,n248);
not (n4,n5);
nand (n5,n6,n211);
xor (n6,n7,n162);
xor (n7,n8,n83);
xor (n8,n9,n57);
xor (n9,n10,n39);
nand (n10,n11,n32);
or (n11,n12,n20);
not (n12,n13);
nand (n13,n14,n18);
or (n14,n15,n16);
not (n16,n17);
or (n18,n19,n17);
not (n19,n15);
not (n20,n21);
and (n21,n22,n29);
not (n22,n23);
nand (n23,n24,n28);
or (n24,n25,n26);
not (n26,n27);
nand (n28,n25,n26);
nand (n29,n30,n31);
or (n30,n25,n19);
nand (n31,n19,n25);
nand (n32,n33,n23);
not (n33,n34);
nor (n34,n35,n37);
and (n35,n19,n36);
and (n37,n15,n38);
not (n38,n36);
nand (n39,n40,n51);
or (n40,n41,n48);
nor (n41,n42,n46);
and (n42,n43,n45);
not (n43,n44);
and (n46,n44,n47);
not (n47,n45);
nand (n48,n44,n49);
not (n49,n50);
or (n51,n52,n49);
nor (n52,n53,n55);
and (n53,n43,n54);
and (n55,n44,n56);
not (n56,n54);
nand (n57,n58,n77);
or (n58,n59,n72);
nand (n59,n60,n67);
nor (n60,n61,n65);
and (n61,n62,n64);
not (n62,n63);
and (n65,n63,n66);
not (n66,n64);
nand (n67,n68,n71);
or (n68,n64,n69);
not (n69,n70);
nand (n71,n69,n64);
nor (n72,n73,n75);
and (n73,n69,n74);
and (n75,n70,n76);
not (n76,n74);
or (n77,n60,n78);
nor (n78,n79,n81);
and (n79,n69,n80);
and (n81,n70,n82);
not (n82,n80);
or (n83,n84,n161);
and (n84,n85,n126);
xor (n85,n86,n94);
nand (n86,n87,n93);
or (n87,n59,n88);
nor (n88,n89,n91);
and (n89,n69,n90);
and (n91,n70,n92);
not (n92,n90);
or (n93,n72,n60);
xor (n94,n95,n103);
and (n95,n96,n15);
nand (n96,n97,n98);
or (n97,n27,n25);
nand (n98,n99,n101);
or (n99,n100,n26);
not (n100,n25);
not (n101,n102);
nand (n103,n104,n119);
or (n104,n105,n109);
not (n105,n106);
nand (n106,n107,n108);
or (n107,n63,n82);
or (n108,n62,n80);
not (n109,n110);
nor (n110,n111,n115);
nand (n111,n112,n114);
or (n112,n43,n113);
nand (n114,n43,n113);
nor (n115,n116,n117);
and (n116,n62,n113);
and (n117,n63,n118);
not (n118,n113);
or (n119,n120,n121);
not (n120,n111);
nor (n121,n122,n125);
and (n122,n123,n63);
not (n123,n124);
and (n125,n124,n62);
or (n126,n127,n160);
and (n127,n128,n142);
xor (n128,n129,n130);
and (n129,n23,n102);
nand (n130,n131,n138);
or (n131,n49,n132);
not (n132,n133);
nor (n133,n134,n137);
and (n134,n135,n43);
not (n135,n136);
and (n137,n44,n136);
or (n138,n139,n48);
nor (n139,n140,n141);
and (n140,n43,n124);
and (n141,n44,n123);
nand (n142,n143,n156);
or (n143,n144,n153);
nand (n144,n145,n149);
nand (n145,n146,n148);
or (n146,n147,n26);
nand (n148,n26,n147);
not (n149,n150);
nand (n150,n151,n152);
or (n151,n69,n147);
nand (n152,n69,n147);
nor (n153,n154,n155);
and (n154,n26,n17);
and (n155,n27,n16);
or (n156,n149,n157);
nor (n157,n158,n159);
and (n158,n38,n27);
and (n159,n36,n26);
and (n160,n129,n130);
and (n161,n86,n94);
xor (n162,n163,n190);
xor (n163,n164,n165);
and (n164,n95,n103);
or (n165,n166,n189);
and (n166,n167,n186);
xor (n167,n168,n179);
nand (n168,n169,n176);
or (n169,n149,n170);
not (n170,n171);
nand (n171,n172,n175);
or (n172,n27,n173);
not (n173,n174);
or (n175,n26,n174);
nand (n176,n177,n178);
not (n177,n157);
not (n178,n144);
nand (n179,n180,n185);
or (n180,n181,n20);
not (n181,n182);
nand (n182,n183,n184);
or (n183,n15,n101);
or (n184,n19,n102);
nand (n185,n13,n23);
nand (n186,n187,n188);
or (n187,n132,n48);
or (n188,n41,n49);
and (n189,n168,n179);
xor (n190,n191,n204);
xor (n191,n192,n198);
nor (n192,n193,n101);
nor (n193,n194,n196);
and (n194,n19,n195);
and (n196,n15,n197);
not (n197,n195);
nand (n198,n199,n200);
or (n199,n121,n109);
nand (n200,n201,n111);
nand (n201,n202,n203);
or (n202,n63,n135);
or (n203,n62,n136);
nand (n204,n205,n206);
or (n205,n170,n144);
nand (n206,n207,n150);
not (n207,n208);
nor (n208,n209,n210);
and (n209,n26,n90);
and (n210,n27,n92);
or (n211,n212,n247);
and (n212,n213,n246);
xor (n213,n214,n215);
xor (n214,n167,n186);
or (n215,n216,n245);
and (n216,n217,n231);
xor (n217,n218,n225);
nand (n218,n219,n224);
or (n219,n220,n109);
not (n220,n221);
nand (n221,n222,n223);
or (n222,n63,n76);
or (n223,n62,n74);
nand (n224,n111,n106);
nand (n225,n226,n230);
or (n226,n59,n227);
nor (n227,n228,n229);
and (n228,n174,n69);
and (n229,n70,n173);
or (n230,n60,n88);
and (n231,n232,n238);
nor (n232,n233,n26);
nor (n233,n234,n236);
and (n234,n235,n101);
nand (n235,n70,n147);
and (n236,n69,n237);
not (n237,n147);
nand (n238,n239,n244);
or (n239,n48,n240);
not (n240,n241);
nor (n241,n242,n243);
and (n242,n44,n80);
and (n243,n82,n43);
or (n244,n139,n49);
and (n245,n218,n225);
xor (n246,n85,n126);
and (n247,n214,n215);
nor (n248,n6,n211);
not (n249,n250);
nor (n250,n251,n449);
and (n251,n252,n432);
or (n252,n253,n431);
and (n253,n254,n322);
xor (n254,n255,n302);
or (n255,n256,n301);
and (n256,n257,n284);
xor (n257,n258,n267);
nand (n258,n259,n263);
or (n259,n59,n260);
nor (n260,n261,n262);
and (n261,n69,n17);
and (n262,n70,n16);
or (n263,n60,n264);
nor (n264,n265,n266);
and (n265,n69,n36);
and (n266,n70,n38);
nor (n267,n268,n279);
not (n268,n269);
nand (n269,n270,n275);
or (n270,n48,n271);
not (n271,n272);
nor (n272,n273,n274);
and (n273,n44,n90);
and (n274,n92,n43);
nand (n275,n276,n50);
nand (n276,n277,n278);
or (n277,n74,n43);
nand (n278,n43,n74);
nand (n279,n280,n70);
nand (n280,n281,n282);
or (n281,n63,n64);
nand (n282,n283,n101);
or (n283,n66,n62);
xor (n284,n285,n291);
xor (n285,n286,n287);
and (n286,n150,n102);
nand (n287,n288,n289);
or (n288,n49,n240);
or (n289,n290,n48);
not (n290,n276);
nand (n291,n292,n297);
or (n292,n293,n109);
not (n293,n294);
nor (n294,n295,n296);
and (n295,n63,n174);
and (n296,n173,n62);
nand (n297,n111,n298);
nand (n298,n299,n300);
or (n299,n63,n92);
or (n300,n62,n90);
and (n301,n258,n267);
xor (n302,n303,n308);
xor (n303,n304,n305);
xor (n304,n232,n238);
or (n305,n306,n307);
and (n306,n285,n291);
and (n307,n286,n287);
xor (n308,n309,n319);
xor (n309,n310,n316);
nand (n310,n311,n315);
or (n311,n144,n312);
nor (n312,n313,n314);
and (n313,n26,n102);
and (n314,n27,n101);
or (n315,n153,n149);
nand (n316,n317,n318);
or (n317,n220,n120);
nand (n318,n110,n298);
nand (n319,n320,n321);
or (n320,n59,n264);
or (n321,n60,n227);
or (n322,n323,n430);
and (n323,n324,n348);
xor (n324,n325,n347);
or (n325,n326,n346);
and (n326,n327,n342);
xor (n327,n328,n335);
nand (n328,n329,n334);
or (n329,n330,n109);
not (n330,n331);
nand (n331,n332,n333);
or (n332,n63,n38);
or (n333,n62,n36);
nand (n334,n111,n294);
nand (n335,n336,n341);
or (n336,n337,n59);
not (n337,n338);
nand (n338,n339,n340);
or (n339,n101,n70);
or (n340,n69,n102);
or (n341,n60,n260);
nand (n342,n343,n345);
or (n343,n344,n268);
not (n344,n279);
or (n345,n269,n279);
and (n346,n328,n335);
xor (n347,n257,n284);
or (n348,n349,n429);
and (n349,n350,n371);
xor (n350,n351,n370);
or (n351,n352,n369);
and (n352,n353,n362);
xor (n353,n354,n355);
nor (n354,n60,n101);
nand (n355,n356,n361);
or (n356,n357,n109);
not (n357,n358);
nor (n358,n359,n360);
and (n359,n16,n62);
and (n360,n63,n17);
nand (n361,n111,n331);
nand (n362,n363,n368);
or (n363,n48,n364);
not (n364,n365);
nor (n365,n366,n367);
and (n366,n173,n43);
and (n367,n44,n174);
or (n368,n271,n49);
and (n369,n354,n355);
xor (n370,n327,n342);
or (n371,n372,n428);
and (n372,n373,n427);
xor (n373,n374,n388);
nor (n374,n375,n383);
not (n375,n376);
nand (n376,n377,n378);
or (n377,n49,n364);
nand (n378,n379,n382);
nor (n379,n380,n381);
and (n380,n38,n43);
and (n381,n44,n36);
not (n382,n48);
nand (n383,n384,n63);
nand (n384,n385,n386);
or (n385,n113,n44);
or (n386,n387,n102);
and (n387,n44,n113);
nand (n388,n389,n426);
or (n389,n390,n414);
not (n390,n391);
nand (n391,n392,n413);
or (n392,n393,n402);
nor (n393,n394,n395);
and (n394,n111,n102);
nand (n395,n396,n398);
or (n396,n49,n397);
not (n397,n379);
nand (n398,n399,n382);
nand (n399,n400,n401);
or (n400,n16,n44);
or (n401,n43,n17);
nand (n402,n403,n406);
not (n403,n404);
nand (n404,n405,n44);
nand (n405,n102,n50);
nand (n406,n407,n409);
or (n407,n49,n408);
not (n408,n399);
nand (n409,n410,n382);
nor (n410,n411,n412);
and (n411,n101,n43);
and (n412,n44,n102);
nand (n413,n394,n395);
not (n414,n415);
nand (n415,n416,n420);
nor (n416,n417,n418);
and (n417,n383,n376);
and (n418,n419,n375);
not (n419,n383);
nor (n420,n421,n425);
and (n421,n110,n422);
nand (n422,n423,n424);
or (n423,n63,n101);
or (n424,n62,n102);
and (n425,n111,n358);
or (n426,n416,n420);
xor (n427,n353,n362);
and (n428,n374,n388);
and (n429,n351,n370);
and (n430,n325,n347);
and (n431,n255,n302);
nor (n432,n433,n444);
nor (n433,n434,n435);
xor (n434,n213,n246);
or (n435,n436,n443);
and (n436,n437,n442);
xor (n437,n438,n441);
or (n438,n439,n440);
and (n439,n309,n319);
and (n440,n310,n316);
xor (n441,n128,n142);
xor (n442,n217,n231);
and (n443,n438,n441);
nor (n444,n445,n446);
xor (n445,n437,n442);
or (n446,n447,n448);
and (n447,n303,n308);
and (n448,n304,n305);
not (n449,n450);
nand (n450,n451,n456);
or (n451,n452,n454);
not (n452,n453);
nand (n453,n445,n446);
not (n454,n455);
nand (n455,n434,n435);
not (n456,n433);
or (n457,n250,n3);
xor (n458,n459,n722);
xor (n459,n460,n719);
xor (n460,n461,n718);
xor (n461,n462,n710);
xor (n462,n463,n709);
xor (n463,n464,n694);
xor (n464,n465,n693);
xor (n465,n466,n673);
xor (n466,n467,n672);
xor (n467,n468,n645);
xor (n468,n469,n644);
xor (n469,n470,n612);
xor (n470,n471,n611);
xor (n471,n472,n574);
xor (n472,n473,n573);
xor (n473,n474,n529);
xor (n474,n475,n528);
xor (n475,n476,n479);
xor (n476,n477,n478);
and (n477,n195,n102);
and (n478,n15,n17);
or (n479,n480,n483);
and (n480,n481,n482);
and (n481,n15,n102);
and (n482,n25,n17);
and (n483,n484,n485);
xor (n484,n481,n482);
or (n485,n486,n489);
and (n486,n487,n488);
and (n487,n25,n102);
and (n488,n27,n17);
and (n489,n490,n491);
xor (n490,n487,n488);
or (n491,n492,n495);
and (n492,n493,n494);
and (n493,n27,n102);
and (n494,n147,n17);
and (n495,n496,n497);
xor (n496,n493,n494);
or (n497,n498,n501);
and (n498,n499,n500);
and (n499,n147,n102);
and (n500,n70,n17);
and (n501,n502,n503);
xor (n502,n499,n500);
or (n503,n504,n507);
and (n504,n505,n506);
and (n505,n70,n102);
and (n506,n64,n17);
and (n507,n508,n509);
xor (n508,n505,n506);
or (n509,n510,n512);
and (n510,n511,n360);
and (n511,n64,n102);
and (n512,n513,n514);
xor (n513,n511,n360);
or (n514,n515,n518);
and (n515,n516,n517);
and (n516,n63,n102);
and (n517,n113,n17);
and (n518,n519,n520);
xor (n519,n516,n517);
or (n520,n521,n524);
and (n521,n522,n523);
and (n522,n113,n102);
and (n523,n44,n17);
and (n524,n525,n526);
xor (n525,n522,n523);
and (n526,n412,n527);
and (n527,n50,n17);
and (n528,n25,n36);
or (n529,n530,n533);
and (n530,n531,n532);
xor (n531,n484,n485);
and (n532,n27,n36);
and (n533,n534,n535);
xor (n534,n531,n532);
or (n535,n536,n539);
and (n536,n537,n538);
xor (n537,n490,n491);
and (n538,n147,n36);
and (n539,n540,n541);
xor (n540,n537,n538);
or (n541,n542,n545);
and (n542,n543,n544);
xor (n543,n496,n497);
and (n544,n70,n36);
and (n545,n546,n547);
xor (n546,n543,n544);
or (n547,n548,n551);
and (n548,n549,n550);
xor (n549,n502,n503);
and (n550,n64,n36);
and (n551,n552,n553);
xor (n552,n549,n550);
or (n553,n554,n557);
and (n554,n555,n556);
xor (n555,n508,n509);
and (n556,n63,n36);
and (n557,n558,n559);
xor (n558,n555,n556);
or (n559,n560,n563);
and (n560,n561,n562);
xor (n561,n513,n514);
and (n562,n113,n36);
and (n563,n564,n565);
xor (n564,n561,n562);
or (n565,n566,n568);
and (n566,n567,n381);
xor (n567,n519,n520);
and (n568,n569,n570);
xor (n569,n567,n381);
and (n570,n571,n572);
xor (n571,n525,n526);
and (n572,n50,n36);
and (n573,n27,n174);
or (n574,n575,n578);
and (n575,n576,n577);
xor (n576,n534,n535);
and (n577,n147,n174);
and (n578,n579,n580);
xor (n579,n576,n577);
or (n580,n581,n584);
and (n581,n582,n583);
xor (n582,n540,n541);
and (n583,n70,n174);
and (n584,n585,n586);
xor (n585,n582,n583);
or (n586,n587,n590);
and (n587,n588,n589);
xor (n588,n546,n547);
and (n589,n64,n174);
and (n590,n591,n592);
xor (n591,n588,n589);
or (n592,n593,n595);
and (n593,n594,n295);
xor (n594,n552,n553);
and (n595,n596,n597);
xor (n596,n594,n295);
or (n597,n598,n601);
and (n598,n599,n600);
xor (n599,n558,n559);
and (n600,n113,n174);
and (n601,n602,n603);
xor (n602,n599,n600);
or (n603,n604,n606);
and (n604,n605,n367);
xor (n605,n564,n565);
and (n606,n607,n608);
xor (n607,n605,n367);
and (n608,n609,n610);
xor (n609,n569,n570);
and (n610,n50,n174);
and (n611,n147,n90);
or (n612,n613,n616);
and (n613,n614,n615);
xor (n614,n579,n580);
and (n615,n70,n90);
and (n616,n617,n618);
xor (n617,n614,n615);
or (n618,n619,n622);
and (n619,n620,n621);
xor (n620,n585,n586);
and (n621,n64,n90);
and (n622,n623,n624);
xor (n623,n620,n621);
or (n624,n625,n628);
and (n625,n626,n627);
xor (n626,n591,n592);
and (n627,n63,n90);
and (n628,n629,n630);
xor (n629,n626,n627);
or (n630,n631,n634);
and (n631,n632,n633);
xor (n632,n596,n597);
and (n633,n113,n90);
and (n634,n635,n636);
xor (n635,n632,n633);
or (n636,n637,n639);
and (n637,n638,n273);
xor (n638,n602,n603);
and (n639,n640,n641);
xor (n640,n638,n273);
and (n641,n642,n643);
xor (n642,n607,n608);
and (n643,n50,n90);
and (n644,n70,n74);
or (n645,n646,n649);
and (n646,n647,n648);
xor (n647,n617,n618);
and (n648,n64,n74);
and (n649,n650,n651);
xor (n650,n647,n648);
or (n651,n652,n655);
and (n652,n653,n654);
xor (n653,n623,n624);
and (n654,n63,n74);
and (n655,n656,n657);
xor (n656,n653,n654);
or (n657,n658,n661);
and (n658,n659,n660);
xor (n659,n629,n630);
and (n660,n113,n74);
and (n661,n662,n663);
xor (n662,n659,n660);
or (n663,n664,n667);
and (n664,n665,n666);
xor (n665,n635,n636);
and (n666,n44,n74);
and (n667,n668,n669);
xor (n668,n665,n666);
and (n669,n670,n671);
xor (n670,n640,n641);
and (n671,n50,n74);
and (n672,n64,n80);
or (n673,n674,n677);
and (n674,n675,n676);
xor (n675,n650,n651);
and (n676,n63,n80);
and (n677,n678,n679);
xor (n678,n675,n676);
or (n679,n680,n683);
and (n680,n681,n682);
xor (n681,n656,n657);
and (n682,n113,n80);
and (n683,n684,n685);
xor (n684,n681,n682);
or (n685,n686,n688);
and (n686,n687,n242);
xor (n687,n662,n663);
and (n688,n689,n690);
xor (n689,n687,n242);
and (n690,n691,n692);
xor (n691,n668,n669);
and (n692,n50,n80);
and (n693,n63,n124);
or (n694,n695,n698);
and (n695,n696,n697);
xor (n696,n678,n679);
and (n697,n113,n124);
and (n698,n699,n700);
xor (n699,n696,n697);
or (n700,n701,n704);
and (n701,n702,n703);
xor (n702,n684,n685);
and (n703,n44,n124);
and (n704,n705,n706);
xor (n705,n702,n703);
and (n706,n707,n708);
xor (n707,n689,n690);
and (n708,n50,n124);
and (n709,n113,n136);
or (n710,n711,n713);
and (n711,n712,n137);
xor (n712,n699,n700);
and (n713,n714,n715);
xor (n714,n712,n137);
and (n715,n716,n717);
xor (n716,n705,n706);
and (n717,n50,n136);
and (n718,n44,n45);
and (n719,n720,n721);
xor (n720,n714,n715);
and (n721,n50,n45);
and (n722,n50,n54);
endmodule
